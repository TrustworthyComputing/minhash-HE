module min_hash(
  input wire [1439:0] set1,
  input wire [1439:0] set2,
  output wire [2887:0] out
);
  wire [15:0] set1_unflattened[90];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  assign set1_unflattened[50] = set1[815:800];
  assign set1_unflattened[51] = set1[831:816];
  assign set1_unflattened[52] = set1[847:832];
  assign set1_unflattened[53] = set1[863:848];
  assign set1_unflattened[54] = set1[879:864];
  assign set1_unflattened[55] = set1[895:880];
  assign set1_unflattened[56] = set1[911:896];
  assign set1_unflattened[57] = set1[927:912];
  assign set1_unflattened[58] = set1[943:928];
  assign set1_unflattened[59] = set1[959:944];
  assign set1_unflattened[60] = set1[975:960];
  assign set1_unflattened[61] = set1[991:976];
  assign set1_unflattened[62] = set1[1007:992];
  assign set1_unflattened[63] = set1[1023:1008];
  assign set1_unflattened[64] = set1[1039:1024];
  assign set1_unflattened[65] = set1[1055:1040];
  assign set1_unflattened[66] = set1[1071:1056];
  assign set1_unflattened[67] = set1[1087:1072];
  assign set1_unflattened[68] = set1[1103:1088];
  assign set1_unflattened[69] = set1[1119:1104];
  assign set1_unflattened[70] = set1[1135:1120];
  assign set1_unflattened[71] = set1[1151:1136];
  assign set1_unflattened[72] = set1[1167:1152];
  assign set1_unflattened[73] = set1[1183:1168];
  assign set1_unflattened[74] = set1[1199:1184];
  assign set1_unflattened[75] = set1[1215:1200];
  assign set1_unflattened[76] = set1[1231:1216];
  assign set1_unflattened[77] = set1[1247:1232];
  assign set1_unflattened[78] = set1[1263:1248];
  assign set1_unflattened[79] = set1[1279:1264];
  assign set1_unflattened[80] = set1[1295:1280];
  assign set1_unflattened[81] = set1[1311:1296];
  assign set1_unflattened[82] = set1[1327:1312];
  assign set1_unflattened[83] = set1[1343:1328];
  assign set1_unflattened[84] = set1[1359:1344];
  assign set1_unflattened[85] = set1[1375:1360];
  assign set1_unflattened[86] = set1[1391:1376];
  assign set1_unflattened[87] = set1[1407:1392];
  assign set1_unflattened[88] = set1[1423:1408];
  assign set1_unflattened[89] = set1[1439:1424];
  wire [15:0] set2_unflattened[90];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  assign set2_unflattened[50] = set2[815:800];
  assign set2_unflattened[51] = set2[831:816];
  assign set2_unflattened[52] = set2[847:832];
  assign set2_unflattened[53] = set2[863:848];
  assign set2_unflattened[54] = set2[879:864];
  assign set2_unflattened[55] = set2[895:880];
  assign set2_unflattened[56] = set2[911:896];
  assign set2_unflattened[57] = set2[927:912];
  assign set2_unflattened[58] = set2[943:928];
  assign set2_unflattened[59] = set2[959:944];
  assign set2_unflattened[60] = set2[975:960];
  assign set2_unflattened[61] = set2[991:976];
  assign set2_unflattened[62] = set2[1007:992];
  assign set2_unflattened[63] = set2[1023:1008];
  assign set2_unflattened[64] = set2[1039:1024];
  assign set2_unflattened[65] = set2[1055:1040];
  assign set2_unflattened[66] = set2[1071:1056];
  assign set2_unflattened[67] = set2[1087:1072];
  assign set2_unflattened[68] = set2[1103:1088];
  assign set2_unflattened[69] = set2[1119:1104];
  assign set2_unflattened[70] = set2[1135:1120];
  assign set2_unflattened[71] = set2[1151:1136];
  assign set2_unflattened[72] = set2[1167:1152];
  assign set2_unflattened[73] = set2[1183:1168];
  assign set2_unflattened[74] = set2[1199:1184];
  assign set2_unflattened[75] = set2[1215:1200];
  assign set2_unflattened[76] = set2[1231:1216];
  assign set2_unflattened[77] = set2[1247:1232];
  assign set2_unflattened[78] = set2[1263:1248];
  assign set2_unflattened[79] = set2[1279:1264];
  assign set2_unflattened[80] = set2[1295:1280];
  assign set2_unflattened[81] = set2[1311:1296];
  assign set2_unflattened[82] = set2[1327:1312];
  assign set2_unflattened[83] = set2[1343:1328];
  assign set2_unflattened[84] = set2[1359:1344];
  assign set2_unflattened[85] = set2[1375:1360];
  assign set2_unflattened[86] = set2[1391:1376];
  assign set2_unflattened[87] = set2[1407:1392];
  assign set2_unflattened[88] = set2[1423:1408];
  assign set2_unflattened[89] = set2[1439:1424];
  wire [15:0] array_index_772631;
  wire [15:0] array_index_772632;
  wire [15:0] array_index_772636;
  wire [1:0] concat_772637;
  wire [1:0] add_772640;
  wire [15:0] array_index_772644;
  wire [2:0] concat_772645;
  wire [2:0] add_772648;
  wire [15:0] array_index_772652;
  wire [3:0] concat_772653;
  wire [3:0] add_772656;
  wire [15:0] array_index_772660;
  wire [4:0] concat_772661;
  wire [4:0] add_772664;
  wire [15:0] array_index_772668;
  wire [5:0] concat_772669;
  wire [5:0] add_772672;
  wire [15:0] array_index_772676;
  wire [6:0] concat_772677;
  wire [6:0] add_772680;
  wire [15:0] array_index_772684;
  wire [7:0] concat_772685;
  wire [7:0] add_772689;
  wire [15:0] array_index_772690;
  wire [7:0] sel_772691;
  wire [7:0] add_772695;
  wire [15:0] array_index_772696;
  wire [7:0] sel_772697;
  wire [7:0] add_772701;
  wire [15:0] array_index_772702;
  wire [7:0] sel_772703;
  wire [7:0] add_772707;
  wire [15:0] array_index_772708;
  wire [7:0] sel_772709;
  wire [7:0] add_772713;
  wire [15:0] array_index_772714;
  wire [7:0] sel_772715;
  wire [7:0] add_772719;
  wire [15:0] array_index_772720;
  wire [7:0] sel_772721;
  wire [7:0] add_772725;
  wire [15:0] array_index_772726;
  wire [7:0] sel_772727;
  wire [7:0] add_772731;
  wire [15:0] array_index_772732;
  wire [7:0] sel_772733;
  wire [7:0] add_772737;
  wire [15:0] array_index_772738;
  wire [7:0] sel_772739;
  wire [7:0] add_772743;
  wire [15:0] array_index_772744;
  wire [7:0] sel_772745;
  wire [7:0] add_772749;
  wire [15:0] array_index_772750;
  wire [7:0] sel_772751;
  wire [7:0] add_772755;
  wire [15:0] array_index_772756;
  wire [7:0] sel_772757;
  wire [7:0] add_772761;
  wire [15:0] array_index_772762;
  wire [7:0] sel_772763;
  wire [7:0] add_772767;
  wire [15:0] array_index_772768;
  wire [7:0] sel_772769;
  wire [7:0] add_772773;
  wire [15:0] array_index_772774;
  wire [7:0] sel_772775;
  wire [7:0] add_772779;
  wire [15:0] array_index_772780;
  wire [7:0] sel_772781;
  wire [7:0] add_772785;
  wire [15:0] array_index_772786;
  wire [7:0] sel_772787;
  wire [7:0] add_772791;
  wire [15:0] array_index_772792;
  wire [7:0] sel_772793;
  wire [7:0] add_772797;
  wire [15:0] array_index_772798;
  wire [7:0] sel_772799;
  wire [7:0] add_772803;
  wire [15:0] array_index_772804;
  wire [7:0] sel_772805;
  wire [7:0] add_772809;
  wire [15:0] array_index_772810;
  wire [7:0] sel_772811;
  wire [7:0] add_772815;
  wire [15:0] array_index_772816;
  wire [7:0] sel_772817;
  wire [7:0] add_772821;
  wire [15:0] array_index_772822;
  wire [7:0] sel_772823;
  wire [7:0] add_772827;
  wire [15:0] array_index_772828;
  wire [7:0] sel_772829;
  wire [7:0] add_772833;
  wire [15:0] array_index_772834;
  wire [7:0] sel_772835;
  wire [7:0] add_772839;
  wire [15:0] array_index_772840;
  wire [7:0] sel_772841;
  wire [7:0] add_772845;
  wire [15:0] array_index_772846;
  wire [7:0] sel_772847;
  wire [7:0] add_772851;
  wire [15:0] array_index_772852;
  wire [7:0] sel_772853;
  wire [7:0] add_772857;
  wire [15:0] array_index_772858;
  wire [7:0] sel_772859;
  wire [7:0] add_772863;
  wire [15:0] array_index_772864;
  wire [7:0] sel_772865;
  wire [7:0] add_772869;
  wire [15:0] array_index_772870;
  wire [7:0] sel_772871;
  wire [7:0] add_772875;
  wire [15:0] array_index_772876;
  wire [7:0] sel_772877;
  wire [7:0] add_772881;
  wire [15:0] array_index_772882;
  wire [7:0] sel_772883;
  wire [7:0] add_772887;
  wire [15:0] array_index_772888;
  wire [7:0] sel_772889;
  wire [7:0] add_772893;
  wire [15:0] array_index_772894;
  wire [7:0] sel_772895;
  wire [7:0] add_772899;
  wire [15:0] array_index_772900;
  wire [7:0] sel_772901;
  wire [7:0] add_772905;
  wire [15:0] array_index_772906;
  wire [7:0] sel_772907;
  wire [7:0] add_772911;
  wire [15:0] array_index_772912;
  wire [7:0] sel_772913;
  wire [7:0] add_772917;
  wire [15:0] array_index_772918;
  wire [7:0] sel_772919;
  wire [7:0] add_772923;
  wire [15:0] array_index_772924;
  wire [7:0] sel_772925;
  wire [7:0] add_772929;
  wire [15:0] array_index_772930;
  wire [7:0] sel_772931;
  wire [7:0] add_772935;
  wire [15:0] array_index_772936;
  wire [7:0] sel_772937;
  wire [7:0] add_772941;
  wire [15:0] array_index_772942;
  wire [7:0] sel_772943;
  wire [7:0] add_772947;
  wire [15:0] array_index_772948;
  wire [7:0] sel_772949;
  wire [7:0] add_772953;
  wire [15:0] array_index_772954;
  wire [7:0] sel_772955;
  wire [7:0] add_772959;
  wire [15:0] array_index_772960;
  wire [7:0] sel_772961;
  wire [7:0] add_772965;
  wire [15:0] array_index_772966;
  wire [7:0] sel_772967;
  wire [7:0] add_772971;
  wire [15:0] array_index_772972;
  wire [7:0] sel_772973;
  wire [7:0] add_772977;
  wire [15:0] array_index_772978;
  wire [7:0] sel_772979;
  wire [7:0] add_772983;
  wire [15:0] array_index_772984;
  wire [7:0] sel_772985;
  wire [7:0] add_772989;
  wire [15:0] array_index_772990;
  wire [7:0] sel_772991;
  wire [7:0] add_772995;
  wire [15:0] array_index_772996;
  wire [7:0] sel_772997;
  wire [7:0] add_773001;
  wire [15:0] array_index_773002;
  wire [7:0] sel_773003;
  wire [7:0] add_773007;
  wire [15:0] array_index_773008;
  wire [7:0] sel_773009;
  wire [7:0] add_773013;
  wire [15:0] array_index_773014;
  wire [7:0] sel_773015;
  wire [7:0] add_773019;
  wire [15:0] array_index_773020;
  wire [7:0] sel_773021;
  wire [7:0] add_773025;
  wire [15:0] array_index_773026;
  wire [7:0] sel_773027;
  wire [7:0] add_773031;
  wire [15:0] array_index_773032;
  wire [7:0] sel_773033;
  wire [7:0] add_773037;
  wire [15:0] array_index_773038;
  wire [7:0] sel_773039;
  wire [7:0] add_773043;
  wire [15:0] array_index_773044;
  wire [7:0] sel_773045;
  wire [7:0] add_773049;
  wire [15:0] array_index_773050;
  wire [7:0] sel_773051;
  wire [7:0] add_773055;
  wire [15:0] array_index_773056;
  wire [7:0] sel_773057;
  wire [7:0] add_773061;
  wire [15:0] array_index_773062;
  wire [7:0] sel_773063;
  wire [7:0] add_773067;
  wire [15:0] array_index_773068;
  wire [7:0] sel_773069;
  wire [7:0] add_773073;
  wire [15:0] array_index_773074;
  wire [7:0] sel_773075;
  wire [7:0] add_773079;
  wire [15:0] array_index_773080;
  wire [7:0] sel_773081;
  wire [7:0] add_773085;
  wire [15:0] array_index_773086;
  wire [7:0] sel_773087;
  wire [7:0] add_773091;
  wire [15:0] array_index_773092;
  wire [7:0] sel_773093;
  wire [7:0] add_773097;
  wire [15:0] array_index_773098;
  wire [7:0] sel_773099;
  wire [7:0] add_773103;
  wire [15:0] array_index_773104;
  wire [7:0] sel_773105;
  wire [7:0] add_773109;
  wire [15:0] array_index_773110;
  wire [7:0] sel_773111;
  wire [7:0] add_773115;
  wire [15:0] array_index_773116;
  wire [7:0] sel_773117;
  wire [7:0] add_773121;
  wire [15:0] array_index_773122;
  wire [7:0] sel_773123;
  wire [7:0] add_773127;
  wire [15:0] array_index_773128;
  wire [7:0] sel_773129;
  wire [7:0] add_773133;
  wire [15:0] array_index_773134;
  wire [7:0] sel_773135;
  wire [7:0] add_773139;
  wire [15:0] array_index_773140;
  wire [7:0] sel_773141;
  wire [7:0] add_773145;
  wire [15:0] array_index_773146;
  wire [7:0] sel_773147;
  wire [7:0] add_773151;
  wire [15:0] array_index_773152;
  wire [7:0] sel_773153;
  wire [7:0] add_773157;
  wire [15:0] array_index_773158;
  wire [7:0] sel_773159;
  wire [7:0] add_773163;
  wire [15:0] array_index_773164;
  wire [7:0] sel_773165;
  wire [7:0] add_773169;
  wire [15:0] array_index_773170;
  wire [7:0] sel_773171;
  wire [7:0] add_773175;
  wire [15:0] array_index_773176;
  wire [7:0] sel_773177;
  wire [7:0] add_773181;
  wire [15:0] array_index_773182;
  wire [7:0] sel_773183;
  wire [7:0] add_773186;
  wire [7:0] sel_773187;
  wire [7:0] add_773190;
  wire [7:0] sel_773191;
  wire [7:0] add_773194;
  wire [7:0] sel_773195;
  wire [7:0] add_773198;
  wire [7:0] sel_773199;
  wire [7:0] add_773202;
  wire [7:0] sel_773203;
  wire [7:0] add_773206;
  wire [7:0] sel_773207;
  wire [7:0] add_773210;
  wire [7:0] sel_773211;
  wire [7:0] add_773214;
  wire [7:0] sel_773215;
  wire [7:0] add_773218;
  wire [7:0] sel_773219;
  wire [7:0] add_773222;
  wire [7:0] sel_773223;
  wire [7:0] add_773226;
  wire [7:0] sel_773227;
  wire [7:0] add_773230;
  wire [7:0] sel_773231;
  wire [7:0] add_773234;
  wire [7:0] sel_773235;
  wire [7:0] add_773238;
  wire [7:0] sel_773239;
  wire [7:0] add_773242;
  wire [7:0] sel_773243;
  wire [7:0] add_773246;
  wire [7:0] sel_773247;
  wire [7:0] add_773250;
  wire [7:0] sel_773251;
  wire [7:0] add_773254;
  wire [7:0] sel_773255;
  wire [7:0] add_773258;
  wire [7:0] sel_773259;
  wire [7:0] add_773262;
  wire [7:0] sel_773263;
  wire [7:0] add_773266;
  wire [7:0] sel_773267;
  wire [7:0] add_773270;
  wire [7:0] sel_773271;
  wire [7:0] add_773274;
  wire [7:0] sel_773275;
  wire [7:0] add_773278;
  wire [7:0] sel_773279;
  wire [7:0] add_773282;
  wire [7:0] sel_773283;
  wire [7:0] add_773286;
  wire [7:0] sel_773287;
  wire [7:0] add_773290;
  wire [7:0] sel_773291;
  wire [7:0] add_773294;
  wire [7:0] sel_773295;
  wire [7:0] add_773298;
  wire [7:0] sel_773299;
  wire [7:0] add_773302;
  wire [7:0] sel_773303;
  wire [7:0] add_773306;
  wire [7:0] sel_773307;
  wire [7:0] add_773310;
  wire [7:0] sel_773311;
  wire [7:0] add_773314;
  wire [7:0] sel_773315;
  wire [7:0] add_773318;
  wire [7:0] sel_773319;
  wire [7:0] add_773322;
  wire [7:0] sel_773323;
  wire [7:0] add_773326;
  wire [7:0] sel_773327;
  wire [7:0] add_773330;
  wire [7:0] sel_773331;
  wire [7:0] add_773334;
  wire [7:0] sel_773335;
  wire [7:0] add_773338;
  wire [7:0] sel_773339;
  wire [7:0] add_773342;
  wire [7:0] sel_773343;
  wire [7:0] add_773346;
  wire [7:0] sel_773347;
  wire [7:0] add_773350;
  wire [7:0] sel_773351;
  wire [7:0] add_773354;
  wire [7:0] sel_773355;
  wire [7:0] add_773358;
  wire [7:0] sel_773359;
  wire [7:0] add_773362;
  wire [7:0] sel_773363;
  wire [7:0] add_773366;
  wire [7:0] sel_773367;
  wire [7:0] add_773370;
  wire [7:0] sel_773371;
  wire [7:0] add_773374;
  wire [7:0] sel_773375;
  wire [7:0] add_773378;
  wire [7:0] sel_773379;
  wire [7:0] add_773382;
  wire [7:0] sel_773383;
  wire [7:0] add_773386;
  wire [7:0] sel_773387;
  wire [7:0] add_773390;
  wire [7:0] sel_773391;
  wire [7:0] add_773394;
  wire [7:0] sel_773395;
  wire [7:0] add_773398;
  wire [7:0] sel_773399;
  wire [7:0] add_773402;
  wire [7:0] sel_773403;
  wire [7:0] add_773406;
  wire [7:0] sel_773407;
  wire [7:0] add_773410;
  wire [7:0] sel_773411;
  wire [7:0] add_773414;
  wire [7:0] sel_773415;
  wire [7:0] add_773418;
  wire [7:0] sel_773419;
  wire [7:0] add_773422;
  wire [7:0] sel_773423;
  wire [7:0] add_773426;
  wire [7:0] sel_773427;
  wire [7:0] add_773430;
  wire [7:0] sel_773431;
  wire [7:0] add_773434;
  wire [7:0] sel_773435;
  wire [7:0] add_773438;
  wire [7:0] sel_773439;
  wire [7:0] add_773442;
  wire [7:0] sel_773443;
  wire [7:0] add_773446;
  wire [7:0] sel_773447;
  wire [7:0] add_773450;
  wire [7:0] sel_773451;
  wire [7:0] add_773454;
  wire [7:0] sel_773455;
  wire [7:0] add_773458;
  wire [7:0] sel_773459;
  wire [7:0] add_773462;
  wire [7:0] sel_773463;
  wire [7:0] add_773466;
  wire [7:0] sel_773467;
  wire [7:0] add_773470;
  wire [7:0] sel_773471;
  wire [7:0] add_773474;
  wire [7:0] sel_773475;
  wire [7:0] add_773478;
  wire [7:0] sel_773479;
  wire [7:0] add_773482;
  wire [7:0] sel_773483;
  wire [7:0] add_773486;
  wire [7:0] sel_773487;
  wire [7:0] add_773490;
  wire [7:0] sel_773491;
  wire [7:0] add_773494;
  wire [7:0] sel_773495;
  wire [7:0] add_773498;
  wire [7:0] sel_773499;
  wire [7:0] add_773502;
  wire [7:0] sel_773503;
  wire [7:0] add_773506;
  wire [7:0] sel_773507;
  wire [7:0] add_773510;
  wire [7:0] sel_773511;
  wire [7:0] add_773514;
  wire [7:0] sel_773515;
  wire [7:0] add_773518;
  wire [7:0] sel_773519;
  wire [7:0] add_773522;
  wire [7:0] sel_773523;
  wire [7:0] add_773526;
  wire [7:0] sel_773527;
  wire [7:0] add_773530;
  wire [7:0] sel_773531;
  wire [7:0] add_773534;
  wire [7:0] sel_773535;
  wire [7:0] add_773538;
  wire [7:0] sel_773539;
  wire [7:0] add_773543;
  wire [15:0] array_index_773544;
  wire [7:0] sel_773545;
  wire [7:0] add_773548;
  wire [7:0] sel_773549;
  wire [7:0] add_773552;
  wire [7:0] sel_773553;
  wire [7:0] add_773556;
  wire [7:0] sel_773557;
  wire [7:0] add_773560;
  wire [7:0] sel_773561;
  wire [7:0] add_773564;
  wire [7:0] sel_773565;
  wire [7:0] add_773568;
  wire [7:0] sel_773569;
  wire [7:0] add_773572;
  wire [7:0] sel_773573;
  wire [7:0] add_773576;
  wire [7:0] sel_773577;
  wire [7:0] add_773580;
  wire [7:0] sel_773581;
  wire [7:0] add_773584;
  wire [7:0] sel_773585;
  wire [7:0] add_773588;
  wire [7:0] sel_773589;
  wire [7:0] add_773592;
  wire [7:0] sel_773593;
  wire [7:0] add_773596;
  wire [7:0] sel_773597;
  wire [7:0] add_773600;
  wire [7:0] sel_773601;
  wire [7:0] add_773604;
  wire [7:0] sel_773605;
  wire [7:0] add_773608;
  wire [7:0] sel_773609;
  wire [7:0] add_773612;
  wire [7:0] sel_773613;
  wire [7:0] add_773616;
  wire [7:0] sel_773617;
  wire [7:0] add_773620;
  wire [7:0] sel_773621;
  wire [7:0] add_773624;
  wire [7:0] sel_773625;
  wire [7:0] add_773628;
  wire [7:0] sel_773629;
  wire [7:0] add_773632;
  wire [7:0] sel_773633;
  wire [7:0] add_773636;
  wire [7:0] sel_773637;
  wire [7:0] add_773640;
  wire [7:0] sel_773641;
  wire [7:0] add_773644;
  wire [7:0] sel_773645;
  wire [7:0] add_773648;
  wire [7:0] sel_773649;
  wire [7:0] add_773652;
  wire [7:0] sel_773653;
  wire [7:0] add_773656;
  wire [7:0] sel_773657;
  wire [7:0] add_773660;
  wire [7:0] sel_773661;
  wire [7:0] add_773664;
  wire [7:0] sel_773665;
  wire [7:0] add_773668;
  wire [7:0] sel_773669;
  wire [7:0] add_773672;
  wire [7:0] sel_773673;
  wire [7:0] add_773676;
  wire [7:0] sel_773677;
  wire [7:0] add_773680;
  wire [7:0] sel_773681;
  wire [7:0] add_773684;
  wire [7:0] sel_773685;
  wire [7:0] add_773688;
  wire [7:0] sel_773689;
  wire [7:0] add_773692;
  wire [7:0] sel_773693;
  wire [7:0] add_773696;
  wire [7:0] sel_773697;
  wire [7:0] add_773700;
  wire [7:0] sel_773701;
  wire [7:0] add_773704;
  wire [7:0] sel_773705;
  wire [7:0] add_773708;
  wire [7:0] sel_773709;
  wire [7:0] add_773712;
  wire [7:0] sel_773713;
  wire [7:0] add_773716;
  wire [7:0] sel_773717;
  wire [7:0] add_773720;
  wire [7:0] sel_773721;
  wire [7:0] add_773724;
  wire [7:0] sel_773725;
  wire [7:0] add_773728;
  wire [7:0] sel_773729;
  wire [7:0] add_773732;
  wire [7:0] sel_773733;
  wire [7:0] add_773736;
  wire [7:0] sel_773737;
  wire [7:0] add_773740;
  wire [7:0] sel_773741;
  wire [7:0] add_773744;
  wire [7:0] sel_773745;
  wire [7:0] add_773748;
  wire [7:0] sel_773749;
  wire [7:0] add_773752;
  wire [7:0] sel_773753;
  wire [7:0] add_773756;
  wire [7:0] sel_773757;
  wire [7:0] add_773760;
  wire [7:0] sel_773761;
  wire [7:0] add_773764;
  wire [7:0] sel_773765;
  wire [7:0] add_773768;
  wire [7:0] sel_773769;
  wire [7:0] add_773772;
  wire [7:0] sel_773773;
  wire [7:0] add_773776;
  wire [7:0] sel_773777;
  wire [7:0] add_773780;
  wire [7:0] sel_773781;
  wire [7:0] add_773784;
  wire [7:0] sel_773785;
  wire [7:0] add_773788;
  wire [7:0] sel_773789;
  wire [7:0] add_773792;
  wire [7:0] sel_773793;
  wire [7:0] add_773796;
  wire [7:0] sel_773797;
  wire [7:0] add_773800;
  wire [7:0] sel_773801;
  wire [7:0] add_773804;
  wire [7:0] sel_773805;
  wire [7:0] add_773808;
  wire [7:0] sel_773809;
  wire [7:0] add_773812;
  wire [7:0] sel_773813;
  wire [7:0] add_773816;
  wire [7:0] sel_773817;
  wire [7:0] add_773820;
  wire [7:0] sel_773821;
  wire [7:0] add_773824;
  wire [7:0] sel_773825;
  wire [7:0] add_773828;
  wire [7:0] sel_773829;
  wire [7:0] add_773832;
  wire [7:0] sel_773833;
  wire [7:0] add_773836;
  wire [7:0] sel_773837;
  wire [7:0] add_773840;
  wire [7:0] sel_773841;
  wire [7:0] add_773844;
  wire [7:0] sel_773845;
  wire [7:0] add_773848;
  wire [7:0] sel_773849;
  wire [7:0] add_773852;
  wire [7:0] sel_773853;
  wire [7:0] add_773856;
  wire [7:0] sel_773857;
  wire [7:0] add_773860;
  wire [7:0] sel_773861;
  wire [7:0] add_773864;
  wire [7:0] sel_773865;
  wire [7:0] add_773868;
  wire [7:0] sel_773869;
  wire [7:0] add_773872;
  wire [7:0] sel_773873;
  wire [7:0] add_773876;
  wire [7:0] sel_773877;
  wire [7:0] add_773880;
  wire [7:0] sel_773881;
  wire [7:0] add_773884;
  wire [7:0] sel_773885;
  wire [7:0] add_773888;
  wire [7:0] sel_773889;
  wire [7:0] add_773892;
  wire [7:0] sel_773893;
  wire [7:0] add_773896;
  wire [7:0] sel_773897;
  wire [7:0] add_773900;
  wire [7:0] sel_773901;
  wire [7:0] add_773905;
  wire [15:0] array_index_773906;
  wire [7:0] sel_773907;
  wire [7:0] add_773910;
  wire [7:0] sel_773911;
  wire [7:0] add_773914;
  wire [7:0] sel_773915;
  wire [7:0] add_773918;
  wire [7:0] sel_773919;
  wire [7:0] add_773922;
  wire [7:0] sel_773923;
  wire [7:0] add_773926;
  wire [7:0] sel_773927;
  wire [7:0] add_773930;
  wire [7:0] sel_773931;
  wire [7:0] add_773934;
  wire [7:0] sel_773935;
  wire [7:0] add_773938;
  wire [7:0] sel_773939;
  wire [7:0] add_773942;
  wire [7:0] sel_773943;
  wire [7:0] add_773946;
  wire [7:0] sel_773947;
  wire [7:0] add_773950;
  wire [7:0] sel_773951;
  wire [7:0] add_773954;
  wire [7:0] sel_773955;
  wire [7:0] add_773958;
  wire [7:0] sel_773959;
  wire [7:0] add_773962;
  wire [7:0] sel_773963;
  wire [7:0] add_773966;
  wire [7:0] sel_773967;
  wire [7:0] add_773970;
  wire [7:0] sel_773971;
  wire [7:0] add_773974;
  wire [7:0] sel_773975;
  wire [7:0] add_773978;
  wire [7:0] sel_773979;
  wire [7:0] add_773982;
  wire [7:0] sel_773983;
  wire [7:0] add_773986;
  wire [7:0] sel_773987;
  wire [7:0] add_773990;
  wire [7:0] sel_773991;
  wire [7:0] add_773994;
  wire [7:0] sel_773995;
  wire [7:0] add_773998;
  wire [7:0] sel_773999;
  wire [7:0] add_774002;
  wire [7:0] sel_774003;
  wire [7:0] add_774006;
  wire [7:0] sel_774007;
  wire [7:0] add_774010;
  wire [7:0] sel_774011;
  wire [7:0] add_774014;
  wire [7:0] sel_774015;
  wire [7:0] add_774018;
  wire [7:0] sel_774019;
  wire [7:0] add_774022;
  wire [7:0] sel_774023;
  wire [7:0] add_774026;
  wire [7:0] sel_774027;
  wire [7:0] add_774030;
  wire [7:0] sel_774031;
  wire [7:0] add_774034;
  wire [7:0] sel_774035;
  wire [7:0] add_774038;
  wire [7:0] sel_774039;
  wire [7:0] add_774042;
  wire [7:0] sel_774043;
  wire [7:0] add_774046;
  wire [7:0] sel_774047;
  wire [7:0] add_774050;
  wire [7:0] sel_774051;
  wire [7:0] add_774054;
  wire [7:0] sel_774055;
  wire [7:0] add_774058;
  wire [7:0] sel_774059;
  wire [7:0] add_774062;
  wire [7:0] sel_774063;
  wire [7:0] add_774066;
  wire [7:0] sel_774067;
  wire [7:0] add_774070;
  wire [7:0] sel_774071;
  wire [7:0] add_774074;
  wire [7:0] sel_774075;
  wire [7:0] add_774078;
  wire [7:0] sel_774079;
  wire [7:0] add_774082;
  wire [7:0] sel_774083;
  wire [7:0] add_774086;
  wire [7:0] sel_774087;
  wire [7:0] add_774090;
  wire [7:0] sel_774091;
  wire [7:0] add_774094;
  wire [7:0] sel_774095;
  wire [7:0] add_774098;
  wire [7:0] sel_774099;
  wire [7:0] add_774102;
  wire [7:0] sel_774103;
  wire [7:0] add_774106;
  wire [7:0] sel_774107;
  wire [7:0] add_774110;
  wire [7:0] sel_774111;
  wire [7:0] add_774114;
  wire [7:0] sel_774115;
  wire [7:0] add_774118;
  wire [7:0] sel_774119;
  wire [7:0] add_774122;
  wire [7:0] sel_774123;
  wire [7:0] add_774126;
  wire [7:0] sel_774127;
  wire [7:0] add_774130;
  wire [7:0] sel_774131;
  wire [7:0] add_774134;
  wire [7:0] sel_774135;
  wire [7:0] add_774138;
  wire [7:0] sel_774139;
  wire [7:0] add_774142;
  wire [7:0] sel_774143;
  wire [7:0] add_774146;
  wire [7:0] sel_774147;
  wire [7:0] add_774150;
  wire [7:0] sel_774151;
  wire [7:0] add_774154;
  wire [7:0] sel_774155;
  wire [7:0] add_774158;
  wire [7:0] sel_774159;
  wire [7:0] add_774162;
  wire [7:0] sel_774163;
  wire [7:0] add_774166;
  wire [7:0] sel_774167;
  wire [7:0] add_774170;
  wire [7:0] sel_774171;
  wire [7:0] add_774174;
  wire [7:0] sel_774175;
  wire [7:0] add_774178;
  wire [7:0] sel_774179;
  wire [7:0] add_774182;
  wire [7:0] sel_774183;
  wire [7:0] add_774186;
  wire [7:0] sel_774187;
  wire [7:0] add_774190;
  wire [7:0] sel_774191;
  wire [7:0] add_774194;
  wire [7:0] sel_774195;
  wire [7:0] add_774198;
  wire [7:0] sel_774199;
  wire [7:0] add_774202;
  wire [7:0] sel_774203;
  wire [7:0] add_774206;
  wire [7:0] sel_774207;
  wire [7:0] add_774210;
  wire [7:0] sel_774211;
  wire [7:0] add_774214;
  wire [7:0] sel_774215;
  wire [7:0] add_774218;
  wire [7:0] sel_774219;
  wire [7:0] add_774222;
  wire [7:0] sel_774223;
  wire [7:0] add_774226;
  wire [7:0] sel_774227;
  wire [7:0] add_774230;
  wire [7:0] sel_774231;
  wire [7:0] add_774234;
  wire [7:0] sel_774235;
  wire [7:0] add_774238;
  wire [7:0] sel_774239;
  wire [7:0] add_774242;
  wire [7:0] sel_774243;
  wire [7:0] add_774246;
  wire [7:0] sel_774247;
  wire [7:0] add_774250;
  wire [7:0] sel_774251;
  wire [7:0] add_774254;
  wire [7:0] sel_774255;
  wire [7:0] add_774258;
  wire [7:0] sel_774259;
  wire [7:0] add_774262;
  wire [7:0] sel_774263;
  wire [7:0] add_774267;
  wire [15:0] array_index_774268;
  wire [7:0] sel_774269;
  wire [7:0] add_774272;
  wire [7:0] sel_774273;
  wire [7:0] add_774276;
  wire [7:0] sel_774277;
  wire [7:0] add_774280;
  wire [7:0] sel_774281;
  wire [7:0] add_774284;
  wire [7:0] sel_774285;
  wire [7:0] add_774288;
  wire [7:0] sel_774289;
  wire [7:0] add_774292;
  wire [7:0] sel_774293;
  wire [7:0] add_774296;
  wire [7:0] sel_774297;
  wire [7:0] add_774300;
  wire [7:0] sel_774301;
  wire [7:0] add_774304;
  wire [7:0] sel_774305;
  wire [7:0] add_774308;
  wire [7:0] sel_774309;
  wire [7:0] add_774312;
  wire [7:0] sel_774313;
  wire [7:0] add_774316;
  wire [7:0] sel_774317;
  wire [7:0] add_774320;
  wire [7:0] sel_774321;
  wire [7:0] add_774324;
  wire [7:0] sel_774325;
  wire [7:0] add_774328;
  wire [7:0] sel_774329;
  wire [7:0] add_774332;
  wire [7:0] sel_774333;
  wire [7:0] add_774336;
  wire [7:0] sel_774337;
  wire [7:0] add_774340;
  wire [7:0] sel_774341;
  wire [7:0] add_774344;
  wire [7:0] sel_774345;
  wire [7:0] add_774348;
  wire [7:0] sel_774349;
  wire [7:0] add_774352;
  wire [7:0] sel_774353;
  wire [7:0] add_774356;
  wire [7:0] sel_774357;
  wire [7:0] add_774360;
  wire [7:0] sel_774361;
  wire [7:0] add_774364;
  wire [7:0] sel_774365;
  wire [7:0] add_774368;
  wire [7:0] sel_774369;
  wire [7:0] add_774372;
  wire [7:0] sel_774373;
  wire [7:0] add_774376;
  wire [7:0] sel_774377;
  wire [7:0] add_774380;
  wire [7:0] sel_774381;
  wire [7:0] add_774384;
  wire [7:0] sel_774385;
  wire [7:0] add_774388;
  wire [7:0] sel_774389;
  wire [7:0] add_774392;
  wire [7:0] sel_774393;
  wire [7:0] add_774396;
  wire [7:0] sel_774397;
  wire [7:0] add_774400;
  wire [7:0] sel_774401;
  wire [7:0] add_774404;
  wire [7:0] sel_774405;
  wire [7:0] add_774408;
  wire [7:0] sel_774409;
  wire [7:0] add_774412;
  wire [7:0] sel_774413;
  wire [7:0] add_774416;
  wire [7:0] sel_774417;
  wire [7:0] add_774420;
  wire [7:0] sel_774421;
  wire [7:0] add_774424;
  wire [7:0] sel_774425;
  wire [7:0] add_774428;
  wire [7:0] sel_774429;
  wire [7:0] add_774432;
  wire [7:0] sel_774433;
  wire [7:0] add_774436;
  wire [7:0] sel_774437;
  wire [7:0] add_774440;
  wire [7:0] sel_774441;
  wire [7:0] add_774444;
  wire [7:0] sel_774445;
  wire [7:0] add_774448;
  wire [7:0] sel_774449;
  wire [7:0] add_774452;
  wire [7:0] sel_774453;
  wire [7:0] add_774456;
  wire [7:0] sel_774457;
  wire [7:0] add_774460;
  wire [7:0] sel_774461;
  wire [7:0] add_774464;
  wire [7:0] sel_774465;
  wire [7:0] add_774468;
  wire [7:0] sel_774469;
  wire [7:0] add_774472;
  wire [7:0] sel_774473;
  wire [7:0] add_774476;
  wire [7:0] sel_774477;
  wire [7:0] add_774480;
  wire [7:0] sel_774481;
  wire [7:0] add_774484;
  wire [7:0] sel_774485;
  wire [7:0] add_774488;
  wire [7:0] sel_774489;
  wire [7:0] add_774492;
  wire [7:0] sel_774493;
  wire [7:0] add_774496;
  wire [7:0] sel_774497;
  wire [7:0] add_774500;
  wire [7:0] sel_774501;
  wire [7:0] add_774504;
  wire [7:0] sel_774505;
  wire [7:0] add_774508;
  wire [7:0] sel_774509;
  wire [7:0] add_774512;
  wire [7:0] sel_774513;
  wire [7:0] add_774516;
  wire [7:0] sel_774517;
  wire [7:0] add_774520;
  wire [7:0] sel_774521;
  wire [7:0] add_774524;
  wire [7:0] sel_774525;
  wire [7:0] add_774528;
  wire [7:0] sel_774529;
  wire [7:0] add_774532;
  wire [7:0] sel_774533;
  wire [7:0] add_774536;
  wire [7:0] sel_774537;
  wire [7:0] add_774540;
  wire [7:0] sel_774541;
  wire [7:0] add_774544;
  wire [7:0] sel_774545;
  wire [7:0] add_774548;
  wire [7:0] sel_774549;
  wire [7:0] add_774552;
  wire [7:0] sel_774553;
  wire [7:0] add_774556;
  wire [7:0] sel_774557;
  wire [7:0] add_774560;
  wire [7:0] sel_774561;
  wire [7:0] add_774564;
  wire [7:0] sel_774565;
  wire [7:0] add_774568;
  wire [7:0] sel_774569;
  wire [7:0] add_774572;
  wire [7:0] sel_774573;
  wire [7:0] add_774576;
  wire [7:0] sel_774577;
  wire [7:0] add_774580;
  wire [7:0] sel_774581;
  wire [7:0] add_774584;
  wire [7:0] sel_774585;
  wire [7:0] add_774588;
  wire [7:0] sel_774589;
  wire [7:0] add_774592;
  wire [7:0] sel_774593;
  wire [7:0] add_774596;
  wire [7:0] sel_774597;
  wire [7:0] add_774600;
  wire [7:0] sel_774601;
  wire [7:0] add_774604;
  wire [7:0] sel_774605;
  wire [7:0] add_774608;
  wire [7:0] sel_774609;
  wire [7:0] add_774612;
  wire [7:0] sel_774613;
  wire [7:0] add_774616;
  wire [7:0] sel_774617;
  wire [7:0] add_774620;
  wire [7:0] sel_774621;
  wire [7:0] add_774624;
  wire [7:0] sel_774625;
  wire [7:0] add_774629;
  wire [15:0] array_index_774630;
  wire [7:0] sel_774631;
  wire [7:0] add_774634;
  wire [7:0] sel_774635;
  wire [7:0] add_774638;
  wire [7:0] sel_774639;
  wire [7:0] add_774642;
  wire [7:0] sel_774643;
  wire [7:0] add_774646;
  wire [7:0] sel_774647;
  wire [7:0] add_774650;
  wire [7:0] sel_774651;
  wire [7:0] add_774654;
  wire [7:0] sel_774655;
  wire [7:0] add_774658;
  wire [7:0] sel_774659;
  wire [7:0] add_774662;
  wire [7:0] sel_774663;
  wire [7:0] add_774666;
  wire [7:0] sel_774667;
  wire [7:0] add_774670;
  wire [7:0] sel_774671;
  wire [7:0] add_774674;
  wire [7:0] sel_774675;
  wire [7:0] add_774678;
  wire [7:0] sel_774679;
  wire [7:0] add_774682;
  wire [7:0] sel_774683;
  wire [7:0] add_774686;
  wire [7:0] sel_774687;
  wire [7:0] add_774690;
  wire [7:0] sel_774691;
  wire [7:0] add_774694;
  wire [7:0] sel_774695;
  wire [7:0] add_774698;
  wire [7:0] sel_774699;
  wire [7:0] add_774702;
  wire [7:0] sel_774703;
  wire [7:0] add_774706;
  wire [7:0] sel_774707;
  wire [7:0] add_774710;
  wire [7:0] sel_774711;
  wire [7:0] add_774714;
  wire [7:0] sel_774715;
  wire [7:0] add_774718;
  wire [7:0] sel_774719;
  wire [7:0] add_774722;
  wire [7:0] sel_774723;
  wire [7:0] add_774726;
  wire [7:0] sel_774727;
  wire [7:0] add_774730;
  wire [7:0] sel_774731;
  wire [7:0] add_774734;
  wire [7:0] sel_774735;
  wire [7:0] add_774738;
  wire [7:0] sel_774739;
  wire [7:0] add_774742;
  wire [7:0] sel_774743;
  wire [7:0] add_774746;
  wire [7:0] sel_774747;
  wire [7:0] add_774750;
  wire [7:0] sel_774751;
  wire [7:0] add_774754;
  wire [7:0] sel_774755;
  wire [7:0] add_774758;
  wire [7:0] sel_774759;
  wire [7:0] add_774762;
  wire [7:0] sel_774763;
  wire [7:0] add_774766;
  wire [7:0] sel_774767;
  wire [7:0] add_774770;
  wire [7:0] sel_774771;
  wire [7:0] add_774774;
  wire [7:0] sel_774775;
  wire [7:0] add_774778;
  wire [7:0] sel_774779;
  wire [7:0] add_774782;
  wire [7:0] sel_774783;
  wire [7:0] add_774786;
  wire [7:0] sel_774787;
  wire [7:0] add_774790;
  wire [7:0] sel_774791;
  wire [7:0] add_774794;
  wire [7:0] sel_774795;
  wire [7:0] add_774798;
  wire [7:0] sel_774799;
  wire [7:0] add_774802;
  wire [7:0] sel_774803;
  wire [7:0] add_774806;
  wire [7:0] sel_774807;
  wire [7:0] add_774810;
  wire [7:0] sel_774811;
  wire [7:0] add_774814;
  wire [7:0] sel_774815;
  wire [7:0] add_774818;
  wire [7:0] sel_774819;
  wire [7:0] add_774822;
  wire [7:0] sel_774823;
  wire [7:0] add_774826;
  wire [7:0] sel_774827;
  wire [7:0] add_774830;
  wire [7:0] sel_774831;
  wire [7:0] add_774834;
  wire [7:0] sel_774835;
  wire [7:0] add_774838;
  wire [7:0] sel_774839;
  wire [7:0] add_774842;
  wire [7:0] sel_774843;
  wire [7:0] add_774846;
  wire [7:0] sel_774847;
  wire [7:0] add_774850;
  wire [7:0] sel_774851;
  wire [7:0] add_774854;
  wire [7:0] sel_774855;
  wire [7:0] add_774858;
  wire [7:0] sel_774859;
  wire [7:0] add_774862;
  wire [7:0] sel_774863;
  wire [7:0] add_774866;
  wire [7:0] sel_774867;
  wire [7:0] add_774870;
  wire [7:0] sel_774871;
  wire [7:0] add_774874;
  wire [7:0] sel_774875;
  wire [7:0] add_774878;
  wire [7:0] sel_774879;
  wire [7:0] add_774882;
  wire [7:0] sel_774883;
  wire [7:0] add_774886;
  wire [7:0] sel_774887;
  wire [7:0] add_774890;
  wire [7:0] sel_774891;
  wire [7:0] add_774894;
  wire [7:0] sel_774895;
  wire [7:0] add_774898;
  wire [7:0] sel_774899;
  wire [7:0] add_774902;
  wire [7:0] sel_774903;
  wire [7:0] add_774906;
  wire [7:0] sel_774907;
  wire [7:0] add_774910;
  wire [7:0] sel_774911;
  wire [7:0] add_774914;
  wire [7:0] sel_774915;
  wire [7:0] add_774918;
  wire [7:0] sel_774919;
  wire [7:0] add_774922;
  wire [7:0] sel_774923;
  wire [7:0] add_774926;
  wire [7:0] sel_774927;
  wire [7:0] add_774930;
  wire [7:0] sel_774931;
  wire [7:0] add_774934;
  wire [7:0] sel_774935;
  wire [7:0] add_774938;
  wire [7:0] sel_774939;
  wire [7:0] add_774942;
  wire [7:0] sel_774943;
  wire [7:0] add_774946;
  wire [7:0] sel_774947;
  wire [7:0] add_774950;
  wire [7:0] sel_774951;
  wire [7:0] add_774954;
  wire [7:0] sel_774955;
  wire [7:0] add_774958;
  wire [7:0] sel_774959;
  wire [7:0] add_774962;
  wire [7:0] sel_774963;
  wire [7:0] add_774966;
  wire [7:0] sel_774967;
  wire [7:0] add_774970;
  wire [7:0] sel_774971;
  wire [7:0] add_774974;
  wire [7:0] sel_774975;
  wire [7:0] add_774978;
  wire [7:0] sel_774979;
  wire [7:0] add_774982;
  wire [7:0] sel_774983;
  wire [7:0] add_774986;
  wire [7:0] sel_774987;
  wire [7:0] add_774991;
  wire [15:0] array_index_774992;
  wire [7:0] sel_774993;
  wire [7:0] add_774996;
  wire [7:0] sel_774997;
  wire [7:0] add_775000;
  wire [7:0] sel_775001;
  wire [7:0] add_775004;
  wire [7:0] sel_775005;
  wire [7:0] add_775008;
  wire [7:0] sel_775009;
  wire [7:0] add_775012;
  wire [7:0] sel_775013;
  wire [7:0] add_775016;
  wire [7:0] sel_775017;
  wire [7:0] add_775020;
  wire [7:0] sel_775021;
  wire [7:0] add_775024;
  wire [7:0] sel_775025;
  wire [7:0] add_775028;
  wire [7:0] sel_775029;
  wire [7:0] add_775032;
  wire [7:0] sel_775033;
  wire [7:0] add_775036;
  wire [7:0] sel_775037;
  wire [7:0] add_775040;
  wire [7:0] sel_775041;
  wire [7:0] add_775044;
  wire [7:0] sel_775045;
  wire [7:0] add_775048;
  wire [7:0] sel_775049;
  wire [7:0] add_775052;
  wire [7:0] sel_775053;
  wire [7:0] add_775056;
  wire [7:0] sel_775057;
  wire [7:0] add_775060;
  wire [7:0] sel_775061;
  wire [7:0] add_775064;
  wire [7:0] sel_775065;
  wire [7:0] add_775068;
  wire [7:0] sel_775069;
  wire [7:0] add_775072;
  wire [7:0] sel_775073;
  wire [7:0] add_775076;
  wire [7:0] sel_775077;
  wire [7:0] add_775080;
  wire [7:0] sel_775081;
  wire [7:0] add_775084;
  wire [7:0] sel_775085;
  wire [7:0] add_775088;
  wire [7:0] sel_775089;
  wire [7:0] add_775092;
  wire [7:0] sel_775093;
  wire [7:0] add_775096;
  wire [7:0] sel_775097;
  wire [7:0] add_775100;
  wire [7:0] sel_775101;
  wire [7:0] add_775104;
  wire [7:0] sel_775105;
  wire [7:0] add_775108;
  wire [7:0] sel_775109;
  wire [7:0] add_775112;
  wire [7:0] sel_775113;
  wire [7:0] add_775116;
  wire [7:0] sel_775117;
  wire [7:0] add_775120;
  wire [7:0] sel_775121;
  wire [7:0] add_775124;
  wire [7:0] sel_775125;
  wire [7:0] add_775128;
  wire [7:0] sel_775129;
  wire [7:0] add_775132;
  wire [7:0] sel_775133;
  wire [7:0] add_775136;
  wire [7:0] sel_775137;
  wire [7:0] add_775140;
  wire [7:0] sel_775141;
  wire [7:0] add_775144;
  wire [7:0] sel_775145;
  wire [7:0] add_775148;
  wire [7:0] sel_775149;
  wire [7:0] add_775152;
  wire [7:0] sel_775153;
  wire [7:0] add_775156;
  wire [7:0] sel_775157;
  wire [7:0] add_775160;
  wire [7:0] sel_775161;
  wire [7:0] add_775164;
  wire [7:0] sel_775165;
  wire [7:0] add_775168;
  wire [7:0] sel_775169;
  wire [7:0] add_775172;
  wire [7:0] sel_775173;
  wire [7:0] add_775176;
  wire [7:0] sel_775177;
  wire [7:0] add_775180;
  wire [7:0] sel_775181;
  wire [7:0] add_775184;
  wire [7:0] sel_775185;
  wire [7:0] add_775188;
  wire [7:0] sel_775189;
  wire [7:0] add_775192;
  wire [7:0] sel_775193;
  wire [7:0] add_775196;
  wire [7:0] sel_775197;
  wire [7:0] add_775200;
  wire [7:0] sel_775201;
  wire [7:0] add_775204;
  wire [7:0] sel_775205;
  wire [7:0] add_775208;
  wire [7:0] sel_775209;
  wire [7:0] add_775212;
  wire [7:0] sel_775213;
  wire [7:0] add_775216;
  wire [7:0] sel_775217;
  wire [7:0] add_775220;
  wire [7:0] sel_775221;
  wire [7:0] add_775224;
  wire [7:0] sel_775225;
  wire [7:0] add_775228;
  wire [7:0] sel_775229;
  wire [7:0] add_775232;
  wire [7:0] sel_775233;
  wire [7:0] add_775236;
  wire [7:0] sel_775237;
  wire [7:0] add_775240;
  wire [7:0] sel_775241;
  wire [7:0] add_775244;
  wire [7:0] sel_775245;
  wire [7:0] add_775248;
  wire [7:0] sel_775249;
  wire [7:0] add_775252;
  wire [7:0] sel_775253;
  wire [7:0] add_775256;
  wire [7:0] sel_775257;
  wire [7:0] add_775260;
  wire [7:0] sel_775261;
  wire [7:0] add_775264;
  wire [7:0] sel_775265;
  wire [7:0] add_775268;
  wire [7:0] sel_775269;
  wire [7:0] add_775272;
  wire [7:0] sel_775273;
  wire [7:0] add_775276;
  wire [7:0] sel_775277;
  wire [7:0] add_775280;
  wire [7:0] sel_775281;
  wire [7:0] add_775284;
  wire [7:0] sel_775285;
  wire [7:0] add_775288;
  wire [7:0] sel_775289;
  wire [7:0] add_775292;
  wire [7:0] sel_775293;
  wire [7:0] add_775296;
  wire [7:0] sel_775297;
  wire [7:0] add_775300;
  wire [7:0] sel_775301;
  wire [7:0] add_775304;
  wire [7:0] sel_775305;
  wire [7:0] add_775308;
  wire [7:0] sel_775309;
  wire [7:0] add_775312;
  wire [7:0] sel_775313;
  wire [7:0] add_775316;
  wire [7:0] sel_775317;
  wire [7:0] add_775320;
  wire [7:0] sel_775321;
  wire [7:0] add_775324;
  wire [7:0] sel_775325;
  wire [7:0] add_775328;
  wire [7:0] sel_775329;
  wire [7:0] add_775332;
  wire [7:0] sel_775333;
  wire [7:0] add_775336;
  wire [7:0] sel_775337;
  wire [7:0] add_775340;
  wire [7:0] sel_775341;
  wire [7:0] add_775344;
  wire [7:0] sel_775345;
  wire [7:0] add_775348;
  wire [7:0] sel_775349;
  wire [7:0] add_775353;
  wire [15:0] array_index_775354;
  wire [7:0] sel_775355;
  wire [7:0] add_775358;
  wire [7:0] sel_775359;
  wire [7:0] add_775362;
  wire [7:0] sel_775363;
  wire [7:0] add_775366;
  wire [7:0] sel_775367;
  wire [7:0] add_775370;
  wire [7:0] sel_775371;
  wire [7:0] add_775374;
  wire [7:0] sel_775375;
  wire [7:0] add_775378;
  wire [7:0] sel_775379;
  wire [7:0] add_775382;
  wire [7:0] sel_775383;
  wire [7:0] add_775386;
  wire [7:0] sel_775387;
  wire [7:0] add_775390;
  wire [7:0] sel_775391;
  wire [7:0] add_775394;
  wire [7:0] sel_775395;
  wire [7:0] add_775398;
  wire [7:0] sel_775399;
  wire [7:0] add_775402;
  wire [7:0] sel_775403;
  wire [7:0] add_775406;
  wire [7:0] sel_775407;
  wire [7:0] add_775410;
  wire [7:0] sel_775411;
  wire [7:0] add_775414;
  wire [7:0] sel_775415;
  wire [7:0] add_775418;
  wire [7:0] sel_775419;
  wire [7:0] add_775422;
  wire [7:0] sel_775423;
  wire [7:0] add_775426;
  wire [7:0] sel_775427;
  wire [7:0] add_775430;
  wire [7:0] sel_775431;
  wire [7:0] add_775434;
  wire [7:0] sel_775435;
  wire [7:0] add_775438;
  wire [7:0] sel_775439;
  wire [7:0] add_775442;
  wire [7:0] sel_775443;
  wire [7:0] add_775446;
  wire [7:0] sel_775447;
  wire [7:0] add_775450;
  wire [7:0] sel_775451;
  wire [7:0] add_775454;
  wire [7:0] sel_775455;
  wire [7:0] add_775458;
  wire [7:0] sel_775459;
  wire [7:0] add_775462;
  wire [7:0] sel_775463;
  wire [7:0] add_775466;
  wire [7:0] sel_775467;
  wire [7:0] add_775470;
  wire [7:0] sel_775471;
  wire [7:0] add_775474;
  wire [7:0] sel_775475;
  wire [7:0] add_775478;
  wire [7:0] sel_775479;
  wire [7:0] add_775482;
  wire [7:0] sel_775483;
  wire [7:0] add_775486;
  wire [7:0] sel_775487;
  wire [7:0] add_775490;
  wire [7:0] sel_775491;
  wire [7:0] add_775494;
  wire [7:0] sel_775495;
  wire [7:0] add_775498;
  wire [7:0] sel_775499;
  wire [7:0] add_775502;
  wire [7:0] sel_775503;
  wire [7:0] add_775506;
  wire [7:0] sel_775507;
  wire [7:0] add_775510;
  wire [7:0] sel_775511;
  wire [7:0] add_775514;
  wire [7:0] sel_775515;
  wire [7:0] add_775518;
  wire [7:0] sel_775519;
  wire [7:0] add_775522;
  wire [7:0] sel_775523;
  wire [7:0] add_775526;
  wire [7:0] sel_775527;
  wire [7:0] add_775530;
  wire [7:0] sel_775531;
  wire [7:0] add_775534;
  wire [7:0] sel_775535;
  wire [7:0] add_775538;
  wire [7:0] sel_775539;
  wire [7:0] add_775542;
  wire [7:0] sel_775543;
  wire [7:0] add_775546;
  wire [7:0] sel_775547;
  wire [7:0] add_775550;
  wire [7:0] sel_775551;
  wire [7:0] add_775554;
  wire [7:0] sel_775555;
  wire [7:0] add_775558;
  wire [7:0] sel_775559;
  wire [7:0] add_775562;
  wire [7:0] sel_775563;
  wire [7:0] add_775566;
  wire [7:0] sel_775567;
  wire [7:0] add_775570;
  wire [7:0] sel_775571;
  wire [7:0] add_775574;
  wire [7:0] sel_775575;
  wire [7:0] add_775578;
  wire [7:0] sel_775579;
  wire [7:0] add_775582;
  wire [7:0] sel_775583;
  wire [7:0] add_775586;
  wire [7:0] sel_775587;
  wire [7:0] add_775590;
  wire [7:0] sel_775591;
  wire [7:0] add_775594;
  wire [7:0] sel_775595;
  wire [7:0] add_775598;
  wire [7:0] sel_775599;
  wire [7:0] add_775602;
  wire [7:0] sel_775603;
  wire [7:0] add_775606;
  wire [7:0] sel_775607;
  wire [7:0] add_775610;
  wire [7:0] sel_775611;
  wire [7:0] add_775614;
  wire [7:0] sel_775615;
  wire [7:0] add_775618;
  wire [7:0] sel_775619;
  wire [7:0] add_775622;
  wire [7:0] sel_775623;
  wire [7:0] add_775626;
  wire [7:0] sel_775627;
  wire [7:0] add_775630;
  wire [7:0] sel_775631;
  wire [7:0] add_775634;
  wire [7:0] sel_775635;
  wire [7:0] add_775638;
  wire [7:0] sel_775639;
  wire [7:0] add_775642;
  wire [7:0] sel_775643;
  wire [7:0] add_775646;
  wire [7:0] sel_775647;
  wire [7:0] add_775650;
  wire [7:0] sel_775651;
  wire [7:0] add_775654;
  wire [7:0] sel_775655;
  wire [7:0] add_775658;
  wire [7:0] sel_775659;
  wire [7:0] add_775662;
  wire [7:0] sel_775663;
  wire [7:0] add_775666;
  wire [7:0] sel_775667;
  wire [7:0] add_775670;
  wire [7:0] sel_775671;
  wire [7:0] add_775674;
  wire [7:0] sel_775675;
  wire [7:0] add_775678;
  wire [7:0] sel_775679;
  wire [7:0] add_775682;
  wire [7:0] sel_775683;
  wire [7:0] add_775686;
  wire [7:0] sel_775687;
  wire [7:0] add_775690;
  wire [7:0] sel_775691;
  wire [7:0] add_775694;
  wire [7:0] sel_775695;
  wire [7:0] add_775698;
  wire [7:0] sel_775699;
  wire [7:0] add_775702;
  wire [7:0] sel_775703;
  wire [7:0] add_775706;
  wire [7:0] sel_775707;
  wire [7:0] add_775710;
  wire [7:0] sel_775711;
  wire [7:0] add_775715;
  wire [15:0] array_index_775716;
  wire [7:0] sel_775717;
  wire [7:0] add_775720;
  wire [7:0] sel_775721;
  wire [7:0] add_775724;
  wire [7:0] sel_775725;
  wire [7:0] add_775728;
  wire [7:0] sel_775729;
  wire [7:0] add_775732;
  wire [7:0] sel_775733;
  wire [7:0] add_775736;
  wire [7:0] sel_775737;
  wire [7:0] add_775740;
  wire [7:0] sel_775741;
  wire [7:0] add_775744;
  wire [7:0] sel_775745;
  wire [7:0] add_775748;
  wire [7:0] sel_775749;
  wire [7:0] add_775752;
  wire [7:0] sel_775753;
  wire [7:0] add_775756;
  wire [7:0] sel_775757;
  wire [7:0] add_775760;
  wire [7:0] sel_775761;
  wire [7:0] add_775764;
  wire [7:0] sel_775765;
  wire [7:0] add_775768;
  wire [7:0] sel_775769;
  wire [7:0] add_775772;
  wire [7:0] sel_775773;
  wire [7:0] add_775776;
  wire [7:0] sel_775777;
  wire [7:0] add_775780;
  wire [7:0] sel_775781;
  wire [7:0] add_775784;
  wire [7:0] sel_775785;
  wire [7:0] add_775788;
  wire [7:0] sel_775789;
  wire [7:0] add_775792;
  wire [7:0] sel_775793;
  wire [7:0] add_775796;
  wire [7:0] sel_775797;
  wire [7:0] add_775800;
  wire [7:0] sel_775801;
  wire [7:0] add_775804;
  wire [7:0] sel_775805;
  wire [7:0] add_775808;
  wire [7:0] sel_775809;
  wire [7:0] add_775812;
  wire [7:0] sel_775813;
  wire [7:0] add_775816;
  wire [7:0] sel_775817;
  wire [7:0] add_775820;
  wire [7:0] sel_775821;
  wire [7:0] add_775824;
  wire [7:0] sel_775825;
  wire [7:0] add_775828;
  wire [7:0] sel_775829;
  wire [7:0] add_775832;
  wire [7:0] sel_775833;
  wire [7:0] add_775836;
  wire [7:0] sel_775837;
  wire [7:0] add_775840;
  wire [7:0] sel_775841;
  wire [7:0] add_775844;
  wire [7:0] sel_775845;
  wire [7:0] add_775848;
  wire [7:0] sel_775849;
  wire [7:0] add_775852;
  wire [7:0] sel_775853;
  wire [7:0] add_775856;
  wire [7:0] sel_775857;
  wire [7:0] add_775860;
  wire [7:0] sel_775861;
  wire [7:0] add_775864;
  wire [7:0] sel_775865;
  wire [7:0] add_775868;
  wire [7:0] sel_775869;
  wire [7:0] add_775872;
  wire [7:0] sel_775873;
  wire [7:0] add_775876;
  wire [7:0] sel_775877;
  wire [7:0] add_775880;
  wire [7:0] sel_775881;
  wire [7:0] add_775884;
  wire [7:0] sel_775885;
  wire [7:0] add_775888;
  wire [7:0] sel_775889;
  wire [7:0] add_775892;
  wire [7:0] sel_775893;
  wire [7:0] add_775896;
  wire [7:0] sel_775897;
  wire [7:0] add_775900;
  wire [7:0] sel_775901;
  wire [7:0] add_775904;
  wire [7:0] sel_775905;
  wire [7:0] add_775908;
  wire [7:0] sel_775909;
  wire [7:0] add_775912;
  wire [7:0] sel_775913;
  wire [7:0] add_775916;
  wire [7:0] sel_775917;
  wire [7:0] add_775920;
  wire [7:0] sel_775921;
  wire [7:0] add_775924;
  wire [7:0] sel_775925;
  wire [7:0] add_775928;
  wire [7:0] sel_775929;
  wire [7:0] add_775932;
  wire [7:0] sel_775933;
  wire [7:0] add_775936;
  wire [7:0] sel_775937;
  wire [7:0] add_775940;
  wire [7:0] sel_775941;
  wire [7:0] add_775944;
  wire [7:0] sel_775945;
  wire [7:0] add_775948;
  wire [7:0] sel_775949;
  wire [7:0] add_775952;
  wire [7:0] sel_775953;
  wire [7:0] add_775956;
  wire [7:0] sel_775957;
  wire [7:0] add_775960;
  wire [7:0] sel_775961;
  wire [7:0] add_775964;
  wire [7:0] sel_775965;
  wire [7:0] add_775968;
  wire [7:0] sel_775969;
  wire [7:0] add_775972;
  wire [7:0] sel_775973;
  wire [7:0] add_775976;
  wire [7:0] sel_775977;
  wire [7:0] add_775980;
  wire [7:0] sel_775981;
  wire [7:0] add_775984;
  wire [7:0] sel_775985;
  wire [7:0] add_775988;
  wire [7:0] sel_775989;
  wire [7:0] add_775992;
  wire [7:0] sel_775993;
  wire [7:0] add_775996;
  wire [7:0] sel_775997;
  wire [7:0] add_776000;
  wire [7:0] sel_776001;
  wire [7:0] add_776004;
  wire [7:0] sel_776005;
  wire [7:0] add_776008;
  wire [7:0] sel_776009;
  wire [7:0] add_776012;
  wire [7:0] sel_776013;
  wire [7:0] add_776016;
  wire [7:0] sel_776017;
  wire [7:0] add_776020;
  wire [7:0] sel_776021;
  wire [7:0] add_776024;
  wire [7:0] sel_776025;
  wire [7:0] add_776028;
  wire [7:0] sel_776029;
  wire [7:0] add_776032;
  wire [7:0] sel_776033;
  wire [7:0] add_776036;
  wire [7:0] sel_776037;
  wire [7:0] add_776040;
  wire [7:0] sel_776041;
  wire [7:0] add_776044;
  wire [7:0] sel_776045;
  wire [7:0] add_776048;
  wire [7:0] sel_776049;
  wire [7:0] add_776052;
  wire [7:0] sel_776053;
  wire [7:0] add_776056;
  wire [7:0] sel_776057;
  wire [7:0] add_776060;
  wire [7:0] sel_776061;
  wire [7:0] add_776064;
  wire [7:0] sel_776065;
  wire [7:0] add_776068;
  wire [7:0] sel_776069;
  wire [7:0] add_776072;
  wire [7:0] sel_776073;
  wire [7:0] add_776077;
  wire [15:0] array_index_776078;
  wire [7:0] sel_776079;
  wire [7:0] add_776082;
  wire [7:0] sel_776083;
  wire [7:0] add_776086;
  wire [7:0] sel_776087;
  wire [7:0] add_776090;
  wire [7:0] sel_776091;
  wire [7:0] add_776094;
  wire [7:0] sel_776095;
  wire [7:0] add_776098;
  wire [7:0] sel_776099;
  wire [7:0] add_776102;
  wire [7:0] sel_776103;
  wire [7:0] add_776106;
  wire [7:0] sel_776107;
  wire [7:0] add_776110;
  wire [7:0] sel_776111;
  wire [7:0] add_776114;
  wire [7:0] sel_776115;
  wire [7:0] add_776118;
  wire [7:0] sel_776119;
  wire [7:0] add_776122;
  wire [7:0] sel_776123;
  wire [7:0] add_776126;
  wire [7:0] sel_776127;
  wire [7:0] add_776130;
  wire [7:0] sel_776131;
  wire [7:0] add_776134;
  wire [7:0] sel_776135;
  wire [7:0] add_776138;
  wire [7:0] sel_776139;
  wire [7:0] add_776142;
  wire [7:0] sel_776143;
  wire [7:0] add_776146;
  wire [7:0] sel_776147;
  wire [7:0] add_776150;
  wire [7:0] sel_776151;
  wire [7:0] add_776154;
  wire [7:0] sel_776155;
  wire [7:0] add_776158;
  wire [7:0] sel_776159;
  wire [7:0] add_776162;
  wire [7:0] sel_776163;
  wire [7:0] add_776166;
  wire [7:0] sel_776167;
  wire [7:0] add_776170;
  wire [7:0] sel_776171;
  wire [7:0] add_776174;
  wire [7:0] sel_776175;
  wire [7:0] add_776178;
  wire [7:0] sel_776179;
  wire [7:0] add_776182;
  wire [7:0] sel_776183;
  wire [7:0] add_776186;
  wire [7:0] sel_776187;
  wire [7:0] add_776190;
  wire [7:0] sel_776191;
  wire [7:0] add_776194;
  wire [7:0] sel_776195;
  wire [7:0] add_776198;
  wire [7:0] sel_776199;
  wire [7:0] add_776202;
  wire [7:0] sel_776203;
  wire [7:0] add_776206;
  wire [7:0] sel_776207;
  wire [7:0] add_776210;
  wire [7:0] sel_776211;
  wire [7:0] add_776214;
  wire [7:0] sel_776215;
  wire [7:0] add_776218;
  wire [7:0] sel_776219;
  wire [7:0] add_776222;
  wire [7:0] sel_776223;
  wire [7:0] add_776226;
  wire [7:0] sel_776227;
  wire [7:0] add_776230;
  wire [7:0] sel_776231;
  wire [7:0] add_776234;
  wire [7:0] sel_776235;
  wire [7:0] add_776238;
  wire [7:0] sel_776239;
  wire [7:0] add_776242;
  wire [7:0] sel_776243;
  wire [7:0] add_776246;
  wire [7:0] sel_776247;
  wire [7:0] add_776250;
  wire [7:0] sel_776251;
  wire [7:0] add_776254;
  wire [7:0] sel_776255;
  wire [7:0] add_776258;
  wire [7:0] sel_776259;
  wire [7:0] add_776262;
  wire [7:0] sel_776263;
  wire [7:0] add_776266;
  wire [7:0] sel_776267;
  wire [7:0] add_776270;
  wire [7:0] sel_776271;
  wire [7:0] add_776274;
  wire [7:0] sel_776275;
  wire [7:0] add_776278;
  wire [7:0] sel_776279;
  wire [7:0] add_776282;
  wire [7:0] sel_776283;
  wire [7:0] add_776286;
  wire [7:0] sel_776287;
  wire [7:0] add_776290;
  wire [7:0] sel_776291;
  wire [7:0] add_776294;
  wire [7:0] sel_776295;
  wire [7:0] add_776298;
  wire [7:0] sel_776299;
  wire [7:0] add_776302;
  wire [7:0] sel_776303;
  wire [7:0] add_776306;
  wire [7:0] sel_776307;
  wire [7:0] add_776310;
  wire [7:0] sel_776311;
  wire [7:0] add_776314;
  wire [7:0] sel_776315;
  wire [7:0] add_776318;
  wire [7:0] sel_776319;
  wire [7:0] add_776322;
  wire [7:0] sel_776323;
  wire [7:0] add_776326;
  wire [7:0] sel_776327;
  wire [7:0] add_776330;
  wire [7:0] sel_776331;
  wire [7:0] add_776334;
  wire [7:0] sel_776335;
  wire [7:0] add_776338;
  wire [7:0] sel_776339;
  wire [7:0] add_776342;
  wire [7:0] sel_776343;
  wire [7:0] add_776346;
  wire [7:0] sel_776347;
  wire [7:0] add_776350;
  wire [7:0] sel_776351;
  wire [7:0] add_776354;
  wire [7:0] sel_776355;
  wire [7:0] add_776358;
  wire [7:0] sel_776359;
  wire [7:0] add_776362;
  wire [7:0] sel_776363;
  wire [7:0] add_776366;
  wire [7:0] sel_776367;
  wire [7:0] add_776370;
  wire [7:0] sel_776371;
  wire [7:0] add_776374;
  wire [7:0] sel_776375;
  wire [7:0] add_776378;
  wire [7:0] sel_776379;
  wire [7:0] add_776382;
  wire [7:0] sel_776383;
  wire [7:0] add_776386;
  wire [7:0] sel_776387;
  wire [7:0] add_776390;
  wire [7:0] sel_776391;
  wire [7:0] add_776394;
  wire [7:0] sel_776395;
  wire [7:0] add_776398;
  wire [7:0] sel_776399;
  wire [7:0] add_776402;
  wire [7:0] sel_776403;
  wire [7:0] add_776406;
  wire [7:0] sel_776407;
  wire [7:0] add_776410;
  wire [7:0] sel_776411;
  wire [7:0] add_776414;
  wire [7:0] sel_776415;
  wire [7:0] add_776418;
  wire [7:0] sel_776419;
  wire [7:0] add_776422;
  wire [7:0] sel_776423;
  wire [7:0] add_776426;
  wire [7:0] sel_776427;
  wire [7:0] add_776430;
  wire [7:0] sel_776431;
  wire [7:0] add_776434;
  wire [7:0] sel_776435;
  wire [7:0] add_776439;
  wire [15:0] array_index_776440;
  wire [7:0] sel_776441;
  wire [7:0] add_776444;
  wire [7:0] sel_776445;
  wire [7:0] add_776448;
  wire [7:0] sel_776449;
  wire [7:0] add_776452;
  wire [7:0] sel_776453;
  wire [7:0] add_776456;
  wire [7:0] sel_776457;
  wire [7:0] add_776460;
  wire [7:0] sel_776461;
  wire [7:0] add_776464;
  wire [7:0] sel_776465;
  wire [7:0] add_776468;
  wire [7:0] sel_776469;
  wire [7:0] add_776472;
  wire [7:0] sel_776473;
  wire [7:0] add_776476;
  wire [7:0] sel_776477;
  wire [7:0] add_776480;
  wire [7:0] sel_776481;
  wire [7:0] add_776484;
  wire [7:0] sel_776485;
  wire [7:0] add_776488;
  wire [7:0] sel_776489;
  wire [7:0] add_776492;
  wire [7:0] sel_776493;
  wire [7:0] add_776496;
  wire [7:0] sel_776497;
  wire [7:0] add_776500;
  wire [7:0] sel_776501;
  wire [7:0] add_776504;
  wire [7:0] sel_776505;
  wire [7:0] add_776508;
  wire [7:0] sel_776509;
  wire [7:0] add_776512;
  wire [7:0] sel_776513;
  wire [7:0] add_776516;
  wire [7:0] sel_776517;
  wire [7:0] add_776520;
  wire [7:0] sel_776521;
  wire [7:0] add_776524;
  wire [7:0] sel_776525;
  wire [7:0] add_776528;
  wire [7:0] sel_776529;
  wire [7:0] add_776532;
  wire [7:0] sel_776533;
  wire [7:0] add_776536;
  wire [7:0] sel_776537;
  wire [7:0] add_776540;
  wire [7:0] sel_776541;
  wire [7:0] add_776544;
  wire [7:0] sel_776545;
  wire [7:0] add_776548;
  wire [7:0] sel_776549;
  wire [7:0] add_776552;
  wire [7:0] sel_776553;
  wire [7:0] add_776556;
  wire [7:0] sel_776557;
  wire [7:0] add_776560;
  wire [7:0] sel_776561;
  wire [7:0] add_776564;
  wire [7:0] sel_776565;
  wire [7:0] add_776568;
  wire [7:0] sel_776569;
  wire [7:0] add_776572;
  wire [7:0] sel_776573;
  wire [7:0] add_776576;
  wire [7:0] sel_776577;
  wire [7:0] add_776580;
  wire [7:0] sel_776581;
  wire [7:0] add_776584;
  wire [7:0] sel_776585;
  wire [7:0] add_776588;
  wire [7:0] sel_776589;
  wire [7:0] add_776592;
  wire [7:0] sel_776593;
  wire [7:0] add_776596;
  wire [7:0] sel_776597;
  wire [7:0] add_776600;
  wire [7:0] sel_776601;
  wire [7:0] add_776604;
  wire [7:0] sel_776605;
  wire [7:0] add_776608;
  wire [7:0] sel_776609;
  wire [7:0] add_776612;
  wire [7:0] sel_776613;
  wire [7:0] add_776616;
  wire [7:0] sel_776617;
  wire [7:0] add_776620;
  wire [7:0] sel_776621;
  wire [7:0] add_776624;
  wire [7:0] sel_776625;
  wire [7:0] add_776628;
  wire [7:0] sel_776629;
  wire [7:0] add_776632;
  wire [7:0] sel_776633;
  wire [7:0] add_776636;
  wire [7:0] sel_776637;
  wire [7:0] add_776640;
  wire [7:0] sel_776641;
  wire [7:0] add_776644;
  wire [7:0] sel_776645;
  wire [7:0] add_776648;
  wire [7:0] sel_776649;
  wire [7:0] add_776652;
  wire [7:0] sel_776653;
  wire [7:0] add_776656;
  wire [7:0] sel_776657;
  wire [7:0] add_776660;
  wire [7:0] sel_776661;
  wire [7:0] add_776664;
  wire [7:0] sel_776665;
  wire [7:0] add_776668;
  wire [7:0] sel_776669;
  wire [7:0] add_776672;
  wire [7:0] sel_776673;
  wire [7:0] add_776676;
  wire [7:0] sel_776677;
  wire [7:0] add_776680;
  wire [7:0] sel_776681;
  wire [7:0] add_776684;
  wire [7:0] sel_776685;
  wire [7:0] add_776688;
  wire [7:0] sel_776689;
  wire [7:0] add_776692;
  wire [7:0] sel_776693;
  wire [7:0] add_776696;
  wire [7:0] sel_776697;
  wire [7:0] add_776700;
  wire [7:0] sel_776701;
  wire [7:0] add_776704;
  wire [7:0] sel_776705;
  wire [7:0] add_776708;
  wire [7:0] sel_776709;
  wire [7:0] add_776712;
  wire [7:0] sel_776713;
  wire [7:0] add_776716;
  wire [7:0] sel_776717;
  wire [7:0] add_776720;
  wire [7:0] sel_776721;
  wire [7:0] add_776724;
  wire [7:0] sel_776725;
  wire [7:0] add_776728;
  wire [7:0] sel_776729;
  wire [7:0] add_776732;
  wire [7:0] sel_776733;
  wire [7:0] add_776736;
  wire [7:0] sel_776737;
  wire [7:0] add_776740;
  wire [7:0] sel_776741;
  wire [7:0] add_776744;
  wire [7:0] sel_776745;
  wire [7:0] add_776748;
  wire [7:0] sel_776749;
  wire [7:0] add_776752;
  wire [7:0] sel_776753;
  wire [7:0] add_776756;
  wire [7:0] sel_776757;
  wire [7:0] add_776760;
  wire [7:0] sel_776761;
  wire [7:0] add_776764;
  wire [7:0] sel_776765;
  wire [7:0] add_776768;
  wire [7:0] sel_776769;
  wire [7:0] add_776772;
  wire [7:0] sel_776773;
  wire [7:0] add_776776;
  wire [7:0] sel_776777;
  wire [7:0] add_776780;
  wire [7:0] sel_776781;
  wire [7:0] add_776784;
  wire [7:0] sel_776785;
  wire [7:0] add_776788;
  wire [7:0] sel_776789;
  wire [7:0] add_776792;
  wire [7:0] sel_776793;
  wire [7:0] add_776796;
  wire [7:0] sel_776797;
  wire [7:0] add_776801;
  wire [15:0] array_index_776802;
  wire [7:0] sel_776803;
  wire [7:0] add_776806;
  wire [7:0] sel_776807;
  wire [7:0] add_776810;
  wire [7:0] sel_776811;
  wire [7:0] add_776814;
  wire [7:0] sel_776815;
  wire [7:0] add_776818;
  wire [7:0] sel_776819;
  wire [7:0] add_776822;
  wire [7:0] sel_776823;
  wire [7:0] add_776826;
  wire [7:0] sel_776827;
  wire [7:0] add_776830;
  wire [7:0] sel_776831;
  wire [7:0] add_776834;
  wire [7:0] sel_776835;
  wire [7:0] add_776838;
  wire [7:0] sel_776839;
  wire [7:0] add_776842;
  wire [7:0] sel_776843;
  wire [7:0] add_776846;
  wire [7:0] sel_776847;
  wire [7:0] add_776850;
  wire [7:0] sel_776851;
  wire [7:0] add_776854;
  wire [7:0] sel_776855;
  wire [7:0] add_776858;
  wire [7:0] sel_776859;
  wire [7:0] add_776862;
  wire [7:0] sel_776863;
  wire [7:0] add_776866;
  wire [7:0] sel_776867;
  wire [7:0] add_776870;
  wire [7:0] sel_776871;
  wire [7:0] add_776874;
  wire [7:0] sel_776875;
  wire [7:0] add_776878;
  wire [7:0] sel_776879;
  wire [7:0] add_776882;
  wire [7:0] sel_776883;
  wire [7:0] add_776886;
  wire [7:0] sel_776887;
  wire [7:0] add_776890;
  wire [7:0] sel_776891;
  wire [7:0] add_776894;
  wire [7:0] sel_776895;
  wire [7:0] add_776898;
  wire [7:0] sel_776899;
  wire [7:0] add_776902;
  wire [7:0] sel_776903;
  wire [7:0] add_776906;
  wire [7:0] sel_776907;
  wire [7:0] add_776910;
  wire [7:0] sel_776911;
  wire [7:0] add_776914;
  wire [7:0] sel_776915;
  wire [7:0] add_776918;
  wire [7:0] sel_776919;
  wire [7:0] add_776922;
  wire [7:0] sel_776923;
  wire [7:0] add_776926;
  wire [7:0] sel_776927;
  wire [7:0] add_776930;
  wire [7:0] sel_776931;
  wire [7:0] add_776934;
  wire [7:0] sel_776935;
  wire [7:0] add_776938;
  wire [7:0] sel_776939;
  wire [7:0] add_776942;
  wire [7:0] sel_776943;
  wire [7:0] add_776946;
  wire [7:0] sel_776947;
  wire [7:0] add_776950;
  wire [7:0] sel_776951;
  wire [7:0] add_776954;
  wire [7:0] sel_776955;
  wire [7:0] add_776958;
  wire [7:0] sel_776959;
  wire [7:0] add_776962;
  wire [7:0] sel_776963;
  wire [7:0] add_776966;
  wire [7:0] sel_776967;
  wire [7:0] add_776970;
  wire [7:0] sel_776971;
  wire [7:0] add_776974;
  wire [7:0] sel_776975;
  wire [7:0] add_776978;
  wire [7:0] sel_776979;
  wire [7:0] add_776982;
  wire [7:0] sel_776983;
  wire [7:0] add_776986;
  wire [7:0] sel_776987;
  wire [7:0] add_776990;
  wire [7:0] sel_776991;
  wire [7:0] add_776994;
  wire [7:0] sel_776995;
  wire [7:0] add_776998;
  wire [7:0] sel_776999;
  wire [7:0] add_777002;
  wire [7:0] sel_777003;
  wire [7:0] add_777006;
  wire [7:0] sel_777007;
  wire [7:0] add_777010;
  wire [7:0] sel_777011;
  wire [7:0] add_777014;
  wire [7:0] sel_777015;
  wire [7:0] add_777018;
  wire [7:0] sel_777019;
  wire [7:0] add_777022;
  wire [7:0] sel_777023;
  wire [7:0] add_777026;
  wire [7:0] sel_777027;
  wire [7:0] add_777030;
  wire [7:0] sel_777031;
  wire [7:0] add_777034;
  wire [7:0] sel_777035;
  wire [7:0] add_777038;
  wire [7:0] sel_777039;
  wire [7:0] add_777042;
  wire [7:0] sel_777043;
  wire [7:0] add_777046;
  wire [7:0] sel_777047;
  wire [7:0] add_777050;
  wire [7:0] sel_777051;
  wire [7:0] add_777054;
  wire [7:0] sel_777055;
  wire [7:0] add_777058;
  wire [7:0] sel_777059;
  wire [7:0] add_777062;
  wire [7:0] sel_777063;
  wire [7:0] add_777066;
  wire [7:0] sel_777067;
  wire [7:0] add_777070;
  wire [7:0] sel_777071;
  wire [7:0] add_777074;
  wire [7:0] sel_777075;
  wire [7:0] add_777078;
  wire [7:0] sel_777079;
  wire [7:0] add_777082;
  wire [7:0] sel_777083;
  wire [7:0] add_777086;
  wire [7:0] sel_777087;
  wire [7:0] add_777090;
  wire [7:0] sel_777091;
  wire [7:0] add_777094;
  wire [7:0] sel_777095;
  wire [7:0] add_777098;
  wire [7:0] sel_777099;
  wire [7:0] add_777102;
  wire [7:0] sel_777103;
  wire [7:0] add_777106;
  wire [7:0] sel_777107;
  wire [7:0] add_777110;
  wire [7:0] sel_777111;
  wire [7:0] add_777114;
  wire [7:0] sel_777115;
  wire [7:0] add_777118;
  wire [7:0] sel_777119;
  wire [7:0] add_777122;
  wire [7:0] sel_777123;
  wire [7:0] add_777126;
  wire [7:0] sel_777127;
  wire [7:0] add_777130;
  wire [7:0] sel_777131;
  wire [7:0] add_777134;
  wire [7:0] sel_777135;
  wire [7:0] add_777138;
  wire [7:0] sel_777139;
  wire [7:0] add_777142;
  wire [7:0] sel_777143;
  wire [7:0] add_777146;
  wire [7:0] sel_777147;
  wire [7:0] add_777150;
  wire [7:0] sel_777151;
  wire [7:0] add_777154;
  wire [7:0] sel_777155;
  wire [7:0] add_777158;
  wire [7:0] sel_777159;
  wire [7:0] add_777163;
  wire [15:0] array_index_777164;
  wire [7:0] sel_777165;
  wire [7:0] add_777168;
  wire [7:0] sel_777169;
  wire [7:0] add_777172;
  wire [7:0] sel_777173;
  wire [7:0] add_777176;
  wire [7:0] sel_777177;
  wire [7:0] add_777180;
  wire [7:0] sel_777181;
  wire [7:0] add_777184;
  wire [7:0] sel_777185;
  wire [7:0] add_777188;
  wire [7:0] sel_777189;
  wire [7:0] add_777192;
  wire [7:0] sel_777193;
  wire [7:0] add_777196;
  wire [7:0] sel_777197;
  wire [7:0] add_777200;
  wire [7:0] sel_777201;
  wire [7:0] add_777204;
  wire [7:0] sel_777205;
  wire [7:0] add_777208;
  wire [7:0] sel_777209;
  wire [7:0] add_777212;
  wire [7:0] sel_777213;
  wire [7:0] add_777216;
  wire [7:0] sel_777217;
  wire [7:0] add_777220;
  wire [7:0] sel_777221;
  wire [7:0] add_777224;
  wire [7:0] sel_777225;
  wire [7:0] add_777228;
  wire [7:0] sel_777229;
  wire [7:0] add_777232;
  wire [7:0] sel_777233;
  wire [7:0] add_777236;
  wire [7:0] sel_777237;
  wire [7:0] add_777240;
  wire [7:0] sel_777241;
  wire [7:0] add_777244;
  wire [7:0] sel_777245;
  wire [7:0] add_777248;
  wire [7:0] sel_777249;
  wire [7:0] add_777252;
  wire [7:0] sel_777253;
  wire [7:0] add_777256;
  wire [7:0] sel_777257;
  wire [7:0] add_777260;
  wire [7:0] sel_777261;
  wire [7:0] add_777264;
  wire [7:0] sel_777265;
  wire [7:0] add_777268;
  wire [7:0] sel_777269;
  wire [7:0] add_777272;
  wire [7:0] sel_777273;
  wire [7:0] add_777276;
  wire [7:0] sel_777277;
  wire [7:0] add_777280;
  wire [7:0] sel_777281;
  wire [7:0] add_777284;
  wire [7:0] sel_777285;
  wire [7:0] add_777288;
  wire [7:0] sel_777289;
  wire [7:0] add_777292;
  wire [7:0] sel_777293;
  wire [7:0] add_777296;
  wire [7:0] sel_777297;
  wire [7:0] add_777300;
  wire [7:0] sel_777301;
  wire [7:0] add_777304;
  wire [7:0] sel_777305;
  wire [7:0] add_777308;
  wire [7:0] sel_777309;
  wire [7:0] add_777312;
  wire [7:0] sel_777313;
  wire [7:0] add_777316;
  wire [7:0] sel_777317;
  wire [7:0] add_777320;
  wire [7:0] sel_777321;
  wire [7:0] add_777324;
  wire [7:0] sel_777325;
  wire [7:0] add_777328;
  wire [7:0] sel_777329;
  wire [7:0] add_777332;
  wire [7:0] sel_777333;
  wire [7:0] add_777336;
  wire [7:0] sel_777337;
  wire [7:0] add_777340;
  wire [7:0] sel_777341;
  wire [7:0] add_777344;
  wire [7:0] sel_777345;
  wire [7:0] add_777348;
  wire [7:0] sel_777349;
  wire [7:0] add_777352;
  wire [7:0] sel_777353;
  wire [7:0] add_777356;
  wire [7:0] sel_777357;
  wire [7:0] add_777360;
  wire [7:0] sel_777361;
  wire [7:0] add_777364;
  wire [7:0] sel_777365;
  wire [7:0] add_777368;
  wire [7:0] sel_777369;
  wire [7:0] add_777372;
  wire [7:0] sel_777373;
  wire [7:0] add_777376;
  wire [7:0] sel_777377;
  wire [7:0] add_777380;
  wire [7:0] sel_777381;
  wire [7:0] add_777384;
  wire [7:0] sel_777385;
  wire [7:0] add_777388;
  wire [7:0] sel_777389;
  wire [7:0] add_777392;
  wire [7:0] sel_777393;
  wire [7:0] add_777396;
  wire [7:0] sel_777397;
  wire [7:0] add_777400;
  wire [7:0] sel_777401;
  wire [7:0] add_777404;
  wire [7:0] sel_777405;
  wire [7:0] add_777408;
  wire [7:0] sel_777409;
  wire [7:0] add_777412;
  wire [7:0] sel_777413;
  wire [7:0] add_777416;
  wire [7:0] sel_777417;
  wire [7:0] add_777420;
  wire [7:0] sel_777421;
  wire [7:0] add_777424;
  wire [7:0] sel_777425;
  wire [7:0] add_777428;
  wire [7:0] sel_777429;
  wire [7:0] add_777432;
  wire [7:0] sel_777433;
  wire [7:0] add_777436;
  wire [7:0] sel_777437;
  wire [7:0] add_777440;
  wire [7:0] sel_777441;
  wire [7:0] add_777444;
  wire [7:0] sel_777445;
  wire [7:0] add_777448;
  wire [7:0] sel_777449;
  wire [7:0] add_777452;
  wire [7:0] sel_777453;
  wire [7:0] add_777456;
  wire [7:0] sel_777457;
  wire [7:0] add_777460;
  wire [7:0] sel_777461;
  wire [7:0] add_777464;
  wire [7:0] sel_777465;
  wire [7:0] add_777468;
  wire [7:0] sel_777469;
  wire [7:0] add_777472;
  wire [7:0] sel_777473;
  wire [7:0] add_777476;
  wire [7:0] sel_777477;
  wire [7:0] add_777480;
  wire [7:0] sel_777481;
  wire [7:0] add_777484;
  wire [7:0] sel_777485;
  wire [7:0] add_777488;
  wire [7:0] sel_777489;
  wire [7:0] add_777492;
  wire [7:0] sel_777493;
  wire [7:0] add_777496;
  wire [7:0] sel_777497;
  wire [7:0] add_777500;
  wire [7:0] sel_777501;
  wire [7:0] add_777504;
  wire [7:0] sel_777505;
  wire [7:0] add_777508;
  wire [7:0] sel_777509;
  wire [7:0] add_777512;
  wire [7:0] sel_777513;
  wire [7:0] add_777516;
  wire [7:0] sel_777517;
  wire [7:0] add_777520;
  wire [7:0] sel_777521;
  wire [7:0] add_777525;
  wire [15:0] array_index_777526;
  wire [7:0] sel_777527;
  wire [7:0] add_777530;
  wire [7:0] sel_777531;
  wire [7:0] add_777534;
  wire [7:0] sel_777535;
  wire [7:0] add_777538;
  wire [7:0] sel_777539;
  wire [7:0] add_777542;
  wire [7:0] sel_777543;
  wire [7:0] add_777546;
  wire [7:0] sel_777547;
  wire [7:0] add_777550;
  wire [7:0] sel_777551;
  wire [7:0] add_777554;
  wire [7:0] sel_777555;
  wire [7:0] add_777558;
  wire [7:0] sel_777559;
  wire [7:0] add_777562;
  wire [7:0] sel_777563;
  wire [7:0] add_777566;
  wire [7:0] sel_777567;
  wire [7:0] add_777570;
  wire [7:0] sel_777571;
  wire [7:0] add_777574;
  wire [7:0] sel_777575;
  wire [7:0] add_777578;
  wire [7:0] sel_777579;
  wire [7:0] add_777582;
  wire [7:0] sel_777583;
  wire [7:0] add_777586;
  wire [7:0] sel_777587;
  wire [7:0] add_777590;
  wire [7:0] sel_777591;
  wire [7:0] add_777594;
  wire [7:0] sel_777595;
  wire [7:0] add_777598;
  wire [7:0] sel_777599;
  wire [7:0] add_777602;
  wire [7:0] sel_777603;
  wire [7:0] add_777606;
  wire [7:0] sel_777607;
  wire [7:0] add_777610;
  wire [7:0] sel_777611;
  wire [7:0] add_777614;
  wire [7:0] sel_777615;
  wire [7:0] add_777618;
  wire [7:0] sel_777619;
  wire [7:0] add_777622;
  wire [7:0] sel_777623;
  wire [7:0] add_777626;
  wire [7:0] sel_777627;
  wire [7:0] add_777630;
  wire [7:0] sel_777631;
  wire [7:0] add_777634;
  wire [7:0] sel_777635;
  wire [7:0] add_777638;
  wire [7:0] sel_777639;
  wire [7:0] add_777642;
  wire [7:0] sel_777643;
  wire [7:0] add_777646;
  wire [7:0] sel_777647;
  wire [7:0] add_777650;
  wire [7:0] sel_777651;
  wire [7:0] add_777654;
  wire [7:0] sel_777655;
  wire [7:0] add_777658;
  wire [7:0] sel_777659;
  wire [7:0] add_777662;
  wire [7:0] sel_777663;
  wire [7:0] add_777666;
  wire [7:0] sel_777667;
  wire [7:0] add_777670;
  wire [7:0] sel_777671;
  wire [7:0] add_777674;
  wire [7:0] sel_777675;
  wire [7:0] add_777678;
  wire [7:0] sel_777679;
  wire [7:0] add_777682;
  wire [7:0] sel_777683;
  wire [7:0] add_777686;
  wire [7:0] sel_777687;
  wire [7:0] add_777690;
  wire [7:0] sel_777691;
  wire [7:0] add_777694;
  wire [7:0] sel_777695;
  wire [7:0] add_777698;
  wire [7:0] sel_777699;
  wire [7:0] add_777702;
  wire [7:0] sel_777703;
  wire [7:0] add_777706;
  wire [7:0] sel_777707;
  wire [7:0] add_777710;
  wire [7:0] sel_777711;
  wire [7:0] add_777714;
  wire [7:0] sel_777715;
  wire [7:0] add_777718;
  wire [7:0] sel_777719;
  wire [7:0] add_777722;
  wire [7:0] sel_777723;
  wire [7:0] add_777726;
  wire [7:0] sel_777727;
  wire [7:0] add_777730;
  wire [7:0] sel_777731;
  wire [7:0] add_777734;
  wire [7:0] sel_777735;
  wire [7:0] add_777738;
  wire [7:0] sel_777739;
  wire [7:0] add_777742;
  wire [7:0] sel_777743;
  wire [7:0] add_777746;
  wire [7:0] sel_777747;
  wire [7:0] add_777750;
  wire [7:0] sel_777751;
  wire [7:0] add_777754;
  wire [7:0] sel_777755;
  wire [7:0] add_777758;
  wire [7:0] sel_777759;
  wire [7:0] add_777762;
  wire [7:0] sel_777763;
  wire [7:0] add_777766;
  wire [7:0] sel_777767;
  wire [7:0] add_777770;
  wire [7:0] sel_777771;
  wire [7:0] add_777774;
  wire [7:0] sel_777775;
  wire [7:0] add_777778;
  wire [7:0] sel_777779;
  wire [7:0] add_777782;
  wire [7:0] sel_777783;
  wire [7:0] add_777786;
  wire [7:0] sel_777787;
  wire [7:0] add_777790;
  wire [7:0] sel_777791;
  wire [7:0] add_777794;
  wire [7:0] sel_777795;
  wire [7:0] add_777798;
  wire [7:0] sel_777799;
  wire [7:0] add_777802;
  wire [7:0] sel_777803;
  wire [7:0] add_777806;
  wire [7:0] sel_777807;
  wire [7:0] add_777810;
  wire [7:0] sel_777811;
  wire [7:0] add_777814;
  wire [7:0] sel_777815;
  wire [7:0] add_777818;
  wire [7:0] sel_777819;
  wire [7:0] add_777822;
  wire [7:0] sel_777823;
  wire [7:0] add_777826;
  wire [7:0] sel_777827;
  wire [7:0] add_777830;
  wire [7:0] sel_777831;
  wire [7:0] add_777834;
  wire [7:0] sel_777835;
  wire [7:0] add_777838;
  wire [7:0] sel_777839;
  wire [7:0] add_777842;
  wire [7:0] sel_777843;
  wire [7:0] add_777846;
  wire [7:0] sel_777847;
  wire [7:0] add_777850;
  wire [7:0] sel_777851;
  wire [7:0] add_777854;
  wire [7:0] sel_777855;
  wire [7:0] add_777858;
  wire [7:0] sel_777859;
  wire [7:0] add_777862;
  wire [7:0] sel_777863;
  wire [7:0] add_777866;
  wire [7:0] sel_777867;
  wire [7:0] add_777870;
  wire [7:0] sel_777871;
  wire [7:0] add_777874;
  wire [7:0] sel_777875;
  wire [7:0] add_777878;
  wire [7:0] sel_777879;
  wire [7:0] add_777882;
  wire [7:0] sel_777883;
  wire [7:0] add_777887;
  wire [15:0] array_index_777888;
  wire [7:0] sel_777889;
  wire [7:0] add_777892;
  wire [7:0] sel_777893;
  wire [7:0] add_777896;
  wire [7:0] sel_777897;
  wire [7:0] add_777900;
  wire [7:0] sel_777901;
  wire [7:0] add_777904;
  wire [7:0] sel_777905;
  wire [7:0] add_777908;
  wire [7:0] sel_777909;
  wire [7:0] add_777912;
  wire [7:0] sel_777913;
  wire [7:0] add_777916;
  wire [7:0] sel_777917;
  wire [7:0] add_777920;
  wire [7:0] sel_777921;
  wire [7:0] add_777924;
  wire [7:0] sel_777925;
  wire [7:0] add_777928;
  wire [7:0] sel_777929;
  wire [7:0] add_777932;
  wire [7:0] sel_777933;
  wire [7:0] add_777936;
  wire [7:0] sel_777937;
  wire [7:0] add_777940;
  wire [7:0] sel_777941;
  wire [7:0] add_777944;
  wire [7:0] sel_777945;
  wire [7:0] add_777948;
  wire [7:0] sel_777949;
  wire [7:0] add_777952;
  wire [7:0] sel_777953;
  wire [7:0] add_777956;
  wire [7:0] sel_777957;
  wire [7:0] add_777960;
  wire [7:0] sel_777961;
  wire [7:0] add_777964;
  wire [7:0] sel_777965;
  wire [7:0] add_777968;
  wire [7:0] sel_777969;
  wire [7:0] add_777972;
  wire [7:0] sel_777973;
  wire [7:0] add_777976;
  wire [7:0] sel_777977;
  wire [7:0] add_777980;
  wire [7:0] sel_777981;
  wire [7:0] add_777984;
  wire [7:0] sel_777985;
  wire [7:0] add_777988;
  wire [7:0] sel_777989;
  wire [7:0] add_777992;
  wire [7:0] sel_777993;
  wire [7:0] add_777996;
  wire [7:0] sel_777997;
  wire [7:0] add_778000;
  wire [7:0] sel_778001;
  wire [7:0] add_778004;
  wire [7:0] sel_778005;
  wire [7:0] add_778008;
  wire [7:0] sel_778009;
  wire [7:0] add_778012;
  wire [7:0] sel_778013;
  wire [7:0] add_778016;
  wire [7:0] sel_778017;
  wire [7:0] add_778020;
  wire [7:0] sel_778021;
  wire [7:0] add_778024;
  wire [7:0] sel_778025;
  wire [7:0] add_778028;
  wire [7:0] sel_778029;
  wire [7:0] add_778032;
  wire [7:0] sel_778033;
  wire [7:0] add_778036;
  wire [7:0] sel_778037;
  wire [7:0] add_778040;
  wire [7:0] sel_778041;
  wire [7:0] add_778044;
  wire [7:0] sel_778045;
  wire [7:0] add_778048;
  wire [7:0] sel_778049;
  wire [7:0] add_778052;
  wire [7:0] sel_778053;
  wire [7:0] add_778056;
  wire [7:0] sel_778057;
  wire [7:0] add_778060;
  wire [7:0] sel_778061;
  wire [7:0] add_778064;
  wire [7:0] sel_778065;
  wire [7:0] add_778068;
  wire [7:0] sel_778069;
  wire [7:0] add_778072;
  wire [7:0] sel_778073;
  wire [7:0] add_778076;
  wire [7:0] sel_778077;
  wire [7:0] add_778080;
  wire [7:0] sel_778081;
  wire [7:0] add_778084;
  wire [7:0] sel_778085;
  wire [7:0] add_778088;
  wire [7:0] sel_778089;
  wire [7:0] add_778092;
  wire [7:0] sel_778093;
  wire [7:0] add_778096;
  wire [7:0] sel_778097;
  wire [7:0] add_778100;
  wire [7:0] sel_778101;
  wire [7:0] add_778104;
  wire [7:0] sel_778105;
  wire [7:0] add_778108;
  wire [7:0] sel_778109;
  wire [7:0] add_778112;
  wire [7:0] sel_778113;
  wire [7:0] add_778116;
  wire [7:0] sel_778117;
  wire [7:0] add_778120;
  wire [7:0] sel_778121;
  wire [7:0] add_778124;
  wire [7:0] sel_778125;
  wire [7:0] add_778128;
  wire [7:0] sel_778129;
  wire [7:0] add_778132;
  wire [7:0] sel_778133;
  wire [7:0] add_778136;
  wire [7:0] sel_778137;
  wire [7:0] add_778140;
  wire [7:0] sel_778141;
  wire [7:0] add_778144;
  wire [7:0] sel_778145;
  wire [7:0] add_778148;
  wire [7:0] sel_778149;
  wire [7:0] add_778152;
  wire [7:0] sel_778153;
  wire [7:0] add_778156;
  wire [7:0] sel_778157;
  wire [7:0] add_778160;
  wire [7:0] sel_778161;
  wire [7:0] add_778164;
  wire [7:0] sel_778165;
  wire [7:0] add_778168;
  wire [7:0] sel_778169;
  wire [7:0] add_778172;
  wire [7:0] sel_778173;
  wire [7:0] add_778176;
  wire [7:0] sel_778177;
  wire [7:0] add_778180;
  wire [7:0] sel_778181;
  wire [7:0] add_778184;
  wire [7:0] sel_778185;
  wire [7:0] add_778188;
  wire [7:0] sel_778189;
  wire [7:0] add_778192;
  wire [7:0] sel_778193;
  wire [7:0] add_778196;
  wire [7:0] sel_778197;
  wire [7:0] add_778200;
  wire [7:0] sel_778201;
  wire [7:0] add_778204;
  wire [7:0] sel_778205;
  wire [7:0] add_778208;
  wire [7:0] sel_778209;
  wire [7:0] add_778212;
  wire [7:0] sel_778213;
  wire [7:0] add_778216;
  wire [7:0] sel_778217;
  wire [7:0] add_778220;
  wire [7:0] sel_778221;
  wire [7:0] add_778224;
  wire [7:0] sel_778225;
  wire [7:0] add_778228;
  wire [7:0] sel_778229;
  wire [7:0] add_778232;
  wire [7:0] sel_778233;
  wire [7:0] add_778236;
  wire [7:0] sel_778237;
  wire [7:0] add_778240;
  wire [7:0] sel_778241;
  wire [7:0] add_778244;
  wire [7:0] sel_778245;
  wire [7:0] add_778249;
  wire [15:0] array_index_778250;
  wire [7:0] sel_778251;
  wire [7:0] add_778254;
  wire [7:0] sel_778255;
  wire [7:0] add_778258;
  wire [7:0] sel_778259;
  wire [7:0] add_778262;
  wire [7:0] sel_778263;
  wire [7:0] add_778266;
  wire [7:0] sel_778267;
  wire [7:0] add_778270;
  wire [7:0] sel_778271;
  wire [7:0] add_778274;
  wire [7:0] sel_778275;
  wire [7:0] add_778278;
  wire [7:0] sel_778279;
  wire [7:0] add_778282;
  wire [7:0] sel_778283;
  wire [7:0] add_778286;
  wire [7:0] sel_778287;
  wire [7:0] add_778290;
  wire [7:0] sel_778291;
  wire [7:0] add_778294;
  wire [7:0] sel_778295;
  wire [7:0] add_778298;
  wire [7:0] sel_778299;
  wire [7:0] add_778302;
  wire [7:0] sel_778303;
  wire [7:0] add_778306;
  wire [7:0] sel_778307;
  wire [7:0] add_778310;
  wire [7:0] sel_778311;
  wire [7:0] add_778314;
  wire [7:0] sel_778315;
  wire [7:0] add_778318;
  wire [7:0] sel_778319;
  wire [7:0] add_778322;
  wire [7:0] sel_778323;
  wire [7:0] add_778326;
  wire [7:0] sel_778327;
  wire [7:0] add_778330;
  wire [7:0] sel_778331;
  wire [7:0] add_778334;
  wire [7:0] sel_778335;
  wire [7:0] add_778338;
  wire [7:0] sel_778339;
  wire [7:0] add_778342;
  wire [7:0] sel_778343;
  wire [7:0] add_778346;
  wire [7:0] sel_778347;
  wire [7:0] add_778350;
  wire [7:0] sel_778351;
  wire [7:0] add_778354;
  wire [7:0] sel_778355;
  wire [7:0] add_778358;
  wire [7:0] sel_778359;
  wire [7:0] add_778362;
  wire [7:0] sel_778363;
  wire [7:0] add_778366;
  wire [7:0] sel_778367;
  wire [7:0] add_778370;
  wire [7:0] sel_778371;
  wire [7:0] add_778374;
  wire [7:0] sel_778375;
  wire [7:0] add_778378;
  wire [7:0] sel_778379;
  wire [7:0] add_778382;
  wire [7:0] sel_778383;
  wire [7:0] add_778386;
  wire [7:0] sel_778387;
  wire [7:0] add_778390;
  wire [7:0] sel_778391;
  wire [7:0] add_778394;
  wire [7:0] sel_778395;
  wire [7:0] add_778398;
  wire [7:0] sel_778399;
  wire [7:0] add_778402;
  wire [7:0] sel_778403;
  wire [7:0] add_778406;
  wire [7:0] sel_778407;
  wire [7:0] add_778410;
  wire [7:0] sel_778411;
  wire [7:0] add_778414;
  wire [7:0] sel_778415;
  wire [7:0] add_778418;
  wire [7:0] sel_778419;
  wire [7:0] add_778422;
  wire [7:0] sel_778423;
  wire [7:0] add_778426;
  wire [7:0] sel_778427;
  wire [7:0] add_778430;
  wire [7:0] sel_778431;
  wire [7:0] add_778434;
  wire [7:0] sel_778435;
  wire [7:0] add_778438;
  wire [7:0] sel_778439;
  wire [7:0] add_778442;
  wire [7:0] sel_778443;
  wire [7:0] add_778446;
  wire [7:0] sel_778447;
  wire [7:0] add_778450;
  wire [7:0] sel_778451;
  wire [7:0] add_778454;
  wire [7:0] sel_778455;
  wire [7:0] add_778458;
  wire [7:0] sel_778459;
  wire [7:0] add_778462;
  wire [7:0] sel_778463;
  wire [7:0] add_778466;
  wire [7:0] sel_778467;
  wire [7:0] add_778470;
  wire [7:0] sel_778471;
  wire [7:0] add_778474;
  wire [7:0] sel_778475;
  wire [7:0] add_778478;
  wire [7:0] sel_778479;
  wire [7:0] add_778482;
  wire [7:0] sel_778483;
  wire [7:0] add_778486;
  wire [7:0] sel_778487;
  wire [7:0] add_778490;
  wire [7:0] sel_778491;
  wire [7:0] add_778494;
  wire [7:0] sel_778495;
  wire [7:0] add_778498;
  wire [7:0] sel_778499;
  wire [7:0] add_778502;
  wire [7:0] sel_778503;
  wire [7:0] add_778506;
  wire [7:0] sel_778507;
  wire [7:0] add_778510;
  wire [7:0] sel_778511;
  wire [7:0] add_778514;
  wire [7:0] sel_778515;
  wire [7:0] add_778518;
  wire [7:0] sel_778519;
  wire [7:0] add_778522;
  wire [7:0] sel_778523;
  wire [7:0] add_778526;
  wire [7:0] sel_778527;
  wire [7:0] add_778530;
  wire [7:0] sel_778531;
  wire [7:0] add_778534;
  wire [7:0] sel_778535;
  wire [7:0] add_778538;
  wire [7:0] sel_778539;
  wire [7:0] add_778542;
  wire [7:0] sel_778543;
  wire [7:0] add_778546;
  wire [7:0] sel_778547;
  wire [7:0] add_778550;
  wire [7:0] sel_778551;
  wire [7:0] add_778554;
  wire [7:0] sel_778555;
  wire [7:0] add_778558;
  wire [7:0] sel_778559;
  wire [7:0] add_778562;
  wire [7:0] sel_778563;
  wire [7:0] add_778566;
  wire [7:0] sel_778567;
  wire [7:0] add_778570;
  wire [7:0] sel_778571;
  wire [7:0] add_778574;
  wire [7:0] sel_778575;
  wire [7:0] add_778578;
  wire [7:0] sel_778579;
  wire [7:0] add_778582;
  wire [7:0] sel_778583;
  wire [7:0] add_778586;
  wire [7:0] sel_778587;
  wire [7:0] add_778590;
  wire [7:0] sel_778591;
  wire [7:0] add_778594;
  wire [7:0] sel_778595;
  wire [7:0] add_778598;
  wire [7:0] sel_778599;
  wire [7:0] add_778602;
  wire [7:0] sel_778603;
  wire [7:0] add_778606;
  wire [7:0] sel_778607;
  wire [7:0] add_778611;
  wire [15:0] array_index_778612;
  wire [7:0] sel_778613;
  wire [7:0] add_778616;
  wire [7:0] sel_778617;
  wire [7:0] add_778620;
  wire [7:0] sel_778621;
  wire [7:0] add_778624;
  wire [7:0] sel_778625;
  wire [7:0] add_778628;
  wire [7:0] sel_778629;
  wire [7:0] add_778632;
  wire [7:0] sel_778633;
  wire [7:0] add_778636;
  wire [7:0] sel_778637;
  wire [7:0] add_778640;
  wire [7:0] sel_778641;
  wire [7:0] add_778644;
  wire [7:0] sel_778645;
  wire [7:0] add_778648;
  wire [7:0] sel_778649;
  wire [7:0] add_778652;
  wire [7:0] sel_778653;
  wire [7:0] add_778656;
  wire [7:0] sel_778657;
  wire [7:0] add_778660;
  wire [7:0] sel_778661;
  wire [7:0] add_778664;
  wire [7:0] sel_778665;
  wire [7:0] add_778668;
  wire [7:0] sel_778669;
  wire [7:0] add_778672;
  wire [7:0] sel_778673;
  wire [7:0] add_778676;
  wire [7:0] sel_778677;
  wire [7:0] add_778680;
  wire [7:0] sel_778681;
  wire [7:0] add_778684;
  wire [7:0] sel_778685;
  wire [7:0] add_778688;
  wire [7:0] sel_778689;
  wire [7:0] add_778692;
  wire [7:0] sel_778693;
  wire [7:0] add_778696;
  wire [7:0] sel_778697;
  wire [7:0] add_778700;
  wire [7:0] sel_778701;
  wire [7:0] add_778704;
  wire [7:0] sel_778705;
  wire [7:0] add_778708;
  wire [7:0] sel_778709;
  wire [7:0] add_778712;
  wire [7:0] sel_778713;
  wire [7:0] add_778716;
  wire [7:0] sel_778717;
  wire [7:0] add_778720;
  wire [7:0] sel_778721;
  wire [7:0] add_778724;
  wire [7:0] sel_778725;
  wire [7:0] add_778728;
  wire [7:0] sel_778729;
  wire [7:0] add_778732;
  wire [7:0] sel_778733;
  wire [7:0] add_778736;
  wire [7:0] sel_778737;
  wire [7:0] add_778740;
  wire [7:0] sel_778741;
  wire [7:0] add_778744;
  wire [7:0] sel_778745;
  wire [7:0] add_778748;
  wire [7:0] sel_778749;
  wire [7:0] add_778752;
  wire [7:0] sel_778753;
  wire [7:0] add_778756;
  wire [7:0] sel_778757;
  wire [7:0] add_778760;
  wire [7:0] sel_778761;
  wire [7:0] add_778764;
  wire [7:0] sel_778765;
  wire [7:0] add_778768;
  wire [7:0] sel_778769;
  wire [7:0] add_778772;
  wire [7:0] sel_778773;
  wire [7:0] add_778776;
  wire [7:0] sel_778777;
  wire [7:0] add_778780;
  wire [7:0] sel_778781;
  wire [7:0] add_778784;
  wire [7:0] sel_778785;
  wire [7:0] add_778788;
  wire [7:0] sel_778789;
  wire [7:0] add_778792;
  wire [7:0] sel_778793;
  wire [7:0] add_778796;
  wire [7:0] sel_778797;
  wire [7:0] add_778800;
  wire [7:0] sel_778801;
  wire [7:0] add_778804;
  wire [7:0] sel_778805;
  wire [7:0] add_778808;
  wire [7:0] sel_778809;
  wire [7:0] add_778812;
  wire [7:0] sel_778813;
  wire [7:0] add_778816;
  wire [7:0] sel_778817;
  wire [7:0] add_778820;
  wire [7:0] sel_778821;
  wire [7:0] add_778824;
  wire [7:0] sel_778825;
  wire [7:0] add_778828;
  wire [7:0] sel_778829;
  wire [7:0] add_778832;
  wire [7:0] sel_778833;
  wire [7:0] add_778836;
  wire [7:0] sel_778837;
  wire [7:0] add_778840;
  wire [7:0] sel_778841;
  wire [7:0] add_778844;
  wire [7:0] sel_778845;
  wire [7:0] add_778848;
  wire [7:0] sel_778849;
  wire [7:0] add_778852;
  wire [7:0] sel_778853;
  wire [7:0] add_778856;
  wire [7:0] sel_778857;
  wire [7:0] add_778860;
  wire [7:0] sel_778861;
  wire [7:0] add_778864;
  wire [7:0] sel_778865;
  wire [7:0] add_778868;
  wire [7:0] sel_778869;
  wire [7:0] add_778872;
  wire [7:0] sel_778873;
  wire [7:0] add_778876;
  wire [7:0] sel_778877;
  wire [7:0] add_778880;
  wire [7:0] sel_778881;
  wire [7:0] add_778884;
  wire [7:0] sel_778885;
  wire [7:0] add_778888;
  wire [7:0] sel_778889;
  wire [7:0] add_778892;
  wire [7:0] sel_778893;
  wire [7:0] add_778896;
  wire [7:0] sel_778897;
  wire [7:0] add_778900;
  wire [7:0] sel_778901;
  wire [7:0] add_778904;
  wire [7:0] sel_778905;
  wire [7:0] add_778908;
  wire [7:0] sel_778909;
  wire [7:0] add_778912;
  wire [7:0] sel_778913;
  wire [7:0] add_778916;
  wire [7:0] sel_778917;
  wire [7:0] add_778920;
  wire [7:0] sel_778921;
  wire [7:0] add_778924;
  wire [7:0] sel_778925;
  wire [7:0] add_778928;
  wire [7:0] sel_778929;
  wire [7:0] add_778932;
  wire [7:0] sel_778933;
  wire [7:0] add_778936;
  wire [7:0] sel_778937;
  wire [7:0] add_778940;
  wire [7:0] sel_778941;
  wire [7:0] add_778944;
  wire [7:0] sel_778945;
  wire [7:0] add_778948;
  wire [7:0] sel_778949;
  wire [7:0] add_778952;
  wire [7:0] sel_778953;
  wire [7:0] add_778956;
  wire [7:0] sel_778957;
  wire [7:0] add_778960;
  wire [7:0] sel_778961;
  wire [7:0] add_778964;
  wire [7:0] sel_778965;
  wire [7:0] add_778968;
  wire [7:0] sel_778969;
  wire [7:0] add_778973;
  wire [15:0] array_index_778974;
  wire [7:0] sel_778975;
  wire [7:0] add_778978;
  wire [7:0] sel_778979;
  wire [7:0] add_778982;
  wire [7:0] sel_778983;
  wire [7:0] add_778986;
  wire [7:0] sel_778987;
  wire [7:0] add_778990;
  wire [7:0] sel_778991;
  wire [7:0] add_778994;
  wire [7:0] sel_778995;
  wire [7:0] add_778998;
  wire [7:0] sel_778999;
  wire [7:0] add_779002;
  wire [7:0] sel_779003;
  wire [7:0] add_779006;
  wire [7:0] sel_779007;
  wire [7:0] add_779010;
  wire [7:0] sel_779011;
  wire [7:0] add_779014;
  wire [7:0] sel_779015;
  wire [7:0] add_779018;
  wire [7:0] sel_779019;
  wire [7:0] add_779022;
  wire [7:0] sel_779023;
  wire [7:0] add_779026;
  wire [7:0] sel_779027;
  wire [7:0] add_779030;
  wire [7:0] sel_779031;
  wire [7:0] add_779034;
  wire [7:0] sel_779035;
  wire [7:0] add_779038;
  wire [7:0] sel_779039;
  wire [7:0] add_779042;
  wire [7:0] sel_779043;
  wire [7:0] add_779046;
  wire [7:0] sel_779047;
  wire [7:0] add_779050;
  wire [7:0] sel_779051;
  wire [7:0] add_779054;
  wire [7:0] sel_779055;
  wire [7:0] add_779058;
  wire [7:0] sel_779059;
  wire [7:0] add_779062;
  wire [7:0] sel_779063;
  wire [7:0] add_779066;
  wire [7:0] sel_779067;
  wire [7:0] add_779070;
  wire [7:0] sel_779071;
  wire [7:0] add_779074;
  wire [7:0] sel_779075;
  wire [7:0] add_779078;
  wire [7:0] sel_779079;
  wire [7:0] add_779082;
  wire [7:0] sel_779083;
  wire [7:0] add_779086;
  wire [7:0] sel_779087;
  wire [7:0] add_779090;
  wire [7:0] sel_779091;
  wire [7:0] add_779094;
  wire [7:0] sel_779095;
  wire [7:0] add_779098;
  wire [7:0] sel_779099;
  wire [7:0] add_779102;
  wire [7:0] sel_779103;
  wire [7:0] add_779106;
  wire [7:0] sel_779107;
  wire [7:0] add_779110;
  wire [7:0] sel_779111;
  wire [7:0] add_779114;
  wire [7:0] sel_779115;
  wire [7:0] add_779118;
  wire [7:0] sel_779119;
  wire [7:0] add_779122;
  wire [7:0] sel_779123;
  wire [7:0] add_779126;
  wire [7:0] sel_779127;
  wire [7:0] add_779130;
  wire [7:0] sel_779131;
  wire [7:0] add_779134;
  wire [7:0] sel_779135;
  wire [7:0] add_779138;
  wire [7:0] sel_779139;
  wire [7:0] add_779142;
  wire [7:0] sel_779143;
  wire [7:0] add_779146;
  wire [7:0] sel_779147;
  wire [7:0] add_779150;
  wire [7:0] sel_779151;
  wire [7:0] add_779154;
  wire [7:0] sel_779155;
  wire [7:0] add_779158;
  wire [7:0] sel_779159;
  wire [7:0] add_779162;
  wire [7:0] sel_779163;
  wire [7:0] add_779166;
  wire [7:0] sel_779167;
  wire [7:0] add_779170;
  wire [7:0] sel_779171;
  wire [7:0] add_779174;
  wire [7:0] sel_779175;
  wire [7:0] add_779178;
  wire [7:0] sel_779179;
  wire [7:0] add_779182;
  wire [7:0] sel_779183;
  wire [7:0] add_779186;
  wire [7:0] sel_779187;
  wire [7:0] add_779190;
  wire [7:0] sel_779191;
  wire [7:0] add_779194;
  wire [7:0] sel_779195;
  wire [7:0] add_779198;
  wire [7:0] sel_779199;
  wire [7:0] add_779202;
  wire [7:0] sel_779203;
  wire [7:0] add_779206;
  wire [7:0] sel_779207;
  wire [7:0] add_779210;
  wire [7:0] sel_779211;
  wire [7:0] add_779214;
  wire [7:0] sel_779215;
  wire [7:0] add_779218;
  wire [7:0] sel_779219;
  wire [7:0] add_779222;
  wire [7:0] sel_779223;
  wire [7:0] add_779226;
  wire [7:0] sel_779227;
  wire [7:0] add_779230;
  wire [7:0] sel_779231;
  wire [7:0] add_779234;
  wire [7:0] sel_779235;
  wire [7:0] add_779238;
  wire [7:0] sel_779239;
  wire [7:0] add_779242;
  wire [7:0] sel_779243;
  wire [7:0] add_779246;
  wire [7:0] sel_779247;
  wire [7:0] add_779250;
  wire [7:0] sel_779251;
  wire [7:0] add_779254;
  wire [7:0] sel_779255;
  wire [7:0] add_779258;
  wire [7:0] sel_779259;
  wire [7:0] add_779262;
  wire [7:0] sel_779263;
  wire [7:0] add_779266;
  wire [7:0] sel_779267;
  wire [7:0] add_779270;
  wire [7:0] sel_779271;
  wire [7:0] add_779274;
  wire [7:0] sel_779275;
  wire [7:0] add_779278;
  wire [7:0] sel_779279;
  wire [7:0] add_779282;
  wire [7:0] sel_779283;
  wire [7:0] add_779286;
  wire [7:0] sel_779287;
  wire [7:0] add_779290;
  wire [7:0] sel_779291;
  wire [7:0] add_779294;
  wire [7:0] sel_779295;
  wire [7:0] add_779298;
  wire [7:0] sel_779299;
  wire [7:0] add_779302;
  wire [7:0] sel_779303;
  wire [7:0] add_779306;
  wire [7:0] sel_779307;
  wire [7:0] add_779310;
  wire [7:0] sel_779311;
  wire [7:0] add_779314;
  wire [7:0] sel_779315;
  wire [7:0] add_779318;
  wire [7:0] sel_779319;
  wire [7:0] add_779322;
  wire [7:0] sel_779323;
  wire [7:0] add_779326;
  wire [7:0] sel_779327;
  wire [7:0] add_779330;
  wire [7:0] sel_779331;
  wire [7:0] add_779335;
  wire [15:0] array_index_779336;
  wire [7:0] sel_779337;
  wire [7:0] add_779340;
  wire [7:0] sel_779341;
  wire [7:0] add_779344;
  wire [7:0] sel_779345;
  wire [7:0] add_779348;
  wire [7:0] sel_779349;
  wire [7:0] add_779352;
  wire [7:0] sel_779353;
  wire [7:0] add_779356;
  wire [7:0] sel_779357;
  wire [7:0] add_779360;
  wire [7:0] sel_779361;
  wire [7:0] add_779364;
  wire [7:0] sel_779365;
  wire [7:0] add_779368;
  wire [7:0] sel_779369;
  wire [7:0] add_779372;
  wire [7:0] sel_779373;
  wire [7:0] add_779376;
  wire [7:0] sel_779377;
  wire [7:0] add_779380;
  wire [7:0] sel_779381;
  wire [7:0] add_779384;
  wire [7:0] sel_779385;
  wire [7:0] add_779388;
  wire [7:0] sel_779389;
  wire [7:0] add_779392;
  wire [7:0] sel_779393;
  wire [7:0] add_779396;
  wire [7:0] sel_779397;
  wire [7:0] add_779400;
  wire [7:0] sel_779401;
  wire [7:0] add_779404;
  wire [7:0] sel_779405;
  wire [7:0] add_779408;
  wire [7:0] sel_779409;
  wire [7:0] add_779412;
  wire [7:0] sel_779413;
  wire [7:0] add_779416;
  wire [7:0] sel_779417;
  wire [7:0] add_779420;
  wire [7:0] sel_779421;
  wire [7:0] add_779424;
  wire [7:0] sel_779425;
  wire [7:0] add_779428;
  wire [7:0] sel_779429;
  wire [7:0] add_779432;
  wire [7:0] sel_779433;
  wire [7:0] add_779436;
  wire [7:0] sel_779437;
  wire [7:0] add_779440;
  wire [7:0] sel_779441;
  wire [7:0] add_779444;
  wire [7:0] sel_779445;
  wire [7:0] add_779448;
  wire [7:0] sel_779449;
  wire [7:0] add_779452;
  wire [7:0] sel_779453;
  wire [7:0] add_779456;
  wire [7:0] sel_779457;
  wire [7:0] add_779460;
  wire [7:0] sel_779461;
  wire [7:0] add_779464;
  wire [7:0] sel_779465;
  wire [7:0] add_779468;
  wire [7:0] sel_779469;
  wire [7:0] add_779472;
  wire [7:0] sel_779473;
  wire [7:0] add_779476;
  wire [7:0] sel_779477;
  wire [7:0] add_779480;
  wire [7:0] sel_779481;
  wire [7:0] add_779484;
  wire [7:0] sel_779485;
  wire [7:0] add_779488;
  wire [7:0] sel_779489;
  wire [7:0] add_779492;
  wire [7:0] sel_779493;
  wire [7:0] add_779496;
  wire [7:0] sel_779497;
  wire [7:0] add_779500;
  wire [7:0] sel_779501;
  wire [7:0] add_779504;
  wire [7:0] sel_779505;
  wire [7:0] add_779508;
  wire [7:0] sel_779509;
  wire [7:0] add_779512;
  wire [7:0] sel_779513;
  wire [7:0] add_779516;
  wire [7:0] sel_779517;
  wire [7:0] add_779520;
  wire [7:0] sel_779521;
  wire [7:0] add_779524;
  wire [7:0] sel_779525;
  wire [7:0] add_779528;
  wire [7:0] sel_779529;
  wire [7:0] add_779532;
  wire [7:0] sel_779533;
  wire [7:0] add_779536;
  wire [7:0] sel_779537;
  wire [7:0] add_779540;
  wire [7:0] sel_779541;
  wire [7:0] add_779544;
  wire [7:0] sel_779545;
  wire [7:0] add_779548;
  wire [7:0] sel_779549;
  wire [7:0] add_779552;
  wire [7:0] sel_779553;
  wire [7:0] add_779556;
  wire [7:0] sel_779557;
  wire [7:0] add_779560;
  wire [7:0] sel_779561;
  wire [7:0] add_779564;
  wire [7:0] sel_779565;
  wire [7:0] add_779568;
  wire [7:0] sel_779569;
  wire [7:0] add_779572;
  wire [7:0] sel_779573;
  wire [7:0] add_779576;
  wire [7:0] sel_779577;
  wire [7:0] add_779580;
  wire [7:0] sel_779581;
  wire [7:0] add_779584;
  wire [7:0] sel_779585;
  wire [7:0] add_779588;
  wire [7:0] sel_779589;
  wire [7:0] add_779592;
  wire [7:0] sel_779593;
  wire [7:0] add_779596;
  wire [7:0] sel_779597;
  wire [7:0] add_779600;
  wire [7:0] sel_779601;
  wire [7:0] add_779604;
  wire [7:0] sel_779605;
  wire [7:0] add_779608;
  wire [7:0] sel_779609;
  wire [7:0] add_779612;
  wire [7:0] sel_779613;
  wire [7:0] add_779616;
  wire [7:0] sel_779617;
  wire [7:0] add_779620;
  wire [7:0] sel_779621;
  wire [7:0] add_779624;
  wire [7:0] sel_779625;
  wire [7:0] add_779628;
  wire [7:0] sel_779629;
  wire [7:0] add_779632;
  wire [7:0] sel_779633;
  wire [7:0] add_779636;
  wire [7:0] sel_779637;
  wire [7:0] add_779640;
  wire [7:0] sel_779641;
  wire [7:0] add_779644;
  wire [7:0] sel_779645;
  wire [7:0] add_779648;
  wire [7:0] sel_779649;
  wire [7:0] add_779652;
  wire [7:0] sel_779653;
  wire [7:0] add_779656;
  wire [7:0] sel_779657;
  wire [7:0] add_779660;
  wire [7:0] sel_779661;
  wire [7:0] add_779664;
  wire [7:0] sel_779665;
  wire [7:0] add_779668;
  wire [7:0] sel_779669;
  wire [7:0] add_779672;
  wire [7:0] sel_779673;
  wire [7:0] add_779676;
  wire [7:0] sel_779677;
  wire [7:0] add_779680;
  wire [7:0] sel_779681;
  wire [7:0] add_779684;
  wire [7:0] sel_779685;
  wire [7:0] add_779688;
  wire [7:0] sel_779689;
  wire [7:0] add_779692;
  wire [7:0] sel_779693;
  wire [7:0] add_779697;
  wire [15:0] array_index_779698;
  wire [7:0] sel_779699;
  wire [7:0] add_779702;
  wire [7:0] sel_779703;
  wire [7:0] add_779706;
  wire [7:0] sel_779707;
  wire [7:0] add_779710;
  wire [7:0] sel_779711;
  wire [7:0] add_779714;
  wire [7:0] sel_779715;
  wire [7:0] add_779718;
  wire [7:0] sel_779719;
  wire [7:0] add_779722;
  wire [7:0] sel_779723;
  wire [7:0] add_779726;
  wire [7:0] sel_779727;
  wire [7:0] add_779730;
  wire [7:0] sel_779731;
  wire [7:0] add_779734;
  wire [7:0] sel_779735;
  wire [7:0] add_779738;
  wire [7:0] sel_779739;
  wire [7:0] add_779742;
  wire [7:0] sel_779743;
  wire [7:0] add_779746;
  wire [7:0] sel_779747;
  wire [7:0] add_779750;
  wire [7:0] sel_779751;
  wire [7:0] add_779754;
  wire [7:0] sel_779755;
  wire [7:0] add_779758;
  wire [7:0] sel_779759;
  wire [7:0] add_779762;
  wire [7:0] sel_779763;
  wire [7:0] add_779766;
  wire [7:0] sel_779767;
  wire [7:0] add_779770;
  wire [7:0] sel_779771;
  wire [7:0] add_779774;
  wire [7:0] sel_779775;
  wire [7:0] add_779778;
  wire [7:0] sel_779779;
  wire [7:0] add_779782;
  wire [7:0] sel_779783;
  wire [7:0] add_779786;
  wire [7:0] sel_779787;
  wire [7:0] add_779790;
  wire [7:0] sel_779791;
  wire [7:0] add_779794;
  wire [7:0] sel_779795;
  wire [7:0] add_779798;
  wire [7:0] sel_779799;
  wire [7:0] add_779802;
  wire [7:0] sel_779803;
  wire [7:0] add_779806;
  wire [7:0] sel_779807;
  wire [7:0] add_779810;
  wire [7:0] sel_779811;
  wire [7:0] add_779814;
  wire [7:0] sel_779815;
  wire [7:0] add_779818;
  wire [7:0] sel_779819;
  wire [7:0] add_779822;
  wire [7:0] sel_779823;
  wire [7:0] add_779826;
  wire [7:0] sel_779827;
  wire [7:0] add_779830;
  wire [7:0] sel_779831;
  wire [7:0] add_779834;
  wire [7:0] sel_779835;
  wire [7:0] add_779838;
  wire [7:0] sel_779839;
  wire [7:0] add_779842;
  wire [7:0] sel_779843;
  wire [7:0] add_779846;
  wire [7:0] sel_779847;
  wire [7:0] add_779850;
  wire [7:0] sel_779851;
  wire [7:0] add_779854;
  wire [7:0] sel_779855;
  wire [7:0] add_779858;
  wire [7:0] sel_779859;
  wire [7:0] add_779862;
  wire [7:0] sel_779863;
  wire [7:0] add_779866;
  wire [7:0] sel_779867;
  wire [7:0] add_779870;
  wire [7:0] sel_779871;
  wire [7:0] add_779874;
  wire [7:0] sel_779875;
  wire [7:0] add_779878;
  wire [7:0] sel_779879;
  wire [7:0] add_779882;
  wire [7:0] sel_779883;
  wire [7:0] add_779886;
  wire [7:0] sel_779887;
  wire [7:0] add_779890;
  wire [7:0] sel_779891;
  wire [7:0] add_779894;
  wire [7:0] sel_779895;
  wire [7:0] add_779898;
  wire [7:0] sel_779899;
  wire [7:0] add_779902;
  wire [7:0] sel_779903;
  wire [7:0] add_779906;
  wire [7:0] sel_779907;
  wire [7:0] add_779910;
  wire [7:0] sel_779911;
  wire [7:0] add_779914;
  wire [7:0] sel_779915;
  wire [7:0] add_779918;
  wire [7:0] sel_779919;
  wire [7:0] add_779922;
  wire [7:0] sel_779923;
  wire [7:0] add_779926;
  wire [7:0] sel_779927;
  wire [7:0] add_779930;
  wire [7:0] sel_779931;
  wire [7:0] add_779934;
  wire [7:0] sel_779935;
  wire [7:0] add_779938;
  wire [7:0] sel_779939;
  wire [7:0] add_779942;
  wire [7:0] sel_779943;
  wire [7:0] add_779946;
  wire [7:0] sel_779947;
  wire [7:0] add_779950;
  wire [7:0] sel_779951;
  wire [7:0] add_779954;
  wire [7:0] sel_779955;
  wire [7:0] add_779958;
  wire [7:0] sel_779959;
  wire [7:0] add_779962;
  wire [7:0] sel_779963;
  wire [7:0] add_779966;
  wire [7:0] sel_779967;
  wire [7:0] add_779970;
  wire [7:0] sel_779971;
  wire [7:0] add_779974;
  wire [7:0] sel_779975;
  wire [7:0] add_779978;
  wire [7:0] sel_779979;
  wire [7:0] add_779982;
  wire [7:0] sel_779983;
  wire [7:0] add_779986;
  wire [7:0] sel_779987;
  wire [7:0] add_779990;
  wire [7:0] sel_779991;
  wire [7:0] add_779994;
  wire [7:0] sel_779995;
  wire [7:0] add_779998;
  wire [7:0] sel_779999;
  wire [7:0] add_780002;
  wire [7:0] sel_780003;
  wire [7:0] add_780006;
  wire [7:0] sel_780007;
  wire [7:0] add_780010;
  wire [7:0] sel_780011;
  wire [7:0] add_780014;
  wire [7:0] sel_780015;
  wire [7:0] add_780018;
  wire [7:0] sel_780019;
  wire [7:0] add_780022;
  wire [7:0] sel_780023;
  wire [7:0] add_780026;
  wire [7:0] sel_780027;
  wire [7:0] add_780030;
  wire [7:0] sel_780031;
  wire [7:0] add_780034;
  wire [7:0] sel_780035;
  wire [7:0] add_780038;
  wire [7:0] sel_780039;
  wire [7:0] add_780042;
  wire [7:0] sel_780043;
  wire [7:0] add_780046;
  wire [7:0] sel_780047;
  wire [7:0] add_780050;
  wire [7:0] sel_780051;
  wire [7:0] add_780054;
  wire [7:0] sel_780055;
  wire [7:0] add_780059;
  wire [15:0] array_index_780060;
  wire [7:0] sel_780061;
  wire [7:0] add_780064;
  wire [7:0] sel_780065;
  wire [7:0] add_780068;
  wire [7:0] sel_780069;
  wire [7:0] add_780072;
  wire [7:0] sel_780073;
  wire [7:0] add_780076;
  wire [7:0] sel_780077;
  wire [7:0] add_780080;
  wire [7:0] sel_780081;
  wire [7:0] add_780084;
  wire [7:0] sel_780085;
  wire [7:0] add_780088;
  wire [7:0] sel_780089;
  wire [7:0] add_780092;
  wire [7:0] sel_780093;
  wire [7:0] add_780096;
  wire [7:0] sel_780097;
  wire [7:0] add_780100;
  wire [7:0] sel_780101;
  wire [7:0] add_780104;
  wire [7:0] sel_780105;
  wire [7:0] add_780108;
  wire [7:0] sel_780109;
  wire [7:0] add_780112;
  wire [7:0] sel_780113;
  wire [7:0] add_780116;
  wire [7:0] sel_780117;
  wire [7:0] add_780120;
  wire [7:0] sel_780121;
  wire [7:0] add_780124;
  wire [7:0] sel_780125;
  wire [7:0] add_780128;
  wire [7:0] sel_780129;
  wire [7:0] add_780132;
  wire [7:0] sel_780133;
  wire [7:0] add_780136;
  wire [7:0] sel_780137;
  wire [7:0] add_780140;
  wire [7:0] sel_780141;
  wire [7:0] add_780144;
  wire [7:0] sel_780145;
  wire [7:0] add_780148;
  wire [7:0] sel_780149;
  wire [7:0] add_780152;
  wire [7:0] sel_780153;
  wire [7:0] add_780156;
  wire [7:0] sel_780157;
  wire [7:0] add_780160;
  wire [7:0] sel_780161;
  wire [7:0] add_780164;
  wire [7:0] sel_780165;
  wire [7:0] add_780168;
  wire [7:0] sel_780169;
  wire [7:0] add_780172;
  wire [7:0] sel_780173;
  wire [7:0] add_780176;
  wire [7:0] sel_780177;
  wire [7:0] add_780180;
  wire [7:0] sel_780181;
  wire [7:0] add_780184;
  wire [7:0] sel_780185;
  wire [7:0] add_780188;
  wire [7:0] sel_780189;
  wire [7:0] add_780192;
  wire [7:0] sel_780193;
  wire [7:0] add_780196;
  wire [7:0] sel_780197;
  wire [7:0] add_780200;
  wire [7:0] sel_780201;
  wire [7:0] add_780204;
  wire [7:0] sel_780205;
  wire [7:0] add_780208;
  wire [7:0] sel_780209;
  wire [7:0] add_780212;
  wire [7:0] sel_780213;
  wire [7:0] add_780216;
  wire [7:0] sel_780217;
  wire [7:0] add_780220;
  wire [7:0] sel_780221;
  wire [7:0] add_780224;
  wire [7:0] sel_780225;
  wire [7:0] add_780228;
  wire [7:0] sel_780229;
  wire [7:0] add_780232;
  wire [7:0] sel_780233;
  wire [7:0] add_780236;
  wire [7:0] sel_780237;
  wire [7:0] add_780240;
  wire [7:0] sel_780241;
  wire [7:0] add_780244;
  wire [7:0] sel_780245;
  wire [7:0] add_780248;
  wire [7:0] sel_780249;
  wire [7:0] add_780252;
  wire [7:0] sel_780253;
  wire [7:0] add_780256;
  wire [7:0] sel_780257;
  wire [7:0] add_780260;
  wire [7:0] sel_780261;
  wire [7:0] add_780264;
  wire [7:0] sel_780265;
  wire [7:0] add_780268;
  wire [7:0] sel_780269;
  wire [7:0] add_780272;
  wire [7:0] sel_780273;
  wire [7:0] add_780276;
  wire [7:0] sel_780277;
  wire [7:0] add_780280;
  wire [7:0] sel_780281;
  wire [7:0] add_780284;
  wire [7:0] sel_780285;
  wire [7:0] add_780288;
  wire [7:0] sel_780289;
  wire [7:0] add_780292;
  wire [7:0] sel_780293;
  wire [7:0] add_780296;
  wire [7:0] sel_780297;
  wire [7:0] add_780300;
  wire [7:0] sel_780301;
  wire [7:0] add_780304;
  wire [7:0] sel_780305;
  wire [7:0] add_780308;
  wire [7:0] sel_780309;
  wire [7:0] add_780312;
  wire [7:0] sel_780313;
  wire [7:0] add_780316;
  wire [7:0] sel_780317;
  wire [7:0] add_780320;
  wire [7:0] sel_780321;
  wire [7:0] add_780324;
  wire [7:0] sel_780325;
  wire [7:0] add_780328;
  wire [7:0] sel_780329;
  wire [7:0] add_780332;
  wire [7:0] sel_780333;
  wire [7:0] add_780336;
  wire [7:0] sel_780337;
  wire [7:0] add_780340;
  wire [7:0] sel_780341;
  wire [7:0] add_780344;
  wire [7:0] sel_780345;
  wire [7:0] add_780348;
  wire [7:0] sel_780349;
  wire [7:0] add_780352;
  wire [7:0] sel_780353;
  wire [7:0] add_780356;
  wire [7:0] sel_780357;
  wire [7:0] add_780360;
  wire [7:0] sel_780361;
  wire [7:0] add_780364;
  wire [7:0] sel_780365;
  wire [7:0] add_780368;
  wire [7:0] sel_780369;
  wire [7:0] add_780372;
  wire [7:0] sel_780373;
  wire [7:0] add_780376;
  wire [7:0] sel_780377;
  wire [7:0] add_780380;
  wire [7:0] sel_780381;
  wire [7:0] add_780384;
  wire [7:0] sel_780385;
  wire [7:0] add_780388;
  wire [7:0] sel_780389;
  wire [7:0] add_780392;
  wire [7:0] sel_780393;
  wire [7:0] add_780396;
  wire [7:0] sel_780397;
  wire [7:0] add_780400;
  wire [7:0] sel_780401;
  wire [7:0] add_780404;
  wire [7:0] sel_780405;
  wire [7:0] add_780408;
  wire [7:0] sel_780409;
  wire [7:0] add_780412;
  wire [7:0] sel_780413;
  wire [7:0] add_780416;
  wire [7:0] sel_780417;
  wire [7:0] add_780421;
  wire [15:0] array_index_780422;
  wire [7:0] sel_780423;
  wire [7:0] add_780426;
  wire [7:0] sel_780427;
  wire [7:0] add_780430;
  wire [7:0] sel_780431;
  wire [7:0] add_780434;
  wire [7:0] sel_780435;
  wire [7:0] add_780438;
  wire [7:0] sel_780439;
  wire [7:0] add_780442;
  wire [7:0] sel_780443;
  wire [7:0] add_780446;
  wire [7:0] sel_780447;
  wire [7:0] add_780450;
  wire [7:0] sel_780451;
  wire [7:0] add_780454;
  wire [7:0] sel_780455;
  wire [7:0] add_780458;
  wire [7:0] sel_780459;
  wire [7:0] add_780462;
  wire [7:0] sel_780463;
  wire [7:0] add_780466;
  wire [7:0] sel_780467;
  wire [7:0] add_780470;
  wire [7:0] sel_780471;
  wire [7:0] add_780474;
  wire [7:0] sel_780475;
  wire [7:0] add_780478;
  wire [7:0] sel_780479;
  wire [7:0] add_780482;
  wire [7:0] sel_780483;
  wire [7:0] add_780486;
  wire [7:0] sel_780487;
  wire [7:0] add_780490;
  wire [7:0] sel_780491;
  wire [7:0] add_780494;
  wire [7:0] sel_780495;
  wire [7:0] add_780498;
  wire [7:0] sel_780499;
  wire [7:0] add_780502;
  wire [7:0] sel_780503;
  wire [7:0] add_780506;
  wire [7:0] sel_780507;
  wire [7:0] add_780510;
  wire [7:0] sel_780511;
  wire [7:0] add_780514;
  wire [7:0] sel_780515;
  wire [7:0] add_780518;
  wire [7:0] sel_780519;
  wire [7:0] add_780522;
  wire [7:0] sel_780523;
  wire [7:0] add_780526;
  wire [7:0] sel_780527;
  wire [7:0] add_780530;
  wire [7:0] sel_780531;
  wire [7:0] add_780534;
  wire [7:0] sel_780535;
  wire [7:0] add_780538;
  wire [7:0] sel_780539;
  wire [7:0] add_780542;
  wire [7:0] sel_780543;
  wire [7:0] add_780546;
  wire [7:0] sel_780547;
  wire [7:0] add_780550;
  wire [7:0] sel_780551;
  wire [7:0] add_780554;
  wire [7:0] sel_780555;
  wire [7:0] add_780558;
  wire [7:0] sel_780559;
  wire [7:0] add_780562;
  wire [7:0] sel_780563;
  wire [7:0] add_780566;
  wire [7:0] sel_780567;
  wire [7:0] add_780570;
  wire [7:0] sel_780571;
  wire [7:0] add_780574;
  wire [7:0] sel_780575;
  wire [7:0] add_780578;
  wire [7:0] sel_780579;
  wire [7:0] add_780582;
  wire [7:0] sel_780583;
  wire [7:0] add_780586;
  wire [7:0] sel_780587;
  wire [7:0] add_780590;
  wire [7:0] sel_780591;
  wire [7:0] add_780594;
  wire [7:0] sel_780595;
  wire [7:0] add_780598;
  wire [7:0] sel_780599;
  wire [7:0] add_780602;
  wire [7:0] sel_780603;
  wire [7:0] add_780606;
  wire [7:0] sel_780607;
  wire [7:0] add_780610;
  wire [7:0] sel_780611;
  wire [7:0] add_780614;
  wire [7:0] sel_780615;
  wire [7:0] add_780618;
  wire [7:0] sel_780619;
  wire [7:0] add_780622;
  wire [7:0] sel_780623;
  wire [7:0] add_780626;
  wire [7:0] sel_780627;
  wire [7:0] add_780630;
  wire [7:0] sel_780631;
  wire [7:0] add_780634;
  wire [7:0] sel_780635;
  wire [7:0] add_780638;
  wire [7:0] sel_780639;
  wire [7:0] add_780642;
  wire [7:0] sel_780643;
  wire [7:0] add_780646;
  wire [7:0] sel_780647;
  wire [7:0] add_780650;
  wire [7:0] sel_780651;
  wire [7:0] add_780654;
  wire [7:0] sel_780655;
  wire [7:0] add_780658;
  wire [7:0] sel_780659;
  wire [7:0] add_780662;
  wire [7:0] sel_780663;
  wire [7:0] add_780666;
  wire [7:0] sel_780667;
  wire [7:0] add_780670;
  wire [7:0] sel_780671;
  wire [7:0] add_780674;
  wire [7:0] sel_780675;
  wire [7:0] add_780678;
  wire [7:0] sel_780679;
  wire [7:0] add_780682;
  wire [7:0] sel_780683;
  wire [7:0] add_780686;
  wire [7:0] sel_780687;
  wire [7:0] add_780690;
  wire [7:0] sel_780691;
  wire [7:0] add_780694;
  wire [7:0] sel_780695;
  wire [7:0] add_780698;
  wire [7:0] sel_780699;
  wire [7:0] add_780702;
  wire [7:0] sel_780703;
  wire [7:0] add_780706;
  wire [7:0] sel_780707;
  wire [7:0] add_780710;
  wire [7:0] sel_780711;
  wire [7:0] add_780714;
  wire [7:0] sel_780715;
  wire [7:0] add_780718;
  wire [7:0] sel_780719;
  wire [7:0] add_780722;
  wire [7:0] sel_780723;
  wire [7:0] add_780726;
  wire [7:0] sel_780727;
  wire [7:0] add_780730;
  wire [7:0] sel_780731;
  wire [7:0] add_780734;
  wire [7:0] sel_780735;
  wire [7:0] add_780738;
  wire [7:0] sel_780739;
  wire [7:0] add_780742;
  wire [7:0] sel_780743;
  wire [7:0] add_780746;
  wire [7:0] sel_780747;
  wire [7:0] add_780750;
  wire [7:0] sel_780751;
  wire [7:0] add_780754;
  wire [7:0] sel_780755;
  wire [7:0] add_780758;
  wire [7:0] sel_780759;
  wire [7:0] add_780762;
  wire [7:0] sel_780763;
  wire [7:0] add_780766;
  wire [7:0] sel_780767;
  wire [7:0] add_780770;
  wire [7:0] sel_780771;
  wire [7:0] add_780774;
  wire [7:0] sel_780775;
  wire [7:0] add_780778;
  wire [7:0] sel_780779;
  wire [7:0] add_780783;
  wire [15:0] array_index_780784;
  wire [7:0] sel_780785;
  wire [7:0] add_780788;
  wire [7:0] sel_780789;
  wire [7:0] add_780792;
  wire [7:0] sel_780793;
  wire [7:0] add_780796;
  wire [7:0] sel_780797;
  wire [7:0] add_780800;
  wire [7:0] sel_780801;
  wire [7:0] add_780804;
  wire [7:0] sel_780805;
  wire [7:0] add_780808;
  wire [7:0] sel_780809;
  wire [7:0] add_780812;
  wire [7:0] sel_780813;
  wire [7:0] add_780816;
  wire [7:0] sel_780817;
  wire [7:0] add_780820;
  wire [7:0] sel_780821;
  wire [7:0] add_780824;
  wire [7:0] sel_780825;
  wire [7:0] add_780828;
  wire [7:0] sel_780829;
  wire [7:0] add_780832;
  wire [7:0] sel_780833;
  wire [7:0] add_780836;
  wire [7:0] sel_780837;
  wire [7:0] add_780840;
  wire [7:0] sel_780841;
  wire [7:0] add_780844;
  wire [7:0] sel_780845;
  wire [7:0] add_780848;
  wire [7:0] sel_780849;
  wire [7:0] add_780852;
  wire [7:0] sel_780853;
  wire [7:0] add_780856;
  wire [7:0] sel_780857;
  wire [7:0] add_780860;
  wire [7:0] sel_780861;
  wire [7:0] add_780864;
  wire [7:0] sel_780865;
  wire [7:0] add_780868;
  wire [7:0] sel_780869;
  wire [7:0] add_780872;
  wire [7:0] sel_780873;
  wire [7:0] add_780876;
  wire [7:0] sel_780877;
  wire [7:0] add_780880;
  wire [7:0] sel_780881;
  wire [7:0] add_780884;
  wire [7:0] sel_780885;
  wire [7:0] add_780888;
  wire [7:0] sel_780889;
  wire [7:0] add_780892;
  wire [7:0] sel_780893;
  wire [7:0] add_780896;
  wire [7:0] sel_780897;
  wire [7:0] add_780900;
  wire [7:0] sel_780901;
  wire [7:0] add_780904;
  wire [7:0] sel_780905;
  wire [7:0] add_780908;
  wire [7:0] sel_780909;
  wire [7:0] add_780912;
  wire [7:0] sel_780913;
  wire [7:0] add_780916;
  wire [7:0] sel_780917;
  wire [7:0] add_780920;
  wire [7:0] sel_780921;
  wire [7:0] add_780924;
  wire [7:0] sel_780925;
  wire [7:0] add_780928;
  wire [7:0] sel_780929;
  wire [7:0] add_780932;
  wire [7:0] sel_780933;
  wire [7:0] add_780936;
  wire [7:0] sel_780937;
  wire [7:0] add_780940;
  wire [7:0] sel_780941;
  wire [7:0] add_780944;
  wire [7:0] sel_780945;
  wire [7:0] add_780948;
  wire [7:0] sel_780949;
  wire [7:0] add_780952;
  wire [7:0] sel_780953;
  wire [7:0] add_780956;
  wire [7:0] sel_780957;
  wire [7:0] add_780960;
  wire [7:0] sel_780961;
  wire [7:0] add_780964;
  wire [7:0] sel_780965;
  wire [7:0] add_780968;
  wire [7:0] sel_780969;
  wire [7:0] add_780972;
  wire [7:0] sel_780973;
  wire [7:0] add_780976;
  wire [7:0] sel_780977;
  wire [7:0] add_780980;
  wire [7:0] sel_780981;
  wire [7:0] add_780984;
  wire [7:0] sel_780985;
  wire [7:0] add_780988;
  wire [7:0] sel_780989;
  wire [7:0] add_780992;
  wire [7:0] sel_780993;
  wire [7:0] add_780996;
  wire [7:0] sel_780997;
  wire [7:0] add_781000;
  wire [7:0] sel_781001;
  wire [7:0] add_781004;
  wire [7:0] sel_781005;
  wire [7:0] add_781008;
  wire [7:0] sel_781009;
  wire [7:0] add_781012;
  wire [7:0] sel_781013;
  wire [7:0] add_781016;
  wire [7:0] sel_781017;
  wire [7:0] add_781020;
  wire [7:0] sel_781021;
  wire [7:0] add_781024;
  wire [7:0] sel_781025;
  wire [7:0] add_781028;
  wire [7:0] sel_781029;
  wire [7:0] add_781032;
  wire [7:0] sel_781033;
  wire [7:0] add_781036;
  wire [7:0] sel_781037;
  wire [7:0] add_781040;
  wire [7:0] sel_781041;
  wire [7:0] add_781044;
  wire [7:0] sel_781045;
  wire [7:0] add_781048;
  wire [7:0] sel_781049;
  wire [7:0] add_781052;
  wire [7:0] sel_781053;
  wire [7:0] add_781056;
  wire [7:0] sel_781057;
  wire [7:0] add_781060;
  wire [7:0] sel_781061;
  wire [7:0] add_781064;
  wire [7:0] sel_781065;
  wire [7:0] add_781068;
  wire [7:0] sel_781069;
  wire [7:0] add_781072;
  wire [7:0] sel_781073;
  wire [7:0] add_781076;
  wire [7:0] sel_781077;
  wire [7:0] add_781080;
  wire [7:0] sel_781081;
  wire [7:0] add_781084;
  wire [7:0] sel_781085;
  wire [7:0] add_781088;
  wire [7:0] sel_781089;
  wire [7:0] add_781092;
  wire [7:0] sel_781093;
  wire [7:0] add_781096;
  wire [7:0] sel_781097;
  wire [7:0] add_781100;
  wire [7:0] sel_781101;
  wire [7:0] add_781104;
  wire [7:0] sel_781105;
  wire [7:0] add_781108;
  wire [7:0] sel_781109;
  wire [7:0] add_781112;
  wire [7:0] sel_781113;
  wire [7:0] add_781116;
  wire [7:0] sel_781117;
  wire [7:0] add_781120;
  wire [7:0] sel_781121;
  wire [7:0] add_781124;
  wire [7:0] sel_781125;
  wire [7:0] add_781128;
  wire [7:0] sel_781129;
  wire [7:0] add_781132;
  wire [7:0] sel_781133;
  wire [7:0] add_781136;
  wire [7:0] sel_781137;
  wire [7:0] add_781140;
  wire [7:0] sel_781141;
  wire [7:0] add_781145;
  wire [15:0] array_index_781146;
  wire [7:0] sel_781147;
  wire [7:0] add_781150;
  wire [7:0] sel_781151;
  wire [7:0] add_781154;
  wire [7:0] sel_781155;
  wire [7:0] add_781158;
  wire [7:0] sel_781159;
  wire [7:0] add_781162;
  wire [7:0] sel_781163;
  wire [7:0] add_781166;
  wire [7:0] sel_781167;
  wire [7:0] add_781170;
  wire [7:0] sel_781171;
  wire [7:0] add_781174;
  wire [7:0] sel_781175;
  wire [7:0] add_781178;
  wire [7:0] sel_781179;
  wire [7:0] add_781182;
  wire [7:0] sel_781183;
  wire [7:0] add_781186;
  wire [7:0] sel_781187;
  wire [7:0] add_781190;
  wire [7:0] sel_781191;
  wire [7:0] add_781194;
  wire [7:0] sel_781195;
  wire [7:0] add_781198;
  wire [7:0] sel_781199;
  wire [7:0] add_781202;
  wire [7:0] sel_781203;
  wire [7:0] add_781206;
  wire [7:0] sel_781207;
  wire [7:0] add_781210;
  wire [7:0] sel_781211;
  wire [7:0] add_781214;
  wire [7:0] sel_781215;
  wire [7:0] add_781218;
  wire [7:0] sel_781219;
  wire [7:0] add_781222;
  wire [7:0] sel_781223;
  wire [7:0] add_781226;
  wire [7:0] sel_781227;
  wire [7:0] add_781230;
  wire [7:0] sel_781231;
  wire [7:0] add_781234;
  wire [7:0] sel_781235;
  wire [7:0] add_781238;
  wire [7:0] sel_781239;
  wire [7:0] add_781242;
  wire [7:0] sel_781243;
  wire [7:0] add_781246;
  wire [7:0] sel_781247;
  wire [7:0] add_781250;
  wire [7:0] sel_781251;
  wire [7:0] add_781254;
  wire [7:0] sel_781255;
  wire [7:0] add_781258;
  wire [7:0] sel_781259;
  wire [7:0] add_781262;
  wire [7:0] sel_781263;
  wire [7:0] add_781266;
  wire [7:0] sel_781267;
  wire [7:0] add_781270;
  wire [7:0] sel_781271;
  wire [7:0] add_781274;
  wire [7:0] sel_781275;
  wire [7:0] add_781278;
  wire [7:0] sel_781279;
  wire [7:0] add_781282;
  wire [7:0] sel_781283;
  wire [7:0] add_781286;
  wire [7:0] sel_781287;
  wire [7:0] add_781290;
  wire [7:0] sel_781291;
  wire [7:0] add_781294;
  wire [7:0] sel_781295;
  wire [7:0] add_781298;
  wire [7:0] sel_781299;
  wire [7:0] add_781302;
  wire [7:0] sel_781303;
  wire [7:0] add_781306;
  wire [7:0] sel_781307;
  wire [7:0] add_781310;
  wire [7:0] sel_781311;
  wire [7:0] add_781314;
  wire [7:0] sel_781315;
  wire [7:0] add_781318;
  wire [7:0] sel_781319;
  wire [7:0] add_781322;
  wire [7:0] sel_781323;
  wire [7:0] add_781326;
  wire [7:0] sel_781327;
  wire [7:0] add_781330;
  wire [7:0] sel_781331;
  wire [7:0] add_781334;
  wire [7:0] sel_781335;
  wire [7:0] add_781338;
  wire [7:0] sel_781339;
  wire [7:0] add_781342;
  wire [7:0] sel_781343;
  wire [7:0] add_781346;
  wire [7:0] sel_781347;
  wire [7:0] add_781350;
  wire [7:0] sel_781351;
  wire [7:0] add_781354;
  wire [7:0] sel_781355;
  wire [7:0] add_781358;
  wire [7:0] sel_781359;
  wire [7:0] add_781362;
  wire [7:0] sel_781363;
  wire [7:0] add_781366;
  wire [7:0] sel_781367;
  wire [7:0] add_781370;
  wire [7:0] sel_781371;
  wire [7:0] add_781374;
  wire [7:0] sel_781375;
  wire [7:0] add_781378;
  wire [7:0] sel_781379;
  wire [7:0] add_781382;
  wire [7:0] sel_781383;
  wire [7:0] add_781386;
  wire [7:0] sel_781387;
  wire [7:0] add_781390;
  wire [7:0] sel_781391;
  wire [7:0] add_781394;
  wire [7:0] sel_781395;
  wire [7:0] add_781398;
  wire [7:0] sel_781399;
  wire [7:0] add_781402;
  wire [7:0] sel_781403;
  wire [7:0] add_781406;
  wire [7:0] sel_781407;
  wire [7:0] add_781410;
  wire [7:0] sel_781411;
  wire [7:0] add_781414;
  wire [7:0] sel_781415;
  wire [7:0] add_781418;
  wire [7:0] sel_781419;
  wire [7:0] add_781422;
  wire [7:0] sel_781423;
  wire [7:0] add_781426;
  wire [7:0] sel_781427;
  wire [7:0] add_781430;
  wire [7:0] sel_781431;
  wire [7:0] add_781434;
  wire [7:0] sel_781435;
  wire [7:0] add_781438;
  wire [7:0] sel_781439;
  wire [7:0] add_781442;
  wire [7:0] sel_781443;
  wire [7:0] add_781446;
  wire [7:0] sel_781447;
  wire [7:0] add_781450;
  wire [7:0] sel_781451;
  wire [7:0] add_781454;
  wire [7:0] sel_781455;
  wire [7:0] add_781458;
  wire [7:0] sel_781459;
  wire [7:0] add_781462;
  wire [7:0] sel_781463;
  wire [7:0] add_781466;
  wire [7:0] sel_781467;
  wire [7:0] add_781470;
  wire [7:0] sel_781471;
  wire [7:0] add_781474;
  wire [7:0] sel_781475;
  wire [7:0] add_781478;
  wire [7:0] sel_781479;
  wire [7:0] add_781482;
  wire [7:0] sel_781483;
  wire [7:0] add_781486;
  wire [7:0] sel_781487;
  wire [7:0] add_781490;
  wire [7:0] sel_781491;
  wire [7:0] add_781494;
  wire [7:0] sel_781495;
  wire [7:0] add_781498;
  wire [7:0] sel_781499;
  wire [7:0] add_781502;
  wire [7:0] sel_781503;
  wire [7:0] add_781507;
  wire [15:0] array_index_781508;
  wire [7:0] sel_781509;
  wire [7:0] add_781512;
  wire [7:0] sel_781513;
  wire [7:0] add_781516;
  wire [7:0] sel_781517;
  wire [7:0] add_781520;
  wire [7:0] sel_781521;
  wire [7:0] add_781524;
  wire [7:0] sel_781525;
  wire [7:0] add_781528;
  wire [7:0] sel_781529;
  wire [7:0] add_781532;
  wire [7:0] sel_781533;
  wire [7:0] add_781536;
  wire [7:0] sel_781537;
  wire [7:0] add_781540;
  wire [7:0] sel_781541;
  wire [7:0] add_781544;
  wire [7:0] sel_781545;
  wire [7:0] add_781548;
  wire [7:0] sel_781549;
  wire [7:0] add_781552;
  wire [7:0] sel_781553;
  wire [7:0] add_781556;
  wire [7:0] sel_781557;
  wire [7:0] add_781560;
  wire [7:0] sel_781561;
  wire [7:0] add_781564;
  wire [7:0] sel_781565;
  wire [7:0] add_781568;
  wire [7:0] sel_781569;
  wire [7:0] add_781572;
  wire [7:0] sel_781573;
  wire [7:0] add_781576;
  wire [7:0] sel_781577;
  wire [7:0] add_781580;
  wire [7:0] sel_781581;
  wire [7:0] add_781584;
  wire [7:0] sel_781585;
  wire [7:0] add_781588;
  wire [7:0] sel_781589;
  wire [7:0] add_781592;
  wire [7:0] sel_781593;
  wire [7:0] add_781596;
  wire [7:0] sel_781597;
  wire [7:0] add_781600;
  wire [7:0] sel_781601;
  wire [7:0] add_781604;
  wire [7:0] sel_781605;
  wire [7:0] add_781608;
  wire [7:0] sel_781609;
  wire [7:0] add_781612;
  wire [7:0] sel_781613;
  wire [7:0] add_781616;
  wire [7:0] sel_781617;
  wire [7:0] add_781620;
  wire [7:0] sel_781621;
  wire [7:0] add_781624;
  wire [7:0] sel_781625;
  wire [7:0] add_781628;
  wire [7:0] sel_781629;
  wire [7:0] add_781632;
  wire [7:0] sel_781633;
  wire [7:0] add_781636;
  wire [7:0] sel_781637;
  wire [7:0] add_781640;
  wire [7:0] sel_781641;
  wire [7:0] add_781644;
  wire [7:0] sel_781645;
  wire [7:0] add_781648;
  wire [7:0] sel_781649;
  wire [7:0] add_781652;
  wire [7:0] sel_781653;
  wire [7:0] add_781656;
  wire [7:0] sel_781657;
  wire [7:0] add_781660;
  wire [7:0] sel_781661;
  wire [7:0] add_781664;
  wire [7:0] sel_781665;
  wire [7:0] add_781668;
  wire [7:0] sel_781669;
  wire [7:0] add_781672;
  wire [7:0] sel_781673;
  wire [7:0] add_781676;
  wire [7:0] sel_781677;
  wire [7:0] add_781680;
  wire [7:0] sel_781681;
  wire [7:0] add_781684;
  wire [7:0] sel_781685;
  wire [7:0] add_781688;
  wire [7:0] sel_781689;
  wire [7:0] add_781692;
  wire [7:0] sel_781693;
  wire [7:0] add_781696;
  wire [7:0] sel_781697;
  wire [7:0] add_781700;
  wire [7:0] sel_781701;
  wire [7:0] add_781704;
  wire [7:0] sel_781705;
  wire [7:0] add_781708;
  wire [7:0] sel_781709;
  wire [7:0] add_781712;
  wire [7:0] sel_781713;
  wire [7:0] add_781716;
  wire [7:0] sel_781717;
  wire [7:0] add_781720;
  wire [7:0] sel_781721;
  wire [7:0] add_781724;
  wire [7:0] sel_781725;
  wire [7:0] add_781728;
  wire [7:0] sel_781729;
  wire [7:0] add_781732;
  wire [7:0] sel_781733;
  wire [7:0] add_781736;
  wire [7:0] sel_781737;
  wire [7:0] add_781740;
  wire [7:0] sel_781741;
  wire [7:0] add_781744;
  wire [7:0] sel_781745;
  wire [7:0] add_781748;
  wire [7:0] sel_781749;
  wire [7:0] add_781752;
  wire [7:0] sel_781753;
  wire [7:0] add_781756;
  wire [7:0] sel_781757;
  wire [7:0] add_781760;
  wire [7:0] sel_781761;
  wire [7:0] add_781764;
  wire [7:0] sel_781765;
  wire [7:0] add_781768;
  wire [7:0] sel_781769;
  wire [7:0] add_781772;
  wire [7:0] sel_781773;
  wire [7:0] add_781776;
  wire [7:0] sel_781777;
  wire [7:0] add_781780;
  wire [7:0] sel_781781;
  wire [7:0] add_781784;
  wire [7:0] sel_781785;
  wire [7:0] add_781788;
  wire [7:0] sel_781789;
  wire [7:0] add_781792;
  wire [7:0] sel_781793;
  wire [7:0] add_781796;
  wire [7:0] sel_781797;
  wire [7:0] add_781800;
  wire [7:0] sel_781801;
  wire [7:0] add_781804;
  wire [7:0] sel_781805;
  wire [7:0] add_781808;
  wire [7:0] sel_781809;
  wire [7:0] add_781812;
  wire [7:0] sel_781813;
  wire [7:0] add_781816;
  wire [7:0] sel_781817;
  wire [7:0] add_781820;
  wire [7:0] sel_781821;
  wire [7:0] add_781824;
  wire [7:0] sel_781825;
  wire [7:0] add_781828;
  wire [7:0] sel_781829;
  wire [7:0] add_781832;
  wire [7:0] sel_781833;
  wire [7:0] add_781836;
  wire [7:0] sel_781837;
  wire [7:0] add_781840;
  wire [7:0] sel_781841;
  wire [7:0] add_781844;
  wire [7:0] sel_781845;
  wire [7:0] add_781848;
  wire [7:0] sel_781849;
  wire [7:0] add_781852;
  wire [7:0] sel_781853;
  wire [7:0] add_781856;
  wire [7:0] sel_781857;
  wire [7:0] add_781860;
  wire [7:0] sel_781861;
  wire [7:0] add_781864;
  wire [7:0] sel_781865;
  wire [7:0] add_781869;
  wire [15:0] array_index_781870;
  wire [7:0] sel_781871;
  wire [7:0] add_781874;
  wire [7:0] sel_781875;
  wire [7:0] add_781878;
  wire [7:0] sel_781879;
  wire [7:0] add_781882;
  wire [7:0] sel_781883;
  wire [7:0] add_781886;
  wire [7:0] sel_781887;
  wire [7:0] add_781890;
  wire [7:0] sel_781891;
  wire [7:0] add_781894;
  wire [7:0] sel_781895;
  wire [7:0] add_781898;
  wire [7:0] sel_781899;
  wire [7:0] add_781902;
  wire [7:0] sel_781903;
  wire [7:0] add_781906;
  wire [7:0] sel_781907;
  wire [7:0] add_781910;
  wire [7:0] sel_781911;
  wire [7:0] add_781914;
  wire [7:0] sel_781915;
  wire [7:0] add_781918;
  wire [7:0] sel_781919;
  wire [7:0] add_781922;
  wire [7:0] sel_781923;
  wire [7:0] add_781926;
  wire [7:0] sel_781927;
  wire [7:0] add_781930;
  wire [7:0] sel_781931;
  wire [7:0] add_781934;
  wire [7:0] sel_781935;
  wire [7:0] add_781938;
  wire [7:0] sel_781939;
  wire [7:0] add_781942;
  wire [7:0] sel_781943;
  wire [7:0] add_781946;
  wire [7:0] sel_781947;
  wire [7:0] add_781950;
  wire [7:0] sel_781951;
  wire [7:0] add_781954;
  wire [7:0] sel_781955;
  wire [7:0] add_781958;
  wire [7:0] sel_781959;
  wire [7:0] add_781962;
  wire [7:0] sel_781963;
  wire [7:0] add_781966;
  wire [7:0] sel_781967;
  wire [7:0] add_781970;
  wire [7:0] sel_781971;
  wire [7:0] add_781974;
  wire [7:0] sel_781975;
  wire [7:0] add_781978;
  wire [7:0] sel_781979;
  wire [7:0] add_781982;
  wire [7:0] sel_781983;
  wire [7:0] add_781986;
  wire [7:0] sel_781987;
  wire [7:0] add_781990;
  wire [7:0] sel_781991;
  wire [7:0] add_781994;
  wire [7:0] sel_781995;
  wire [7:0] add_781998;
  wire [7:0] sel_781999;
  wire [7:0] add_782002;
  wire [7:0] sel_782003;
  wire [7:0] add_782006;
  wire [7:0] sel_782007;
  wire [7:0] add_782010;
  wire [7:0] sel_782011;
  wire [7:0] add_782014;
  wire [7:0] sel_782015;
  wire [7:0] add_782018;
  wire [7:0] sel_782019;
  wire [7:0] add_782022;
  wire [7:0] sel_782023;
  wire [7:0] add_782026;
  wire [7:0] sel_782027;
  wire [7:0] add_782030;
  wire [7:0] sel_782031;
  wire [7:0] add_782034;
  wire [7:0] sel_782035;
  wire [7:0] add_782038;
  wire [7:0] sel_782039;
  wire [7:0] add_782042;
  wire [7:0] sel_782043;
  wire [7:0] add_782046;
  wire [7:0] sel_782047;
  wire [7:0] add_782050;
  wire [7:0] sel_782051;
  wire [7:0] add_782054;
  wire [7:0] sel_782055;
  wire [7:0] add_782058;
  wire [7:0] sel_782059;
  wire [7:0] add_782062;
  wire [7:0] sel_782063;
  wire [7:0] add_782066;
  wire [7:0] sel_782067;
  wire [7:0] add_782070;
  wire [7:0] sel_782071;
  wire [7:0] add_782074;
  wire [7:0] sel_782075;
  wire [7:0] add_782078;
  wire [7:0] sel_782079;
  wire [7:0] add_782082;
  wire [7:0] sel_782083;
  wire [7:0] add_782086;
  wire [7:0] sel_782087;
  wire [7:0] add_782090;
  wire [7:0] sel_782091;
  wire [7:0] add_782094;
  wire [7:0] sel_782095;
  wire [7:0] add_782098;
  wire [7:0] sel_782099;
  wire [7:0] add_782102;
  wire [7:0] sel_782103;
  wire [7:0] add_782106;
  wire [7:0] sel_782107;
  wire [7:0] add_782110;
  wire [7:0] sel_782111;
  wire [7:0] add_782114;
  wire [7:0] sel_782115;
  wire [7:0] add_782118;
  wire [7:0] sel_782119;
  wire [7:0] add_782122;
  wire [7:0] sel_782123;
  wire [7:0] add_782126;
  wire [7:0] sel_782127;
  wire [7:0] add_782130;
  wire [7:0] sel_782131;
  wire [7:0] add_782134;
  wire [7:0] sel_782135;
  wire [7:0] add_782138;
  wire [7:0] sel_782139;
  wire [7:0] add_782142;
  wire [7:0] sel_782143;
  wire [7:0] add_782146;
  wire [7:0] sel_782147;
  wire [7:0] add_782150;
  wire [7:0] sel_782151;
  wire [7:0] add_782154;
  wire [7:0] sel_782155;
  wire [7:0] add_782158;
  wire [7:0] sel_782159;
  wire [7:0] add_782162;
  wire [7:0] sel_782163;
  wire [7:0] add_782166;
  wire [7:0] sel_782167;
  wire [7:0] add_782170;
  wire [7:0] sel_782171;
  wire [7:0] add_782174;
  wire [7:0] sel_782175;
  wire [7:0] add_782178;
  wire [7:0] sel_782179;
  wire [7:0] add_782182;
  wire [7:0] sel_782183;
  wire [7:0] add_782186;
  wire [7:0] sel_782187;
  wire [7:0] add_782190;
  wire [7:0] sel_782191;
  wire [7:0] add_782194;
  wire [7:0] sel_782195;
  wire [7:0] add_782198;
  wire [7:0] sel_782199;
  wire [7:0] add_782202;
  wire [7:0] sel_782203;
  wire [7:0] add_782206;
  wire [7:0] sel_782207;
  wire [7:0] add_782210;
  wire [7:0] sel_782211;
  wire [7:0] add_782214;
  wire [7:0] sel_782215;
  wire [7:0] add_782218;
  wire [7:0] sel_782219;
  wire [7:0] add_782222;
  wire [7:0] sel_782223;
  wire [7:0] add_782226;
  wire [7:0] sel_782227;
  wire [7:0] add_782231;
  wire [15:0] array_index_782232;
  wire [7:0] sel_782233;
  wire [7:0] add_782236;
  wire [7:0] sel_782237;
  wire [7:0] add_782240;
  wire [7:0] sel_782241;
  wire [7:0] add_782244;
  wire [7:0] sel_782245;
  wire [7:0] add_782248;
  wire [7:0] sel_782249;
  wire [7:0] add_782252;
  wire [7:0] sel_782253;
  wire [7:0] add_782256;
  wire [7:0] sel_782257;
  wire [7:0] add_782260;
  wire [7:0] sel_782261;
  wire [7:0] add_782264;
  wire [7:0] sel_782265;
  wire [7:0] add_782268;
  wire [7:0] sel_782269;
  wire [7:0] add_782272;
  wire [7:0] sel_782273;
  wire [7:0] add_782276;
  wire [7:0] sel_782277;
  wire [7:0] add_782280;
  wire [7:0] sel_782281;
  wire [7:0] add_782284;
  wire [7:0] sel_782285;
  wire [7:0] add_782288;
  wire [7:0] sel_782289;
  wire [7:0] add_782292;
  wire [7:0] sel_782293;
  wire [7:0] add_782296;
  wire [7:0] sel_782297;
  wire [7:0] add_782300;
  wire [7:0] sel_782301;
  wire [7:0] add_782304;
  wire [7:0] sel_782305;
  wire [7:0] add_782308;
  wire [7:0] sel_782309;
  wire [7:0] add_782312;
  wire [7:0] sel_782313;
  wire [7:0] add_782316;
  wire [7:0] sel_782317;
  wire [7:0] add_782320;
  wire [7:0] sel_782321;
  wire [7:0] add_782324;
  wire [7:0] sel_782325;
  wire [7:0] add_782328;
  wire [7:0] sel_782329;
  wire [7:0] add_782332;
  wire [7:0] sel_782333;
  wire [7:0] add_782336;
  wire [7:0] sel_782337;
  wire [7:0] add_782340;
  wire [7:0] sel_782341;
  wire [7:0] add_782344;
  wire [7:0] sel_782345;
  wire [7:0] add_782348;
  wire [7:0] sel_782349;
  wire [7:0] add_782352;
  wire [7:0] sel_782353;
  wire [7:0] add_782356;
  wire [7:0] sel_782357;
  wire [7:0] add_782360;
  wire [7:0] sel_782361;
  wire [7:0] add_782364;
  wire [7:0] sel_782365;
  wire [7:0] add_782368;
  wire [7:0] sel_782369;
  wire [7:0] add_782372;
  wire [7:0] sel_782373;
  wire [7:0] add_782376;
  wire [7:0] sel_782377;
  wire [7:0] add_782380;
  wire [7:0] sel_782381;
  wire [7:0] add_782384;
  wire [7:0] sel_782385;
  wire [7:0] add_782388;
  wire [7:0] sel_782389;
  wire [7:0] add_782392;
  wire [7:0] sel_782393;
  wire [7:0] add_782396;
  wire [7:0] sel_782397;
  wire [7:0] add_782400;
  wire [7:0] sel_782401;
  wire [7:0] add_782404;
  wire [7:0] sel_782405;
  wire [7:0] add_782408;
  wire [7:0] sel_782409;
  wire [7:0] add_782412;
  wire [7:0] sel_782413;
  wire [7:0] add_782416;
  wire [7:0] sel_782417;
  wire [7:0] add_782420;
  wire [7:0] sel_782421;
  wire [7:0] add_782424;
  wire [7:0] sel_782425;
  wire [7:0] add_782428;
  wire [7:0] sel_782429;
  wire [7:0] add_782432;
  wire [7:0] sel_782433;
  wire [7:0] add_782436;
  wire [7:0] sel_782437;
  wire [7:0] add_782440;
  wire [7:0] sel_782441;
  wire [7:0] add_782444;
  wire [7:0] sel_782445;
  wire [7:0] add_782448;
  wire [7:0] sel_782449;
  wire [7:0] add_782452;
  wire [7:0] sel_782453;
  wire [7:0] add_782456;
  wire [7:0] sel_782457;
  wire [7:0] add_782460;
  wire [7:0] sel_782461;
  wire [7:0] add_782464;
  wire [7:0] sel_782465;
  wire [7:0] add_782468;
  wire [7:0] sel_782469;
  wire [7:0] add_782472;
  wire [7:0] sel_782473;
  wire [7:0] add_782476;
  wire [7:0] sel_782477;
  wire [7:0] add_782480;
  wire [7:0] sel_782481;
  wire [7:0] add_782484;
  wire [7:0] sel_782485;
  wire [7:0] add_782488;
  wire [7:0] sel_782489;
  wire [7:0] add_782492;
  wire [7:0] sel_782493;
  wire [7:0] add_782496;
  wire [7:0] sel_782497;
  wire [7:0] add_782500;
  wire [7:0] sel_782501;
  wire [7:0] add_782504;
  wire [7:0] sel_782505;
  wire [7:0] add_782508;
  wire [7:0] sel_782509;
  wire [7:0] add_782512;
  wire [7:0] sel_782513;
  wire [7:0] add_782516;
  wire [7:0] sel_782517;
  wire [7:0] add_782520;
  wire [7:0] sel_782521;
  wire [7:0] add_782524;
  wire [7:0] sel_782525;
  wire [7:0] add_782528;
  wire [7:0] sel_782529;
  wire [7:0] add_782532;
  wire [7:0] sel_782533;
  wire [7:0] add_782536;
  wire [7:0] sel_782537;
  wire [7:0] add_782540;
  wire [7:0] sel_782541;
  wire [7:0] add_782544;
  wire [7:0] sel_782545;
  wire [7:0] add_782548;
  wire [7:0] sel_782549;
  wire [7:0] add_782552;
  wire [7:0] sel_782553;
  wire [7:0] add_782556;
  wire [7:0] sel_782557;
  wire [7:0] add_782560;
  wire [7:0] sel_782561;
  wire [7:0] add_782564;
  wire [7:0] sel_782565;
  wire [7:0] add_782568;
  wire [7:0] sel_782569;
  wire [7:0] add_782572;
  wire [7:0] sel_782573;
  wire [7:0] add_782576;
  wire [7:0] sel_782577;
  wire [7:0] add_782580;
  wire [7:0] sel_782581;
  wire [7:0] add_782584;
  wire [7:0] sel_782585;
  wire [7:0] add_782588;
  wire [7:0] sel_782589;
  wire [7:0] add_782593;
  wire [15:0] array_index_782594;
  wire [7:0] sel_782595;
  wire [7:0] add_782598;
  wire [7:0] sel_782599;
  wire [7:0] add_782602;
  wire [7:0] sel_782603;
  wire [7:0] add_782606;
  wire [7:0] sel_782607;
  wire [7:0] add_782610;
  wire [7:0] sel_782611;
  wire [7:0] add_782614;
  wire [7:0] sel_782615;
  wire [7:0] add_782618;
  wire [7:0] sel_782619;
  wire [7:0] add_782622;
  wire [7:0] sel_782623;
  wire [7:0] add_782626;
  wire [7:0] sel_782627;
  wire [7:0] add_782630;
  wire [7:0] sel_782631;
  wire [7:0] add_782634;
  wire [7:0] sel_782635;
  wire [7:0] add_782638;
  wire [7:0] sel_782639;
  wire [7:0] add_782642;
  wire [7:0] sel_782643;
  wire [7:0] add_782646;
  wire [7:0] sel_782647;
  wire [7:0] add_782650;
  wire [7:0] sel_782651;
  wire [7:0] add_782654;
  wire [7:0] sel_782655;
  wire [7:0] add_782658;
  wire [7:0] sel_782659;
  wire [7:0] add_782662;
  wire [7:0] sel_782663;
  wire [7:0] add_782666;
  wire [7:0] sel_782667;
  wire [7:0] add_782670;
  wire [7:0] sel_782671;
  wire [7:0] add_782674;
  wire [7:0] sel_782675;
  wire [7:0] add_782678;
  wire [7:0] sel_782679;
  wire [7:0] add_782682;
  wire [7:0] sel_782683;
  wire [7:0] add_782686;
  wire [7:0] sel_782687;
  wire [7:0] add_782690;
  wire [7:0] sel_782691;
  wire [7:0] add_782694;
  wire [7:0] sel_782695;
  wire [7:0] add_782698;
  wire [7:0] sel_782699;
  wire [7:0] add_782702;
  wire [7:0] sel_782703;
  wire [7:0] add_782706;
  wire [7:0] sel_782707;
  wire [7:0] add_782710;
  wire [7:0] sel_782711;
  wire [7:0] add_782714;
  wire [7:0] sel_782715;
  wire [7:0] add_782718;
  wire [7:0] sel_782719;
  wire [7:0] add_782722;
  wire [7:0] sel_782723;
  wire [7:0] add_782726;
  wire [7:0] sel_782727;
  wire [7:0] add_782730;
  wire [7:0] sel_782731;
  wire [7:0] add_782734;
  wire [7:0] sel_782735;
  wire [7:0] add_782738;
  wire [7:0] sel_782739;
  wire [7:0] add_782742;
  wire [7:0] sel_782743;
  wire [7:0] add_782746;
  wire [7:0] sel_782747;
  wire [7:0] add_782750;
  wire [7:0] sel_782751;
  wire [7:0] add_782754;
  wire [7:0] sel_782755;
  wire [7:0] add_782758;
  wire [7:0] sel_782759;
  wire [7:0] add_782762;
  wire [7:0] sel_782763;
  wire [7:0] add_782766;
  wire [7:0] sel_782767;
  wire [7:0] add_782770;
  wire [7:0] sel_782771;
  wire [7:0] add_782774;
  wire [7:0] sel_782775;
  wire [7:0] add_782778;
  wire [7:0] sel_782779;
  wire [7:0] add_782782;
  wire [7:0] sel_782783;
  wire [7:0] add_782786;
  wire [7:0] sel_782787;
  wire [7:0] add_782790;
  wire [7:0] sel_782791;
  wire [7:0] add_782794;
  wire [7:0] sel_782795;
  wire [7:0] add_782798;
  wire [7:0] sel_782799;
  wire [7:0] add_782802;
  wire [7:0] sel_782803;
  wire [7:0] add_782806;
  wire [7:0] sel_782807;
  wire [7:0] add_782810;
  wire [7:0] sel_782811;
  wire [7:0] add_782814;
  wire [7:0] sel_782815;
  wire [7:0] add_782818;
  wire [7:0] sel_782819;
  wire [7:0] add_782822;
  wire [7:0] sel_782823;
  wire [7:0] add_782826;
  wire [7:0] sel_782827;
  wire [7:0] add_782830;
  wire [7:0] sel_782831;
  wire [7:0] add_782834;
  wire [7:0] sel_782835;
  wire [7:0] add_782838;
  wire [7:0] sel_782839;
  wire [7:0] add_782842;
  wire [7:0] sel_782843;
  wire [7:0] add_782846;
  wire [7:0] sel_782847;
  wire [7:0] add_782850;
  wire [7:0] sel_782851;
  wire [7:0] add_782854;
  wire [7:0] sel_782855;
  wire [7:0] add_782858;
  wire [7:0] sel_782859;
  wire [7:0] add_782862;
  wire [7:0] sel_782863;
  wire [7:0] add_782866;
  wire [7:0] sel_782867;
  wire [7:0] add_782870;
  wire [7:0] sel_782871;
  wire [7:0] add_782874;
  wire [7:0] sel_782875;
  wire [7:0] add_782878;
  wire [7:0] sel_782879;
  wire [7:0] add_782882;
  wire [7:0] sel_782883;
  wire [7:0] add_782886;
  wire [7:0] sel_782887;
  wire [7:0] add_782890;
  wire [7:0] sel_782891;
  wire [7:0] add_782894;
  wire [7:0] sel_782895;
  wire [7:0] add_782898;
  wire [7:0] sel_782899;
  wire [7:0] add_782902;
  wire [7:0] sel_782903;
  wire [7:0] add_782906;
  wire [7:0] sel_782907;
  wire [7:0] add_782910;
  wire [7:0] sel_782911;
  wire [7:0] add_782914;
  wire [7:0] sel_782915;
  wire [7:0] add_782918;
  wire [7:0] sel_782919;
  wire [7:0] add_782922;
  wire [7:0] sel_782923;
  wire [7:0] add_782926;
  wire [7:0] sel_782927;
  wire [7:0] add_782930;
  wire [7:0] sel_782931;
  wire [7:0] add_782934;
  wire [7:0] sel_782935;
  wire [7:0] add_782938;
  wire [7:0] sel_782939;
  wire [7:0] add_782942;
  wire [7:0] sel_782943;
  wire [7:0] add_782946;
  wire [7:0] sel_782947;
  wire [7:0] add_782950;
  wire [7:0] sel_782951;
  wire [7:0] add_782955;
  wire [15:0] array_index_782956;
  wire [7:0] sel_782957;
  wire [7:0] add_782960;
  wire [7:0] sel_782961;
  wire [7:0] add_782964;
  wire [7:0] sel_782965;
  wire [7:0] add_782968;
  wire [7:0] sel_782969;
  wire [7:0] add_782972;
  wire [7:0] sel_782973;
  wire [7:0] add_782976;
  wire [7:0] sel_782977;
  wire [7:0] add_782980;
  wire [7:0] sel_782981;
  wire [7:0] add_782984;
  wire [7:0] sel_782985;
  wire [7:0] add_782988;
  wire [7:0] sel_782989;
  wire [7:0] add_782992;
  wire [7:0] sel_782993;
  wire [7:0] add_782996;
  wire [7:0] sel_782997;
  wire [7:0] add_783000;
  wire [7:0] sel_783001;
  wire [7:0] add_783004;
  wire [7:0] sel_783005;
  wire [7:0] add_783008;
  wire [7:0] sel_783009;
  wire [7:0] add_783012;
  wire [7:0] sel_783013;
  wire [7:0] add_783016;
  wire [7:0] sel_783017;
  wire [7:0] add_783020;
  wire [7:0] sel_783021;
  wire [7:0] add_783024;
  wire [7:0] sel_783025;
  wire [7:0] add_783028;
  wire [7:0] sel_783029;
  wire [7:0] add_783032;
  wire [7:0] sel_783033;
  wire [7:0] add_783036;
  wire [7:0] sel_783037;
  wire [7:0] add_783040;
  wire [7:0] sel_783041;
  wire [7:0] add_783044;
  wire [7:0] sel_783045;
  wire [7:0] add_783048;
  wire [7:0] sel_783049;
  wire [7:0] add_783052;
  wire [7:0] sel_783053;
  wire [7:0] add_783056;
  wire [7:0] sel_783057;
  wire [7:0] add_783060;
  wire [7:0] sel_783061;
  wire [7:0] add_783064;
  wire [7:0] sel_783065;
  wire [7:0] add_783068;
  wire [7:0] sel_783069;
  wire [7:0] add_783072;
  wire [7:0] sel_783073;
  wire [7:0] add_783076;
  wire [7:0] sel_783077;
  wire [7:0] add_783080;
  wire [7:0] sel_783081;
  wire [7:0] add_783084;
  wire [7:0] sel_783085;
  wire [7:0] add_783088;
  wire [7:0] sel_783089;
  wire [7:0] add_783092;
  wire [7:0] sel_783093;
  wire [7:0] add_783096;
  wire [7:0] sel_783097;
  wire [7:0] add_783100;
  wire [7:0] sel_783101;
  wire [7:0] add_783104;
  wire [7:0] sel_783105;
  wire [7:0] add_783108;
  wire [7:0] sel_783109;
  wire [7:0] add_783112;
  wire [7:0] sel_783113;
  wire [7:0] add_783116;
  wire [7:0] sel_783117;
  wire [7:0] add_783120;
  wire [7:0] sel_783121;
  wire [7:0] add_783124;
  wire [7:0] sel_783125;
  wire [7:0] add_783128;
  wire [7:0] sel_783129;
  wire [7:0] add_783132;
  wire [7:0] sel_783133;
  wire [7:0] add_783136;
  wire [7:0] sel_783137;
  wire [7:0] add_783140;
  wire [7:0] sel_783141;
  wire [7:0] add_783144;
  wire [7:0] sel_783145;
  wire [7:0] add_783148;
  wire [7:0] sel_783149;
  wire [7:0] add_783152;
  wire [7:0] sel_783153;
  wire [7:0] add_783156;
  wire [7:0] sel_783157;
  wire [7:0] add_783160;
  wire [7:0] sel_783161;
  wire [7:0] add_783164;
  wire [7:0] sel_783165;
  wire [7:0] add_783168;
  wire [7:0] sel_783169;
  wire [7:0] add_783172;
  wire [7:0] sel_783173;
  wire [7:0] add_783176;
  wire [7:0] sel_783177;
  wire [7:0] add_783180;
  wire [7:0] sel_783181;
  wire [7:0] add_783184;
  wire [7:0] sel_783185;
  wire [7:0] add_783188;
  wire [7:0] sel_783189;
  wire [7:0] add_783192;
  wire [7:0] sel_783193;
  wire [7:0] add_783196;
  wire [7:0] sel_783197;
  wire [7:0] add_783200;
  wire [7:0] sel_783201;
  wire [7:0] add_783204;
  wire [7:0] sel_783205;
  wire [7:0] add_783208;
  wire [7:0] sel_783209;
  wire [7:0] add_783212;
  wire [7:0] sel_783213;
  wire [7:0] add_783216;
  wire [7:0] sel_783217;
  wire [7:0] add_783220;
  wire [7:0] sel_783221;
  wire [7:0] add_783224;
  wire [7:0] sel_783225;
  wire [7:0] add_783228;
  wire [7:0] sel_783229;
  wire [7:0] add_783232;
  wire [7:0] sel_783233;
  wire [7:0] add_783236;
  wire [7:0] sel_783237;
  wire [7:0] add_783240;
  wire [7:0] sel_783241;
  wire [7:0] add_783244;
  wire [7:0] sel_783245;
  wire [7:0] add_783248;
  wire [7:0] sel_783249;
  wire [7:0] add_783252;
  wire [7:0] sel_783253;
  wire [7:0] add_783256;
  wire [7:0] sel_783257;
  wire [7:0] add_783260;
  wire [7:0] sel_783261;
  wire [7:0] add_783264;
  wire [7:0] sel_783265;
  wire [7:0] add_783268;
  wire [7:0] sel_783269;
  wire [7:0] add_783272;
  wire [7:0] sel_783273;
  wire [7:0] add_783276;
  wire [7:0] sel_783277;
  wire [7:0] add_783280;
  wire [7:0] sel_783281;
  wire [7:0] add_783284;
  wire [7:0] sel_783285;
  wire [7:0] add_783288;
  wire [7:0] sel_783289;
  wire [7:0] add_783292;
  wire [7:0] sel_783293;
  wire [7:0] add_783296;
  wire [7:0] sel_783297;
  wire [7:0] add_783300;
  wire [7:0] sel_783301;
  wire [7:0] add_783304;
  wire [7:0] sel_783305;
  wire [7:0] add_783308;
  wire [7:0] sel_783309;
  wire [7:0] add_783312;
  wire [7:0] sel_783313;
  wire [7:0] add_783317;
  wire [15:0] array_index_783318;
  wire [7:0] sel_783319;
  wire [7:0] add_783322;
  wire [7:0] sel_783323;
  wire [7:0] add_783326;
  wire [7:0] sel_783327;
  wire [7:0] add_783330;
  wire [7:0] sel_783331;
  wire [7:0] add_783334;
  wire [7:0] sel_783335;
  wire [7:0] add_783338;
  wire [7:0] sel_783339;
  wire [7:0] add_783342;
  wire [7:0] sel_783343;
  wire [7:0] add_783346;
  wire [7:0] sel_783347;
  wire [7:0] add_783350;
  wire [7:0] sel_783351;
  wire [7:0] add_783354;
  wire [7:0] sel_783355;
  wire [7:0] add_783358;
  wire [7:0] sel_783359;
  wire [7:0] add_783362;
  wire [7:0] sel_783363;
  wire [7:0] add_783366;
  wire [7:0] sel_783367;
  wire [7:0] add_783370;
  wire [7:0] sel_783371;
  wire [7:0] add_783374;
  wire [7:0] sel_783375;
  wire [7:0] add_783378;
  wire [7:0] sel_783379;
  wire [7:0] add_783382;
  wire [7:0] sel_783383;
  wire [7:0] add_783386;
  wire [7:0] sel_783387;
  wire [7:0] add_783390;
  wire [7:0] sel_783391;
  wire [7:0] add_783394;
  wire [7:0] sel_783395;
  wire [7:0] add_783398;
  wire [7:0] sel_783399;
  wire [7:0] add_783402;
  wire [7:0] sel_783403;
  wire [7:0] add_783406;
  wire [7:0] sel_783407;
  wire [7:0] add_783410;
  wire [7:0] sel_783411;
  wire [7:0] add_783414;
  wire [7:0] sel_783415;
  wire [7:0] add_783418;
  wire [7:0] sel_783419;
  wire [7:0] add_783422;
  wire [7:0] sel_783423;
  wire [7:0] add_783426;
  wire [7:0] sel_783427;
  wire [7:0] add_783430;
  wire [7:0] sel_783431;
  wire [7:0] add_783434;
  wire [7:0] sel_783435;
  wire [7:0] add_783438;
  wire [7:0] sel_783439;
  wire [7:0] add_783442;
  wire [7:0] sel_783443;
  wire [7:0] add_783446;
  wire [7:0] sel_783447;
  wire [7:0] add_783450;
  wire [7:0] sel_783451;
  wire [7:0] add_783454;
  wire [7:0] sel_783455;
  wire [7:0] add_783458;
  wire [7:0] sel_783459;
  wire [7:0] add_783462;
  wire [7:0] sel_783463;
  wire [7:0] add_783466;
  wire [7:0] sel_783467;
  wire [7:0] add_783470;
  wire [7:0] sel_783471;
  wire [7:0] add_783474;
  wire [7:0] sel_783475;
  wire [7:0] add_783478;
  wire [7:0] sel_783479;
  wire [7:0] add_783482;
  wire [7:0] sel_783483;
  wire [7:0] add_783486;
  wire [7:0] sel_783487;
  wire [7:0] add_783490;
  wire [7:0] sel_783491;
  wire [7:0] add_783494;
  wire [7:0] sel_783495;
  wire [7:0] add_783498;
  wire [7:0] sel_783499;
  wire [7:0] add_783502;
  wire [7:0] sel_783503;
  wire [7:0] add_783506;
  wire [7:0] sel_783507;
  wire [7:0] add_783510;
  wire [7:0] sel_783511;
  wire [7:0] add_783514;
  wire [7:0] sel_783515;
  wire [7:0] add_783518;
  wire [7:0] sel_783519;
  wire [7:0] add_783522;
  wire [7:0] sel_783523;
  wire [7:0] add_783526;
  wire [7:0] sel_783527;
  wire [7:0] add_783530;
  wire [7:0] sel_783531;
  wire [7:0] add_783534;
  wire [7:0] sel_783535;
  wire [7:0] add_783538;
  wire [7:0] sel_783539;
  wire [7:0] add_783542;
  wire [7:0] sel_783543;
  wire [7:0] add_783546;
  wire [7:0] sel_783547;
  wire [7:0] add_783550;
  wire [7:0] sel_783551;
  wire [7:0] add_783554;
  wire [7:0] sel_783555;
  wire [7:0] add_783558;
  wire [7:0] sel_783559;
  wire [7:0] add_783562;
  wire [7:0] sel_783563;
  wire [7:0] add_783566;
  wire [7:0] sel_783567;
  wire [7:0] add_783570;
  wire [7:0] sel_783571;
  wire [7:0] add_783574;
  wire [7:0] sel_783575;
  wire [7:0] add_783578;
  wire [7:0] sel_783579;
  wire [7:0] add_783582;
  wire [7:0] sel_783583;
  wire [7:0] add_783586;
  wire [7:0] sel_783587;
  wire [7:0] add_783590;
  wire [7:0] sel_783591;
  wire [7:0] add_783594;
  wire [7:0] sel_783595;
  wire [7:0] add_783598;
  wire [7:0] sel_783599;
  wire [7:0] add_783602;
  wire [7:0] sel_783603;
  wire [7:0] add_783606;
  wire [7:0] sel_783607;
  wire [7:0] add_783610;
  wire [7:0] sel_783611;
  wire [7:0] add_783614;
  wire [7:0] sel_783615;
  wire [7:0] add_783618;
  wire [7:0] sel_783619;
  wire [7:0] add_783622;
  wire [7:0] sel_783623;
  wire [7:0] add_783626;
  wire [7:0] sel_783627;
  wire [7:0] add_783630;
  wire [7:0] sel_783631;
  wire [7:0] add_783634;
  wire [7:0] sel_783635;
  wire [7:0] add_783638;
  wire [7:0] sel_783639;
  wire [7:0] add_783642;
  wire [7:0] sel_783643;
  wire [7:0] add_783646;
  wire [7:0] sel_783647;
  wire [7:0] add_783650;
  wire [7:0] sel_783651;
  wire [7:0] add_783654;
  wire [7:0] sel_783655;
  wire [7:0] add_783658;
  wire [7:0] sel_783659;
  wire [7:0] add_783662;
  wire [7:0] sel_783663;
  wire [7:0] add_783666;
  wire [7:0] sel_783667;
  wire [7:0] add_783670;
  wire [7:0] sel_783671;
  wire [7:0] add_783674;
  wire [7:0] sel_783675;
  wire [7:0] add_783679;
  wire [15:0] array_index_783680;
  wire [7:0] sel_783681;
  wire [7:0] add_783684;
  wire [7:0] sel_783685;
  wire [7:0] add_783688;
  wire [7:0] sel_783689;
  wire [7:0] add_783692;
  wire [7:0] sel_783693;
  wire [7:0] add_783696;
  wire [7:0] sel_783697;
  wire [7:0] add_783700;
  wire [7:0] sel_783701;
  wire [7:0] add_783704;
  wire [7:0] sel_783705;
  wire [7:0] add_783708;
  wire [7:0] sel_783709;
  wire [7:0] add_783712;
  wire [7:0] sel_783713;
  wire [7:0] add_783716;
  wire [7:0] sel_783717;
  wire [7:0] add_783720;
  wire [7:0] sel_783721;
  wire [7:0] add_783724;
  wire [7:0] sel_783725;
  wire [7:0] add_783728;
  wire [7:0] sel_783729;
  wire [7:0] add_783732;
  wire [7:0] sel_783733;
  wire [7:0] add_783736;
  wire [7:0] sel_783737;
  wire [7:0] add_783740;
  wire [7:0] sel_783741;
  wire [7:0] add_783744;
  wire [7:0] sel_783745;
  wire [7:0] add_783748;
  wire [7:0] sel_783749;
  wire [7:0] add_783752;
  wire [7:0] sel_783753;
  wire [7:0] add_783756;
  wire [7:0] sel_783757;
  wire [7:0] add_783760;
  wire [7:0] sel_783761;
  wire [7:0] add_783764;
  wire [7:0] sel_783765;
  wire [7:0] add_783768;
  wire [7:0] sel_783769;
  wire [7:0] add_783772;
  wire [7:0] sel_783773;
  wire [7:0] add_783776;
  wire [7:0] sel_783777;
  wire [7:0] add_783780;
  wire [7:0] sel_783781;
  wire [7:0] add_783784;
  wire [7:0] sel_783785;
  wire [7:0] add_783788;
  wire [7:0] sel_783789;
  wire [7:0] add_783792;
  wire [7:0] sel_783793;
  wire [7:0] add_783796;
  wire [7:0] sel_783797;
  wire [7:0] add_783800;
  wire [7:0] sel_783801;
  wire [7:0] add_783804;
  wire [7:0] sel_783805;
  wire [7:0] add_783808;
  wire [7:0] sel_783809;
  wire [7:0] add_783812;
  wire [7:0] sel_783813;
  wire [7:0] add_783816;
  wire [7:0] sel_783817;
  wire [7:0] add_783820;
  wire [7:0] sel_783821;
  wire [7:0] add_783824;
  wire [7:0] sel_783825;
  wire [7:0] add_783828;
  wire [7:0] sel_783829;
  wire [7:0] add_783832;
  wire [7:0] sel_783833;
  wire [7:0] add_783836;
  wire [7:0] sel_783837;
  wire [7:0] add_783840;
  wire [7:0] sel_783841;
  wire [7:0] add_783844;
  wire [7:0] sel_783845;
  wire [7:0] add_783848;
  wire [7:0] sel_783849;
  wire [7:0] add_783852;
  wire [7:0] sel_783853;
  wire [7:0] add_783856;
  wire [7:0] sel_783857;
  wire [7:0] add_783860;
  wire [7:0] sel_783861;
  wire [7:0] add_783864;
  wire [7:0] sel_783865;
  wire [7:0] add_783868;
  wire [7:0] sel_783869;
  wire [7:0] add_783872;
  wire [7:0] sel_783873;
  wire [7:0] add_783876;
  wire [7:0] sel_783877;
  wire [7:0] add_783880;
  wire [7:0] sel_783881;
  wire [7:0] add_783884;
  wire [7:0] sel_783885;
  wire [7:0] add_783888;
  wire [7:0] sel_783889;
  wire [7:0] add_783892;
  wire [7:0] sel_783893;
  wire [7:0] add_783896;
  wire [7:0] sel_783897;
  wire [7:0] add_783900;
  wire [7:0] sel_783901;
  wire [7:0] add_783904;
  wire [7:0] sel_783905;
  wire [7:0] add_783908;
  wire [7:0] sel_783909;
  wire [7:0] add_783912;
  wire [7:0] sel_783913;
  wire [7:0] add_783916;
  wire [7:0] sel_783917;
  wire [7:0] add_783920;
  wire [7:0] sel_783921;
  wire [7:0] add_783924;
  wire [7:0] sel_783925;
  wire [7:0] add_783928;
  wire [7:0] sel_783929;
  wire [7:0] add_783932;
  wire [7:0] sel_783933;
  wire [7:0] add_783936;
  wire [7:0] sel_783937;
  wire [7:0] add_783940;
  wire [7:0] sel_783941;
  wire [7:0] add_783944;
  wire [7:0] sel_783945;
  wire [7:0] add_783948;
  wire [7:0] sel_783949;
  wire [7:0] add_783952;
  wire [7:0] sel_783953;
  wire [7:0] add_783956;
  wire [7:0] sel_783957;
  wire [7:0] add_783960;
  wire [7:0] sel_783961;
  wire [7:0] add_783964;
  wire [7:0] sel_783965;
  wire [7:0] add_783968;
  wire [7:0] sel_783969;
  wire [7:0] add_783972;
  wire [7:0] sel_783973;
  wire [7:0] add_783976;
  wire [7:0] sel_783977;
  wire [7:0] add_783980;
  wire [7:0] sel_783981;
  wire [7:0] add_783984;
  wire [7:0] sel_783985;
  wire [7:0] add_783988;
  wire [7:0] sel_783989;
  wire [7:0] add_783992;
  wire [7:0] sel_783993;
  wire [7:0] add_783996;
  wire [7:0] sel_783997;
  wire [7:0] add_784000;
  wire [7:0] sel_784001;
  wire [7:0] add_784004;
  wire [7:0] sel_784005;
  wire [7:0] add_784008;
  wire [7:0] sel_784009;
  wire [7:0] add_784012;
  wire [7:0] sel_784013;
  wire [7:0] add_784016;
  wire [7:0] sel_784017;
  wire [7:0] add_784020;
  wire [7:0] sel_784021;
  wire [7:0] add_784024;
  wire [7:0] sel_784025;
  wire [7:0] add_784028;
  wire [7:0] sel_784029;
  wire [7:0] add_784032;
  wire [7:0] sel_784033;
  wire [7:0] add_784036;
  wire [7:0] sel_784037;
  wire [7:0] add_784041;
  wire [15:0] array_index_784042;
  wire [7:0] sel_784043;
  wire [7:0] add_784046;
  wire [7:0] sel_784047;
  wire [7:0] add_784050;
  wire [7:0] sel_784051;
  wire [7:0] add_784054;
  wire [7:0] sel_784055;
  wire [7:0] add_784058;
  wire [7:0] sel_784059;
  wire [7:0] add_784062;
  wire [7:0] sel_784063;
  wire [7:0] add_784066;
  wire [7:0] sel_784067;
  wire [7:0] add_784070;
  wire [7:0] sel_784071;
  wire [7:0] add_784074;
  wire [7:0] sel_784075;
  wire [7:0] add_784078;
  wire [7:0] sel_784079;
  wire [7:0] add_784082;
  wire [7:0] sel_784083;
  wire [7:0] add_784086;
  wire [7:0] sel_784087;
  wire [7:0] add_784090;
  wire [7:0] sel_784091;
  wire [7:0] add_784094;
  wire [7:0] sel_784095;
  wire [7:0] add_784098;
  wire [7:0] sel_784099;
  wire [7:0] add_784102;
  wire [7:0] sel_784103;
  wire [7:0] add_784106;
  wire [7:0] sel_784107;
  wire [7:0] add_784110;
  wire [7:0] sel_784111;
  wire [7:0] add_784114;
  wire [7:0] sel_784115;
  wire [7:0] add_784118;
  wire [7:0] sel_784119;
  wire [7:0] add_784122;
  wire [7:0] sel_784123;
  wire [7:0] add_784126;
  wire [7:0] sel_784127;
  wire [7:0] add_784130;
  wire [7:0] sel_784131;
  wire [7:0] add_784134;
  wire [7:0] sel_784135;
  wire [7:0] add_784138;
  wire [7:0] sel_784139;
  wire [7:0] add_784142;
  wire [7:0] sel_784143;
  wire [7:0] add_784146;
  wire [7:0] sel_784147;
  wire [7:0] add_784150;
  wire [7:0] sel_784151;
  wire [7:0] add_784154;
  wire [7:0] sel_784155;
  wire [7:0] add_784158;
  wire [7:0] sel_784159;
  wire [7:0] add_784162;
  wire [7:0] sel_784163;
  wire [7:0] add_784166;
  wire [7:0] sel_784167;
  wire [7:0] add_784170;
  wire [7:0] sel_784171;
  wire [7:0] add_784174;
  wire [7:0] sel_784175;
  wire [7:0] add_784178;
  wire [7:0] sel_784179;
  wire [7:0] add_784182;
  wire [7:0] sel_784183;
  wire [7:0] add_784186;
  wire [7:0] sel_784187;
  wire [7:0] add_784190;
  wire [7:0] sel_784191;
  wire [7:0] add_784194;
  wire [7:0] sel_784195;
  wire [7:0] add_784198;
  wire [7:0] sel_784199;
  wire [7:0] add_784202;
  wire [7:0] sel_784203;
  wire [7:0] add_784206;
  wire [7:0] sel_784207;
  wire [7:0] add_784210;
  wire [7:0] sel_784211;
  wire [7:0] add_784214;
  wire [7:0] sel_784215;
  wire [7:0] add_784218;
  wire [7:0] sel_784219;
  wire [7:0] add_784222;
  wire [7:0] sel_784223;
  wire [7:0] add_784226;
  wire [7:0] sel_784227;
  wire [7:0] add_784230;
  wire [7:0] sel_784231;
  wire [7:0] add_784234;
  wire [7:0] sel_784235;
  wire [7:0] add_784238;
  wire [7:0] sel_784239;
  wire [7:0] add_784242;
  wire [7:0] sel_784243;
  wire [7:0] add_784246;
  wire [7:0] sel_784247;
  wire [7:0] add_784250;
  wire [7:0] sel_784251;
  wire [7:0] add_784254;
  wire [7:0] sel_784255;
  wire [7:0] add_784258;
  wire [7:0] sel_784259;
  wire [7:0] add_784262;
  wire [7:0] sel_784263;
  wire [7:0] add_784266;
  wire [7:0] sel_784267;
  wire [7:0] add_784270;
  wire [7:0] sel_784271;
  wire [7:0] add_784274;
  wire [7:0] sel_784275;
  wire [7:0] add_784278;
  wire [7:0] sel_784279;
  wire [7:0] add_784282;
  wire [7:0] sel_784283;
  wire [7:0] add_784286;
  wire [7:0] sel_784287;
  wire [7:0] add_784290;
  wire [7:0] sel_784291;
  wire [7:0] add_784294;
  wire [7:0] sel_784295;
  wire [7:0] add_784298;
  wire [7:0] sel_784299;
  wire [7:0] add_784302;
  wire [7:0] sel_784303;
  wire [7:0] add_784306;
  wire [7:0] sel_784307;
  wire [7:0] add_784310;
  wire [7:0] sel_784311;
  wire [7:0] add_784314;
  wire [7:0] sel_784315;
  wire [7:0] add_784318;
  wire [7:0] sel_784319;
  wire [7:0] add_784322;
  wire [7:0] sel_784323;
  wire [7:0] add_784326;
  wire [7:0] sel_784327;
  wire [7:0] add_784330;
  wire [7:0] sel_784331;
  wire [7:0] add_784334;
  wire [7:0] sel_784335;
  wire [7:0] add_784338;
  wire [7:0] sel_784339;
  wire [7:0] add_784342;
  wire [7:0] sel_784343;
  wire [7:0] add_784346;
  wire [7:0] sel_784347;
  wire [7:0] add_784350;
  wire [7:0] sel_784351;
  wire [7:0] add_784354;
  wire [7:0] sel_784355;
  wire [7:0] add_784358;
  wire [7:0] sel_784359;
  wire [7:0] add_784362;
  wire [7:0] sel_784363;
  wire [7:0] add_784366;
  wire [7:0] sel_784367;
  wire [7:0] add_784370;
  wire [7:0] sel_784371;
  wire [7:0] add_784374;
  wire [7:0] sel_784375;
  wire [7:0] add_784378;
  wire [7:0] sel_784379;
  wire [7:0] add_784382;
  wire [7:0] sel_784383;
  wire [7:0] add_784386;
  wire [7:0] sel_784387;
  wire [7:0] add_784390;
  wire [7:0] sel_784391;
  wire [7:0] add_784394;
  wire [7:0] sel_784395;
  wire [7:0] add_784398;
  wire [7:0] sel_784399;
  wire [7:0] add_784403;
  wire [15:0] array_index_784404;
  wire [7:0] sel_784405;
  wire [7:0] add_784408;
  wire [7:0] sel_784409;
  wire [7:0] add_784412;
  wire [7:0] sel_784413;
  wire [7:0] add_784416;
  wire [7:0] sel_784417;
  wire [7:0] add_784420;
  wire [7:0] sel_784421;
  wire [7:0] add_784424;
  wire [7:0] sel_784425;
  wire [7:0] add_784428;
  wire [7:0] sel_784429;
  wire [7:0] add_784432;
  wire [7:0] sel_784433;
  wire [7:0] add_784436;
  wire [7:0] sel_784437;
  wire [7:0] add_784440;
  wire [7:0] sel_784441;
  wire [7:0] add_784444;
  wire [7:0] sel_784445;
  wire [7:0] add_784448;
  wire [7:0] sel_784449;
  wire [7:0] add_784452;
  wire [7:0] sel_784453;
  wire [7:0] add_784456;
  wire [7:0] sel_784457;
  wire [7:0] add_784460;
  wire [7:0] sel_784461;
  wire [7:0] add_784464;
  wire [7:0] sel_784465;
  wire [7:0] add_784468;
  wire [7:0] sel_784469;
  wire [7:0] add_784472;
  wire [7:0] sel_784473;
  wire [7:0] add_784476;
  wire [7:0] sel_784477;
  wire [7:0] add_784480;
  wire [7:0] sel_784481;
  wire [7:0] add_784484;
  wire [7:0] sel_784485;
  wire [7:0] add_784488;
  wire [7:0] sel_784489;
  wire [7:0] add_784492;
  wire [7:0] sel_784493;
  wire [7:0] add_784496;
  wire [7:0] sel_784497;
  wire [7:0] add_784500;
  wire [7:0] sel_784501;
  wire [7:0] add_784504;
  wire [7:0] sel_784505;
  wire [7:0] add_784508;
  wire [7:0] sel_784509;
  wire [7:0] add_784512;
  wire [7:0] sel_784513;
  wire [7:0] add_784516;
  wire [7:0] sel_784517;
  wire [7:0] add_784520;
  wire [7:0] sel_784521;
  wire [7:0] add_784524;
  wire [7:0] sel_784525;
  wire [7:0] add_784528;
  wire [7:0] sel_784529;
  wire [7:0] add_784532;
  wire [7:0] sel_784533;
  wire [7:0] add_784536;
  wire [7:0] sel_784537;
  wire [7:0] add_784540;
  wire [7:0] sel_784541;
  wire [7:0] add_784544;
  wire [7:0] sel_784545;
  wire [7:0] add_784548;
  wire [7:0] sel_784549;
  wire [7:0] add_784552;
  wire [7:0] sel_784553;
  wire [7:0] add_784556;
  wire [7:0] sel_784557;
  wire [7:0] add_784560;
  wire [7:0] sel_784561;
  wire [7:0] add_784564;
  wire [7:0] sel_784565;
  wire [7:0] add_784568;
  wire [7:0] sel_784569;
  wire [7:0] add_784572;
  wire [7:0] sel_784573;
  wire [7:0] add_784576;
  wire [7:0] sel_784577;
  wire [7:0] add_784580;
  wire [7:0] sel_784581;
  wire [7:0] add_784584;
  wire [7:0] sel_784585;
  wire [7:0] add_784588;
  wire [7:0] sel_784589;
  wire [7:0] add_784592;
  wire [7:0] sel_784593;
  wire [7:0] add_784596;
  wire [7:0] sel_784597;
  wire [7:0] add_784600;
  wire [7:0] sel_784601;
  wire [7:0] add_784604;
  wire [7:0] sel_784605;
  wire [7:0] add_784608;
  wire [7:0] sel_784609;
  wire [7:0] add_784612;
  wire [7:0] sel_784613;
  wire [7:0] add_784616;
  wire [7:0] sel_784617;
  wire [7:0] add_784620;
  wire [7:0] sel_784621;
  wire [7:0] add_784624;
  wire [7:0] sel_784625;
  wire [7:0] add_784628;
  wire [7:0] sel_784629;
  wire [7:0] add_784632;
  wire [7:0] sel_784633;
  wire [7:0] add_784636;
  wire [7:0] sel_784637;
  wire [7:0] add_784640;
  wire [7:0] sel_784641;
  wire [7:0] add_784644;
  wire [7:0] sel_784645;
  wire [7:0] add_784648;
  wire [7:0] sel_784649;
  wire [7:0] add_784652;
  wire [7:0] sel_784653;
  wire [7:0] add_784656;
  wire [7:0] sel_784657;
  wire [7:0] add_784660;
  wire [7:0] sel_784661;
  wire [7:0] add_784664;
  wire [7:0] sel_784665;
  wire [7:0] add_784668;
  wire [7:0] sel_784669;
  wire [7:0] add_784672;
  wire [7:0] sel_784673;
  wire [7:0] add_784676;
  wire [7:0] sel_784677;
  wire [7:0] add_784680;
  wire [7:0] sel_784681;
  wire [7:0] add_784684;
  wire [7:0] sel_784685;
  wire [7:0] add_784688;
  wire [7:0] sel_784689;
  wire [7:0] add_784692;
  wire [7:0] sel_784693;
  wire [7:0] add_784696;
  wire [7:0] sel_784697;
  wire [7:0] add_784700;
  wire [7:0] sel_784701;
  wire [7:0] add_784704;
  wire [7:0] sel_784705;
  wire [7:0] add_784708;
  wire [7:0] sel_784709;
  wire [7:0] add_784712;
  wire [7:0] sel_784713;
  wire [7:0] add_784716;
  wire [7:0] sel_784717;
  wire [7:0] add_784720;
  wire [7:0] sel_784721;
  wire [7:0] add_784724;
  wire [7:0] sel_784725;
  wire [7:0] add_784728;
  wire [7:0] sel_784729;
  wire [7:0] add_784732;
  wire [7:0] sel_784733;
  wire [7:0] add_784736;
  wire [7:0] sel_784737;
  wire [7:0] add_784740;
  wire [7:0] sel_784741;
  wire [7:0] add_784744;
  wire [7:0] sel_784745;
  wire [7:0] add_784748;
  wire [7:0] sel_784749;
  wire [7:0] add_784752;
  wire [7:0] sel_784753;
  wire [7:0] add_784756;
  wire [7:0] sel_784757;
  wire [7:0] add_784760;
  wire [7:0] sel_784761;
  wire [7:0] add_784765;
  wire [15:0] array_index_784766;
  wire [7:0] sel_784767;
  wire [7:0] add_784770;
  wire [7:0] sel_784771;
  wire [7:0] add_784774;
  wire [7:0] sel_784775;
  wire [7:0] add_784778;
  wire [7:0] sel_784779;
  wire [7:0] add_784782;
  wire [7:0] sel_784783;
  wire [7:0] add_784786;
  wire [7:0] sel_784787;
  wire [7:0] add_784790;
  wire [7:0] sel_784791;
  wire [7:0] add_784794;
  wire [7:0] sel_784795;
  wire [7:0] add_784798;
  wire [7:0] sel_784799;
  wire [7:0] add_784802;
  wire [7:0] sel_784803;
  wire [7:0] add_784806;
  wire [7:0] sel_784807;
  wire [7:0] add_784810;
  wire [7:0] sel_784811;
  wire [7:0] add_784814;
  wire [7:0] sel_784815;
  wire [7:0] add_784818;
  wire [7:0] sel_784819;
  wire [7:0] add_784822;
  wire [7:0] sel_784823;
  wire [7:0] add_784826;
  wire [7:0] sel_784827;
  wire [7:0] add_784830;
  wire [7:0] sel_784831;
  wire [7:0] add_784834;
  wire [7:0] sel_784835;
  wire [7:0] add_784838;
  wire [7:0] sel_784839;
  wire [7:0] add_784842;
  wire [7:0] sel_784843;
  wire [7:0] add_784846;
  wire [7:0] sel_784847;
  wire [7:0] add_784850;
  wire [7:0] sel_784851;
  wire [7:0] add_784854;
  wire [7:0] sel_784855;
  wire [7:0] add_784858;
  wire [7:0] sel_784859;
  wire [7:0] add_784862;
  wire [7:0] sel_784863;
  wire [7:0] add_784866;
  wire [7:0] sel_784867;
  wire [7:0] add_784870;
  wire [7:0] sel_784871;
  wire [7:0] add_784874;
  wire [7:0] sel_784875;
  wire [7:0] add_784878;
  wire [7:0] sel_784879;
  wire [7:0] add_784882;
  wire [7:0] sel_784883;
  wire [7:0] add_784886;
  wire [7:0] sel_784887;
  wire [7:0] add_784890;
  wire [7:0] sel_784891;
  wire [7:0] add_784894;
  wire [7:0] sel_784895;
  wire [7:0] add_784898;
  wire [7:0] sel_784899;
  wire [7:0] add_784902;
  wire [7:0] sel_784903;
  wire [7:0] add_784906;
  wire [7:0] sel_784907;
  wire [7:0] add_784910;
  wire [7:0] sel_784911;
  wire [7:0] add_784914;
  wire [7:0] sel_784915;
  wire [7:0] add_784918;
  wire [7:0] sel_784919;
  wire [7:0] add_784922;
  wire [7:0] sel_784923;
  wire [7:0] add_784926;
  wire [7:0] sel_784927;
  wire [7:0] add_784930;
  wire [7:0] sel_784931;
  wire [7:0] add_784934;
  wire [7:0] sel_784935;
  wire [7:0] add_784938;
  wire [7:0] sel_784939;
  wire [7:0] add_784942;
  wire [7:0] sel_784943;
  wire [7:0] add_784946;
  wire [7:0] sel_784947;
  wire [7:0] add_784950;
  wire [7:0] sel_784951;
  wire [7:0] add_784954;
  wire [7:0] sel_784955;
  wire [7:0] add_784958;
  wire [7:0] sel_784959;
  wire [7:0] add_784962;
  wire [7:0] sel_784963;
  wire [7:0] add_784966;
  wire [7:0] sel_784967;
  wire [7:0] add_784970;
  wire [7:0] sel_784971;
  wire [7:0] add_784974;
  wire [7:0] sel_784975;
  wire [7:0] add_784978;
  wire [7:0] sel_784979;
  wire [7:0] add_784982;
  wire [7:0] sel_784983;
  wire [7:0] add_784986;
  wire [7:0] sel_784987;
  wire [7:0] add_784990;
  wire [7:0] sel_784991;
  wire [7:0] add_784994;
  wire [7:0] sel_784995;
  wire [7:0] add_784998;
  wire [7:0] sel_784999;
  wire [7:0] add_785002;
  wire [7:0] sel_785003;
  wire [7:0] add_785006;
  wire [7:0] sel_785007;
  wire [7:0] add_785010;
  wire [7:0] sel_785011;
  wire [7:0] add_785014;
  wire [7:0] sel_785015;
  wire [7:0] add_785018;
  wire [7:0] sel_785019;
  wire [7:0] add_785022;
  wire [7:0] sel_785023;
  wire [7:0] add_785026;
  wire [7:0] sel_785027;
  wire [7:0] add_785030;
  wire [7:0] sel_785031;
  wire [7:0] add_785034;
  wire [7:0] sel_785035;
  wire [7:0] add_785038;
  wire [7:0] sel_785039;
  wire [7:0] add_785042;
  wire [7:0] sel_785043;
  wire [7:0] add_785046;
  wire [7:0] sel_785047;
  wire [7:0] add_785050;
  wire [7:0] sel_785051;
  wire [7:0] add_785054;
  wire [7:0] sel_785055;
  wire [7:0] add_785058;
  wire [7:0] sel_785059;
  wire [7:0] add_785062;
  wire [7:0] sel_785063;
  wire [7:0] add_785066;
  wire [7:0] sel_785067;
  wire [7:0] add_785070;
  wire [7:0] sel_785071;
  wire [7:0] add_785074;
  wire [7:0] sel_785075;
  wire [7:0] add_785078;
  wire [7:0] sel_785079;
  wire [7:0] add_785082;
  wire [7:0] sel_785083;
  wire [7:0] add_785086;
  wire [7:0] sel_785087;
  wire [7:0] add_785090;
  wire [7:0] sel_785091;
  wire [7:0] add_785094;
  wire [7:0] sel_785095;
  wire [7:0] add_785098;
  wire [7:0] sel_785099;
  wire [7:0] add_785102;
  wire [7:0] sel_785103;
  wire [7:0] add_785106;
  wire [7:0] sel_785107;
  wire [7:0] add_785110;
  wire [7:0] sel_785111;
  wire [7:0] add_785114;
  wire [7:0] sel_785115;
  wire [7:0] add_785118;
  wire [7:0] sel_785119;
  wire [7:0] add_785122;
  wire [7:0] sel_785123;
  wire [7:0] add_785127;
  wire [15:0] array_index_785128;
  wire [7:0] sel_785129;
  wire [7:0] add_785132;
  wire [7:0] sel_785133;
  wire [7:0] add_785136;
  wire [7:0] sel_785137;
  wire [7:0] add_785140;
  wire [7:0] sel_785141;
  wire [7:0] add_785144;
  wire [7:0] sel_785145;
  wire [7:0] add_785148;
  wire [7:0] sel_785149;
  wire [7:0] add_785152;
  wire [7:0] sel_785153;
  wire [7:0] add_785156;
  wire [7:0] sel_785157;
  wire [7:0] add_785160;
  wire [7:0] sel_785161;
  wire [7:0] add_785164;
  wire [7:0] sel_785165;
  wire [7:0] add_785168;
  wire [7:0] sel_785169;
  wire [7:0] add_785172;
  wire [7:0] sel_785173;
  wire [7:0] add_785176;
  wire [7:0] sel_785177;
  wire [7:0] add_785180;
  wire [7:0] sel_785181;
  wire [7:0] add_785184;
  wire [7:0] sel_785185;
  wire [7:0] add_785188;
  wire [7:0] sel_785189;
  wire [7:0] add_785192;
  wire [7:0] sel_785193;
  wire [7:0] add_785196;
  wire [7:0] sel_785197;
  wire [7:0] add_785200;
  wire [7:0] sel_785201;
  wire [7:0] add_785204;
  wire [7:0] sel_785205;
  wire [7:0] add_785208;
  wire [7:0] sel_785209;
  wire [7:0] add_785212;
  wire [7:0] sel_785213;
  wire [7:0] add_785216;
  wire [7:0] sel_785217;
  wire [7:0] add_785220;
  wire [7:0] sel_785221;
  wire [7:0] add_785224;
  wire [7:0] sel_785225;
  wire [7:0] add_785228;
  wire [7:0] sel_785229;
  wire [7:0] add_785232;
  wire [7:0] sel_785233;
  wire [7:0] add_785236;
  wire [7:0] sel_785237;
  wire [7:0] add_785240;
  wire [7:0] sel_785241;
  wire [7:0] add_785244;
  wire [7:0] sel_785245;
  wire [7:0] add_785248;
  wire [7:0] sel_785249;
  wire [7:0] add_785252;
  wire [7:0] sel_785253;
  wire [7:0] add_785256;
  wire [7:0] sel_785257;
  wire [7:0] add_785260;
  wire [7:0] sel_785261;
  wire [7:0] add_785264;
  wire [7:0] sel_785265;
  wire [7:0] add_785268;
  wire [7:0] sel_785269;
  wire [7:0] add_785272;
  wire [7:0] sel_785273;
  wire [7:0] add_785276;
  wire [7:0] sel_785277;
  wire [7:0] add_785280;
  wire [7:0] sel_785281;
  wire [7:0] add_785284;
  wire [7:0] sel_785285;
  wire [7:0] add_785288;
  wire [7:0] sel_785289;
  wire [7:0] add_785292;
  wire [7:0] sel_785293;
  wire [7:0] add_785296;
  wire [7:0] sel_785297;
  wire [7:0] add_785300;
  wire [7:0] sel_785301;
  wire [7:0] add_785304;
  wire [7:0] sel_785305;
  wire [7:0] add_785308;
  wire [7:0] sel_785309;
  wire [7:0] add_785312;
  wire [7:0] sel_785313;
  wire [7:0] add_785316;
  wire [7:0] sel_785317;
  wire [7:0] add_785320;
  wire [7:0] sel_785321;
  wire [7:0] add_785324;
  wire [7:0] sel_785325;
  wire [7:0] add_785328;
  wire [7:0] sel_785329;
  wire [7:0] add_785332;
  wire [7:0] sel_785333;
  wire [7:0] add_785336;
  wire [7:0] sel_785337;
  wire [7:0] add_785340;
  wire [7:0] sel_785341;
  wire [7:0] add_785344;
  wire [7:0] sel_785345;
  wire [7:0] add_785348;
  wire [7:0] sel_785349;
  wire [7:0] add_785352;
  wire [7:0] sel_785353;
  wire [7:0] add_785356;
  wire [7:0] sel_785357;
  wire [7:0] add_785360;
  wire [7:0] sel_785361;
  wire [7:0] add_785364;
  wire [7:0] sel_785365;
  wire [7:0] add_785368;
  wire [7:0] sel_785369;
  wire [7:0] add_785372;
  wire [7:0] sel_785373;
  wire [7:0] add_785376;
  wire [7:0] sel_785377;
  wire [7:0] add_785380;
  wire [7:0] sel_785381;
  wire [7:0] add_785384;
  wire [7:0] sel_785385;
  wire [7:0] add_785388;
  wire [7:0] sel_785389;
  wire [7:0] add_785392;
  wire [7:0] sel_785393;
  wire [7:0] add_785396;
  wire [7:0] sel_785397;
  wire [7:0] add_785400;
  wire [7:0] sel_785401;
  wire [7:0] add_785404;
  wire [7:0] sel_785405;
  wire [7:0] add_785408;
  wire [7:0] sel_785409;
  wire [7:0] add_785412;
  wire [7:0] sel_785413;
  wire [7:0] add_785416;
  wire [7:0] sel_785417;
  wire [7:0] add_785420;
  wire [7:0] sel_785421;
  wire [7:0] add_785424;
  wire [7:0] sel_785425;
  wire [7:0] add_785428;
  wire [7:0] sel_785429;
  wire [7:0] add_785432;
  wire [7:0] sel_785433;
  wire [7:0] add_785436;
  wire [7:0] sel_785437;
  wire [7:0] add_785440;
  wire [7:0] sel_785441;
  wire [7:0] add_785444;
  wire [7:0] sel_785445;
  wire [7:0] add_785448;
  wire [7:0] sel_785449;
  wire [7:0] add_785452;
  wire [7:0] sel_785453;
  wire [7:0] add_785456;
  wire [7:0] sel_785457;
  wire [7:0] add_785460;
  wire [7:0] sel_785461;
  wire [7:0] add_785464;
  wire [7:0] sel_785465;
  wire [7:0] add_785468;
  wire [7:0] sel_785469;
  wire [7:0] add_785472;
  wire [7:0] sel_785473;
  wire [7:0] add_785476;
  wire [7:0] sel_785477;
  wire [7:0] add_785480;
  wire [7:0] sel_785481;
  wire [7:0] add_785484;
  wire [7:0] sel_785485;
  wire [7:0] add_785489;
  wire [15:0] array_index_785490;
  wire [7:0] sel_785491;
  wire [7:0] add_785494;
  wire [7:0] sel_785495;
  wire [7:0] add_785498;
  wire [7:0] sel_785499;
  wire [7:0] add_785502;
  wire [7:0] sel_785503;
  wire [7:0] add_785506;
  wire [7:0] sel_785507;
  wire [7:0] add_785510;
  wire [7:0] sel_785511;
  wire [7:0] add_785514;
  wire [7:0] sel_785515;
  wire [7:0] add_785518;
  wire [7:0] sel_785519;
  wire [7:0] add_785522;
  wire [7:0] sel_785523;
  wire [7:0] add_785526;
  wire [7:0] sel_785527;
  wire [7:0] add_785530;
  wire [7:0] sel_785531;
  wire [7:0] add_785534;
  wire [7:0] sel_785535;
  wire [7:0] add_785538;
  wire [7:0] sel_785539;
  wire [7:0] add_785542;
  wire [7:0] sel_785543;
  wire [7:0] add_785546;
  wire [7:0] sel_785547;
  wire [7:0] add_785550;
  wire [7:0] sel_785551;
  wire [7:0] add_785554;
  wire [7:0] sel_785555;
  wire [7:0] add_785558;
  wire [7:0] sel_785559;
  wire [7:0] add_785562;
  wire [7:0] sel_785563;
  wire [7:0] add_785566;
  wire [7:0] sel_785567;
  wire [7:0] add_785570;
  wire [7:0] sel_785571;
  wire [7:0] add_785574;
  wire [7:0] sel_785575;
  wire [7:0] add_785578;
  wire [7:0] sel_785579;
  wire [7:0] add_785582;
  wire [7:0] sel_785583;
  wire [7:0] add_785586;
  wire [7:0] sel_785587;
  wire [7:0] add_785590;
  wire [7:0] sel_785591;
  wire [7:0] add_785594;
  wire [7:0] sel_785595;
  wire [7:0] add_785598;
  wire [7:0] sel_785599;
  wire [7:0] add_785602;
  wire [7:0] sel_785603;
  wire [7:0] add_785606;
  wire [7:0] sel_785607;
  wire [7:0] add_785610;
  wire [7:0] sel_785611;
  wire [7:0] add_785614;
  wire [7:0] sel_785615;
  wire [7:0] add_785618;
  wire [7:0] sel_785619;
  wire [7:0] add_785622;
  wire [7:0] sel_785623;
  wire [7:0] add_785626;
  wire [7:0] sel_785627;
  wire [7:0] add_785630;
  wire [7:0] sel_785631;
  wire [7:0] add_785634;
  wire [7:0] sel_785635;
  wire [7:0] add_785638;
  wire [7:0] sel_785639;
  wire [7:0] add_785642;
  wire [7:0] sel_785643;
  wire [7:0] add_785646;
  wire [7:0] sel_785647;
  wire [7:0] add_785650;
  wire [7:0] sel_785651;
  wire [7:0] add_785654;
  wire [7:0] sel_785655;
  wire [7:0] add_785658;
  wire [7:0] sel_785659;
  wire [7:0] add_785662;
  wire [7:0] sel_785663;
  wire [7:0] add_785666;
  wire [7:0] sel_785667;
  wire [7:0] add_785670;
  wire [7:0] sel_785671;
  wire [7:0] add_785674;
  wire [7:0] sel_785675;
  wire [7:0] add_785678;
  wire [7:0] sel_785679;
  wire [7:0] add_785682;
  wire [7:0] sel_785683;
  wire [7:0] add_785686;
  wire [7:0] sel_785687;
  wire [7:0] add_785690;
  wire [7:0] sel_785691;
  wire [7:0] add_785694;
  wire [7:0] sel_785695;
  wire [7:0] add_785698;
  wire [7:0] sel_785699;
  wire [7:0] add_785702;
  wire [7:0] sel_785703;
  wire [7:0] add_785706;
  wire [7:0] sel_785707;
  wire [7:0] add_785710;
  wire [7:0] sel_785711;
  wire [7:0] add_785714;
  wire [7:0] sel_785715;
  wire [7:0] add_785718;
  wire [7:0] sel_785719;
  wire [7:0] add_785722;
  wire [7:0] sel_785723;
  wire [7:0] add_785726;
  wire [7:0] sel_785727;
  wire [7:0] add_785730;
  wire [7:0] sel_785731;
  wire [7:0] add_785734;
  wire [7:0] sel_785735;
  wire [7:0] add_785738;
  wire [7:0] sel_785739;
  wire [7:0] add_785742;
  wire [7:0] sel_785743;
  wire [7:0] add_785746;
  wire [7:0] sel_785747;
  wire [7:0] add_785750;
  wire [7:0] sel_785751;
  wire [7:0] add_785754;
  wire [7:0] sel_785755;
  wire [7:0] add_785758;
  wire [7:0] sel_785759;
  wire [7:0] add_785762;
  wire [7:0] sel_785763;
  wire [7:0] add_785766;
  wire [7:0] sel_785767;
  wire [7:0] add_785770;
  wire [7:0] sel_785771;
  wire [7:0] add_785774;
  wire [7:0] sel_785775;
  wire [7:0] add_785778;
  wire [7:0] sel_785779;
  wire [7:0] add_785782;
  wire [7:0] sel_785783;
  wire [7:0] add_785786;
  wire [7:0] sel_785787;
  wire [7:0] add_785790;
  wire [7:0] sel_785791;
  wire [7:0] add_785794;
  wire [7:0] sel_785795;
  wire [7:0] add_785798;
  wire [7:0] sel_785799;
  wire [7:0] add_785802;
  wire [7:0] sel_785803;
  wire [7:0] add_785806;
  wire [7:0] sel_785807;
  wire [7:0] add_785810;
  wire [7:0] sel_785811;
  wire [7:0] add_785814;
  wire [7:0] sel_785815;
  wire [7:0] add_785818;
  wire [7:0] sel_785819;
  wire [7:0] add_785822;
  wire [7:0] sel_785823;
  wire [7:0] add_785826;
  wire [7:0] sel_785827;
  wire [7:0] add_785830;
  wire [7:0] sel_785831;
  wire [7:0] add_785834;
  wire [7:0] sel_785835;
  wire [7:0] add_785838;
  wire [7:0] sel_785839;
  wire [7:0] add_785842;
  wire [7:0] sel_785843;
  wire [7:0] add_785846;
  wire [7:0] sel_785847;
  wire [7:0] add_785851;
  wire [15:0] array_index_785852;
  wire [7:0] sel_785853;
  wire [7:0] add_785856;
  wire [7:0] sel_785857;
  wire [7:0] add_785860;
  wire [7:0] sel_785861;
  wire [7:0] add_785864;
  wire [7:0] sel_785865;
  wire [7:0] add_785868;
  wire [7:0] sel_785869;
  wire [7:0] add_785872;
  wire [7:0] sel_785873;
  wire [7:0] add_785876;
  wire [7:0] sel_785877;
  wire [7:0] add_785880;
  wire [7:0] sel_785881;
  wire [7:0] add_785884;
  wire [7:0] sel_785885;
  wire [7:0] add_785888;
  wire [7:0] sel_785889;
  wire [7:0] add_785892;
  wire [7:0] sel_785893;
  wire [7:0] add_785896;
  wire [7:0] sel_785897;
  wire [7:0] add_785900;
  wire [7:0] sel_785901;
  wire [7:0] add_785904;
  wire [7:0] sel_785905;
  wire [7:0] add_785908;
  wire [7:0] sel_785909;
  wire [7:0] add_785912;
  wire [7:0] sel_785913;
  wire [7:0] add_785916;
  wire [7:0] sel_785917;
  wire [7:0] add_785920;
  wire [7:0] sel_785921;
  wire [7:0] add_785924;
  wire [7:0] sel_785925;
  wire [7:0] add_785928;
  wire [7:0] sel_785929;
  wire [7:0] add_785932;
  wire [7:0] sel_785933;
  wire [7:0] add_785936;
  wire [7:0] sel_785937;
  wire [7:0] add_785940;
  wire [7:0] sel_785941;
  wire [7:0] add_785944;
  wire [7:0] sel_785945;
  wire [7:0] add_785948;
  wire [7:0] sel_785949;
  wire [7:0] add_785952;
  wire [7:0] sel_785953;
  wire [7:0] add_785956;
  wire [7:0] sel_785957;
  wire [7:0] add_785960;
  wire [7:0] sel_785961;
  wire [7:0] add_785964;
  wire [7:0] sel_785965;
  wire [7:0] add_785968;
  wire [7:0] sel_785969;
  wire [7:0] add_785972;
  wire [7:0] sel_785973;
  wire [7:0] add_785976;
  wire [7:0] sel_785977;
  wire [7:0] add_785980;
  wire [7:0] sel_785981;
  wire [7:0] add_785984;
  wire [7:0] sel_785985;
  wire [7:0] add_785988;
  wire [7:0] sel_785989;
  wire [7:0] add_785992;
  wire [7:0] sel_785993;
  wire [7:0] add_785996;
  wire [7:0] sel_785997;
  wire [7:0] add_786000;
  wire [7:0] sel_786001;
  wire [7:0] add_786004;
  wire [7:0] sel_786005;
  wire [7:0] add_786008;
  wire [7:0] sel_786009;
  wire [7:0] add_786012;
  wire [7:0] sel_786013;
  wire [7:0] add_786016;
  wire [7:0] sel_786017;
  wire [7:0] add_786020;
  wire [7:0] sel_786021;
  wire [7:0] add_786024;
  wire [7:0] sel_786025;
  wire [7:0] add_786028;
  wire [7:0] sel_786029;
  wire [7:0] add_786032;
  wire [7:0] sel_786033;
  wire [7:0] add_786036;
  wire [7:0] sel_786037;
  wire [7:0] add_786040;
  wire [7:0] sel_786041;
  wire [7:0] add_786044;
  wire [7:0] sel_786045;
  wire [7:0] add_786048;
  wire [7:0] sel_786049;
  wire [7:0] add_786052;
  wire [7:0] sel_786053;
  wire [7:0] add_786056;
  wire [7:0] sel_786057;
  wire [7:0] add_786060;
  wire [7:0] sel_786061;
  wire [7:0] add_786064;
  wire [7:0] sel_786065;
  wire [7:0] add_786068;
  wire [7:0] sel_786069;
  wire [7:0] add_786072;
  wire [7:0] sel_786073;
  wire [7:0] add_786076;
  wire [7:0] sel_786077;
  wire [7:0] add_786080;
  wire [7:0] sel_786081;
  wire [7:0] add_786084;
  wire [7:0] sel_786085;
  wire [7:0] add_786088;
  wire [7:0] sel_786089;
  wire [7:0] add_786092;
  wire [7:0] sel_786093;
  wire [7:0] add_786096;
  wire [7:0] sel_786097;
  wire [7:0] add_786100;
  wire [7:0] sel_786101;
  wire [7:0] add_786104;
  wire [7:0] sel_786105;
  wire [7:0] add_786108;
  wire [7:0] sel_786109;
  wire [7:0] add_786112;
  wire [7:0] sel_786113;
  wire [7:0] add_786116;
  wire [7:0] sel_786117;
  wire [7:0] add_786120;
  wire [7:0] sel_786121;
  wire [7:0] add_786124;
  wire [7:0] sel_786125;
  wire [7:0] add_786128;
  wire [7:0] sel_786129;
  wire [7:0] add_786132;
  wire [7:0] sel_786133;
  wire [7:0] add_786136;
  wire [7:0] sel_786137;
  wire [7:0] add_786140;
  wire [7:0] sel_786141;
  wire [7:0] add_786144;
  wire [7:0] sel_786145;
  wire [7:0] add_786148;
  wire [7:0] sel_786149;
  wire [7:0] add_786152;
  wire [7:0] sel_786153;
  wire [7:0] add_786156;
  wire [7:0] sel_786157;
  wire [7:0] add_786160;
  wire [7:0] sel_786161;
  wire [7:0] add_786164;
  wire [7:0] sel_786165;
  wire [7:0] add_786168;
  wire [7:0] sel_786169;
  wire [7:0] add_786172;
  wire [7:0] sel_786173;
  wire [7:0] add_786176;
  wire [7:0] sel_786177;
  wire [7:0] add_786180;
  wire [7:0] sel_786181;
  wire [7:0] add_786184;
  wire [7:0] sel_786185;
  wire [7:0] add_786188;
  wire [7:0] sel_786189;
  wire [7:0] add_786192;
  wire [7:0] sel_786193;
  wire [7:0] add_786196;
  wire [7:0] sel_786197;
  wire [7:0] add_786200;
  wire [7:0] sel_786201;
  wire [7:0] add_786204;
  wire [7:0] sel_786205;
  wire [7:0] add_786208;
  wire [7:0] sel_786209;
  wire [7:0] add_786213;
  wire [15:0] array_index_786214;
  wire [7:0] sel_786215;
  wire [7:0] add_786218;
  wire [7:0] sel_786219;
  wire [7:0] add_786222;
  wire [7:0] sel_786223;
  wire [7:0] add_786226;
  wire [7:0] sel_786227;
  wire [7:0] add_786230;
  wire [7:0] sel_786231;
  wire [7:0] add_786234;
  wire [7:0] sel_786235;
  wire [7:0] add_786238;
  wire [7:0] sel_786239;
  wire [7:0] add_786242;
  wire [7:0] sel_786243;
  wire [7:0] add_786246;
  wire [7:0] sel_786247;
  wire [7:0] add_786250;
  wire [7:0] sel_786251;
  wire [7:0] add_786254;
  wire [7:0] sel_786255;
  wire [7:0] add_786258;
  wire [7:0] sel_786259;
  wire [7:0] add_786262;
  wire [7:0] sel_786263;
  wire [7:0] add_786266;
  wire [7:0] sel_786267;
  wire [7:0] add_786270;
  wire [7:0] sel_786271;
  wire [7:0] add_786274;
  wire [7:0] sel_786275;
  wire [7:0] add_786278;
  wire [7:0] sel_786279;
  wire [7:0] add_786282;
  wire [7:0] sel_786283;
  wire [7:0] add_786286;
  wire [7:0] sel_786287;
  wire [7:0] add_786290;
  wire [7:0] sel_786291;
  wire [7:0] add_786294;
  wire [7:0] sel_786295;
  wire [7:0] add_786298;
  wire [7:0] sel_786299;
  wire [7:0] add_786302;
  wire [7:0] sel_786303;
  wire [7:0] add_786306;
  wire [7:0] sel_786307;
  wire [7:0] add_786310;
  wire [7:0] sel_786311;
  wire [7:0] add_786314;
  wire [7:0] sel_786315;
  wire [7:0] add_786318;
  wire [7:0] sel_786319;
  wire [7:0] add_786322;
  wire [7:0] sel_786323;
  wire [7:0] add_786326;
  wire [7:0] sel_786327;
  wire [7:0] add_786330;
  wire [7:0] sel_786331;
  wire [7:0] add_786334;
  wire [7:0] sel_786335;
  wire [7:0] add_786338;
  wire [7:0] sel_786339;
  wire [7:0] add_786342;
  wire [7:0] sel_786343;
  wire [7:0] add_786346;
  wire [7:0] sel_786347;
  wire [7:0] add_786350;
  wire [7:0] sel_786351;
  wire [7:0] add_786354;
  wire [7:0] sel_786355;
  wire [7:0] add_786358;
  wire [7:0] sel_786359;
  wire [7:0] add_786362;
  wire [7:0] sel_786363;
  wire [7:0] add_786366;
  wire [7:0] sel_786367;
  wire [7:0] add_786370;
  wire [7:0] sel_786371;
  wire [7:0] add_786374;
  wire [7:0] sel_786375;
  wire [7:0] add_786378;
  wire [7:0] sel_786379;
  wire [7:0] add_786382;
  wire [7:0] sel_786383;
  wire [7:0] add_786386;
  wire [7:0] sel_786387;
  wire [7:0] add_786390;
  wire [7:0] sel_786391;
  wire [7:0] add_786394;
  wire [7:0] sel_786395;
  wire [7:0] add_786398;
  wire [7:0] sel_786399;
  wire [7:0] add_786402;
  wire [7:0] sel_786403;
  wire [7:0] add_786406;
  wire [7:0] sel_786407;
  wire [7:0] add_786410;
  wire [7:0] sel_786411;
  wire [7:0] add_786414;
  wire [7:0] sel_786415;
  wire [7:0] add_786418;
  wire [7:0] sel_786419;
  wire [7:0] add_786422;
  wire [7:0] sel_786423;
  wire [7:0] add_786426;
  wire [7:0] sel_786427;
  wire [7:0] add_786430;
  wire [7:0] sel_786431;
  wire [7:0] add_786434;
  wire [7:0] sel_786435;
  wire [7:0] add_786438;
  wire [7:0] sel_786439;
  wire [7:0] add_786442;
  wire [7:0] sel_786443;
  wire [7:0] add_786446;
  wire [7:0] sel_786447;
  wire [7:0] add_786450;
  wire [7:0] sel_786451;
  wire [7:0] add_786454;
  wire [7:0] sel_786455;
  wire [7:0] add_786458;
  wire [7:0] sel_786459;
  wire [7:0] add_786462;
  wire [7:0] sel_786463;
  wire [7:0] add_786466;
  wire [7:0] sel_786467;
  wire [7:0] add_786470;
  wire [7:0] sel_786471;
  wire [7:0] add_786474;
  wire [7:0] sel_786475;
  wire [7:0] add_786478;
  wire [7:0] sel_786479;
  wire [7:0] add_786482;
  wire [7:0] sel_786483;
  wire [7:0] add_786486;
  wire [7:0] sel_786487;
  wire [7:0] add_786490;
  wire [7:0] sel_786491;
  wire [7:0] add_786494;
  wire [7:0] sel_786495;
  wire [7:0] add_786498;
  wire [7:0] sel_786499;
  wire [7:0] add_786502;
  wire [7:0] sel_786503;
  wire [7:0] add_786506;
  wire [7:0] sel_786507;
  wire [7:0] add_786510;
  wire [7:0] sel_786511;
  wire [7:0] add_786514;
  wire [7:0] sel_786515;
  wire [7:0] add_786518;
  wire [7:0] sel_786519;
  wire [7:0] add_786522;
  wire [7:0] sel_786523;
  wire [7:0] add_786526;
  wire [7:0] sel_786527;
  wire [7:0] add_786530;
  wire [7:0] sel_786531;
  wire [7:0] add_786534;
  wire [7:0] sel_786535;
  wire [7:0] add_786538;
  wire [7:0] sel_786539;
  wire [7:0] add_786542;
  wire [7:0] sel_786543;
  wire [7:0] add_786546;
  wire [7:0] sel_786547;
  wire [7:0] add_786550;
  wire [7:0] sel_786551;
  wire [7:0] add_786554;
  wire [7:0] sel_786555;
  wire [7:0] add_786558;
  wire [7:0] sel_786559;
  wire [7:0] add_786562;
  wire [7:0] sel_786563;
  wire [7:0] add_786566;
  wire [7:0] sel_786567;
  wire [7:0] add_786570;
  wire [7:0] sel_786571;
  wire [7:0] add_786575;
  wire [15:0] array_index_786576;
  wire [7:0] sel_786577;
  wire [7:0] add_786580;
  wire [7:0] sel_786581;
  wire [7:0] add_786584;
  wire [7:0] sel_786585;
  wire [7:0] add_786588;
  wire [7:0] sel_786589;
  wire [7:0] add_786592;
  wire [7:0] sel_786593;
  wire [7:0] add_786596;
  wire [7:0] sel_786597;
  wire [7:0] add_786600;
  wire [7:0] sel_786601;
  wire [7:0] add_786604;
  wire [7:0] sel_786605;
  wire [7:0] add_786608;
  wire [7:0] sel_786609;
  wire [7:0] add_786612;
  wire [7:0] sel_786613;
  wire [7:0] add_786616;
  wire [7:0] sel_786617;
  wire [7:0] add_786620;
  wire [7:0] sel_786621;
  wire [7:0] add_786624;
  wire [7:0] sel_786625;
  wire [7:0] add_786628;
  wire [7:0] sel_786629;
  wire [7:0] add_786632;
  wire [7:0] sel_786633;
  wire [7:0] add_786636;
  wire [7:0] sel_786637;
  wire [7:0] add_786640;
  wire [7:0] sel_786641;
  wire [7:0] add_786644;
  wire [7:0] sel_786645;
  wire [7:0] add_786648;
  wire [7:0] sel_786649;
  wire [7:0] add_786652;
  wire [7:0] sel_786653;
  wire [7:0] add_786656;
  wire [7:0] sel_786657;
  wire [7:0] add_786660;
  wire [7:0] sel_786661;
  wire [7:0] add_786664;
  wire [7:0] sel_786665;
  wire [7:0] add_786668;
  wire [7:0] sel_786669;
  wire [7:0] add_786672;
  wire [7:0] sel_786673;
  wire [7:0] add_786676;
  wire [7:0] sel_786677;
  wire [7:0] add_786680;
  wire [7:0] sel_786681;
  wire [7:0] add_786684;
  wire [7:0] sel_786685;
  wire [7:0] add_786688;
  wire [7:0] sel_786689;
  wire [7:0] add_786692;
  wire [7:0] sel_786693;
  wire [7:0] add_786696;
  wire [7:0] sel_786697;
  wire [7:0] add_786700;
  wire [7:0] sel_786701;
  wire [7:0] add_786704;
  wire [7:0] sel_786705;
  wire [7:0] add_786708;
  wire [7:0] sel_786709;
  wire [7:0] add_786712;
  wire [7:0] sel_786713;
  wire [7:0] add_786716;
  wire [7:0] sel_786717;
  wire [7:0] add_786720;
  wire [7:0] sel_786721;
  wire [7:0] add_786724;
  wire [7:0] sel_786725;
  wire [7:0] add_786728;
  wire [7:0] sel_786729;
  wire [7:0] add_786732;
  wire [7:0] sel_786733;
  wire [7:0] add_786736;
  wire [7:0] sel_786737;
  wire [7:0] add_786740;
  wire [7:0] sel_786741;
  wire [7:0] add_786744;
  wire [7:0] sel_786745;
  wire [7:0] add_786748;
  wire [7:0] sel_786749;
  wire [7:0] add_786752;
  wire [7:0] sel_786753;
  wire [7:0] add_786756;
  wire [7:0] sel_786757;
  wire [7:0] add_786760;
  wire [7:0] sel_786761;
  wire [7:0] add_786764;
  wire [7:0] sel_786765;
  wire [7:0] add_786768;
  wire [7:0] sel_786769;
  wire [7:0] add_786772;
  wire [7:0] sel_786773;
  wire [7:0] add_786776;
  wire [7:0] sel_786777;
  wire [7:0] add_786780;
  wire [7:0] sel_786781;
  wire [7:0] add_786784;
  wire [7:0] sel_786785;
  wire [7:0] add_786788;
  wire [7:0] sel_786789;
  wire [7:0] add_786792;
  wire [7:0] sel_786793;
  wire [7:0] add_786796;
  wire [7:0] sel_786797;
  wire [7:0] add_786800;
  wire [7:0] sel_786801;
  wire [7:0] add_786804;
  wire [7:0] sel_786805;
  wire [7:0] add_786808;
  wire [7:0] sel_786809;
  wire [7:0] add_786812;
  wire [7:0] sel_786813;
  wire [7:0] add_786816;
  wire [7:0] sel_786817;
  wire [7:0] add_786820;
  wire [7:0] sel_786821;
  wire [7:0] add_786824;
  wire [7:0] sel_786825;
  wire [7:0] add_786828;
  wire [7:0] sel_786829;
  wire [7:0] add_786832;
  wire [7:0] sel_786833;
  wire [7:0] add_786836;
  wire [7:0] sel_786837;
  wire [7:0] add_786840;
  wire [7:0] sel_786841;
  wire [7:0] add_786844;
  wire [7:0] sel_786845;
  wire [7:0] add_786848;
  wire [7:0] sel_786849;
  wire [7:0] add_786852;
  wire [7:0] sel_786853;
  wire [7:0] add_786856;
  wire [7:0] sel_786857;
  wire [7:0] add_786860;
  wire [7:0] sel_786861;
  wire [7:0] add_786864;
  wire [7:0] sel_786865;
  wire [7:0] add_786868;
  wire [7:0] sel_786869;
  wire [7:0] add_786872;
  wire [7:0] sel_786873;
  wire [7:0] add_786876;
  wire [7:0] sel_786877;
  wire [7:0] add_786880;
  wire [7:0] sel_786881;
  wire [7:0] add_786884;
  wire [7:0] sel_786885;
  wire [7:0] add_786888;
  wire [7:0] sel_786889;
  wire [7:0] add_786892;
  wire [7:0] sel_786893;
  wire [7:0] add_786896;
  wire [7:0] sel_786897;
  wire [7:0] add_786900;
  wire [7:0] sel_786901;
  wire [7:0] add_786904;
  wire [7:0] sel_786905;
  wire [7:0] add_786908;
  wire [7:0] sel_786909;
  wire [7:0] add_786912;
  wire [7:0] sel_786913;
  wire [7:0] add_786916;
  wire [7:0] sel_786917;
  wire [7:0] add_786920;
  wire [7:0] sel_786921;
  wire [7:0] add_786924;
  wire [7:0] sel_786925;
  wire [7:0] add_786928;
  wire [7:0] sel_786929;
  wire [7:0] add_786932;
  wire [7:0] sel_786933;
  wire [7:0] add_786937;
  wire [15:0] array_index_786938;
  wire [7:0] sel_786939;
  wire [7:0] add_786942;
  wire [7:0] sel_786943;
  wire [7:0] add_786946;
  wire [7:0] sel_786947;
  wire [7:0] add_786950;
  wire [7:0] sel_786951;
  wire [7:0] add_786954;
  wire [7:0] sel_786955;
  wire [7:0] add_786958;
  wire [7:0] sel_786959;
  wire [7:0] add_786962;
  wire [7:0] sel_786963;
  wire [7:0] add_786966;
  wire [7:0] sel_786967;
  wire [7:0] add_786970;
  wire [7:0] sel_786971;
  wire [7:0] add_786974;
  wire [7:0] sel_786975;
  wire [7:0] add_786978;
  wire [7:0] sel_786979;
  wire [7:0] add_786982;
  wire [7:0] sel_786983;
  wire [7:0] add_786986;
  wire [7:0] sel_786987;
  wire [7:0] add_786990;
  wire [7:0] sel_786991;
  wire [7:0] add_786994;
  wire [7:0] sel_786995;
  wire [7:0] add_786998;
  wire [7:0] sel_786999;
  wire [7:0] add_787002;
  wire [7:0] sel_787003;
  wire [7:0] add_787006;
  wire [7:0] sel_787007;
  wire [7:0] add_787010;
  wire [7:0] sel_787011;
  wire [7:0] add_787014;
  wire [7:0] sel_787015;
  wire [7:0] add_787018;
  wire [7:0] sel_787019;
  wire [7:0] add_787022;
  wire [7:0] sel_787023;
  wire [7:0] add_787026;
  wire [7:0] sel_787027;
  wire [7:0] add_787030;
  wire [7:0] sel_787031;
  wire [7:0] add_787034;
  wire [7:0] sel_787035;
  wire [7:0] add_787038;
  wire [7:0] sel_787039;
  wire [7:0] add_787042;
  wire [7:0] sel_787043;
  wire [7:0] add_787046;
  wire [7:0] sel_787047;
  wire [7:0] add_787050;
  wire [7:0] sel_787051;
  wire [7:0] add_787054;
  wire [7:0] sel_787055;
  wire [7:0] add_787058;
  wire [7:0] sel_787059;
  wire [7:0] add_787062;
  wire [7:0] sel_787063;
  wire [7:0] add_787066;
  wire [7:0] sel_787067;
  wire [7:0] add_787070;
  wire [7:0] sel_787071;
  wire [7:0] add_787074;
  wire [7:0] sel_787075;
  wire [7:0] add_787078;
  wire [7:0] sel_787079;
  wire [7:0] add_787082;
  wire [7:0] sel_787083;
  wire [7:0] add_787086;
  wire [7:0] sel_787087;
  wire [7:0] add_787090;
  wire [7:0] sel_787091;
  wire [7:0] add_787094;
  wire [7:0] sel_787095;
  wire [7:0] add_787098;
  wire [7:0] sel_787099;
  wire [7:0] add_787102;
  wire [7:0] sel_787103;
  wire [7:0] add_787106;
  wire [7:0] sel_787107;
  wire [7:0] add_787110;
  wire [7:0] sel_787111;
  wire [7:0] add_787114;
  wire [7:0] sel_787115;
  wire [7:0] add_787118;
  wire [7:0] sel_787119;
  wire [7:0] add_787122;
  wire [7:0] sel_787123;
  wire [7:0] add_787126;
  wire [7:0] sel_787127;
  wire [7:0] add_787130;
  wire [7:0] sel_787131;
  wire [7:0] add_787134;
  wire [7:0] sel_787135;
  wire [7:0] add_787138;
  wire [7:0] sel_787139;
  wire [7:0] add_787142;
  wire [7:0] sel_787143;
  wire [7:0] add_787146;
  wire [7:0] sel_787147;
  wire [7:0] add_787150;
  wire [7:0] sel_787151;
  wire [7:0] add_787154;
  wire [7:0] sel_787155;
  wire [7:0] add_787158;
  wire [7:0] sel_787159;
  wire [7:0] add_787162;
  wire [7:0] sel_787163;
  wire [7:0] add_787166;
  wire [7:0] sel_787167;
  wire [7:0] add_787170;
  wire [7:0] sel_787171;
  wire [7:0] add_787174;
  wire [7:0] sel_787175;
  wire [7:0] add_787178;
  wire [7:0] sel_787179;
  wire [7:0] add_787182;
  wire [7:0] sel_787183;
  wire [7:0] add_787186;
  wire [7:0] sel_787187;
  wire [7:0] add_787190;
  wire [7:0] sel_787191;
  wire [7:0] add_787194;
  wire [7:0] sel_787195;
  wire [7:0] add_787198;
  wire [7:0] sel_787199;
  wire [7:0] add_787202;
  wire [7:0] sel_787203;
  wire [7:0] add_787206;
  wire [7:0] sel_787207;
  wire [7:0] add_787210;
  wire [7:0] sel_787211;
  wire [7:0] add_787214;
  wire [7:0] sel_787215;
  wire [7:0] add_787218;
  wire [7:0] sel_787219;
  wire [7:0] add_787222;
  wire [7:0] sel_787223;
  wire [7:0] add_787226;
  wire [7:0] sel_787227;
  wire [7:0] add_787230;
  wire [7:0] sel_787231;
  wire [7:0] add_787234;
  wire [7:0] sel_787235;
  wire [7:0] add_787238;
  wire [7:0] sel_787239;
  wire [7:0] add_787242;
  wire [7:0] sel_787243;
  wire [7:0] add_787246;
  wire [7:0] sel_787247;
  wire [7:0] add_787250;
  wire [7:0] sel_787251;
  wire [7:0] add_787254;
  wire [7:0] sel_787255;
  wire [7:0] add_787258;
  wire [7:0] sel_787259;
  wire [7:0] add_787262;
  wire [7:0] sel_787263;
  wire [7:0] add_787266;
  wire [7:0] sel_787267;
  wire [7:0] add_787270;
  wire [7:0] sel_787271;
  wire [7:0] add_787274;
  wire [7:0] sel_787275;
  wire [7:0] add_787278;
  wire [7:0] sel_787279;
  wire [7:0] add_787282;
  wire [7:0] sel_787283;
  wire [7:0] add_787286;
  wire [7:0] sel_787287;
  wire [7:0] add_787290;
  wire [7:0] sel_787291;
  wire [7:0] add_787294;
  wire [7:0] sel_787295;
  wire [7:0] add_787299;
  wire [15:0] array_index_787300;
  wire [7:0] sel_787301;
  wire [7:0] add_787304;
  wire [7:0] sel_787305;
  wire [7:0] add_787308;
  wire [7:0] sel_787309;
  wire [7:0] add_787312;
  wire [7:0] sel_787313;
  wire [7:0] add_787316;
  wire [7:0] sel_787317;
  wire [7:0] add_787320;
  wire [7:0] sel_787321;
  wire [7:0] add_787324;
  wire [7:0] sel_787325;
  wire [7:0] add_787328;
  wire [7:0] sel_787329;
  wire [7:0] add_787332;
  wire [7:0] sel_787333;
  wire [7:0] add_787336;
  wire [7:0] sel_787337;
  wire [7:0] add_787340;
  wire [7:0] sel_787341;
  wire [7:0] add_787344;
  wire [7:0] sel_787345;
  wire [7:0] add_787348;
  wire [7:0] sel_787349;
  wire [7:0] add_787352;
  wire [7:0] sel_787353;
  wire [7:0] add_787356;
  wire [7:0] sel_787357;
  wire [7:0] add_787360;
  wire [7:0] sel_787361;
  wire [7:0] add_787364;
  wire [7:0] sel_787365;
  wire [7:0] add_787368;
  wire [7:0] sel_787369;
  wire [7:0] add_787372;
  wire [7:0] sel_787373;
  wire [7:0] add_787376;
  wire [7:0] sel_787377;
  wire [7:0] add_787380;
  wire [7:0] sel_787381;
  wire [7:0] add_787384;
  wire [7:0] sel_787385;
  wire [7:0] add_787388;
  wire [7:0] sel_787389;
  wire [7:0] add_787392;
  wire [7:0] sel_787393;
  wire [7:0] add_787396;
  wire [7:0] sel_787397;
  wire [7:0] add_787400;
  wire [7:0] sel_787401;
  wire [7:0] add_787404;
  wire [7:0] sel_787405;
  wire [7:0] add_787408;
  wire [7:0] sel_787409;
  wire [7:0] add_787412;
  wire [7:0] sel_787413;
  wire [7:0] add_787416;
  wire [7:0] sel_787417;
  wire [7:0] add_787420;
  wire [7:0] sel_787421;
  wire [7:0] add_787424;
  wire [7:0] sel_787425;
  wire [7:0] add_787428;
  wire [7:0] sel_787429;
  wire [7:0] add_787432;
  wire [7:0] sel_787433;
  wire [7:0] add_787436;
  wire [7:0] sel_787437;
  wire [7:0] add_787440;
  wire [7:0] sel_787441;
  wire [7:0] add_787444;
  wire [7:0] sel_787445;
  wire [7:0] add_787448;
  wire [7:0] sel_787449;
  wire [7:0] add_787452;
  wire [7:0] sel_787453;
  wire [7:0] add_787456;
  wire [7:0] sel_787457;
  wire [7:0] add_787460;
  wire [7:0] sel_787461;
  wire [7:0] add_787464;
  wire [7:0] sel_787465;
  wire [7:0] add_787468;
  wire [7:0] sel_787469;
  wire [7:0] add_787472;
  wire [7:0] sel_787473;
  wire [7:0] add_787476;
  wire [7:0] sel_787477;
  wire [7:0] add_787480;
  wire [7:0] sel_787481;
  wire [7:0] add_787484;
  wire [7:0] sel_787485;
  wire [7:0] add_787488;
  wire [7:0] sel_787489;
  wire [7:0] add_787492;
  wire [7:0] sel_787493;
  wire [7:0] add_787496;
  wire [7:0] sel_787497;
  wire [7:0] add_787500;
  wire [7:0] sel_787501;
  wire [7:0] add_787504;
  wire [7:0] sel_787505;
  wire [7:0] add_787508;
  wire [7:0] sel_787509;
  wire [7:0] add_787512;
  wire [7:0] sel_787513;
  wire [7:0] add_787516;
  wire [7:0] sel_787517;
  wire [7:0] add_787520;
  wire [7:0] sel_787521;
  wire [7:0] add_787524;
  wire [7:0] sel_787525;
  wire [7:0] add_787528;
  wire [7:0] sel_787529;
  wire [7:0] add_787532;
  wire [7:0] sel_787533;
  wire [7:0] add_787536;
  wire [7:0] sel_787537;
  wire [7:0] add_787540;
  wire [7:0] sel_787541;
  wire [7:0] add_787544;
  wire [7:0] sel_787545;
  wire [7:0] add_787548;
  wire [7:0] sel_787549;
  wire [7:0] add_787552;
  wire [7:0] sel_787553;
  wire [7:0] add_787556;
  wire [7:0] sel_787557;
  wire [7:0] add_787560;
  wire [7:0] sel_787561;
  wire [7:0] add_787564;
  wire [7:0] sel_787565;
  wire [7:0] add_787568;
  wire [7:0] sel_787569;
  wire [7:0] add_787572;
  wire [7:0] sel_787573;
  wire [7:0] add_787576;
  wire [7:0] sel_787577;
  wire [7:0] add_787580;
  wire [7:0] sel_787581;
  wire [7:0] add_787584;
  wire [7:0] sel_787585;
  wire [7:0] add_787588;
  wire [7:0] sel_787589;
  wire [7:0] add_787592;
  wire [7:0] sel_787593;
  wire [7:0] add_787596;
  wire [7:0] sel_787597;
  wire [7:0] add_787600;
  wire [7:0] sel_787601;
  wire [7:0] add_787604;
  wire [7:0] sel_787605;
  wire [7:0] add_787608;
  wire [7:0] sel_787609;
  wire [7:0] add_787612;
  wire [7:0] sel_787613;
  wire [7:0] add_787616;
  wire [7:0] sel_787617;
  wire [7:0] add_787620;
  wire [7:0] sel_787621;
  wire [7:0] add_787624;
  wire [7:0] sel_787625;
  wire [7:0] add_787628;
  wire [7:0] sel_787629;
  wire [7:0] add_787632;
  wire [7:0] sel_787633;
  wire [7:0] add_787636;
  wire [7:0] sel_787637;
  wire [7:0] add_787640;
  wire [7:0] sel_787641;
  wire [7:0] add_787644;
  wire [7:0] sel_787645;
  wire [7:0] add_787648;
  wire [7:0] sel_787649;
  wire [7:0] add_787652;
  wire [7:0] sel_787653;
  wire [7:0] add_787656;
  wire [7:0] sel_787657;
  wire [7:0] add_787661;
  wire [15:0] array_index_787662;
  wire [7:0] sel_787663;
  wire [7:0] add_787666;
  wire [7:0] sel_787667;
  wire [7:0] add_787670;
  wire [7:0] sel_787671;
  wire [7:0] add_787674;
  wire [7:0] sel_787675;
  wire [7:0] add_787678;
  wire [7:0] sel_787679;
  wire [7:0] add_787682;
  wire [7:0] sel_787683;
  wire [7:0] add_787686;
  wire [7:0] sel_787687;
  wire [7:0] add_787690;
  wire [7:0] sel_787691;
  wire [7:0] add_787694;
  wire [7:0] sel_787695;
  wire [7:0] add_787698;
  wire [7:0] sel_787699;
  wire [7:0] add_787702;
  wire [7:0] sel_787703;
  wire [7:0] add_787706;
  wire [7:0] sel_787707;
  wire [7:0] add_787710;
  wire [7:0] sel_787711;
  wire [7:0] add_787714;
  wire [7:0] sel_787715;
  wire [7:0] add_787718;
  wire [7:0] sel_787719;
  wire [7:0] add_787722;
  wire [7:0] sel_787723;
  wire [7:0] add_787726;
  wire [7:0] sel_787727;
  wire [7:0] add_787730;
  wire [7:0] sel_787731;
  wire [7:0] add_787734;
  wire [7:0] sel_787735;
  wire [7:0] add_787738;
  wire [7:0] sel_787739;
  wire [7:0] add_787742;
  wire [7:0] sel_787743;
  wire [7:0] add_787746;
  wire [7:0] sel_787747;
  wire [7:0] add_787750;
  wire [7:0] sel_787751;
  wire [7:0] add_787754;
  wire [7:0] sel_787755;
  wire [7:0] add_787758;
  wire [7:0] sel_787759;
  wire [7:0] add_787762;
  wire [7:0] sel_787763;
  wire [7:0] add_787766;
  wire [7:0] sel_787767;
  wire [7:0] add_787770;
  wire [7:0] sel_787771;
  wire [7:0] add_787774;
  wire [7:0] sel_787775;
  wire [7:0] add_787778;
  wire [7:0] sel_787779;
  wire [7:0] add_787782;
  wire [7:0] sel_787783;
  wire [7:0] add_787786;
  wire [7:0] sel_787787;
  wire [7:0] add_787790;
  wire [7:0] sel_787791;
  wire [7:0] add_787794;
  wire [7:0] sel_787795;
  wire [7:0] add_787798;
  wire [7:0] sel_787799;
  wire [7:0] add_787802;
  wire [7:0] sel_787803;
  wire [7:0] add_787806;
  wire [7:0] sel_787807;
  wire [7:0] add_787810;
  wire [7:0] sel_787811;
  wire [7:0] add_787814;
  wire [7:0] sel_787815;
  wire [7:0] add_787818;
  wire [7:0] sel_787819;
  wire [7:0] add_787822;
  wire [7:0] sel_787823;
  wire [7:0] add_787826;
  wire [7:0] sel_787827;
  wire [7:0] add_787830;
  wire [7:0] sel_787831;
  wire [7:0] add_787834;
  wire [7:0] sel_787835;
  wire [7:0] add_787838;
  wire [7:0] sel_787839;
  wire [7:0] add_787842;
  wire [7:0] sel_787843;
  wire [7:0] add_787846;
  wire [7:0] sel_787847;
  wire [7:0] add_787850;
  wire [7:0] sel_787851;
  wire [7:0] add_787854;
  wire [7:0] sel_787855;
  wire [7:0] add_787858;
  wire [7:0] sel_787859;
  wire [7:0] add_787862;
  wire [7:0] sel_787863;
  wire [7:0] add_787866;
  wire [7:0] sel_787867;
  wire [7:0] add_787870;
  wire [7:0] sel_787871;
  wire [7:0] add_787874;
  wire [7:0] sel_787875;
  wire [7:0] add_787878;
  wire [7:0] sel_787879;
  wire [7:0] add_787882;
  wire [7:0] sel_787883;
  wire [7:0] add_787886;
  wire [7:0] sel_787887;
  wire [7:0] add_787890;
  wire [7:0] sel_787891;
  wire [7:0] add_787894;
  wire [7:0] sel_787895;
  wire [7:0] add_787898;
  wire [7:0] sel_787899;
  wire [7:0] add_787902;
  wire [7:0] sel_787903;
  wire [7:0] add_787906;
  wire [7:0] sel_787907;
  wire [7:0] add_787910;
  wire [7:0] sel_787911;
  wire [7:0] add_787914;
  wire [7:0] sel_787915;
  wire [7:0] add_787918;
  wire [7:0] sel_787919;
  wire [7:0] add_787922;
  wire [7:0] sel_787923;
  wire [7:0] add_787926;
  wire [7:0] sel_787927;
  wire [7:0] add_787930;
  wire [7:0] sel_787931;
  wire [7:0] add_787934;
  wire [7:0] sel_787935;
  wire [7:0] add_787938;
  wire [7:0] sel_787939;
  wire [7:0] add_787942;
  wire [7:0] sel_787943;
  wire [7:0] add_787946;
  wire [7:0] sel_787947;
  wire [7:0] add_787950;
  wire [7:0] sel_787951;
  wire [7:0] add_787954;
  wire [7:0] sel_787955;
  wire [7:0] add_787958;
  wire [7:0] sel_787959;
  wire [7:0] add_787962;
  wire [7:0] sel_787963;
  wire [7:0] add_787966;
  wire [7:0] sel_787967;
  wire [7:0] add_787970;
  wire [7:0] sel_787971;
  wire [7:0] add_787974;
  wire [7:0] sel_787975;
  wire [7:0] add_787978;
  wire [7:0] sel_787979;
  wire [7:0] add_787982;
  wire [7:0] sel_787983;
  wire [7:0] add_787986;
  wire [7:0] sel_787987;
  wire [7:0] add_787990;
  wire [7:0] sel_787991;
  wire [7:0] add_787994;
  wire [7:0] sel_787995;
  wire [7:0] add_787998;
  wire [7:0] sel_787999;
  wire [7:0] add_788002;
  wire [7:0] sel_788003;
  wire [7:0] add_788006;
  wire [7:0] sel_788007;
  wire [7:0] add_788010;
  wire [7:0] sel_788011;
  wire [7:0] add_788014;
  wire [7:0] sel_788015;
  wire [7:0] add_788018;
  wire [7:0] sel_788019;
  wire [7:0] add_788023;
  wire [15:0] array_index_788024;
  wire [7:0] sel_788025;
  wire [7:0] add_788028;
  wire [7:0] sel_788029;
  wire [7:0] add_788032;
  wire [7:0] sel_788033;
  wire [7:0] add_788036;
  wire [7:0] sel_788037;
  wire [7:0] add_788040;
  wire [7:0] sel_788041;
  wire [7:0] add_788044;
  wire [7:0] sel_788045;
  wire [7:0] add_788048;
  wire [7:0] sel_788049;
  wire [7:0] add_788052;
  wire [7:0] sel_788053;
  wire [7:0] add_788056;
  wire [7:0] sel_788057;
  wire [7:0] add_788060;
  wire [7:0] sel_788061;
  wire [7:0] add_788064;
  wire [7:0] sel_788065;
  wire [7:0] add_788068;
  wire [7:0] sel_788069;
  wire [7:0] add_788072;
  wire [7:0] sel_788073;
  wire [7:0] add_788076;
  wire [7:0] sel_788077;
  wire [7:0] add_788080;
  wire [7:0] sel_788081;
  wire [7:0] add_788084;
  wire [7:0] sel_788085;
  wire [7:0] add_788088;
  wire [7:0] sel_788089;
  wire [7:0] add_788092;
  wire [7:0] sel_788093;
  wire [7:0] add_788096;
  wire [7:0] sel_788097;
  wire [7:0] add_788100;
  wire [7:0] sel_788101;
  wire [7:0] add_788104;
  wire [7:0] sel_788105;
  wire [7:0] add_788108;
  wire [7:0] sel_788109;
  wire [7:0] add_788112;
  wire [7:0] sel_788113;
  wire [7:0] add_788116;
  wire [7:0] sel_788117;
  wire [7:0] add_788120;
  wire [7:0] sel_788121;
  wire [7:0] add_788124;
  wire [7:0] sel_788125;
  wire [7:0] add_788128;
  wire [7:0] sel_788129;
  wire [7:0] add_788132;
  wire [7:0] sel_788133;
  wire [7:0] add_788136;
  wire [7:0] sel_788137;
  wire [7:0] add_788140;
  wire [7:0] sel_788141;
  wire [7:0] add_788144;
  wire [7:0] sel_788145;
  wire [7:0] add_788148;
  wire [7:0] sel_788149;
  wire [7:0] add_788152;
  wire [7:0] sel_788153;
  wire [7:0] add_788156;
  wire [7:0] sel_788157;
  wire [7:0] add_788160;
  wire [7:0] sel_788161;
  wire [7:0] add_788164;
  wire [7:0] sel_788165;
  wire [7:0] add_788168;
  wire [7:0] sel_788169;
  wire [7:0] add_788172;
  wire [7:0] sel_788173;
  wire [7:0] add_788176;
  wire [7:0] sel_788177;
  wire [7:0] add_788180;
  wire [7:0] sel_788181;
  wire [7:0] add_788184;
  wire [7:0] sel_788185;
  wire [7:0] add_788188;
  wire [7:0] sel_788189;
  wire [7:0] add_788192;
  wire [7:0] sel_788193;
  wire [7:0] add_788196;
  wire [7:0] sel_788197;
  wire [7:0] add_788200;
  wire [7:0] sel_788201;
  wire [7:0] add_788204;
  wire [7:0] sel_788205;
  wire [7:0] add_788208;
  wire [7:0] sel_788209;
  wire [7:0] add_788212;
  wire [7:0] sel_788213;
  wire [7:0] add_788216;
  wire [7:0] sel_788217;
  wire [7:0] add_788220;
  wire [7:0] sel_788221;
  wire [7:0] add_788224;
  wire [7:0] sel_788225;
  wire [7:0] add_788228;
  wire [7:0] sel_788229;
  wire [7:0] add_788232;
  wire [7:0] sel_788233;
  wire [7:0] add_788236;
  wire [7:0] sel_788237;
  wire [7:0] add_788240;
  wire [7:0] sel_788241;
  wire [7:0] add_788244;
  wire [7:0] sel_788245;
  wire [7:0] add_788248;
  wire [7:0] sel_788249;
  wire [7:0] add_788252;
  wire [7:0] sel_788253;
  wire [7:0] add_788256;
  wire [7:0] sel_788257;
  wire [7:0] add_788260;
  wire [7:0] sel_788261;
  wire [7:0] add_788264;
  wire [7:0] sel_788265;
  wire [7:0] add_788268;
  wire [7:0] sel_788269;
  wire [7:0] add_788272;
  wire [7:0] sel_788273;
  wire [7:0] add_788276;
  wire [7:0] sel_788277;
  wire [7:0] add_788280;
  wire [7:0] sel_788281;
  wire [7:0] add_788284;
  wire [7:0] sel_788285;
  wire [7:0] add_788288;
  wire [7:0] sel_788289;
  wire [7:0] add_788292;
  wire [7:0] sel_788293;
  wire [7:0] add_788296;
  wire [7:0] sel_788297;
  wire [7:0] add_788300;
  wire [7:0] sel_788301;
  wire [7:0] add_788304;
  wire [7:0] sel_788305;
  wire [7:0] add_788308;
  wire [7:0] sel_788309;
  wire [7:0] add_788312;
  wire [7:0] sel_788313;
  wire [7:0] add_788316;
  wire [7:0] sel_788317;
  wire [7:0] add_788320;
  wire [7:0] sel_788321;
  wire [7:0] add_788324;
  wire [7:0] sel_788325;
  wire [7:0] add_788328;
  wire [7:0] sel_788329;
  wire [7:0] add_788332;
  wire [7:0] sel_788333;
  wire [7:0] add_788336;
  wire [7:0] sel_788337;
  wire [7:0] add_788340;
  wire [7:0] sel_788341;
  wire [7:0] add_788344;
  wire [7:0] sel_788345;
  wire [7:0] add_788348;
  wire [7:0] sel_788349;
  wire [7:0] add_788352;
  wire [7:0] sel_788353;
  wire [7:0] add_788356;
  wire [7:0] sel_788357;
  wire [7:0] add_788360;
  wire [7:0] sel_788361;
  wire [7:0] add_788364;
  wire [7:0] sel_788365;
  wire [7:0] add_788368;
  wire [7:0] sel_788369;
  wire [7:0] add_788372;
  wire [7:0] sel_788373;
  wire [7:0] add_788376;
  wire [7:0] sel_788377;
  wire [7:0] add_788380;
  wire [7:0] sel_788381;
  wire [7:0] add_788385;
  wire [15:0] array_index_788386;
  wire [7:0] sel_788387;
  wire [7:0] add_788390;
  wire [7:0] sel_788391;
  wire [7:0] add_788394;
  wire [7:0] sel_788395;
  wire [7:0] add_788398;
  wire [7:0] sel_788399;
  wire [7:0] add_788402;
  wire [7:0] sel_788403;
  wire [7:0] add_788406;
  wire [7:0] sel_788407;
  wire [7:0] add_788410;
  wire [7:0] sel_788411;
  wire [7:0] add_788414;
  wire [7:0] sel_788415;
  wire [7:0] add_788418;
  wire [7:0] sel_788419;
  wire [7:0] add_788422;
  wire [7:0] sel_788423;
  wire [7:0] add_788426;
  wire [7:0] sel_788427;
  wire [7:0] add_788430;
  wire [7:0] sel_788431;
  wire [7:0] add_788434;
  wire [7:0] sel_788435;
  wire [7:0] add_788438;
  wire [7:0] sel_788439;
  wire [7:0] add_788442;
  wire [7:0] sel_788443;
  wire [7:0] add_788446;
  wire [7:0] sel_788447;
  wire [7:0] add_788450;
  wire [7:0] sel_788451;
  wire [7:0] add_788454;
  wire [7:0] sel_788455;
  wire [7:0] add_788458;
  wire [7:0] sel_788459;
  wire [7:0] add_788462;
  wire [7:0] sel_788463;
  wire [7:0] add_788466;
  wire [7:0] sel_788467;
  wire [7:0] add_788470;
  wire [7:0] sel_788471;
  wire [7:0] add_788474;
  wire [7:0] sel_788475;
  wire [7:0] add_788478;
  wire [7:0] sel_788479;
  wire [7:0] add_788482;
  wire [7:0] sel_788483;
  wire [7:0] add_788486;
  wire [7:0] sel_788487;
  wire [7:0] add_788490;
  wire [7:0] sel_788491;
  wire [7:0] add_788494;
  wire [7:0] sel_788495;
  wire [7:0] add_788498;
  wire [7:0] sel_788499;
  wire [7:0] add_788502;
  wire [7:0] sel_788503;
  wire [7:0] add_788506;
  wire [7:0] sel_788507;
  wire [7:0] add_788510;
  wire [7:0] sel_788511;
  wire [7:0] add_788514;
  wire [7:0] sel_788515;
  wire [7:0] add_788518;
  wire [7:0] sel_788519;
  wire [7:0] add_788522;
  wire [7:0] sel_788523;
  wire [7:0] add_788526;
  wire [7:0] sel_788527;
  wire [7:0] add_788530;
  wire [7:0] sel_788531;
  wire [7:0] add_788534;
  wire [7:0] sel_788535;
  wire [7:0] add_788538;
  wire [7:0] sel_788539;
  wire [7:0] add_788542;
  wire [7:0] sel_788543;
  wire [7:0] add_788546;
  wire [7:0] sel_788547;
  wire [7:0] add_788550;
  wire [7:0] sel_788551;
  wire [7:0] add_788554;
  wire [7:0] sel_788555;
  wire [7:0] add_788558;
  wire [7:0] sel_788559;
  wire [7:0] add_788562;
  wire [7:0] sel_788563;
  wire [7:0] add_788566;
  wire [7:0] sel_788567;
  wire [7:0] add_788570;
  wire [7:0] sel_788571;
  wire [7:0] add_788574;
  wire [7:0] sel_788575;
  wire [7:0] add_788578;
  wire [7:0] sel_788579;
  wire [7:0] add_788582;
  wire [7:0] sel_788583;
  wire [7:0] add_788586;
  wire [7:0] sel_788587;
  wire [7:0] add_788590;
  wire [7:0] sel_788591;
  wire [7:0] add_788594;
  wire [7:0] sel_788595;
  wire [7:0] add_788598;
  wire [7:0] sel_788599;
  wire [7:0] add_788602;
  wire [7:0] sel_788603;
  wire [7:0] add_788606;
  wire [7:0] sel_788607;
  wire [7:0] add_788610;
  wire [7:0] sel_788611;
  wire [7:0] add_788614;
  wire [7:0] sel_788615;
  wire [7:0] add_788618;
  wire [7:0] sel_788619;
  wire [7:0] add_788622;
  wire [7:0] sel_788623;
  wire [7:0] add_788626;
  wire [7:0] sel_788627;
  wire [7:0] add_788630;
  wire [7:0] sel_788631;
  wire [7:0] add_788634;
  wire [7:0] sel_788635;
  wire [7:0] add_788638;
  wire [7:0] sel_788639;
  wire [7:0] add_788642;
  wire [7:0] sel_788643;
  wire [7:0] add_788646;
  wire [7:0] sel_788647;
  wire [7:0] add_788650;
  wire [7:0] sel_788651;
  wire [7:0] add_788654;
  wire [7:0] sel_788655;
  wire [7:0] add_788658;
  wire [7:0] sel_788659;
  wire [7:0] add_788662;
  wire [7:0] sel_788663;
  wire [7:0] add_788666;
  wire [7:0] sel_788667;
  wire [7:0] add_788670;
  wire [7:0] sel_788671;
  wire [7:0] add_788674;
  wire [7:0] sel_788675;
  wire [7:0] add_788678;
  wire [7:0] sel_788679;
  wire [7:0] add_788682;
  wire [7:0] sel_788683;
  wire [7:0] add_788686;
  wire [7:0] sel_788687;
  wire [7:0] add_788690;
  wire [7:0] sel_788691;
  wire [7:0] add_788694;
  wire [7:0] sel_788695;
  wire [7:0] add_788698;
  wire [7:0] sel_788699;
  wire [7:0] add_788702;
  wire [7:0] sel_788703;
  wire [7:0] add_788706;
  wire [7:0] sel_788707;
  wire [7:0] add_788710;
  wire [7:0] sel_788711;
  wire [7:0] add_788714;
  wire [7:0] sel_788715;
  wire [7:0] add_788718;
  wire [7:0] sel_788719;
  wire [7:0] add_788722;
  wire [7:0] sel_788723;
  wire [7:0] add_788726;
  wire [7:0] sel_788727;
  wire [7:0] add_788730;
  wire [7:0] sel_788731;
  wire [7:0] add_788734;
  wire [7:0] sel_788735;
  wire [7:0] add_788738;
  wire [7:0] sel_788739;
  wire [7:0] add_788742;
  wire [7:0] sel_788743;
  wire [7:0] add_788747;
  wire [15:0] array_index_788748;
  wire [7:0] sel_788749;
  wire [7:0] add_788752;
  wire [7:0] sel_788753;
  wire [7:0] add_788756;
  wire [7:0] sel_788757;
  wire [7:0] add_788760;
  wire [7:0] sel_788761;
  wire [7:0] add_788764;
  wire [7:0] sel_788765;
  wire [7:0] add_788768;
  wire [7:0] sel_788769;
  wire [7:0] add_788772;
  wire [7:0] sel_788773;
  wire [7:0] add_788776;
  wire [7:0] sel_788777;
  wire [7:0] add_788780;
  wire [7:0] sel_788781;
  wire [7:0] add_788784;
  wire [7:0] sel_788785;
  wire [7:0] add_788788;
  wire [7:0] sel_788789;
  wire [7:0] add_788792;
  wire [7:0] sel_788793;
  wire [7:0] add_788796;
  wire [7:0] sel_788797;
  wire [7:0] add_788800;
  wire [7:0] sel_788801;
  wire [7:0] add_788804;
  wire [7:0] sel_788805;
  wire [7:0] add_788808;
  wire [7:0] sel_788809;
  wire [7:0] add_788812;
  wire [7:0] sel_788813;
  wire [7:0] add_788816;
  wire [7:0] sel_788817;
  wire [7:0] add_788820;
  wire [7:0] sel_788821;
  wire [7:0] add_788824;
  wire [7:0] sel_788825;
  wire [7:0] add_788828;
  wire [7:0] sel_788829;
  wire [7:0] add_788832;
  wire [7:0] sel_788833;
  wire [7:0] add_788836;
  wire [7:0] sel_788837;
  wire [7:0] add_788840;
  wire [7:0] sel_788841;
  wire [7:0] add_788844;
  wire [7:0] sel_788845;
  wire [7:0] add_788848;
  wire [7:0] sel_788849;
  wire [7:0] add_788852;
  wire [7:0] sel_788853;
  wire [7:0] add_788856;
  wire [7:0] sel_788857;
  wire [7:0] add_788860;
  wire [7:0] sel_788861;
  wire [7:0] add_788864;
  wire [7:0] sel_788865;
  wire [7:0] add_788868;
  wire [7:0] sel_788869;
  wire [7:0] add_788872;
  wire [7:0] sel_788873;
  wire [7:0] add_788876;
  wire [7:0] sel_788877;
  wire [7:0] add_788880;
  wire [7:0] sel_788881;
  wire [7:0] add_788884;
  wire [7:0] sel_788885;
  wire [7:0] add_788888;
  wire [7:0] sel_788889;
  wire [7:0] add_788892;
  wire [7:0] sel_788893;
  wire [7:0] add_788896;
  wire [7:0] sel_788897;
  wire [7:0] add_788900;
  wire [7:0] sel_788901;
  wire [7:0] add_788904;
  wire [7:0] sel_788905;
  wire [7:0] add_788908;
  wire [7:0] sel_788909;
  wire [7:0] add_788912;
  wire [7:0] sel_788913;
  wire [7:0] add_788916;
  wire [7:0] sel_788917;
  wire [7:0] add_788920;
  wire [7:0] sel_788921;
  wire [7:0] add_788924;
  wire [7:0] sel_788925;
  wire [7:0] add_788928;
  wire [7:0] sel_788929;
  wire [7:0] add_788932;
  wire [7:0] sel_788933;
  wire [7:0] add_788936;
  wire [7:0] sel_788937;
  wire [7:0] add_788940;
  wire [7:0] sel_788941;
  wire [7:0] add_788944;
  wire [7:0] sel_788945;
  wire [7:0] add_788948;
  wire [7:0] sel_788949;
  wire [7:0] add_788952;
  wire [7:0] sel_788953;
  wire [7:0] add_788956;
  wire [7:0] sel_788957;
  wire [7:0] add_788960;
  wire [7:0] sel_788961;
  wire [7:0] add_788964;
  wire [7:0] sel_788965;
  wire [7:0] add_788968;
  wire [7:0] sel_788969;
  wire [7:0] add_788972;
  wire [7:0] sel_788973;
  wire [7:0] add_788976;
  wire [7:0] sel_788977;
  wire [7:0] add_788980;
  wire [7:0] sel_788981;
  wire [7:0] add_788984;
  wire [7:0] sel_788985;
  wire [7:0] add_788988;
  wire [7:0] sel_788989;
  wire [7:0] add_788992;
  wire [7:0] sel_788993;
  wire [7:0] add_788996;
  wire [7:0] sel_788997;
  wire [7:0] add_789000;
  wire [7:0] sel_789001;
  wire [7:0] add_789004;
  wire [7:0] sel_789005;
  wire [7:0] add_789008;
  wire [7:0] sel_789009;
  wire [7:0] add_789012;
  wire [7:0] sel_789013;
  wire [7:0] add_789016;
  wire [7:0] sel_789017;
  wire [7:0] add_789020;
  wire [7:0] sel_789021;
  wire [7:0] add_789024;
  wire [7:0] sel_789025;
  wire [7:0] add_789028;
  wire [7:0] sel_789029;
  wire [7:0] add_789032;
  wire [7:0] sel_789033;
  wire [7:0] add_789036;
  wire [7:0] sel_789037;
  wire [7:0] add_789040;
  wire [7:0] sel_789041;
  wire [7:0] add_789044;
  wire [7:0] sel_789045;
  wire [7:0] add_789048;
  wire [7:0] sel_789049;
  wire [7:0] add_789052;
  wire [7:0] sel_789053;
  wire [7:0] add_789056;
  wire [7:0] sel_789057;
  wire [7:0] add_789060;
  wire [7:0] sel_789061;
  wire [7:0] add_789064;
  wire [7:0] sel_789065;
  wire [7:0] add_789068;
  wire [7:0] sel_789069;
  wire [7:0] add_789072;
  wire [7:0] sel_789073;
  wire [7:0] add_789076;
  wire [7:0] sel_789077;
  wire [7:0] add_789080;
  wire [7:0] sel_789081;
  wire [7:0] add_789084;
  wire [7:0] sel_789085;
  wire [7:0] add_789088;
  wire [7:0] sel_789089;
  wire [7:0] add_789092;
  wire [7:0] sel_789093;
  wire [7:0] add_789096;
  wire [7:0] sel_789097;
  wire [7:0] add_789100;
  wire [7:0] sel_789101;
  wire [7:0] add_789104;
  wire [7:0] sel_789105;
  wire [7:0] add_789109;
  wire [15:0] array_index_789110;
  wire [7:0] sel_789111;
  wire [7:0] add_789114;
  wire [7:0] sel_789115;
  wire [7:0] add_789118;
  wire [7:0] sel_789119;
  wire [7:0] add_789122;
  wire [7:0] sel_789123;
  wire [7:0] add_789126;
  wire [7:0] sel_789127;
  wire [7:0] add_789130;
  wire [7:0] sel_789131;
  wire [7:0] add_789134;
  wire [7:0] sel_789135;
  wire [7:0] add_789138;
  wire [7:0] sel_789139;
  wire [7:0] add_789142;
  wire [7:0] sel_789143;
  wire [7:0] add_789146;
  wire [7:0] sel_789147;
  wire [7:0] add_789150;
  wire [7:0] sel_789151;
  wire [7:0] add_789154;
  wire [7:0] sel_789155;
  wire [7:0] add_789158;
  wire [7:0] sel_789159;
  wire [7:0] add_789162;
  wire [7:0] sel_789163;
  wire [7:0] add_789166;
  wire [7:0] sel_789167;
  wire [7:0] add_789170;
  wire [7:0] sel_789171;
  wire [7:0] add_789174;
  wire [7:0] sel_789175;
  wire [7:0] add_789178;
  wire [7:0] sel_789179;
  wire [7:0] add_789182;
  wire [7:0] sel_789183;
  wire [7:0] add_789186;
  wire [7:0] sel_789187;
  wire [7:0] add_789190;
  wire [7:0] sel_789191;
  wire [7:0] add_789194;
  wire [7:0] sel_789195;
  wire [7:0] add_789198;
  wire [7:0] sel_789199;
  wire [7:0] add_789202;
  wire [7:0] sel_789203;
  wire [7:0] add_789206;
  wire [7:0] sel_789207;
  wire [7:0] add_789210;
  wire [7:0] sel_789211;
  wire [7:0] add_789214;
  wire [7:0] sel_789215;
  wire [7:0] add_789218;
  wire [7:0] sel_789219;
  wire [7:0] add_789222;
  wire [7:0] sel_789223;
  wire [7:0] add_789226;
  wire [7:0] sel_789227;
  wire [7:0] add_789230;
  wire [7:0] sel_789231;
  wire [7:0] add_789234;
  wire [7:0] sel_789235;
  wire [7:0] add_789238;
  wire [7:0] sel_789239;
  wire [7:0] add_789242;
  wire [7:0] sel_789243;
  wire [7:0] add_789246;
  wire [7:0] sel_789247;
  wire [7:0] add_789250;
  wire [7:0] sel_789251;
  wire [7:0] add_789254;
  wire [7:0] sel_789255;
  wire [7:0] add_789258;
  wire [7:0] sel_789259;
  wire [7:0] add_789262;
  wire [7:0] sel_789263;
  wire [7:0] add_789266;
  wire [7:0] sel_789267;
  wire [7:0] add_789270;
  wire [7:0] sel_789271;
  wire [7:0] add_789274;
  wire [7:0] sel_789275;
  wire [7:0] add_789278;
  wire [7:0] sel_789279;
  wire [7:0] add_789282;
  wire [7:0] sel_789283;
  wire [7:0] add_789286;
  wire [7:0] sel_789287;
  wire [7:0] add_789290;
  wire [7:0] sel_789291;
  wire [7:0] add_789294;
  wire [7:0] sel_789295;
  wire [7:0] add_789298;
  wire [7:0] sel_789299;
  wire [7:0] add_789302;
  wire [7:0] sel_789303;
  wire [7:0] add_789306;
  wire [7:0] sel_789307;
  wire [7:0] add_789310;
  wire [7:0] sel_789311;
  wire [7:0] add_789314;
  wire [7:0] sel_789315;
  wire [7:0] add_789318;
  wire [7:0] sel_789319;
  wire [7:0] add_789322;
  wire [7:0] sel_789323;
  wire [7:0] add_789326;
  wire [7:0] sel_789327;
  wire [7:0] add_789330;
  wire [7:0] sel_789331;
  wire [7:0] add_789334;
  wire [7:0] sel_789335;
  wire [7:0] add_789338;
  wire [7:0] sel_789339;
  wire [7:0] add_789342;
  wire [7:0] sel_789343;
  wire [7:0] add_789346;
  wire [7:0] sel_789347;
  wire [7:0] add_789350;
  wire [7:0] sel_789351;
  wire [7:0] add_789354;
  wire [7:0] sel_789355;
  wire [7:0] add_789358;
  wire [7:0] sel_789359;
  wire [7:0] add_789362;
  wire [7:0] sel_789363;
  wire [7:0] add_789366;
  wire [7:0] sel_789367;
  wire [7:0] add_789370;
  wire [7:0] sel_789371;
  wire [7:0] add_789374;
  wire [7:0] sel_789375;
  wire [7:0] add_789378;
  wire [7:0] sel_789379;
  wire [7:0] add_789382;
  wire [7:0] sel_789383;
  wire [7:0] add_789386;
  wire [7:0] sel_789387;
  wire [7:0] add_789390;
  wire [7:0] sel_789391;
  wire [7:0] add_789394;
  wire [7:0] sel_789395;
  wire [7:0] add_789398;
  wire [7:0] sel_789399;
  wire [7:0] add_789402;
  wire [7:0] sel_789403;
  wire [7:0] add_789406;
  wire [7:0] sel_789407;
  wire [7:0] add_789410;
  wire [7:0] sel_789411;
  wire [7:0] add_789414;
  wire [7:0] sel_789415;
  wire [7:0] add_789418;
  wire [7:0] sel_789419;
  wire [7:0] add_789422;
  wire [7:0] sel_789423;
  wire [7:0] add_789426;
  wire [7:0] sel_789427;
  wire [7:0] add_789430;
  wire [7:0] sel_789431;
  wire [7:0] add_789434;
  wire [7:0] sel_789435;
  wire [7:0] add_789438;
  wire [7:0] sel_789439;
  wire [7:0] add_789442;
  wire [7:0] sel_789443;
  wire [7:0] add_789446;
  wire [7:0] sel_789447;
  wire [7:0] add_789450;
  wire [7:0] sel_789451;
  wire [7:0] add_789454;
  wire [7:0] sel_789455;
  wire [7:0] add_789458;
  wire [7:0] sel_789459;
  wire [7:0] add_789462;
  wire [7:0] sel_789463;
  wire [7:0] add_789466;
  wire [7:0] sel_789467;
  wire [7:0] add_789471;
  wire [15:0] array_index_789472;
  wire [7:0] sel_789473;
  wire [7:0] add_789476;
  wire [7:0] sel_789477;
  wire [7:0] add_789480;
  wire [7:0] sel_789481;
  wire [7:0] add_789484;
  wire [7:0] sel_789485;
  wire [7:0] add_789488;
  wire [7:0] sel_789489;
  wire [7:0] add_789492;
  wire [7:0] sel_789493;
  wire [7:0] add_789496;
  wire [7:0] sel_789497;
  wire [7:0] add_789500;
  wire [7:0] sel_789501;
  wire [7:0] add_789504;
  wire [7:0] sel_789505;
  wire [7:0] add_789508;
  wire [7:0] sel_789509;
  wire [7:0] add_789512;
  wire [7:0] sel_789513;
  wire [7:0] add_789516;
  wire [7:0] sel_789517;
  wire [7:0] add_789520;
  wire [7:0] sel_789521;
  wire [7:0] add_789524;
  wire [7:0] sel_789525;
  wire [7:0] add_789528;
  wire [7:0] sel_789529;
  wire [7:0] add_789532;
  wire [7:0] sel_789533;
  wire [7:0] add_789536;
  wire [7:0] sel_789537;
  wire [7:0] add_789540;
  wire [7:0] sel_789541;
  wire [7:0] add_789544;
  wire [7:0] sel_789545;
  wire [7:0] add_789548;
  wire [7:0] sel_789549;
  wire [7:0] add_789552;
  wire [7:0] sel_789553;
  wire [7:0] add_789556;
  wire [7:0] sel_789557;
  wire [7:0] add_789560;
  wire [7:0] sel_789561;
  wire [7:0] add_789564;
  wire [7:0] sel_789565;
  wire [7:0] add_789568;
  wire [7:0] sel_789569;
  wire [7:0] add_789572;
  wire [7:0] sel_789573;
  wire [7:0] add_789576;
  wire [7:0] sel_789577;
  wire [7:0] add_789580;
  wire [7:0] sel_789581;
  wire [7:0] add_789584;
  wire [7:0] sel_789585;
  wire [7:0] add_789588;
  wire [7:0] sel_789589;
  wire [7:0] add_789592;
  wire [7:0] sel_789593;
  wire [7:0] add_789596;
  wire [7:0] sel_789597;
  wire [7:0] add_789600;
  wire [7:0] sel_789601;
  wire [7:0] add_789604;
  wire [7:0] sel_789605;
  wire [7:0] add_789608;
  wire [7:0] sel_789609;
  wire [7:0] add_789612;
  wire [7:0] sel_789613;
  wire [7:0] add_789616;
  wire [7:0] sel_789617;
  wire [7:0] add_789620;
  wire [7:0] sel_789621;
  wire [7:0] add_789624;
  wire [7:0] sel_789625;
  wire [7:0] add_789628;
  wire [7:0] sel_789629;
  wire [7:0] add_789632;
  wire [7:0] sel_789633;
  wire [7:0] add_789636;
  wire [7:0] sel_789637;
  wire [7:0] add_789640;
  wire [7:0] sel_789641;
  wire [7:0] add_789644;
  wire [7:0] sel_789645;
  wire [7:0] add_789648;
  wire [7:0] sel_789649;
  wire [7:0] add_789652;
  wire [7:0] sel_789653;
  wire [7:0] add_789656;
  wire [7:0] sel_789657;
  wire [7:0] add_789660;
  wire [7:0] sel_789661;
  wire [7:0] add_789664;
  wire [7:0] sel_789665;
  wire [7:0] add_789668;
  wire [7:0] sel_789669;
  wire [7:0] add_789672;
  wire [7:0] sel_789673;
  wire [7:0] add_789676;
  wire [7:0] sel_789677;
  wire [7:0] add_789680;
  wire [7:0] sel_789681;
  wire [7:0] add_789684;
  wire [7:0] sel_789685;
  wire [7:0] add_789688;
  wire [7:0] sel_789689;
  wire [7:0] add_789692;
  wire [7:0] sel_789693;
  wire [7:0] add_789696;
  wire [7:0] sel_789697;
  wire [7:0] add_789700;
  wire [7:0] sel_789701;
  wire [7:0] add_789704;
  wire [7:0] sel_789705;
  wire [7:0] add_789708;
  wire [7:0] sel_789709;
  wire [7:0] add_789712;
  wire [7:0] sel_789713;
  wire [7:0] add_789716;
  wire [7:0] sel_789717;
  wire [7:0] add_789720;
  wire [7:0] sel_789721;
  wire [7:0] add_789724;
  wire [7:0] sel_789725;
  wire [7:0] add_789728;
  wire [7:0] sel_789729;
  wire [7:0] add_789732;
  wire [7:0] sel_789733;
  wire [7:0] add_789736;
  wire [7:0] sel_789737;
  wire [7:0] add_789740;
  wire [7:0] sel_789741;
  wire [7:0] add_789744;
  wire [7:0] sel_789745;
  wire [7:0] add_789748;
  wire [7:0] sel_789749;
  wire [7:0] add_789752;
  wire [7:0] sel_789753;
  wire [7:0] add_789756;
  wire [7:0] sel_789757;
  wire [7:0] add_789760;
  wire [7:0] sel_789761;
  wire [7:0] add_789764;
  wire [7:0] sel_789765;
  wire [7:0] add_789768;
  wire [7:0] sel_789769;
  wire [7:0] add_789772;
  wire [7:0] sel_789773;
  wire [7:0] add_789776;
  wire [7:0] sel_789777;
  wire [7:0] add_789780;
  wire [7:0] sel_789781;
  wire [7:0] add_789784;
  wire [7:0] sel_789785;
  wire [7:0] add_789788;
  wire [7:0] sel_789789;
  wire [7:0] add_789792;
  wire [7:0] sel_789793;
  wire [7:0] add_789796;
  wire [7:0] sel_789797;
  wire [7:0] add_789800;
  wire [7:0] sel_789801;
  wire [7:0] add_789804;
  wire [7:0] sel_789805;
  wire [7:0] add_789808;
  wire [7:0] sel_789809;
  wire [7:0] add_789812;
  wire [7:0] sel_789813;
  wire [7:0] add_789816;
  wire [7:0] sel_789817;
  wire [7:0] add_789820;
  wire [7:0] sel_789821;
  wire [7:0] add_789824;
  wire [7:0] sel_789825;
  wire [7:0] add_789828;
  wire [7:0] sel_789829;
  wire [7:0] add_789833;
  wire [15:0] array_index_789834;
  wire [7:0] sel_789835;
  wire [7:0] add_789838;
  wire [7:0] sel_789839;
  wire [7:0] add_789842;
  wire [7:0] sel_789843;
  wire [7:0] add_789846;
  wire [7:0] sel_789847;
  wire [7:0] add_789850;
  wire [7:0] sel_789851;
  wire [7:0] add_789854;
  wire [7:0] sel_789855;
  wire [7:0] add_789858;
  wire [7:0] sel_789859;
  wire [7:0] add_789862;
  wire [7:0] sel_789863;
  wire [7:0] add_789866;
  wire [7:0] sel_789867;
  wire [7:0] add_789870;
  wire [7:0] sel_789871;
  wire [7:0] add_789874;
  wire [7:0] sel_789875;
  wire [7:0] add_789878;
  wire [7:0] sel_789879;
  wire [7:0] add_789882;
  wire [7:0] sel_789883;
  wire [7:0] add_789886;
  wire [7:0] sel_789887;
  wire [7:0] add_789890;
  wire [7:0] sel_789891;
  wire [7:0] add_789894;
  wire [7:0] sel_789895;
  wire [7:0] add_789898;
  wire [7:0] sel_789899;
  wire [7:0] add_789902;
  wire [7:0] sel_789903;
  wire [7:0] add_789906;
  wire [7:0] sel_789907;
  wire [7:0] add_789910;
  wire [7:0] sel_789911;
  wire [7:0] add_789914;
  wire [7:0] sel_789915;
  wire [7:0] add_789918;
  wire [7:0] sel_789919;
  wire [7:0] add_789922;
  wire [7:0] sel_789923;
  wire [7:0] add_789926;
  wire [7:0] sel_789927;
  wire [7:0] add_789930;
  wire [7:0] sel_789931;
  wire [7:0] add_789934;
  wire [7:0] sel_789935;
  wire [7:0] add_789938;
  wire [7:0] sel_789939;
  wire [7:0] add_789942;
  wire [7:0] sel_789943;
  wire [7:0] add_789946;
  wire [7:0] sel_789947;
  wire [7:0] add_789950;
  wire [7:0] sel_789951;
  wire [7:0] add_789954;
  wire [7:0] sel_789955;
  wire [7:0] add_789958;
  wire [7:0] sel_789959;
  wire [7:0] add_789962;
  wire [7:0] sel_789963;
  wire [7:0] add_789966;
  wire [7:0] sel_789967;
  wire [7:0] add_789970;
  wire [7:0] sel_789971;
  wire [7:0] add_789974;
  wire [7:0] sel_789975;
  wire [7:0] add_789978;
  wire [7:0] sel_789979;
  wire [7:0] add_789982;
  wire [7:0] sel_789983;
  wire [7:0] add_789986;
  wire [7:0] sel_789987;
  wire [7:0] add_789990;
  wire [7:0] sel_789991;
  wire [7:0] add_789994;
  wire [7:0] sel_789995;
  wire [7:0] add_789998;
  wire [7:0] sel_789999;
  wire [7:0] add_790002;
  wire [7:0] sel_790003;
  wire [7:0] add_790006;
  wire [7:0] sel_790007;
  wire [7:0] add_790010;
  wire [7:0] sel_790011;
  wire [7:0] add_790014;
  wire [7:0] sel_790015;
  wire [7:0] add_790018;
  wire [7:0] sel_790019;
  wire [7:0] add_790022;
  wire [7:0] sel_790023;
  wire [7:0] add_790026;
  wire [7:0] sel_790027;
  wire [7:0] add_790030;
  wire [7:0] sel_790031;
  wire [7:0] add_790034;
  wire [7:0] sel_790035;
  wire [7:0] add_790038;
  wire [7:0] sel_790039;
  wire [7:0] add_790042;
  wire [7:0] sel_790043;
  wire [7:0] add_790046;
  wire [7:0] sel_790047;
  wire [7:0] add_790050;
  wire [7:0] sel_790051;
  wire [7:0] add_790054;
  wire [7:0] sel_790055;
  wire [7:0] add_790058;
  wire [7:0] sel_790059;
  wire [7:0] add_790062;
  wire [7:0] sel_790063;
  wire [7:0] add_790066;
  wire [7:0] sel_790067;
  wire [7:0] add_790070;
  wire [7:0] sel_790071;
  wire [7:0] add_790074;
  wire [7:0] sel_790075;
  wire [7:0] add_790078;
  wire [7:0] sel_790079;
  wire [7:0] add_790082;
  wire [7:0] sel_790083;
  wire [7:0] add_790086;
  wire [7:0] sel_790087;
  wire [7:0] add_790090;
  wire [7:0] sel_790091;
  wire [7:0] add_790094;
  wire [7:0] sel_790095;
  wire [7:0] add_790098;
  wire [7:0] sel_790099;
  wire [7:0] add_790102;
  wire [7:0] sel_790103;
  wire [7:0] add_790106;
  wire [7:0] sel_790107;
  wire [7:0] add_790110;
  wire [7:0] sel_790111;
  wire [7:0] add_790114;
  wire [7:0] sel_790115;
  wire [7:0] add_790118;
  wire [7:0] sel_790119;
  wire [7:0] add_790122;
  wire [7:0] sel_790123;
  wire [7:0] add_790126;
  wire [7:0] sel_790127;
  wire [7:0] add_790130;
  wire [7:0] sel_790131;
  wire [7:0] add_790134;
  wire [7:0] sel_790135;
  wire [7:0] add_790138;
  wire [7:0] sel_790139;
  wire [7:0] add_790142;
  wire [7:0] sel_790143;
  wire [7:0] add_790146;
  wire [7:0] sel_790147;
  wire [7:0] add_790150;
  wire [7:0] sel_790151;
  wire [7:0] add_790154;
  wire [7:0] sel_790155;
  wire [7:0] add_790158;
  wire [7:0] sel_790159;
  wire [7:0] add_790162;
  wire [7:0] sel_790163;
  wire [7:0] add_790166;
  wire [7:0] sel_790167;
  wire [7:0] add_790170;
  wire [7:0] sel_790171;
  wire [7:0] add_790174;
  wire [7:0] sel_790175;
  wire [7:0] add_790178;
  wire [7:0] sel_790179;
  wire [7:0] add_790182;
  wire [7:0] sel_790183;
  wire [7:0] add_790186;
  wire [7:0] sel_790187;
  wire [7:0] add_790190;
  wire [7:0] sel_790191;
  wire [7:0] add_790195;
  wire [15:0] array_index_790196;
  wire [7:0] sel_790197;
  wire [7:0] add_790200;
  wire [7:0] sel_790201;
  wire [7:0] add_790204;
  wire [7:0] sel_790205;
  wire [7:0] add_790208;
  wire [7:0] sel_790209;
  wire [7:0] add_790212;
  wire [7:0] sel_790213;
  wire [7:0] add_790216;
  wire [7:0] sel_790217;
  wire [7:0] add_790220;
  wire [7:0] sel_790221;
  wire [7:0] add_790224;
  wire [7:0] sel_790225;
  wire [7:0] add_790228;
  wire [7:0] sel_790229;
  wire [7:0] add_790232;
  wire [7:0] sel_790233;
  wire [7:0] add_790236;
  wire [7:0] sel_790237;
  wire [7:0] add_790240;
  wire [7:0] sel_790241;
  wire [7:0] add_790244;
  wire [7:0] sel_790245;
  wire [7:0] add_790248;
  wire [7:0] sel_790249;
  wire [7:0] add_790252;
  wire [7:0] sel_790253;
  wire [7:0] add_790256;
  wire [7:0] sel_790257;
  wire [7:0] add_790260;
  wire [7:0] sel_790261;
  wire [7:0] add_790264;
  wire [7:0] sel_790265;
  wire [7:0] add_790268;
  wire [7:0] sel_790269;
  wire [7:0] add_790272;
  wire [7:0] sel_790273;
  wire [7:0] add_790276;
  wire [7:0] sel_790277;
  wire [7:0] add_790280;
  wire [7:0] sel_790281;
  wire [7:0] add_790284;
  wire [7:0] sel_790285;
  wire [7:0] add_790288;
  wire [7:0] sel_790289;
  wire [7:0] add_790292;
  wire [7:0] sel_790293;
  wire [7:0] add_790296;
  wire [7:0] sel_790297;
  wire [7:0] add_790300;
  wire [7:0] sel_790301;
  wire [7:0] add_790304;
  wire [7:0] sel_790305;
  wire [7:0] add_790308;
  wire [7:0] sel_790309;
  wire [7:0] add_790312;
  wire [7:0] sel_790313;
  wire [7:0] add_790316;
  wire [7:0] sel_790317;
  wire [7:0] add_790320;
  wire [7:0] sel_790321;
  wire [7:0] add_790324;
  wire [7:0] sel_790325;
  wire [7:0] add_790328;
  wire [7:0] sel_790329;
  wire [7:0] add_790332;
  wire [7:0] sel_790333;
  wire [7:0] add_790336;
  wire [7:0] sel_790337;
  wire [7:0] add_790340;
  wire [7:0] sel_790341;
  wire [7:0] add_790344;
  wire [7:0] sel_790345;
  wire [7:0] add_790348;
  wire [7:0] sel_790349;
  wire [7:0] add_790352;
  wire [7:0] sel_790353;
  wire [7:0] add_790356;
  wire [7:0] sel_790357;
  wire [7:0] add_790360;
  wire [7:0] sel_790361;
  wire [7:0] add_790364;
  wire [7:0] sel_790365;
  wire [7:0] add_790368;
  wire [7:0] sel_790369;
  wire [7:0] add_790372;
  wire [7:0] sel_790373;
  wire [7:0] add_790376;
  wire [7:0] sel_790377;
  wire [7:0] add_790380;
  wire [7:0] sel_790381;
  wire [7:0] add_790384;
  wire [7:0] sel_790385;
  wire [7:0] add_790388;
  wire [7:0] sel_790389;
  wire [7:0] add_790392;
  wire [7:0] sel_790393;
  wire [7:0] add_790396;
  wire [7:0] sel_790397;
  wire [7:0] add_790400;
  wire [7:0] sel_790401;
  wire [7:0] add_790404;
  wire [7:0] sel_790405;
  wire [7:0] add_790408;
  wire [7:0] sel_790409;
  wire [7:0] add_790412;
  wire [7:0] sel_790413;
  wire [7:0] add_790416;
  wire [7:0] sel_790417;
  wire [7:0] add_790420;
  wire [7:0] sel_790421;
  wire [7:0] add_790424;
  wire [7:0] sel_790425;
  wire [7:0] add_790428;
  wire [7:0] sel_790429;
  wire [7:0] add_790432;
  wire [7:0] sel_790433;
  wire [7:0] add_790436;
  wire [7:0] sel_790437;
  wire [7:0] add_790440;
  wire [7:0] sel_790441;
  wire [7:0] add_790444;
  wire [7:0] sel_790445;
  wire [7:0] add_790448;
  wire [7:0] sel_790449;
  wire [7:0] add_790452;
  wire [7:0] sel_790453;
  wire [7:0] add_790456;
  wire [7:0] sel_790457;
  wire [7:0] add_790460;
  wire [7:0] sel_790461;
  wire [7:0] add_790464;
  wire [7:0] sel_790465;
  wire [7:0] add_790468;
  wire [7:0] sel_790469;
  wire [7:0] add_790472;
  wire [7:0] sel_790473;
  wire [7:0] add_790476;
  wire [7:0] sel_790477;
  wire [7:0] add_790480;
  wire [7:0] sel_790481;
  wire [7:0] add_790484;
  wire [7:0] sel_790485;
  wire [7:0] add_790488;
  wire [7:0] sel_790489;
  wire [7:0] add_790492;
  wire [7:0] sel_790493;
  wire [7:0] add_790496;
  wire [7:0] sel_790497;
  wire [7:0] add_790500;
  wire [7:0] sel_790501;
  wire [7:0] add_790504;
  wire [7:0] sel_790505;
  wire [7:0] add_790508;
  wire [7:0] sel_790509;
  wire [7:0] add_790512;
  wire [7:0] sel_790513;
  wire [7:0] add_790516;
  wire [7:0] sel_790517;
  wire [7:0] add_790520;
  wire [7:0] sel_790521;
  wire [7:0] add_790524;
  wire [7:0] sel_790525;
  wire [7:0] add_790528;
  wire [7:0] sel_790529;
  wire [7:0] add_790532;
  wire [7:0] sel_790533;
  wire [7:0] add_790536;
  wire [7:0] sel_790537;
  wire [7:0] add_790540;
  wire [7:0] sel_790541;
  wire [7:0] add_790544;
  wire [7:0] sel_790545;
  wire [7:0] add_790548;
  wire [7:0] sel_790549;
  wire [7:0] add_790552;
  wire [7:0] sel_790553;
  wire [7:0] add_790557;
  wire [15:0] array_index_790558;
  wire [7:0] sel_790559;
  wire [7:0] add_790562;
  wire [7:0] sel_790563;
  wire [7:0] add_790566;
  wire [7:0] sel_790567;
  wire [7:0] add_790570;
  wire [7:0] sel_790571;
  wire [7:0] add_790574;
  wire [7:0] sel_790575;
  wire [7:0] add_790578;
  wire [7:0] sel_790579;
  wire [7:0] add_790582;
  wire [7:0] sel_790583;
  wire [7:0] add_790586;
  wire [7:0] sel_790587;
  wire [7:0] add_790590;
  wire [7:0] sel_790591;
  wire [7:0] add_790594;
  wire [7:0] sel_790595;
  wire [7:0] add_790598;
  wire [7:0] sel_790599;
  wire [7:0] add_790602;
  wire [7:0] sel_790603;
  wire [7:0] add_790606;
  wire [7:0] sel_790607;
  wire [7:0] add_790610;
  wire [7:0] sel_790611;
  wire [7:0] add_790614;
  wire [7:0] sel_790615;
  wire [7:0] add_790618;
  wire [7:0] sel_790619;
  wire [7:0] add_790622;
  wire [7:0] sel_790623;
  wire [7:0] add_790626;
  wire [7:0] sel_790627;
  wire [7:0] add_790630;
  wire [7:0] sel_790631;
  wire [7:0] add_790634;
  wire [7:0] sel_790635;
  wire [7:0] add_790638;
  wire [7:0] sel_790639;
  wire [7:0] add_790642;
  wire [7:0] sel_790643;
  wire [7:0] add_790646;
  wire [7:0] sel_790647;
  wire [7:0] add_790650;
  wire [7:0] sel_790651;
  wire [7:0] add_790654;
  wire [7:0] sel_790655;
  wire [7:0] add_790658;
  wire [7:0] sel_790659;
  wire [7:0] add_790662;
  wire [7:0] sel_790663;
  wire [7:0] add_790666;
  wire [7:0] sel_790667;
  wire [7:0] add_790670;
  wire [7:0] sel_790671;
  wire [7:0] add_790674;
  wire [7:0] sel_790675;
  wire [7:0] add_790678;
  wire [7:0] sel_790679;
  wire [7:0] add_790682;
  wire [7:0] sel_790683;
  wire [7:0] add_790686;
  wire [7:0] sel_790687;
  wire [7:0] add_790690;
  wire [7:0] sel_790691;
  wire [7:0] add_790694;
  wire [7:0] sel_790695;
  wire [7:0] add_790698;
  wire [7:0] sel_790699;
  wire [7:0] add_790702;
  wire [7:0] sel_790703;
  wire [7:0] add_790706;
  wire [7:0] sel_790707;
  wire [7:0] add_790710;
  wire [7:0] sel_790711;
  wire [7:0] add_790714;
  wire [7:0] sel_790715;
  wire [7:0] add_790718;
  wire [7:0] sel_790719;
  wire [7:0] add_790722;
  wire [7:0] sel_790723;
  wire [7:0] add_790726;
  wire [7:0] sel_790727;
  wire [7:0] add_790730;
  wire [7:0] sel_790731;
  wire [7:0] add_790734;
  wire [7:0] sel_790735;
  wire [7:0] add_790738;
  wire [7:0] sel_790739;
  wire [7:0] add_790742;
  wire [7:0] sel_790743;
  wire [7:0] add_790746;
  wire [7:0] sel_790747;
  wire [7:0] add_790750;
  wire [7:0] sel_790751;
  wire [7:0] add_790754;
  wire [7:0] sel_790755;
  wire [7:0] add_790758;
  wire [7:0] sel_790759;
  wire [7:0] add_790762;
  wire [7:0] sel_790763;
  wire [7:0] add_790766;
  wire [7:0] sel_790767;
  wire [7:0] add_790770;
  wire [7:0] sel_790771;
  wire [7:0] add_790774;
  wire [7:0] sel_790775;
  wire [7:0] add_790778;
  wire [7:0] sel_790779;
  wire [7:0] add_790782;
  wire [7:0] sel_790783;
  wire [7:0] add_790786;
  wire [7:0] sel_790787;
  wire [7:0] add_790790;
  wire [7:0] sel_790791;
  wire [7:0] add_790794;
  wire [7:0] sel_790795;
  wire [7:0] add_790798;
  wire [7:0] sel_790799;
  wire [7:0] add_790802;
  wire [7:0] sel_790803;
  wire [7:0] add_790806;
  wire [7:0] sel_790807;
  wire [7:0] add_790810;
  wire [7:0] sel_790811;
  wire [7:0] add_790814;
  wire [7:0] sel_790815;
  wire [7:0] add_790818;
  wire [7:0] sel_790819;
  wire [7:0] add_790822;
  wire [7:0] sel_790823;
  wire [7:0] add_790826;
  wire [7:0] sel_790827;
  wire [7:0] add_790830;
  wire [7:0] sel_790831;
  wire [7:0] add_790834;
  wire [7:0] sel_790835;
  wire [7:0] add_790838;
  wire [7:0] sel_790839;
  wire [7:0] add_790842;
  wire [7:0] sel_790843;
  wire [7:0] add_790846;
  wire [7:0] sel_790847;
  wire [7:0] add_790850;
  wire [7:0] sel_790851;
  wire [7:0] add_790854;
  wire [7:0] sel_790855;
  wire [7:0] add_790858;
  wire [7:0] sel_790859;
  wire [7:0] add_790862;
  wire [7:0] sel_790863;
  wire [7:0] add_790866;
  wire [7:0] sel_790867;
  wire [7:0] add_790870;
  wire [7:0] sel_790871;
  wire [7:0] add_790874;
  wire [7:0] sel_790875;
  wire [7:0] add_790878;
  wire [7:0] sel_790879;
  wire [7:0] add_790882;
  wire [7:0] sel_790883;
  wire [7:0] add_790886;
  wire [7:0] sel_790887;
  wire [7:0] add_790890;
  wire [7:0] sel_790891;
  wire [7:0] add_790894;
  wire [7:0] sel_790895;
  wire [7:0] add_790898;
  wire [7:0] sel_790899;
  wire [7:0] add_790902;
  wire [7:0] sel_790903;
  wire [7:0] add_790906;
  wire [7:0] sel_790907;
  wire [7:0] add_790910;
  wire [7:0] sel_790911;
  wire [7:0] add_790914;
  wire [7:0] sel_790915;
  wire [7:0] add_790919;
  wire [15:0] array_index_790920;
  wire [7:0] sel_790921;
  wire [7:0] add_790924;
  wire [7:0] sel_790925;
  wire [7:0] add_790928;
  wire [7:0] sel_790929;
  wire [7:0] add_790932;
  wire [7:0] sel_790933;
  wire [7:0] add_790936;
  wire [7:0] sel_790937;
  wire [7:0] add_790940;
  wire [7:0] sel_790941;
  wire [7:0] add_790944;
  wire [7:0] sel_790945;
  wire [7:0] add_790948;
  wire [7:0] sel_790949;
  wire [7:0] add_790952;
  wire [7:0] sel_790953;
  wire [7:0] add_790956;
  wire [7:0] sel_790957;
  wire [7:0] add_790960;
  wire [7:0] sel_790961;
  wire [7:0] add_790964;
  wire [7:0] sel_790965;
  wire [7:0] add_790968;
  wire [7:0] sel_790969;
  wire [7:0] add_790972;
  wire [7:0] sel_790973;
  wire [7:0] add_790976;
  wire [7:0] sel_790977;
  wire [7:0] add_790980;
  wire [7:0] sel_790981;
  wire [7:0] add_790984;
  wire [7:0] sel_790985;
  wire [7:0] add_790988;
  wire [7:0] sel_790989;
  wire [7:0] add_790992;
  wire [7:0] sel_790993;
  wire [7:0] add_790996;
  wire [7:0] sel_790997;
  wire [7:0] add_791000;
  wire [7:0] sel_791001;
  wire [7:0] add_791004;
  wire [7:0] sel_791005;
  wire [7:0] add_791008;
  wire [7:0] sel_791009;
  wire [7:0] add_791012;
  wire [7:0] sel_791013;
  wire [7:0] add_791016;
  wire [7:0] sel_791017;
  wire [7:0] add_791020;
  wire [7:0] sel_791021;
  wire [7:0] add_791024;
  wire [7:0] sel_791025;
  wire [7:0] add_791028;
  wire [7:0] sel_791029;
  wire [7:0] add_791032;
  wire [7:0] sel_791033;
  wire [7:0] add_791036;
  wire [7:0] sel_791037;
  wire [7:0] add_791040;
  wire [7:0] sel_791041;
  wire [7:0] add_791044;
  wire [7:0] sel_791045;
  wire [7:0] add_791048;
  wire [7:0] sel_791049;
  wire [7:0] add_791052;
  wire [7:0] sel_791053;
  wire [7:0] add_791056;
  wire [7:0] sel_791057;
  wire [7:0] add_791060;
  wire [7:0] sel_791061;
  wire [7:0] add_791064;
  wire [7:0] sel_791065;
  wire [7:0] add_791068;
  wire [7:0] sel_791069;
  wire [7:0] add_791072;
  wire [7:0] sel_791073;
  wire [7:0] add_791076;
  wire [7:0] sel_791077;
  wire [7:0] add_791080;
  wire [7:0] sel_791081;
  wire [7:0] add_791084;
  wire [7:0] sel_791085;
  wire [7:0] add_791088;
  wire [7:0] sel_791089;
  wire [7:0] add_791092;
  wire [7:0] sel_791093;
  wire [7:0] add_791096;
  wire [7:0] sel_791097;
  wire [7:0] add_791100;
  wire [7:0] sel_791101;
  wire [7:0] add_791104;
  wire [7:0] sel_791105;
  wire [7:0] add_791108;
  wire [7:0] sel_791109;
  wire [7:0] add_791112;
  wire [7:0] sel_791113;
  wire [7:0] add_791116;
  wire [7:0] sel_791117;
  wire [7:0] add_791120;
  wire [7:0] sel_791121;
  wire [7:0] add_791124;
  wire [7:0] sel_791125;
  wire [7:0] add_791128;
  wire [7:0] sel_791129;
  wire [7:0] add_791132;
  wire [7:0] sel_791133;
  wire [7:0] add_791136;
  wire [7:0] sel_791137;
  wire [7:0] add_791140;
  wire [7:0] sel_791141;
  wire [7:0] add_791144;
  wire [7:0] sel_791145;
  wire [7:0] add_791148;
  wire [7:0] sel_791149;
  wire [7:0] add_791152;
  wire [7:0] sel_791153;
  wire [7:0] add_791156;
  wire [7:0] sel_791157;
  wire [7:0] add_791160;
  wire [7:0] sel_791161;
  wire [7:0] add_791164;
  wire [7:0] sel_791165;
  wire [7:0] add_791168;
  wire [7:0] sel_791169;
  wire [7:0] add_791172;
  wire [7:0] sel_791173;
  wire [7:0] add_791176;
  wire [7:0] sel_791177;
  wire [7:0] add_791180;
  wire [7:0] sel_791181;
  wire [7:0] add_791184;
  wire [7:0] sel_791185;
  wire [7:0] add_791188;
  wire [7:0] sel_791189;
  wire [7:0] add_791192;
  wire [7:0] sel_791193;
  wire [7:0] add_791196;
  wire [7:0] sel_791197;
  wire [7:0] add_791200;
  wire [7:0] sel_791201;
  wire [7:0] add_791204;
  wire [7:0] sel_791205;
  wire [7:0] add_791208;
  wire [7:0] sel_791209;
  wire [7:0] add_791212;
  wire [7:0] sel_791213;
  wire [7:0] add_791216;
  wire [7:0] sel_791217;
  wire [7:0] add_791220;
  wire [7:0] sel_791221;
  wire [7:0] add_791224;
  wire [7:0] sel_791225;
  wire [7:0] add_791228;
  wire [7:0] sel_791229;
  wire [7:0] add_791232;
  wire [7:0] sel_791233;
  wire [7:0] add_791236;
  wire [7:0] sel_791237;
  wire [7:0] add_791240;
  wire [7:0] sel_791241;
  wire [7:0] add_791244;
  wire [7:0] sel_791245;
  wire [7:0] add_791248;
  wire [7:0] sel_791249;
  wire [7:0] add_791252;
  wire [7:0] sel_791253;
  wire [7:0] add_791256;
  wire [7:0] sel_791257;
  wire [7:0] add_791260;
  wire [7:0] sel_791261;
  wire [7:0] add_791264;
  wire [7:0] sel_791265;
  wire [7:0] add_791268;
  wire [7:0] sel_791269;
  wire [7:0] add_791272;
  wire [7:0] sel_791273;
  wire [7:0] add_791276;
  wire [7:0] sel_791277;
  wire [7:0] add_791281;
  wire [15:0] array_index_791282;
  wire [7:0] sel_791283;
  wire [7:0] add_791286;
  wire [7:0] sel_791287;
  wire [7:0] add_791290;
  wire [7:0] sel_791291;
  wire [7:0] add_791294;
  wire [7:0] sel_791295;
  wire [7:0] add_791298;
  wire [7:0] sel_791299;
  wire [7:0] add_791302;
  wire [7:0] sel_791303;
  wire [7:0] add_791306;
  wire [7:0] sel_791307;
  wire [7:0] add_791310;
  wire [7:0] sel_791311;
  wire [7:0] add_791314;
  wire [7:0] sel_791315;
  wire [7:0] add_791318;
  wire [7:0] sel_791319;
  wire [7:0] add_791322;
  wire [7:0] sel_791323;
  wire [7:0] add_791326;
  wire [7:0] sel_791327;
  wire [7:0] add_791330;
  wire [7:0] sel_791331;
  wire [7:0] add_791334;
  wire [7:0] sel_791335;
  wire [7:0] add_791338;
  wire [7:0] sel_791339;
  wire [7:0] add_791342;
  wire [7:0] sel_791343;
  wire [7:0] add_791346;
  wire [7:0] sel_791347;
  wire [7:0] add_791350;
  wire [7:0] sel_791351;
  wire [7:0] add_791354;
  wire [7:0] sel_791355;
  wire [7:0] add_791358;
  wire [7:0] sel_791359;
  wire [7:0] add_791362;
  wire [7:0] sel_791363;
  wire [7:0] add_791366;
  wire [7:0] sel_791367;
  wire [7:0] add_791370;
  wire [7:0] sel_791371;
  wire [7:0] add_791374;
  wire [7:0] sel_791375;
  wire [7:0] add_791378;
  wire [7:0] sel_791379;
  wire [7:0] add_791382;
  wire [7:0] sel_791383;
  wire [7:0] add_791386;
  wire [7:0] sel_791387;
  wire [7:0] add_791390;
  wire [7:0] sel_791391;
  wire [7:0] add_791394;
  wire [7:0] sel_791395;
  wire [7:0] add_791398;
  wire [7:0] sel_791399;
  wire [7:0] add_791402;
  wire [7:0] sel_791403;
  wire [7:0] add_791406;
  wire [7:0] sel_791407;
  wire [7:0] add_791410;
  wire [7:0] sel_791411;
  wire [7:0] add_791414;
  wire [7:0] sel_791415;
  wire [7:0] add_791418;
  wire [7:0] sel_791419;
  wire [7:0] add_791422;
  wire [7:0] sel_791423;
  wire [7:0] add_791426;
  wire [7:0] sel_791427;
  wire [7:0] add_791430;
  wire [7:0] sel_791431;
  wire [7:0] add_791434;
  wire [7:0] sel_791435;
  wire [7:0] add_791438;
  wire [7:0] sel_791439;
  wire [7:0] add_791442;
  wire [7:0] sel_791443;
  wire [7:0] add_791446;
  wire [7:0] sel_791447;
  wire [7:0] add_791450;
  wire [7:0] sel_791451;
  wire [7:0] add_791454;
  wire [7:0] sel_791455;
  wire [7:0] add_791458;
  wire [7:0] sel_791459;
  wire [7:0] add_791462;
  wire [7:0] sel_791463;
  wire [7:0] add_791466;
  wire [7:0] sel_791467;
  wire [7:0] add_791470;
  wire [7:0] sel_791471;
  wire [7:0] add_791474;
  wire [7:0] sel_791475;
  wire [7:0] add_791478;
  wire [7:0] sel_791479;
  wire [7:0] add_791482;
  wire [7:0] sel_791483;
  wire [7:0] add_791486;
  wire [7:0] sel_791487;
  wire [7:0] add_791490;
  wire [7:0] sel_791491;
  wire [7:0] add_791494;
  wire [7:0] sel_791495;
  wire [7:0] add_791498;
  wire [7:0] sel_791499;
  wire [7:0] add_791502;
  wire [7:0] sel_791503;
  wire [7:0] add_791506;
  wire [7:0] sel_791507;
  wire [7:0] add_791510;
  wire [7:0] sel_791511;
  wire [7:0] add_791514;
  wire [7:0] sel_791515;
  wire [7:0] add_791518;
  wire [7:0] sel_791519;
  wire [7:0] add_791522;
  wire [7:0] sel_791523;
  wire [7:0] add_791526;
  wire [7:0] sel_791527;
  wire [7:0] add_791530;
  wire [7:0] sel_791531;
  wire [7:0] add_791534;
  wire [7:0] sel_791535;
  wire [7:0] add_791538;
  wire [7:0] sel_791539;
  wire [7:0] add_791542;
  wire [7:0] sel_791543;
  wire [7:0] add_791546;
  wire [7:0] sel_791547;
  wire [7:0] add_791550;
  wire [7:0] sel_791551;
  wire [7:0] add_791554;
  wire [7:0] sel_791555;
  wire [7:0] add_791558;
  wire [7:0] sel_791559;
  wire [7:0] add_791562;
  wire [7:0] sel_791563;
  wire [7:0] add_791566;
  wire [7:0] sel_791567;
  wire [7:0] add_791570;
  wire [7:0] sel_791571;
  wire [7:0] add_791574;
  wire [7:0] sel_791575;
  wire [7:0] add_791578;
  wire [7:0] sel_791579;
  wire [7:0] add_791582;
  wire [7:0] sel_791583;
  wire [7:0] add_791586;
  wire [7:0] sel_791587;
  wire [7:0] add_791590;
  wire [7:0] sel_791591;
  wire [7:0] add_791594;
  wire [7:0] sel_791595;
  wire [7:0] add_791598;
  wire [7:0] sel_791599;
  wire [7:0] add_791602;
  wire [7:0] sel_791603;
  wire [7:0] add_791606;
  wire [7:0] sel_791607;
  wire [7:0] add_791610;
  wire [7:0] sel_791611;
  wire [7:0] add_791614;
  wire [7:0] sel_791615;
  wire [7:0] add_791618;
  wire [7:0] sel_791619;
  wire [7:0] add_791622;
  wire [7:0] sel_791623;
  wire [7:0] add_791626;
  wire [7:0] sel_791627;
  wire [7:0] add_791630;
  wire [7:0] sel_791631;
  wire [7:0] add_791634;
  wire [7:0] sel_791635;
  wire [7:0] add_791638;
  wire [7:0] sel_791639;
  wire [7:0] add_791643;
  wire [15:0] array_index_791644;
  wire [7:0] sel_791645;
  wire [7:0] add_791648;
  wire [7:0] sel_791649;
  wire [7:0] add_791652;
  wire [7:0] sel_791653;
  wire [7:0] add_791656;
  wire [7:0] sel_791657;
  wire [7:0] add_791660;
  wire [7:0] sel_791661;
  wire [7:0] add_791664;
  wire [7:0] sel_791665;
  wire [7:0] add_791668;
  wire [7:0] sel_791669;
  wire [7:0] add_791672;
  wire [7:0] sel_791673;
  wire [7:0] add_791676;
  wire [7:0] sel_791677;
  wire [7:0] add_791680;
  wire [7:0] sel_791681;
  wire [7:0] add_791684;
  wire [7:0] sel_791685;
  wire [7:0] add_791688;
  wire [7:0] sel_791689;
  wire [7:0] add_791692;
  wire [7:0] sel_791693;
  wire [7:0] add_791696;
  wire [7:0] sel_791697;
  wire [7:0] add_791700;
  wire [7:0] sel_791701;
  wire [7:0] add_791704;
  wire [7:0] sel_791705;
  wire [7:0] add_791708;
  wire [7:0] sel_791709;
  wire [7:0] add_791712;
  wire [7:0] sel_791713;
  wire [7:0] add_791716;
  wire [7:0] sel_791717;
  wire [7:0] add_791720;
  wire [7:0] sel_791721;
  wire [7:0] add_791724;
  wire [7:0] sel_791725;
  wire [7:0] add_791728;
  wire [7:0] sel_791729;
  wire [7:0] add_791732;
  wire [7:0] sel_791733;
  wire [7:0] add_791736;
  wire [7:0] sel_791737;
  wire [7:0] add_791740;
  wire [7:0] sel_791741;
  wire [7:0] add_791744;
  wire [7:0] sel_791745;
  wire [7:0] add_791748;
  wire [7:0] sel_791749;
  wire [7:0] add_791752;
  wire [7:0] sel_791753;
  wire [7:0] add_791756;
  wire [7:0] sel_791757;
  wire [7:0] add_791760;
  wire [7:0] sel_791761;
  wire [7:0] add_791764;
  wire [7:0] sel_791765;
  wire [7:0] add_791768;
  wire [7:0] sel_791769;
  wire [7:0] add_791772;
  wire [7:0] sel_791773;
  wire [7:0] add_791776;
  wire [7:0] sel_791777;
  wire [7:0] add_791780;
  wire [7:0] sel_791781;
  wire [7:0] add_791784;
  wire [7:0] sel_791785;
  wire [7:0] add_791788;
  wire [7:0] sel_791789;
  wire [7:0] add_791792;
  wire [7:0] sel_791793;
  wire [7:0] add_791796;
  wire [7:0] sel_791797;
  wire [7:0] add_791800;
  wire [7:0] sel_791801;
  wire [7:0] add_791804;
  wire [7:0] sel_791805;
  wire [7:0] add_791808;
  wire [7:0] sel_791809;
  wire [7:0] add_791812;
  wire [7:0] sel_791813;
  wire [7:0] add_791816;
  wire [7:0] sel_791817;
  wire [7:0] add_791820;
  wire [7:0] sel_791821;
  wire [7:0] add_791824;
  wire [7:0] sel_791825;
  wire [7:0] add_791828;
  wire [7:0] sel_791829;
  wire [7:0] add_791832;
  wire [7:0] sel_791833;
  wire [7:0] add_791836;
  wire [7:0] sel_791837;
  wire [7:0] add_791840;
  wire [7:0] sel_791841;
  wire [7:0] add_791844;
  wire [7:0] sel_791845;
  wire [7:0] add_791848;
  wire [7:0] sel_791849;
  wire [7:0] add_791852;
  wire [7:0] sel_791853;
  wire [7:0] add_791856;
  wire [7:0] sel_791857;
  wire [7:0] add_791860;
  wire [7:0] sel_791861;
  wire [7:0] add_791864;
  wire [7:0] sel_791865;
  wire [7:0] add_791868;
  wire [7:0] sel_791869;
  wire [7:0] add_791872;
  wire [7:0] sel_791873;
  wire [7:0] add_791876;
  wire [7:0] sel_791877;
  wire [7:0] add_791880;
  wire [7:0] sel_791881;
  wire [7:0] add_791884;
  wire [7:0] sel_791885;
  wire [7:0] add_791888;
  wire [7:0] sel_791889;
  wire [7:0] add_791892;
  wire [7:0] sel_791893;
  wire [7:0] add_791896;
  wire [7:0] sel_791897;
  wire [7:0] add_791900;
  wire [7:0] sel_791901;
  wire [7:0] add_791904;
  wire [7:0] sel_791905;
  wire [7:0] add_791908;
  wire [7:0] sel_791909;
  wire [7:0] add_791912;
  wire [7:0] sel_791913;
  wire [7:0] add_791916;
  wire [7:0] sel_791917;
  wire [7:0] add_791920;
  wire [7:0] sel_791921;
  wire [7:0] add_791924;
  wire [7:0] sel_791925;
  wire [7:0] add_791928;
  wire [7:0] sel_791929;
  wire [7:0] add_791932;
  wire [7:0] sel_791933;
  wire [7:0] add_791936;
  wire [7:0] sel_791937;
  wire [7:0] add_791940;
  wire [7:0] sel_791941;
  wire [7:0] add_791944;
  wire [7:0] sel_791945;
  wire [7:0] add_791948;
  wire [7:0] sel_791949;
  wire [7:0] add_791952;
  wire [7:0] sel_791953;
  wire [7:0] add_791956;
  wire [7:0] sel_791957;
  wire [7:0] add_791960;
  wire [7:0] sel_791961;
  wire [7:0] add_791964;
  wire [7:0] sel_791965;
  wire [7:0] add_791968;
  wire [7:0] sel_791969;
  wire [7:0] add_791972;
  wire [7:0] sel_791973;
  wire [7:0] add_791976;
  wire [7:0] sel_791977;
  wire [7:0] add_791980;
  wire [7:0] sel_791981;
  wire [7:0] add_791984;
  wire [7:0] sel_791985;
  wire [7:0] add_791988;
  wire [7:0] sel_791989;
  wire [7:0] add_791992;
  wire [7:0] sel_791993;
  wire [7:0] add_791996;
  wire [7:0] sel_791997;
  wire [7:0] add_792000;
  wire [7:0] sel_792001;
  wire [7:0] add_792005;
  wire [15:0] array_index_792006;
  wire [7:0] sel_792007;
  wire [7:0] add_792010;
  wire [7:0] sel_792011;
  wire [7:0] add_792014;
  wire [7:0] sel_792015;
  wire [7:0] add_792018;
  wire [7:0] sel_792019;
  wire [7:0] add_792022;
  wire [7:0] sel_792023;
  wire [7:0] add_792026;
  wire [7:0] sel_792027;
  wire [7:0] add_792030;
  wire [7:0] sel_792031;
  wire [7:0] add_792034;
  wire [7:0] sel_792035;
  wire [7:0] add_792038;
  wire [7:0] sel_792039;
  wire [7:0] add_792042;
  wire [7:0] sel_792043;
  wire [7:0] add_792046;
  wire [7:0] sel_792047;
  wire [7:0] add_792050;
  wire [7:0] sel_792051;
  wire [7:0] add_792054;
  wire [7:0] sel_792055;
  wire [7:0] add_792058;
  wire [7:0] sel_792059;
  wire [7:0] add_792062;
  wire [7:0] sel_792063;
  wire [7:0] add_792066;
  wire [7:0] sel_792067;
  wire [7:0] add_792070;
  wire [7:0] sel_792071;
  wire [7:0] add_792074;
  wire [7:0] sel_792075;
  wire [7:0] add_792078;
  wire [7:0] sel_792079;
  wire [7:0] add_792082;
  wire [7:0] sel_792083;
  wire [7:0] add_792086;
  wire [7:0] sel_792087;
  wire [7:0] add_792090;
  wire [7:0] sel_792091;
  wire [7:0] add_792094;
  wire [7:0] sel_792095;
  wire [7:0] add_792098;
  wire [7:0] sel_792099;
  wire [7:0] add_792102;
  wire [7:0] sel_792103;
  wire [7:0] add_792106;
  wire [7:0] sel_792107;
  wire [7:0] add_792110;
  wire [7:0] sel_792111;
  wire [7:0] add_792114;
  wire [7:0] sel_792115;
  wire [7:0] add_792118;
  wire [7:0] sel_792119;
  wire [7:0] add_792122;
  wire [7:0] sel_792123;
  wire [7:0] add_792126;
  wire [7:0] sel_792127;
  wire [7:0] add_792130;
  wire [7:0] sel_792131;
  wire [7:0] add_792134;
  wire [7:0] sel_792135;
  wire [7:0] add_792138;
  wire [7:0] sel_792139;
  wire [7:0] add_792142;
  wire [7:0] sel_792143;
  wire [7:0] add_792146;
  wire [7:0] sel_792147;
  wire [7:0] add_792150;
  wire [7:0] sel_792151;
  wire [7:0] add_792154;
  wire [7:0] sel_792155;
  wire [7:0] add_792158;
  wire [7:0] sel_792159;
  wire [7:0] add_792162;
  wire [7:0] sel_792163;
  wire [7:0] add_792166;
  wire [7:0] sel_792167;
  wire [7:0] add_792170;
  wire [7:0] sel_792171;
  wire [7:0] add_792174;
  wire [7:0] sel_792175;
  wire [7:0] add_792178;
  wire [7:0] sel_792179;
  wire [7:0] add_792182;
  wire [7:0] sel_792183;
  wire [7:0] add_792186;
  wire [7:0] sel_792187;
  wire [7:0] add_792190;
  wire [7:0] sel_792191;
  wire [7:0] add_792194;
  wire [7:0] sel_792195;
  wire [7:0] add_792198;
  wire [7:0] sel_792199;
  wire [7:0] add_792202;
  wire [7:0] sel_792203;
  wire [7:0] add_792206;
  wire [7:0] sel_792207;
  wire [7:0] add_792210;
  wire [7:0] sel_792211;
  wire [7:0] add_792214;
  wire [7:0] sel_792215;
  wire [7:0] add_792218;
  wire [7:0] sel_792219;
  wire [7:0] add_792222;
  wire [7:0] sel_792223;
  wire [7:0] add_792226;
  wire [7:0] sel_792227;
  wire [7:0] add_792230;
  wire [7:0] sel_792231;
  wire [7:0] add_792234;
  wire [7:0] sel_792235;
  wire [7:0] add_792238;
  wire [7:0] sel_792239;
  wire [7:0] add_792242;
  wire [7:0] sel_792243;
  wire [7:0] add_792246;
  wire [7:0] sel_792247;
  wire [7:0] add_792250;
  wire [7:0] sel_792251;
  wire [7:0] add_792254;
  wire [7:0] sel_792255;
  wire [7:0] add_792258;
  wire [7:0] sel_792259;
  wire [7:0] add_792262;
  wire [7:0] sel_792263;
  wire [7:0] add_792266;
  wire [7:0] sel_792267;
  wire [7:0] add_792270;
  wire [7:0] sel_792271;
  wire [7:0] add_792274;
  wire [7:0] sel_792275;
  wire [7:0] add_792278;
  wire [7:0] sel_792279;
  wire [7:0] add_792282;
  wire [7:0] sel_792283;
  wire [7:0] add_792286;
  wire [7:0] sel_792287;
  wire [7:0] add_792290;
  wire [7:0] sel_792291;
  wire [7:0] add_792294;
  wire [7:0] sel_792295;
  wire [7:0] add_792298;
  wire [7:0] sel_792299;
  wire [7:0] add_792302;
  wire [7:0] sel_792303;
  wire [7:0] add_792306;
  wire [7:0] sel_792307;
  wire [7:0] add_792310;
  wire [7:0] sel_792311;
  wire [7:0] add_792314;
  wire [7:0] sel_792315;
  wire [7:0] add_792318;
  wire [7:0] sel_792319;
  wire [7:0] add_792322;
  wire [7:0] sel_792323;
  wire [7:0] add_792326;
  wire [7:0] sel_792327;
  wire [7:0] add_792330;
  wire [7:0] sel_792331;
  wire [7:0] add_792334;
  wire [7:0] sel_792335;
  wire [7:0] add_792338;
  wire [7:0] sel_792339;
  wire [7:0] add_792342;
  wire [7:0] sel_792343;
  wire [7:0] add_792346;
  wire [7:0] sel_792347;
  wire [7:0] add_792350;
  wire [7:0] sel_792351;
  wire [7:0] add_792354;
  wire [7:0] sel_792355;
  wire [7:0] add_792358;
  wire [7:0] sel_792359;
  wire [7:0] add_792362;
  wire [7:0] sel_792363;
  wire [7:0] add_792367;
  wire [15:0] array_index_792368;
  wire [7:0] sel_792369;
  wire [7:0] add_792372;
  wire [7:0] sel_792373;
  wire [7:0] add_792376;
  wire [7:0] sel_792377;
  wire [7:0] add_792380;
  wire [7:0] sel_792381;
  wire [7:0] add_792384;
  wire [7:0] sel_792385;
  wire [7:0] add_792388;
  wire [7:0] sel_792389;
  wire [7:0] add_792392;
  wire [7:0] sel_792393;
  wire [7:0] add_792396;
  wire [7:0] sel_792397;
  wire [7:0] add_792400;
  wire [7:0] sel_792401;
  wire [7:0] add_792404;
  wire [7:0] sel_792405;
  wire [7:0] add_792408;
  wire [7:0] sel_792409;
  wire [7:0] add_792412;
  wire [7:0] sel_792413;
  wire [7:0] add_792416;
  wire [7:0] sel_792417;
  wire [7:0] add_792420;
  wire [7:0] sel_792421;
  wire [7:0] add_792424;
  wire [7:0] sel_792425;
  wire [7:0] add_792428;
  wire [7:0] sel_792429;
  wire [7:0] add_792432;
  wire [7:0] sel_792433;
  wire [7:0] add_792436;
  wire [7:0] sel_792437;
  wire [7:0] add_792440;
  wire [7:0] sel_792441;
  wire [7:0] add_792444;
  wire [7:0] sel_792445;
  wire [7:0] add_792448;
  wire [7:0] sel_792449;
  wire [7:0] add_792452;
  wire [7:0] sel_792453;
  wire [7:0] add_792456;
  wire [7:0] sel_792457;
  wire [7:0] add_792460;
  wire [7:0] sel_792461;
  wire [7:0] add_792464;
  wire [7:0] sel_792465;
  wire [7:0] add_792468;
  wire [7:0] sel_792469;
  wire [7:0] add_792472;
  wire [7:0] sel_792473;
  wire [7:0] add_792476;
  wire [7:0] sel_792477;
  wire [7:0] add_792480;
  wire [7:0] sel_792481;
  wire [7:0] add_792484;
  wire [7:0] sel_792485;
  wire [7:0] add_792488;
  wire [7:0] sel_792489;
  wire [7:0] add_792492;
  wire [7:0] sel_792493;
  wire [7:0] add_792496;
  wire [7:0] sel_792497;
  wire [7:0] add_792500;
  wire [7:0] sel_792501;
  wire [7:0] add_792504;
  wire [7:0] sel_792505;
  wire [7:0] add_792508;
  wire [7:0] sel_792509;
  wire [7:0] add_792512;
  wire [7:0] sel_792513;
  wire [7:0] add_792516;
  wire [7:0] sel_792517;
  wire [7:0] add_792520;
  wire [7:0] sel_792521;
  wire [7:0] add_792524;
  wire [7:0] sel_792525;
  wire [7:0] add_792528;
  wire [7:0] sel_792529;
  wire [7:0] add_792532;
  wire [7:0] sel_792533;
  wire [7:0] add_792536;
  wire [7:0] sel_792537;
  wire [7:0] add_792540;
  wire [7:0] sel_792541;
  wire [7:0] add_792544;
  wire [7:0] sel_792545;
  wire [7:0] add_792548;
  wire [7:0] sel_792549;
  wire [7:0] add_792552;
  wire [7:0] sel_792553;
  wire [7:0] add_792556;
  wire [7:0] sel_792557;
  wire [7:0] add_792560;
  wire [7:0] sel_792561;
  wire [7:0] add_792564;
  wire [7:0] sel_792565;
  wire [7:0] add_792568;
  wire [7:0] sel_792569;
  wire [7:0] add_792572;
  wire [7:0] sel_792573;
  wire [7:0] add_792576;
  wire [7:0] sel_792577;
  wire [7:0] add_792580;
  wire [7:0] sel_792581;
  wire [7:0] add_792584;
  wire [7:0] sel_792585;
  wire [7:0] add_792588;
  wire [7:0] sel_792589;
  wire [7:0] add_792592;
  wire [7:0] sel_792593;
  wire [7:0] add_792596;
  wire [7:0] sel_792597;
  wire [7:0] add_792600;
  wire [7:0] sel_792601;
  wire [7:0] add_792604;
  wire [7:0] sel_792605;
  wire [7:0] add_792608;
  wire [7:0] sel_792609;
  wire [7:0] add_792612;
  wire [7:0] sel_792613;
  wire [7:0] add_792616;
  wire [7:0] sel_792617;
  wire [7:0] add_792620;
  wire [7:0] sel_792621;
  wire [7:0] add_792624;
  wire [7:0] sel_792625;
  wire [7:0] add_792628;
  wire [7:0] sel_792629;
  wire [7:0] add_792632;
  wire [7:0] sel_792633;
  wire [7:0] add_792636;
  wire [7:0] sel_792637;
  wire [7:0] add_792640;
  wire [7:0] sel_792641;
  wire [7:0] add_792644;
  wire [7:0] sel_792645;
  wire [7:0] add_792648;
  wire [7:0] sel_792649;
  wire [7:0] add_792652;
  wire [7:0] sel_792653;
  wire [7:0] add_792656;
  wire [7:0] sel_792657;
  wire [7:0] add_792660;
  wire [7:0] sel_792661;
  wire [7:0] add_792664;
  wire [7:0] sel_792665;
  wire [7:0] add_792668;
  wire [7:0] sel_792669;
  wire [7:0] add_792672;
  wire [7:0] sel_792673;
  wire [7:0] add_792676;
  wire [7:0] sel_792677;
  wire [7:0] add_792680;
  wire [7:0] sel_792681;
  wire [7:0] add_792684;
  wire [7:0] sel_792685;
  wire [7:0] add_792688;
  wire [7:0] sel_792689;
  wire [7:0] add_792692;
  wire [7:0] sel_792693;
  wire [7:0] add_792696;
  wire [7:0] sel_792697;
  wire [7:0] add_792700;
  wire [7:0] sel_792701;
  wire [7:0] add_792704;
  wire [7:0] sel_792705;
  wire [7:0] add_792708;
  wire [7:0] sel_792709;
  wire [7:0] add_792712;
  wire [7:0] sel_792713;
  wire [7:0] add_792716;
  wire [7:0] sel_792717;
  wire [7:0] add_792720;
  wire [7:0] sel_792721;
  wire [7:0] add_792724;
  wire [7:0] sel_792725;
  wire [7:0] add_792729;
  wire [15:0] array_index_792730;
  wire [7:0] sel_792731;
  wire [7:0] add_792734;
  wire [7:0] sel_792735;
  wire [7:0] add_792738;
  wire [7:0] sel_792739;
  wire [7:0] add_792742;
  wire [7:0] sel_792743;
  wire [7:0] add_792746;
  wire [7:0] sel_792747;
  wire [7:0] add_792750;
  wire [7:0] sel_792751;
  wire [7:0] add_792754;
  wire [7:0] sel_792755;
  wire [7:0] add_792758;
  wire [7:0] sel_792759;
  wire [7:0] add_792762;
  wire [7:0] sel_792763;
  wire [7:0] add_792766;
  wire [7:0] sel_792767;
  wire [7:0] add_792770;
  wire [7:0] sel_792771;
  wire [7:0] add_792774;
  wire [7:0] sel_792775;
  wire [7:0] add_792778;
  wire [7:0] sel_792779;
  wire [7:0] add_792782;
  wire [7:0] sel_792783;
  wire [7:0] add_792786;
  wire [7:0] sel_792787;
  wire [7:0] add_792790;
  wire [7:0] sel_792791;
  wire [7:0] add_792794;
  wire [7:0] sel_792795;
  wire [7:0] add_792798;
  wire [7:0] sel_792799;
  wire [7:0] add_792802;
  wire [7:0] sel_792803;
  wire [7:0] add_792806;
  wire [7:0] sel_792807;
  wire [7:0] add_792810;
  wire [7:0] sel_792811;
  wire [7:0] add_792814;
  wire [7:0] sel_792815;
  wire [7:0] add_792818;
  wire [7:0] sel_792819;
  wire [7:0] add_792822;
  wire [7:0] sel_792823;
  wire [7:0] add_792826;
  wire [7:0] sel_792827;
  wire [7:0] add_792830;
  wire [7:0] sel_792831;
  wire [7:0] add_792834;
  wire [7:0] sel_792835;
  wire [7:0] add_792838;
  wire [7:0] sel_792839;
  wire [7:0] add_792842;
  wire [7:0] sel_792843;
  wire [7:0] add_792846;
  wire [7:0] sel_792847;
  wire [7:0] add_792850;
  wire [7:0] sel_792851;
  wire [7:0] add_792854;
  wire [7:0] sel_792855;
  wire [7:0] add_792858;
  wire [7:0] sel_792859;
  wire [7:0] add_792862;
  wire [7:0] sel_792863;
  wire [7:0] add_792866;
  wire [7:0] sel_792867;
  wire [7:0] add_792870;
  wire [7:0] sel_792871;
  wire [7:0] add_792874;
  wire [7:0] sel_792875;
  wire [7:0] add_792878;
  wire [7:0] sel_792879;
  wire [7:0] add_792882;
  wire [7:0] sel_792883;
  wire [7:0] add_792886;
  wire [7:0] sel_792887;
  wire [7:0] add_792890;
  wire [7:0] sel_792891;
  wire [7:0] add_792894;
  wire [7:0] sel_792895;
  wire [7:0] add_792898;
  wire [7:0] sel_792899;
  wire [7:0] add_792902;
  wire [7:0] sel_792903;
  wire [7:0] add_792906;
  wire [7:0] sel_792907;
  wire [7:0] add_792910;
  wire [7:0] sel_792911;
  wire [7:0] add_792914;
  wire [7:0] sel_792915;
  wire [7:0] add_792918;
  wire [7:0] sel_792919;
  wire [7:0] add_792922;
  wire [7:0] sel_792923;
  wire [7:0] add_792926;
  wire [7:0] sel_792927;
  wire [7:0] add_792930;
  wire [7:0] sel_792931;
  wire [7:0] add_792934;
  wire [7:0] sel_792935;
  wire [7:0] add_792938;
  wire [7:0] sel_792939;
  wire [7:0] add_792942;
  wire [7:0] sel_792943;
  wire [7:0] add_792946;
  wire [7:0] sel_792947;
  wire [7:0] add_792950;
  wire [7:0] sel_792951;
  wire [7:0] add_792954;
  wire [7:0] sel_792955;
  wire [7:0] add_792958;
  wire [7:0] sel_792959;
  wire [7:0] add_792962;
  wire [7:0] sel_792963;
  wire [7:0] add_792966;
  wire [7:0] sel_792967;
  wire [7:0] add_792970;
  wire [7:0] sel_792971;
  wire [7:0] add_792974;
  wire [7:0] sel_792975;
  wire [7:0] add_792978;
  wire [7:0] sel_792979;
  wire [7:0] add_792982;
  wire [7:0] sel_792983;
  wire [7:0] add_792986;
  wire [7:0] sel_792987;
  wire [7:0] add_792990;
  wire [7:0] sel_792991;
  wire [7:0] add_792994;
  wire [7:0] sel_792995;
  wire [7:0] add_792998;
  wire [7:0] sel_792999;
  wire [7:0] add_793002;
  wire [7:0] sel_793003;
  wire [7:0] add_793006;
  wire [7:0] sel_793007;
  wire [7:0] add_793010;
  wire [7:0] sel_793011;
  wire [7:0] add_793014;
  wire [7:0] sel_793015;
  wire [7:0] add_793018;
  wire [7:0] sel_793019;
  wire [7:0] add_793022;
  wire [7:0] sel_793023;
  wire [7:0] add_793026;
  wire [7:0] sel_793027;
  wire [7:0] add_793030;
  wire [7:0] sel_793031;
  wire [7:0] add_793034;
  wire [7:0] sel_793035;
  wire [7:0] add_793038;
  wire [7:0] sel_793039;
  wire [7:0] add_793042;
  wire [7:0] sel_793043;
  wire [7:0] add_793046;
  wire [7:0] sel_793047;
  wire [7:0] add_793050;
  wire [7:0] sel_793051;
  wire [7:0] add_793054;
  wire [7:0] sel_793055;
  wire [7:0] add_793058;
  wire [7:0] sel_793059;
  wire [7:0] add_793062;
  wire [7:0] sel_793063;
  wire [7:0] add_793066;
  wire [7:0] sel_793067;
  wire [7:0] add_793070;
  wire [7:0] sel_793071;
  wire [7:0] add_793074;
  wire [7:0] sel_793075;
  wire [7:0] add_793078;
  wire [7:0] sel_793079;
  wire [7:0] add_793082;
  wire [7:0] sel_793083;
  wire [7:0] add_793086;
  wire [7:0] sel_793087;
  wire [7:0] add_793091;
  wire [15:0] array_index_793092;
  wire [7:0] sel_793093;
  wire [7:0] add_793096;
  wire [7:0] sel_793097;
  wire [7:0] add_793100;
  wire [7:0] sel_793101;
  wire [7:0] add_793104;
  wire [7:0] sel_793105;
  wire [7:0] add_793108;
  wire [7:0] sel_793109;
  wire [7:0] add_793112;
  wire [7:0] sel_793113;
  wire [7:0] add_793116;
  wire [7:0] sel_793117;
  wire [7:0] add_793120;
  wire [7:0] sel_793121;
  wire [7:0] add_793124;
  wire [7:0] sel_793125;
  wire [7:0] add_793128;
  wire [7:0] sel_793129;
  wire [7:0] add_793132;
  wire [7:0] sel_793133;
  wire [7:0] add_793136;
  wire [7:0] sel_793137;
  wire [7:0] add_793140;
  wire [7:0] sel_793141;
  wire [7:0] add_793144;
  wire [7:0] sel_793145;
  wire [7:0] add_793148;
  wire [7:0] sel_793149;
  wire [7:0] add_793152;
  wire [7:0] sel_793153;
  wire [7:0] add_793156;
  wire [7:0] sel_793157;
  wire [7:0] add_793160;
  wire [7:0] sel_793161;
  wire [7:0] add_793164;
  wire [7:0] sel_793165;
  wire [7:0] add_793168;
  wire [7:0] sel_793169;
  wire [7:0] add_793172;
  wire [7:0] sel_793173;
  wire [7:0] add_793176;
  wire [7:0] sel_793177;
  wire [7:0] add_793180;
  wire [7:0] sel_793181;
  wire [7:0] add_793184;
  wire [7:0] sel_793185;
  wire [7:0] add_793188;
  wire [7:0] sel_793189;
  wire [7:0] add_793192;
  wire [7:0] sel_793193;
  wire [7:0] add_793196;
  wire [7:0] sel_793197;
  wire [7:0] add_793200;
  wire [7:0] sel_793201;
  wire [7:0] add_793204;
  wire [7:0] sel_793205;
  wire [7:0] add_793208;
  wire [7:0] sel_793209;
  wire [7:0] add_793212;
  wire [7:0] sel_793213;
  wire [7:0] add_793216;
  wire [7:0] sel_793217;
  wire [7:0] add_793220;
  wire [7:0] sel_793221;
  wire [7:0] add_793224;
  wire [7:0] sel_793225;
  wire [7:0] add_793228;
  wire [7:0] sel_793229;
  wire [7:0] add_793232;
  wire [7:0] sel_793233;
  wire [7:0] add_793236;
  wire [7:0] sel_793237;
  wire [7:0] add_793240;
  wire [7:0] sel_793241;
  wire [7:0] add_793244;
  wire [7:0] sel_793245;
  wire [7:0] add_793248;
  wire [7:0] sel_793249;
  wire [7:0] add_793252;
  wire [7:0] sel_793253;
  wire [7:0] add_793256;
  wire [7:0] sel_793257;
  wire [7:0] add_793260;
  wire [7:0] sel_793261;
  wire [7:0] add_793264;
  wire [7:0] sel_793265;
  wire [7:0] add_793268;
  wire [7:0] sel_793269;
  wire [7:0] add_793272;
  wire [7:0] sel_793273;
  wire [7:0] add_793276;
  wire [7:0] sel_793277;
  wire [7:0] add_793280;
  wire [7:0] sel_793281;
  wire [7:0] add_793284;
  wire [7:0] sel_793285;
  wire [7:0] add_793288;
  wire [7:0] sel_793289;
  wire [7:0] add_793292;
  wire [7:0] sel_793293;
  wire [7:0] add_793296;
  wire [7:0] sel_793297;
  wire [7:0] add_793300;
  wire [7:0] sel_793301;
  wire [7:0] add_793304;
  wire [7:0] sel_793305;
  wire [7:0] add_793308;
  wire [7:0] sel_793309;
  wire [7:0] add_793312;
  wire [7:0] sel_793313;
  wire [7:0] add_793316;
  wire [7:0] sel_793317;
  wire [7:0] add_793320;
  wire [7:0] sel_793321;
  wire [7:0] add_793324;
  wire [7:0] sel_793325;
  wire [7:0] add_793328;
  wire [7:0] sel_793329;
  wire [7:0] add_793332;
  wire [7:0] sel_793333;
  wire [7:0] add_793336;
  wire [7:0] sel_793337;
  wire [7:0] add_793340;
  wire [7:0] sel_793341;
  wire [7:0] add_793344;
  wire [7:0] sel_793345;
  wire [7:0] add_793348;
  wire [7:0] sel_793349;
  wire [7:0] add_793352;
  wire [7:0] sel_793353;
  wire [7:0] add_793356;
  wire [7:0] sel_793357;
  wire [7:0] add_793360;
  wire [7:0] sel_793361;
  wire [7:0] add_793364;
  wire [7:0] sel_793365;
  wire [7:0] add_793368;
  wire [7:0] sel_793369;
  wire [7:0] add_793372;
  wire [7:0] sel_793373;
  wire [7:0] add_793376;
  wire [7:0] sel_793377;
  wire [7:0] add_793380;
  wire [7:0] sel_793381;
  wire [7:0] add_793384;
  wire [7:0] sel_793385;
  wire [7:0] add_793388;
  wire [7:0] sel_793389;
  wire [7:0] add_793392;
  wire [7:0] sel_793393;
  wire [7:0] add_793396;
  wire [7:0] sel_793397;
  wire [7:0] add_793400;
  wire [7:0] sel_793401;
  wire [7:0] add_793404;
  wire [7:0] sel_793405;
  wire [7:0] add_793408;
  wire [7:0] sel_793409;
  wire [7:0] add_793412;
  wire [7:0] sel_793413;
  wire [7:0] add_793416;
  wire [7:0] sel_793417;
  wire [7:0] add_793420;
  wire [7:0] sel_793421;
  wire [7:0] add_793424;
  wire [7:0] sel_793425;
  wire [7:0] add_793428;
  wire [7:0] sel_793429;
  wire [7:0] add_793432;
  wire [7:0] sel_793433;
  wire [7:0] add_793436;
  wire [7:0] sel_793437;
  wire [7:0] add_793440;
  wire [7:0] sel_793441;
  wire [7:0] add_793444;
  wire [7:0] sel_793445;
  wire [7:0] add_793448;
  wire [7:0] sel_793449;
  wire [7:0] add_793453;
  wire [15:0] array_index_793454;
  wire [7:0] sel_793455;
  wire [7:0] add_793458;
  wire [7:0] sel_793459;
  wire [7:0] add_793462;
  wire [7:0] sel_793463;
  wire [7:0] add_793466;
  wire [7:0] sel_793467;
  wire [7:0] add_793470;
  wire [7:0] sel_793471;
  wire [7:0] add_793474;
  wire [7:0] sel_793475;
  wire [7:0] add_793478;
  wire [7:0] sel_793479;
  wire [7:0] add_793482;
  wire [7:0] sel_793483;
  wire [7:0] add_793486;
  wire [7:0] sel_793487;
  wire [7:0] add_793490;
  wire [7:0] sel_793491;
  wire [7:0] add_793494;
  wire [7:0] sel_793495;
  wire [7:0] add_793498;
  wire [7:0] sel_793499;
  wire [7:0] add_793502;
  wire [7:0] sel_793503;
  wire [7:0] add_793506;
  wire [7:0] sel_793507;
  wire [7:0] add_793510;
  wire [7:0] sel_793511;
  wire [7:0] add_793514;
  wire [7:0] sel_793515;
  wire [7:0] add_793518;
  wire [7:0] sel_793519;
  wire [7:0] add_793522;
  wire [7:0] sel_793523;
  wire [7:0] add_793526;
  wire [7:0] sel_793527;
  wire [7:0] add_793530;
  wire [7:0] sel_793531;
  wire [7:0] add_793534;
  wire [7:0] sel_793535;
  wire [7:0] add_793538;
  wire [7:0] sel_793539;
  wire [7:0] add_793542;
  wire [7:0] sel_793543;
  wire [7:0] add_793546;
  wire [7:0] sel_793547;
  wire [7:0] add_793550;
  wire [7:0] sel_793551;
  wire [7:0] add_793554;
  wire [7:0] sel_793555;
  wire [7:0] add_793558;
  wire [7:0] sel_793559;
  wire [7:0] add_793562;
  wire [7:0] sel_793563;
  wire [7:0] add_793566;
  wire [7:0] sel_793567;
  wire [7:0] add_793570;
  wire [7:0] sel_793571;
  wire [7:0] add_793574;
  wire [7:0] sel_793575;
  wire [7:0] add_793578;
  wire [7:0] sel_793579;
  wire [7:0] add_793582;
  wire [7:0] sel_793583;
  wire [7:0] add_793586;
  wire [7:0] sel_793587;
  wire [7:0] add_793590;
  wire [7:0] sel_793591;
  wire [7:0] add_793594;
  wire [7:0] sel_793595;
  wire [7:0] add_793598;
  wire [7:0] sel_793599;
  wire [7:0] add_793602;
  wire [7:0] sel_793603;
  wire [7:0] add_793606;
  wire [7:0] sel_793607;
  wire [7:0] add_793610;
  wire [7:0] sel_793611;
  wire [7:0] add_793614;
  wire [7:0] sel_793615;
  wire [7:0] add_793618;
  wire [7:0] sel_793619;
  wire [7:0] add_793622;
  wire [7:0] sel_793623;
  wire [7:0] add_793626;
  wire [7:0] sel_793627;
  wire [7:0] add_793630;
  wire [7:0] sel_793631;
  wire [7:0] add_793634;
  wire [7:0] sel_793635;
  wire [7:0] add_793638;
  wire [7:0] sel_793639;
  wire [7:0] add_793642;
  wire [7:0] sel_793643;
  wire [7:0] add_793646;
  wire [7:0] sel_793647;
  wire [7:0] add_793650;
  wire [7:0] sel_793651;
  wire [7:0] add_793654;
  wire [7:0] sel_793655;
  wire [7:0] add_793658;
  wire [7:0] sel_793659;
  wire [7:0] add_793662;
  wire [7:0] sel_793663;
  wire [7:0] add_793666;
  wire [7:0] sel_793667;
  wire [7:0] add_793670;
  wire [7:0] sel_793671;
  wire [7:0] add_793674;
  wire [7:0] sel_793675;
  wire [7:0] add_793678;
  wire [7:0] sel_793679;
  wire [7:0] add_793682;
  wire [7:0] sel_793683;
  wire [7:0] add_793686;
  wire [7:0] sel_793687;
  wire [7:0] add_793690;
  wire [7:0] sel_793691;
  wire [7:0] add_793694;
  wire [7:0] sel_793695;
  wire [7:0] add_793698;
  wire [7:0] sel_793699;
  wire [7:0] add_793702;
  wire [7:0] sel_793703;
  wire [7:0] add_793706;
  wire [7:0] sel_793707;
  wire [7:0] add_793710;
  wire [7:0] sel_793711;
  wire [7:0] add_793714;
  wire [7:0] sel_793715;
  wire [7:0] add_793718;
  wire [7:0] sel_793719;
  wire [7:0] add_793722;
  wire [7:0] sel_793723;
  wire [7:0] add_793726;
  wire [7:0] sel_793727;
  wire [7:0] add_793730;
  wire [7:0] sel_793731;
  wire [7:0] add_793734;
  wire [7:0] sel_793735;
  wire [7:0] add_793738;
  wire [7:0] sel_793739;
  wire [7:0] add_793742;
  wire [7:0] sel_793743;
  wire [7:0] add_793746;
  wire [7:0] sel_793747;
  wire [7:0] add_793750;
  wire [7:0] sel_793751;
  wire [7:0] add_793754;
  wire [7:0] sel_793755;
  wire [7:0] add_793758;
  wire [7:0] sel_793759;
  wire [7:0] add_793762;
  wire [7:0] sel_793763;
  wire [7:0] add_793766;
  wire [7:0] sel_793767;
  wire [7:0] add_793770;
  wire [7:0] sel_793771;
  wire [7:0] add_793774;
  wire [7:0] sel_793775;
  wire [7:0] add_793778;
  wire [7:0] sel_793779;
  wire [7:0] add_793782;
  wire [7:0] sel_793783;
  wire [7:0] add_793786;
  wire [7:0] sel_793787;
  wire [7:0] add_793790;
  wire [7:0] sel_793791;
  wire [7:0] add_793794;
  wire [7:0] sel_793795;
  wire [7:0] add_793798;
  wire [7:0] sel_793799;
  wire [7:0] add_793802;
  wire [7:0] sel_793803;
  wire [7:0] add_793806;
  wire [7:0] sel_793807;
  wire [7:0] add_793810;
  wire [7:0] sel_793811;
  wire [7:0] add_793815;
  wire [15:0] array_index_793816;
  wire [7:0] sel_793817;
  wire [7:0] add_793820;
  wire [7:0] sel_793821;
  wire [7:0] add_793824;
  wire [7:0] sel_793825;
  wire [7:0] add_793828;
  wire [7:0] sel_793829;
  wire [7:0] add_793832;
  wire [7:0] sel_793833;
  wire [7:0] add_793836;
  wire [7:0] sel_793837;
  wire [7:0] add_793840;
  wire [7:0] sel_793841;
  wire [7:0] add_793844;
  wire [7:0] sel_793845;
  wire [7:0] add_793848;
  wire [7:0] sel_793849;
  wire [7:0] add_793852;
  wire [7:0] sel_793853;
  wire [7:0] add_793856;
  wire [7:0] sel_793857;
  wire [7:0] add_793860;
  wire [7:0] sel_793861;
  wire [7:0] add_793864;
  wire [7:0] sel_793865;
  wire [7:0] add_793868;
  wire [7:0] sel_793869;
  wire [7:0] add_793872;
  wire [7:0] sel_793873;
  wire [7:0] add_793876;
  wire [7:0] sel_793877;
  wire [7:0] add_793880;
  wire [7:0] sel_793881;
  wire [7:0] add_793884;
  wire [7:0] sel_793885;
  wire [7:0] add_793888;
  wire [7:0] sel_793889;
  wire [7:0] add_793892;
  wire [7:0] sel_793893;
  wire [7:0] add_793896;
  wire [7:0] sel_793897;
  wire [7:0] add_793900;
  wire [7:0] sel_793901;
  wire [7:0] add_793904;
  wire [7:0] sel_793905;
  wire [7:0] add_793908;
  wire [7:0] sel_793909;
  wire [7:0] add_793912;
  wire [7:0] sel_793913;
  wire [7:0] add_793916;
  wire [7:0] sel_793917;
  wire [7:0] add_793920;
  wire [7:0] sel_793921;
  wire [7:0] add_793924;
  wire [7:0] sel_793925;
  wire [7:0] add_793928;
  wire [7:0] sel_793929;
  wire [7:0] add_793932;
  wire [7:0] sel_793933;
  wire [7:0] add_793936;
  wire [7:0] sel_793937;
  wire [7:0] add_793940;
  wire [7:0] sel_793941;
  wire [7:0] add_793944;
  wire [7:0] sel_793945;
  wire [7:0] add_793948;
  wire [7:0] sel_793949;
  wire [7:0] add_793952;
  wire [7:0] sel_793953;
  wire [7:0] add_793956;
  wire [7:0] sel_793957;
  wire [7:0] add_793960;
  wire [7:0] sel_793961;
  wire [7:0] add_793964;
  wire [7:0] sel_793965;
  wire [7:0] add_793968;
  wire [7:0] sel_793969;
  wire [7:0] add_793972;
  wire [7:0] sel_793973;
  wire [7:0] add_793976;
  wire [7:0] sel_793977;
  wire [7:0] add_793980;
  wire [7:0] sel_793981;
  wire [7:0] add_793984;
  wire [7:0] sel_793985;
  wire [7:0] add_793988;
  wire [7:0] sel_793989;
  wire [7:0] add_793992;
  wire [7:0] sel_793993;
  wire [7:0] add_793996;
  wire [7:0] sel_793997;
  wire [7:0] add_794000;
  wire [7:0] sel_794001;
  wire [7:0] add_794004;
  wire [7:0] sel_794005;
  wire [7:0] add_794008;
  wire [7:0] sel_794009;
  wire [7:0] add_794012;
  wire [7:0] sel_794013;
  wire [7:0] add_794016;
  wire [7:0] sel_794017;
  wire [7:0] add_794020;
  wire [7:0] sel_794021;
  wire [7:0] add_794024;
  wire [7:0] sel_794025;
  wire [7:0] add_794028;
  wire [7:0] sel_794029;
  wire [7:0] add_794032;
  wire [7:0] sel_794033;
  wire [7:0] add_794036;
  wire [7:0] sel_794037;
  wire [7:0] add_794040;
  wire [7:0] sel_794041;
  wire [7:0] add_794044;
  wire [7:0] sel_794045;
  wire [7:0] add_794048;
  wire [7:0] sel_794049;
  wire [7:0] add_794052;
  wire [7:0] sel_794053;
  wire [7:0] add_794056;
  wire [7:0] sel_794057;
  wire [7:0] add_794060;
  wire [7:0] sel_794061;
  wire [7:0] add_794064;
  wire [7:0] sel_794065;
  wire [7:0] add_794068;
  wire [7:0] sel_794069;
  wire [7:0] add_794072;
  wire [7:0] sel_794073;
  wire [7:0] add_794076;
  wire [7:0] sel_794077;
  wire [7:0] add_794080;
  wire [7:0] sel_794081;
  wire [7:0] add_794084;
  wire [7:0] sel_794085;
  wire [7:0] add_794088;
  wire [7:0] sel_794089;
  wire [7:0] add_794092;
  wire [7:0] sel_794093;
  wire [7:0] add_794096;
  wire [7:0] sel_794097;
  wire [7:0] add_794100;
  wire [7:0] sel_794101;
  wire [7:0] add_794104;
  wire [7:0] sel_794105;
  wire [7:0] add_794108;
  wire [7:0] sel_794109;
  wire [7:0] add_794112;
  wire [7:0] sel_794113;
  wire [7:0] add_794116;
  wire [7:0] sel_794117;
  wire [7:0] add_794120;
  wire [7:0] sel_794121;
  wire [7:0] add_794124;
  wire [7:0] sel_794125;
  wire [7:0] add_794128;
  wire [7:0] sel_794129;
  wire [7:0] add_794132;
  wire [7:0] sel_794133;
  wire [7:0] add_794136;
  wire [7:0] sel_794137;
  wire [7:0] add_794140;
  wire [7:0] sel_794141;
  wire [7:0] add_794144;
  wire [7:0] sel_794145;
  wire [7:0] add_794148;
  wire [7:0] sel_794149;
  wire [7:0] add_794152;
  wire [7:0] sel_794153;
  wire [7:0] add_794156;
  wire [7:0] sel_794157;
  wire [7:0] add_794160;
  wire [7:0] sel_794161;
  wire [7:0] add_794164;
  wire [7:0] sel_794165;
  wire [7:0] add_794168;
  wire [7:0] sel_794169;
  wire [7:0] add_794172;
  wire [7:0] sel_794173;
  wire [7:0] add_794177;
  wire [15:0] array_index_794178;
  wire [7:0] sel_794179;
  wire [7:0] add_794182;
  wire [7:0] sel_794183;
  wire [7:0] add_794186;
  wire [7:0] sel_794187;
  wire [7:0] add_794190;
  wire [7:0] sel_794191;
  wire [7:0] add_794194;
  wire [7:0] sel_794195;
  wire [7:0] add_794198;
  wire [7:0] sel_794199;
  wire [7:0] add_794202;
  wire [7:0] sel_794203;
  wire [7:0] add_794206;
  wire [7:0] sel_794207;
  wire [7:0] add_794210;
  wire [7:0] sel_794211;
  wire [7:0] add_794214;
  wire [7:0] sel_794215;
  wire [7:0] add_794218;
  wire [7:0] sel_794219;
  wire [7:0] add_794222;
  wire [7:0] sel_794223;
  wire [7:0] add_794226;
  wire [7:0] sel_794227;
  wire [7:0] add_794230;
  wire [7:0] sel_794231;
  wire [7:0] add_794234;
  wire [7:0] sel_794235;
  wire [7:0] add_794238;
  wire [7:0] sel_794239;
  wire [7:0] add_794242;
  wire [7:0] sel_794243;
  wire [7:0] add_794246;
  wire [7:0] sel_794247;
  wire [7:0] add_794250;
  wire [7:0] sel_794251;
  wire [7:0] add_794254;
  wire [7:0] sel_794255;
  wire [7:0] add_794258;
  wire [7:0] sel_794259;
  wire [7:0] add_794262;
  wire [7:0] sel_794263;
  wire [7:0] add_794266;
  wire [7:0] sel_794267;
  wire [7:0] add_794270;
  wire [7:0] sel_794271;
  wire [7:0] add_794274;
  wire [7:0] sel_794275;
  wire [7:0] add_794278;
  wire [7:0] sel_794279;
  wire [7:0] add_794282;
  wire [7:0] sel_794283;
  wire [7:0] add_794286;
  wire [7:0] sel_794287;
  wire [7:0] add_794290;
  wire [7:0] sel_794291;
  wire [7:0] add_794294;
  wire [7:0] sel_794295;
  wire [7:0] add_794298;
  wire [7:0] sel_794299;
  wire [7:0] add_794302;
  wire [7:0] sel_794303;
  wire [7:0] add_794306;
  wire [7:0] sel_794307;
  wire [7:0] add_794310;
  wire [7:0] sel_794311;
  wire [7:0] add_794314;
  wire [7:0] sel_794315;
  wire [7:0] add_794318;
  wire [7:0] sel_794319;
  wire [7:0] add_794322;
  wire [7:0] sel_794323;
  wire [7:0] add_794326;
  wire [7:0] sel_794327;
  wire [7:0] add_794330;
  wire [7:0] sel_794331;
  wire [7:0] add_794334;
  wire [7:0] sel_794335;
  wire [7:0] add_794338;
  wire [7:0] sel_794339;
  wire [7:0] add_794342;
  wire [7:0] sel_794343;
  wire [7:0] add_794346;
  wire [7:0] sel_794347;
  wire [7:0] add_794350;
  wire [7:0] sel_794351;
  wire [7:0] add_794354;
  wire [7:0] sel_794355;
  wire [7:0] add_794358;
  wire [7:0] sel_794359;
  wire [7:0] add_794362;
  wire [7:0] sel_794363;
  wire [7:0] add_794366;
  wire [7:0] sel_794367;
  wire [7:0] add_794370;
  wire [7:0] sel_794371;
  wire [7:0] add_794374;
  wire [7:0] sel_794375;
  wire [7:0] add_794378;
  wire [7:0] sel_794379;
  wire [7:0] add_794382;
  wire [7:0] sel_794383;
  wire [7:0] add_794386;
  wire [7:0] sel_794387;
  wire [7:0] add_794390;
  wire [7:0] sel_794391;
  wire [7:0] add_794394;
  wire [7:0] sel_794395;
  wire [7:0] add_794398;
  wire [7:0] sel_794399;
  wire [7:0] add_794402;
  wire [7:0] sel_794403;
  wire [7:0] add_794406;
  wire [7:0] sel_794407;
  wire [7:0] add_794410;
  wire [7:0] sel_794411;
  wire [7:0] add_794414;
  wire [7:0] sel_794415;
  wire [7:0] add_794418;
  wire [7:0] sel_794419;
  wire [7:0] add_794422;
  wire [7:0] sel_794423;
  wire [7:0] add_794426;
  wire [7:0] sel_794427;
  wire [7:0] add_794430;
  wire [7:0] sel_794431;
  wire [7:0] add_794434;
  wire [7:0] sel_794435;
  wire [7:0] add_794438;
  wire [7:0] sel_794439;
  wire [7:0] add_794442;
  wire [7:0] sel_794443;
  wire [7:0] add_794446;
  wire [7:0] sel_794447;
  wire [7:0] add_794450;
  wire [7:0] sel_794451;
  wire [7:0] add_794454;
  wire [7:0] sel_794455;
  wire [7:0] add_794458;
  wire [7:0] sel_794459;
  wire [7:0] add_794462;
  wire [7:0] sel_794463;
  wire [7:0] add_794466;
  wire [7:0] sel_794467;
  wire [7:0] add_794470;
  wire [7:0] sel_794471;
  wire [7:0] add_794474;
  wire [7:0] sel_794475;
  wire [7:0] add_794478;
  wire [7:0] sel_794479;
  wire [7:0] add_794482;
  wire [7:0] sel_794483;
  wire [7:0] add_794486;
  wire [7:0] sel_794487;
  wire [7:0] add_794490;
  wire [7:0] sel_794491;
  wire [7:0] add_794494;
  wire [7:0] sel_794495;
  wire [7:0] add_794498;
  wire [7:0] sel_794499;
  wire [7:0] add_794502;
  wire [7:0] sel_794503;
  wire [7:0] add_794506;
  wire [7:0] sel_794507;
  wire [7:0] add_794510;
  wire [7:0] sel_794511;
  wire [7:0] add_794514;
  wire [7:0] sel_794515;
  wire [7:0] add_794518;
  wire [7:0] sel_794519;
  wire [7:0] add_794522;
  wire [7:0] sel_794523;
  wire [7:0] add_794526;
  wire [7:0] sel_794527;
  wire [7:0] add_794530;
  wire [7:0] sel_794531;
  wire [7:0] add_794534;
  wire [7:0] sel_794535;
  wire [7:0] add_794539;
  wire [15:0] array_index_794540;
  wire [7:0] sel_794541;
  wire [7:0] add_794544;
  wire [7:0] sel_794545;
  wire [7:0] add_794548;
  wire [7:0] sel_794549;
  wire [7:0] add_794552;
  wire [7:0] sel_794553;
  wire [7:0] add_794556;
  wire [7:0] sel_794557;
  wire [7:0] add_794560;
  wire [7:0] sel_794561;
  wire [7:0] add_794564;
  wire [7:0] sel_794565;
  wire [7:0] add_794568;
  wire [7:0] sel_794569;
  wire [7:0] add_794572;
  wire [7:0] sel_794573;
  wire [7:0] add_794576;
  wire [7:0] sel_794577;
  wire [7:0] add_794580;
  wire [7:0] sel_794581;
  wire [7:0] add_794584;
  wire [7:0] sel_794585;
  wire [7:0] add_794588;
  wire [7:0] sel_794589;
  wire [7:0] add_794592;
  wire [7:0] sel_794593;
  wire [7:0] add_794596;
  wire [7:0] sel_794597;
  wire [7:0] add_794600;
  wire [7:0] sel_794601;
  wire [7:0] add_794604;
  wire [7:0] sel_794605;
  wire [7:0] add_794608;
  wire [7:0] sel_794609;
  wire [7:0] add_794612;
  wire [7:0] sel_794613;
  wire [7:0] add_794616;
  wire [7:0] sel_794617;
  wire [7:0] add_794620;
  wire [7:0] sel_794621;
  wire [7:0] add_794624;
  wire [7:0] sel_794625;
  wire [7:0] add_794628;
  wire [7:0] sel_794629;
  wire [7:0] add_794632;
  wire [7:0] sel_794633;
  wire [7:0] add_794636;
  wire [7:0] sel_794637;
  wire [7:0] add_794640;
  wire [7:0] sel_794641;
  wire [7:0] add_794644;
  wire [7:0] sel_794645;
  wire [7:0] add_794648;
  wire [7:0] sel_794649;
  wire [7:0] add_794652;
  wire [7:0] sel_794653;
  wire [7:0] add_794656;
  wire [7:0] sel_794657;
  wire [7:0] add_794660;
  wire [7:0] sel_794661;
  wire [7:0] add_794664;
  wire [7:0] sel_794665;
  wire [7:0] add_794668;
  wire [7:0] sel_794669;
  wire [7:0] add_794672;
  wire [7:0] sel_794673;
  wire [7:0] add_794676;
  wire [7:0] sel_794677;
  wire [7:0] add_794680;
  wire [7:0] sel_794681;
  wire [7:0] add_794684;
  wire [7:0] sel_794685;
  wire [7:0] add_794688;
  wire [7:0] sel_794689;
  wire [7:0] add_794692;
  wire [7:0] sel_794693;
  wire [7:0] add_794696;
  wire [7:0] sel_794697;
  wire [7:0] add_794700;
  wire [7:0] sel_794701;
  wire [7:0] add_794704;
  wire [7:0] sel_794705;
  wire [7:0] add_794708;
  wire [7:0] sel_794709;
  wire [7:0] add_794712;
  wire [7:0] sel_794713;
  wire [7:0] add_794716;
  wire [7:0] sel_794717;
  wire [7:0] add_794720;
  wire [7:0] sel_794721;
  wire [7:0] add_794724;
  wire [7:0] sel_794725;
  wire [7:0] add_794728;
  wire [7:0] sel_794729;
  wire [7:0] add_794732;
  wire [7:0] sel_794733;
  wire [7:0] add_794736;
  wire [7:0] sel_794737;
  wire [7:0] add_794740;
  wire [7:0] sel_794741;
  wire [7:0] add_794744;
  wire [7:0] sel_794745;
  wire [7:0] add_794748;
  wire [7:0] sel_794749;
  wire [7:0] add_794752;
  wire [7:0] sel_794753;
  wire [7:0] add_794756;
  wire [7:0] sel_794757;
  wire [7:0] add_794760;
  wire [7:0] sel_794761;
  wire [7:0] add_794764;
  wire [7:0] sel_794765;
  wire [7:0] add_794768;
  wire [7:0] sel_794769;
  wire [7:0] add_794772;
  wire [7:0] sel_794773;
  wire [7:0] add_794776;
  wire [7:0] sel_794777;
  wire [7:0] add_794780;
  wire [7:0] sel_794781;
  wire [7:0] add_794784;
  wire [7:0] sel_794785;
  wire [7:0] add_794788;
  wire [7:0] sel_794789;
  wire [7:0] add_794792;
  wire [7:0] sel_794793;
  wire [7:0] add_794796;
  wire [7:0] sel_794797;
  wire [7:0] add_794800;
  wire [7:0] sel_794801;
  wire [7:0] add_794804;
  wire [7:0] sel_794805;
  wire [7:0] add_794808;
  wire [7:0] sel_794809;
  wire [7:0] add_794812;
  wire [7:0] sel_794813;
  wire [7:0] add_794816;
  wire [7:0] sel_794817;
  wire [7:0] add_794820;
  wire [7:0] sel_794821;
  wire [7:0] add_794824;
  wire [7:0] sel_794825;
  wire [7:0] add_794828;
  wire [7:0] sel_794829;
  wire [7:0] add_794832;
  wire [7:0] sel_794833;
  wire [7:0] add_794836;
  wire [7:0] sel_794837;
  wire [7:0] add_794840;
  wire [7:0] sel_794841;
  wire [7:0] add_794844;
  wire [7:0] sel_794845;
  wire [7:0] add_794848;
  wire [7:0] sel_794849;
  wire [7:0] add_794852;
  wire [7:0] sel_794853;
  wire [7:0] add_794856;
  wire [7:0] sel_794857;
  wire [7:0] add_794860;
  wire [7:0] sel_794861;
  wire [7:0] add_794864;
  wire [7:0] sel_794865;
  wire [7:0] add_794868;
  wire [7:0] sel_794869;
  wire [7:0] add_794872;
  wire [7:0] sel_794873;
  wire [7:0] add_794876;
  wire [7:0] sel_794877;
  wire [7:0] add_794880;
  wire [7:0] sel_794881;
  wire [7:0] add_794884;
  wire [7:0] sel_794885;
  wire [7:0] add_794888;
  wire [7:0] sel_794889;
  wire [7:0] add_794892;
  wire [7:0] sel_794893;
  wire [7:0] add_794896;
  wire [7:0] sel_794897;
  wire [7:0] add_794901;
  wire [15:0] array_index_794902;
  wire [7:0] sel_794903;
  wire [7:0] add_794906;
  wire [7:0] sel_794907;
  wire [7:0] add_794910;
  wire [7:0] sel_794911;
  wire [7:0] add_794914;
  wire [7:0] sel_794915;
  wire [7:0] add_794918;
  wire [7:0] sel_794919;
  wire [7:0] add_794922;
  wire [7:0] sel_794923;
  wire [7:0] add_794926;
  wire [7:0] sel_794927;
  wire [7:0] add_794930;
  wire [7:0] sel_794931;
  wire [7:0] add_794934;
  wire [7:0] sel_794935;
  wire [7:0] add_794938;
  wire [7:0] sel_794939;
  wire [7:0] add_794942;
  wire [7:0] sel_794943;
  wire [7:0] add_794946;
  wire [7:0] sel_794947;
  wire [7:0] add_794950;
  wire [7:0] sel_794951;
  wire [7:0] add_794954;
  wire [7:0] sel_794955;
  wire [7:0] add_794958;
  wire [7:0] sel_794959;
  wire [7:0] add_794962;
  wire [7:0] sel_794963;
  wire [7:0] add_794966;
  wire [7:0] sel_794967;
  wire [7:0] add_794970;
  wire [7:0] sel_794971;
  wire [7:0] add_794974;
  wire [7:0] sel_794975;
  wire [7:0] add_794978;
  wire [7:0] sel_794979;
  wire [7:0] add_794982;
  wire [7:0] sel_794983;
  wire [7:0] add_794986;
  wire [7:0] sel_794987;
  wire [7:0] add_794990;
  wire [7:0] sel_794991;
  wire [7:0] add_794994;
  wire [7:0] sel_794995;
  wire [7:0] add_794998;
  wire [7:0] sel_794999;
  wire [7:0] add_795002;
  wire [7:0] sel_795003;
  wire [7:0] add_795006;
  wire [7:0] sel_795007;
  wire [7:0] add_795010;
  wire [7:0] sel_795011;
  wire [7:0] add_795014;
  wire [7:0] sel_795015;
  wire [7:0] add_795018;
  wire [7:0] sel_795019;
  wire [7:0] add_795022;
  wire [7:0] sel_795023;
  wire [7:0] add_795026;
  wire [7:0] sel_795027;
  wire [7:0] add_795030;
  wire [7:0] sel_795031;
  wire [7:0] add_795034;
  wire [7:0] sel_795035;
  wire [7:0] add_795038;
  wire [7:0] sel_795039;
  wire [7:0] add_795042;
  wire [7:0] sel_795043;
  wire [7:0] add_795046;
  wire [7:0] sel_795047;
  wire [7:0] add_795050;
  wire [7:0] sel_795051;
  wire [7:0] add_795054;
  wire [7:0] sel_795055;
  wire [7:0] add_795058;
  wire [7:0] sel_795059;
  wire [7:0] add_795062;
  wire [7:0] sel_795063;
  wire [7:0] add_795066;
  wire [7:0] sel_795067;
  wire [7:0] add_795070;
  wire [7:0] sel_795071;
  wire [7:0] add_795074;
  wire [7:0] sel_795075;
  wire [7:0] add_795078;
  wire [7:0] sel_795079;
  wire [7:0] add_795082;
  wire [7:0] sel_795083;
  wire [7:0] add_795086;
  wire [7:0] sel_795087;
  wire [7:0] add_795090;
  wire [7:0] sel_795091;
  wire [7:0] add_795094;
  wire [7:0] sel_795095;
  wire [7:0] add_795098;
  wire [7:0] sel_795099;
  wire [7:0] add_795102;
  wire [7:0] sel_795103;
  wire [7:0] add_795106;
  wire [7:0] sel_795107;
  wire [7:0] add_795110;
  wire [7:0] sel_795111;
  wire [7:0] add_795114;
  wire [7:0] sel_795115;
  wire [7:0] add_795118;
  wire [7:0] sel_795119;
  wire [7:0] add_795122;
  wire [7:0] sel_795123;
  wire [7:0] add_795126;
  wire [7:0] sel_795127;
  wire [7:0] add_795130;
  wire [7:0] sel_795131;
  wire [7:0] add_795134;
  wire [7:0] sel_795135;
  wire [7:0] add_795138;
  wire [7:0] sel_795139;
  wire [7:0] add_795142;
  wire [7:0] sel_795143;
  wire [7:0] add_795146;
  wire [7:0] sel_795147;
  wire [7:0] add_795150;
  wire [7:0] sel_795151;
  wire [7:0] add_795154;
  wire [7:0] sel_795155;
  wire [7:0] add_795158;
  wire [7:0] sel_795159;
  wire [7:0] add_795162;
  wire [7:0] sel_795163;
  wire [7:0] add_795166;
  wire [7:0] sel_795167;
  wire [7:0] add_795170;
  wire [7:0] sel_795171;
  wire [7:0] add_795174;
  wire [7:0] sel_795175;
  wire [7:0] add_795178;
  wire [7:0] sel_795179;
  wire [7:0] add_795182;
  wire [7:0] sel_795183;
  wire [7:0] add_795186;
  wire [7:0] sel_795187;
  wire [7:0] add_795190;
  wire [7:0] sel_795191;
  wire [7:0] add_795194;
  wire [7:0] sel_795195;
  wire [7:0] add_795198;
  wire [7:0] sel_795199;
  wire [7:0] add_795202;
  wire [7:0] sel_795203;
  wire [7:0] add_795206;
  wire [7:0] sel_795207;
  wire [7:0] add_795210;
  wire [7:0] sel_795211;
  wire [7:0] add_795214;
  wire [7:0] sel_795215;
  wire [7:0] add_795218;
  wire [7:0] sel_795219;
  wire [7:0] add_795222;
  wire [7:0] sel_795223;
  wire [7:0] add_795226;
  wire [7:0] sel_795227;
  wire [7:0] add_795230;
  wire [7:0] sel_795231;
  wire [7:0] add_795234;
  wire [7:0] sel_795235;
  wire [7:0] add_795238;
  wire [7:0] sel_795239;
  wire [7:0] add_795242;
  wire [7:0] sel_795243;
  wire [7:0] add_795246;
  wire [7:0] sel_795247;
  wire [7:0] add_795250;
  wire [7:0] sel_795251;
  wire [7:0] add_795254;
  wire [7:0] sel_795255;
  wire [7:0] add_795258;
  wire [7:0] sel_795259;
  wire [7:0] add_795263;
  wire [15:0] array_index_795264;
  wire [7:0] sel_795265;
  wire [7:0] add_795268;
  wire [7:0] sel_795269;
  wire [7:0] add_795272;
  wire [7:0] sel_795273;
  wire [7:0] add_795276;
  wire [7:0] sel_795277;
  wire [7:0] add_795280;
  wire [7:0] sel_795281;
  wire [7:0] add_795284;
  wire [7:0] sel_795285;
  wire [7:0] add_795288;
  wire [7:0] sel_795289;
  wire [7:0] add_795292;
  wire [7:0] sel_795293;
  wire [7:0] add_795296;
  wire [7:0] sel_795297;
  wire [7:0] add_795300;
  wire [7:0] sel_795301;
  wire [7:0] add_795304;
  wire [7:0] sel_795305;
  wire [7:0] add_795308;
  wire [7:0] sel_795309;
  wire [7:0] add_795312;
  wire [7:0] sel_795313;
  wire [7:0] add_795316;
  wire [7:0] sel_795317;
  wire [7:0] add_795320;
  wire [7:0] sel_795321;
  wire [7:0] add_795324;
  wire [7:0] sel_795325;
  wire [7:0] add_795328;
  wire [7:0] sel_795329;
  wire [7:0] add_795332;
  wire [7:0] sel_795333;
  wire [7:0] add_795336;
  wire [7:0] sel_795337;
  wire [7:0] add_795340;
  wire [7:0] sel_795341;
  wire [7:0] add_795344;
  wire [7:0] sel_795345;
  wire [7:0] add_795348;
  wire [7:0] sel_795349;
  wire [7:0] add_795352;
  wire [7:0] sel_795353;
  wire [7:0] add_795356;
  wire [7:0] sel_795357;
  wire [7:0] add_795360;
  wire [7:0] sel_795361;
  wire [7:0] add_795364;
  wire [7:0] sel_795365;
  wire [7:0] add_795368;
  wire [7:0] sel_795369;
  wire [7:0] add_795372;
  wire [7:0] sel_795373;
  wire [7:0] add_795376;
  wire [7:0] sel_795377;
  wire [7:0] add_795380;
  wire [7:0] sel_795381;
  wire [7:0] add_795384;
  wire [7:0] sel_795385;
  wire [7:0] add_795388;
  wire [7:0] sel_795389;
  wire [7:0] add_795392;
  wire [7:0] sel_795393;
  wire [7:0] add_795396;
  wire [7:0] sel_795397;
  wire [7:0] add_795400;
  wire [7:0] sel_795401;
  wire [7:0] add_795404;
  wire [7:0] sel_795405;
  wire [7:0] add_795408;
  wire [7:0] sel_795409;
  wire [7:0] add_795412;
  wire [7:0] sel_795413;
  wire [7:0] add_795416;
  wire [7:0] sel_795417;
  wire [7:0] add_795420;
  wire [7:0] sel_795421;
  wire [7:0] add_795424;
  wire [7:0] sel_795425;
  wire [7:0] add_795428;
  wire [7:0] sel_795429;
  wire [7:0] add_795432;
  wire [7:0] sel_795433;
  wire [7:0] add_795436;
  wire [7:0] sel_795437;
  wire [7:0] add_795440;
  wire [7:0] sel_795441;
  wire [7:0] add_795444;
  wire [7:0] sel_795445;
  wire [7:0] add_795448;
  wire [7:0] sel_795449;
  wire [7:0] add_795452;
  wire [7:0] sel_795453;
  wire [7:0] add_795456;
  wire [7:0] sel_795457;
  wire [7:0] add_795460;
  wire [7:0] sel_795461;
  wire [7:0] add_795464;
  wire [7:0] sel_795465;
  wire [7:0] add_795468;
  wire [7:0] sel_795469;
  wire [7:0] add_795472;
  wire [7:0] sel_795473;
  wire [7:0] add_795476;
  wire [7:0] sel_795477;
  wire [7:0] add_795480;
  wire [7:0] sel_795481;
  wire [7:0] add_795484;
  wire [7:0] sel_795485;
  wire [7:0] add_795488;
  wire [7:0] sel_795489;
  wire [7:0] add_795492;
  wire [7:0] sel_795493;
  wire [7:0] add_795496;
  wire [7:0] sel_795497;
  wire [7:0] add_795500;
  wire [7:0] sel_795501;
  wire [7:0] add_795504;
  wire [7:0] sel_795505;
  wire [7:0] add_795508;
  wire [7:0] sel_795509;
  wire [7:0] add_795512;
  wire [7:0] sel_795513;
  wire [7:0] add_795516;
  wire [7:0] sel_795517;
  wire [7:0] add_795520;
  wire [7:0] sel_795521;
  wire [7:0] add_795524;
  wire [7:0] sel_795525;
  wire [7:0] add_795528;
  wire [7:0] sel_795529;
  wire [7:0] add_795532;
  wire [7:0] sel_795533;
  wire [7:0] add_795536;
  wire [7:0] sel_795537;
  wire [7:0] add_795540;
  wire [7:0] sel_795541;
  wire [7:0] add_795544;
  wire [7:0] sel_795545;
  wire [7:0] add_795548;
  wire [7:0] sel_795549;
  wire [7:0] add_795552;
  wire [7:0] sel_795553;
  wire [7:0] add_795556;
  wire [7:0] sel_795557;
  wire [7:0] add_795560;
  wire [7:0] sel_795561;
  wire [7:0] add_795564;
  wire [7:0] sel_795565;
  wire [7:0] add_795568;
  wire [7:0] sel_795569;
  wire [7:0] add_795572;
  wire [7:0] sel_795573;
  wire [7:0] add_795576;
  wire [7:0] sel_795577;
  wire [7:0] add_795580;
  wire [7:0] sel_795581;
  wire [7:0] add_795584;
  wire [7:0] sel_795585;
  wire [7:0] add_795588;
  wire [7:0] sel_795589;
  wire [7:0] add_795592;
  wire [7:0] sel_795593;
  wire [7:0] add_795596;
  wire [7:0] sel_795597;
  wire [7:0] add_795600;
  wire [7:0] sel_795601;
  wire [7:0] add_795604;
  wire [7:0] sel_795605;
  wire [7:0] add_795608;
  wire [7:0] sel_795609;
  wire [7:0] add_795612;
  wire [7:0] sel_795613;
  wire [7:0] add_795616;
  wire [7:0] sel_795617;
  wire [7:0] add_795620;
  wire [7:0] sel_795621;
  wire [7:0] add_795625;
  wire [15:0] array_index_795626;
  wire [7:0] sel_795627;
  wire [7:0] add_795630;
  wire [7:0] sel_795631;
  wire [7:0] add_795634;
  wire [7:0] sel_795635;
  wire [7:0] add_795638;
  wire [7:0] sel_795639;
  wire [7:0] add_795642;
  wire [7:0] sel_795643;
  wire [7:0] add_795646;
  wire [7:0] sel_795647;
  wire [7:0] add_795650;
  wire [7:0] sel_795651;
  wire [7:0] add_795654;
  wire [7:0] sel_795655;
  wire [7:0] add_795658;
  wire [7:0] sel_795659;
  wire [7:0] add_795662;
  wire [7:0] sel_795663;
  wire [7:0] add_795666;
  wire [7:0] sel_795667;
  wire [7:0] add_795670;
  wire [7:0] sel_795671;
  wire [7:0] add_795674;
  wire [7:0] sel_795675;
  wire [7:0] add_795678;
  wire [7:0] sel_795679;
  wire [7:0] add_795682;
  wire [7:0] sel_795683;
  wire [7:0] add_795686;
  wire [7:0] sel_795687;
  wire [7:0] add_795690;
  wire [7:0] sel_795691;
  wire [7:0] add_795694;
  wire [7:0] sel_795695;
  wire [7:0] add_795698;
  wire [7:0] sel_795699;
  wire [7:0] add_795702;
  wire [7:0] sel_795703;
  wire [7:0] add_795706;
  wire [7:0] sel_795707;
  wire [7:0] add_795710;
  wire [7:0] sel_795711;
  wire [7:0] add_795714;
  wire [7:0] sel_795715;
  wire [7:0] add_795718;
  wire [7:0] sel_795719;
  wire [7:0] add_795722;
  wire [7:0] sel_795723;
  wire [7:0] add_795726;
  wire [7:0] sel_795727;
  wire [7:0] add_795730;
  wire [7:0] sel_795731;
  wire [7:0] add_795734;
  wire [7:0] sel_795735;
  wire [7:0] add_795738;
  wire [7:0] sel_795739;
  wire [7:0] add_795742;
  wire [7:0] sel_795743;
  wire [7:0] add_795746;
  wire [7:0] sel_795747;
  wire [7:0] add_795750;
  wire [7:0] sel_795751;
  wire [7:0] add_795754;
  wire [7:0] sel_795755;
  wire [7:0] add_795758;
  wire [7:0] sel_795759;
  wire [7:0] add_795762;
  wire [7:0] sel_795763;
  wire [7:0] add_795766;
  wire [7:0] sel_795767;
  wire [7:0] add_795770;
  wire [7:0] sel_795771;
  wire [7:0] add_795774;
  wire [7:0] sel_795775;
  wire [7:0] add_795778;
  wire [7:0] sel_795779;
  wire [7:0] add_795782;
  wire [7:0] sel_795783;
  wire [7:0] add_795786;
  wire [7:0] sel_795787;
  wire [7:0] add_795790;
  wire [7:0] sel_795791;
  wire [7:0] add_795794;
  wire [7:0] sel_795795;
  wire [7:0] add_795798;
  wire [7:0] sel_795799;
  wire [7:0] add_795802;
  wire [7:0] sel_795803;
  wire [7:0] add_795806;
  wire [7:0] sel_795807;
  wire [7:0] add_795810;
  wire [7:0] sel_795811;
  wire [7:0] add_795814;
  wire [7:0] sel_795815;
  wire [7:0] add_795818;
  wire [7:0] sel_795819;
  wire [7:0] add_795822;
  wire [7:0] sel_795823;
  wire [7:0] add_795826;
  wire [7:0] sel_795827;
  wire [7:0] add_795830;
  wire [7:0] sel_795831;
  wire [7:0] add_795834;
  wire [7:0] sel_795835;
  wire [7:0] add_795838;
  wire [7:0] sel_795839;
  wire [7:0] add_795842;
  wire [7:0] sel_795843;
  wire [7:0] add_795846;
  wire [7:0] sel_795847;
  wire [7:0] add_795850;
  wire [7:0] sel_795851;
  wire [7:0] add_795854;
  wire [7:0] sel_795855;
  wire [7:0] add_795858;
  wire [7:0] sel_795859;
  wire [7:0] add_795862;
  wire [7:0] sel_795863;
  wire [7:0] add_795866;
  wire [7:0] sel_795867;
  wire [7:0] add_795870;
  wire [7:0] sel_795871;
  wire [7:0] add_795874;
  wire [7:0] sel_795875;
  wire [7:0] add_795878;
  wire [7:0] sel_795879;
  wire [7:0] add_795882;
  wire [7:0] sel_795883;
  wire [7:0] add_795886;
  wire [7:0] sel_795887;
  wire [7:0] add_795890;
  wire [7:0] sel_795891;
  wire [7:0] add_795894;
  wire [7:0] sel_795895;
  wire [7:0] add_795898;
  wire [7:0] sel_795899;
  wire [7:0] add_795902;
  wire [7:0] sel_795903;
  wire [7:0] add_795906;
  wire [7:0] sel_795907;
  wire [7:0] add_795910;
  wire [7:0] sel_795911;
  wire [7:0] add_795914;
  wire [7:0] sel_795915;
  wire [7:0] add_795918;
  wire [7:0] sel_795919;
  wire [7:0] add_795922;
  wire [7:0] sel_795923;
  wire [7:0] add_795926;
  wire [7:0] sel_795927;
  wire [7:0] add_795930;
  wire [7:0] sel_795931;
  wire [7:0] add_795934;
  wire [7:0] sel_795935;
  wire [7:0] add_795938;
  wire [7:0] sel_795939;
  wire [7:0] add_795942;
  wire [7:0] sel_795943;
  wire [7:0] add_795946;
  wire [7:0] sel_795947;
  wire [7:0] add_795950;
  wire [7:0] sel_795951;
  wire [7:0] add_795954;
  wire [7:0] sel_795955;
  wire [7:0] add_795958;
  wire [7:0] sel_795959;
  wire [7:0] add_795962;
  wire [7:0] sel_795963;
  wire [7:0] add_795966;
  wire [7:0] sel_795967;
  wire [7:0] add_795970;
  wire [7:0] sel_795971;
  wire [7:0] add_795974;
  wire [7:0] sel_795975;
  wire [7:0] add_795978;
  wire [7:0] sel_795979;
  wire [7:0] add_795982;
  wire [7:0] sel_795983;
  wire [7:0] add_795987;
  wire [15:0] array_index_795988;
  wire [7:0] sel_795989;
  wire [7:0] add_795992;
  wire [7:0] sel_795993;
  wire [7:0] add_795996;
  wire [7:0] sel_795997;
  wire [7:0] add_796000;
  wire [7:0] sel_796001;
  wire [7:0] add_796004;
  wire [7:0] sel_796005;
  wire [7:0] add_796008;
  wire [7:0] sel_796009;
  wire [7:0] add_796012;
  wire [7:0] sel_796013;
  wire [7:0] add_796016;
  wire [7:0] sel_796017;
  wire [7:0] add_796020;
  wire [7:0] sel_796021;
  wire [7:0] add_796024;
  wire [7:0] sel_796025;
  wire [7:0] add_796028;
  wire [7:0] sel_796029;
  wire [7:0] add_796032;
  wire [7:0] sel_796033;
  wire [7:0] add_796036;
  wire [7:0] sel_796037;
  wire [7:0] add_796040;
  wire [7:0] sel_796041;
  wire [7:0] add_796044;
  wire [7:0] sel_796045;
  wire [7:0] add_796048;
  wire [7:0] sel_796049;
  wire [7:0] add_796052;
  wire [7:0] sel_796053;
  wire [7:0] add_796056;
  wire [7:0] sel_796057;
  wire [7:0] add_796060;
  wire [7:0] sel_796061;
  wire [7:0] add_796064;
  wire [7:0] sel_796065;
  wire [7:0] add_796068;
  wire [7:0] sel_796069;
  wire [7:0] add_796072;
  wire [7:0] sel_796073;
  wire [7:0] add_796076;
  wire [7:0] sel_796077;
  wire [7:0] add_796080;
  wire [7:0] sel_796081;
  wire [7:0] add_796084;
  wire [7:0] sel_796085;
  wire [7:0] add_796088;
  wire [7:0] sel_796089;
  wire [7:0] add_796092;
  wire [7:0] sel_796093;
  wire [7:0] add_796096;
  wire [7:0] sel_796097;
  wire [7:0] add_796100;
  wire [7:0] sel_796101;
  wire [7:0] add_796104;
  wire [7:0] sel_796105;
  wire [7:0] add_796108;
  wire [7:0] sel_796109;
  wire [7:0] add_796112;
  wire [7:0] sel_796113;
  wire [7:0] add_796116;
  wire [7:0] sel_796117;
  wire [7:0] add_796120;
  wire [7:0] sel_796121;
  wire [7:0] add_796124;
  wire [7:0] sel_796125;
  wire [7:0] add_796128;
  wire [7:0] sel_796129;
  wire [7:0] add_796132;
  wire [7:0] sel_796133;
  wire [7:0] add_796136;
  wire [7:0] sel_796137;
  wire [7:0] add_796140;
  wire [7:0] sel_796141;
  wire [7:0] add_796144;
  wire [7:0] sel_796145;
  wire [7:0] add_796148;
  wire [7:0] sel_796149;
  wire [7:0] add_796152;
  wire [7:0] sel_796153;
  wire [7:0] add_796156;
  wire [7:0] sel_796157;
  wire [7:0] add_796160;
  wire [7:0] sel_796161;
  wire [7:0] add_796164;
  wire [7:0] sel_796165;
  wire [7:0] add_796168;
  wire [7:0] sel_796169;
  wire [7:0] add_796172;
  wire [7:0] sel_796173;
  wire [7:0] add_796176;
  wire [7:0] sel_796177;
  wire [7:0] add_796180;
  wire [7:0] sel_796181;
  wire [7:0] add_796184;
  wire [7:0] sel_796185;
  wire [7:0] add_796188;
  wire [7:0] sel_796189;
  wire [7:0] add_796192;
  wire [7:0] sel_796193;
  wire [7:0] add_796196;
  wire [7:0] sel_796197;
  wire [7:0] add_796200;
  wire [7:0] sel_796201;
  wire [7:0] add_796204;
  wire [7:0] sel_796205;
  wire [7:0] add_796208;
  wire [7:0] sel_796209;
  wire [7:0] add_796212;
  wire [7:0] sel_796213;
  wire [7:0] add_796216;
  wire [7:0] sel_796217;
  wire [7:0] add_796220;
  wire [7:0] sel_796221;
  wire [7:0] add_796224;
  wire [7:0] sel_796225;
  wire [7:0] add_796228;
  wire [7:0] sel_796229;
  wire [7:0] add_796232;
  wire [7:0] sel_796233;
  wire [7:0] add_796236;
  wire [7:0] sel_796237;
  wire [7:0] add_796240;
  wire [7:0] sel_796241;
  wire [7:0] add_796244;
  wire [7:0] sel_796245;
  wire [7:0] add_796248;
  wire [7:0] sel_796249;
  wire [7:0] add_796252;
  wire [7:0] sel_796253;
  wire [7:0] add_796256;
  wire [7:0] sel_796257;
  wire [7:0] add_796260;
  wire [7:0] sel_796261;
  wire [7:0] add_796264;
  wire [7:0] sel_796265;
  wire [7:0] add_796268;
  wire [7:0] sel_796269;
  wire [7:0] add_796272;
  wire [7:0] sel_796273;
  wire [7:0] add_796276;
  wire [7:0] sel_796277;
  wire [7:0] add_796280;
  wire [7:0] sel_796281;
  wire [7:0] add_796284;
  wire [7:0] sel_796285;
  wire [7:0] add_796288;
  wire [7:0] sel_796289;
  wire [7:0] add_796292;
  wire [7:0] sel_796293;
  wire [7:0] add_796296;
  wire [7:0] sel_796297;
  wire [7:0] add_796300;
  wire [7:0] sel_796301;
  wire [7:0] add_796304;
  wire [7:0] sel_796305;
  wire [7:0] add_796308;
  wire [7:0] sel_796309;
  wire [7:0] add_796312;
  wire [7:0] sel_796313;
  wire [7:0] add_796316;
  wire [7:0] sel_796317;
  wire [7:0] add_796320;
  wire [7:0] sel_796321;
  wire [7:0] add_796324;
  wire [7:0] sel_796325;
  wire [7:0] add_796328;
  wire [7:0] sel_796329;
  wire [7:0] add_796332;
  wire [7:0] sel_796333;
  wire [7:0] add_796336;
  wire [7:0] sel_796337;
  wire [7:0] add_796340;
  wire [7:0] sel_796341;
  wire [7:0] add_796344;
  wire [7:0] sel_796345;
  wire [7:0] add_796349;
  wire [15:0] array_index_796350;
  wire [7:0] sel_796351;
  wire [7:0] add_796354;
  wire [7:0] sel_796355;
  wire [7:0] add_796358;
  wire [7:0] sel_796359;
  wire [7:0] add_796362;
  wire [7:0] sel_796363;
  wire [7:0] add_796366;
  wire [7:0] sel_796367;
  wire [7:0] add_796370;
  wire [7:0] sel_796371;
  wire [7:0] add_796374;
  wire [7:0] sel_796375;
  wire [7:0] add_796378;
  wire [7:0] sel_796379;
  wire [7:0] add_796382;
  wire [7:0] sel_796383;
  wire [7:0] add_796386;
  wire [7:0] sel_796387;
  wire [7:0] add_796390;
  wire [7:0] sel_796391;
  wire [7:0] add_796394;
  wire [7:0] sel_796395;
  wire [7:0] add_796398;
  wire [7:0] sel_796399;
  wire [7:0] add_796402;
  wire [7:0] sel_796403;
  wire [7:0] add_796406;
  wire [7:0] sel_796407;
  wire [7:0] add_796410;
  wire [7:0] sel_796411;
  wire [7:0] add_796414;
  wire [7:0] sel_796415;
  wire [7:0] add_796418;
  wire [7:0] sel_796419;
  wire [7:0] add_796422;
  wire [7:0] sel_796423;
  wire [7:0] add_796426;
  wire [7:0] sel_796427;
  wire [7:0] add_796430;
  wire [7:0] sel_796431;
  wire [7:0] add_796434;
  wire [7:0] sel_796435;
  wire [7:0] add_796438;
  wire [7:0] sel_796439;
  wire [7:0] add_796442;
  wire [7:0] sel_796443;
  wire [7:0] add_796446;
  wire [7:0] sel_796447;
  wire [7:0] add_796450;
  wire [7:0] sel_796451;
  wire [7:0] add_796454;
  wire [7:0] sel_796455;
  wire [7:0] add_796458;
  wire [7:0] sel_796459;
  wire [7:0] add_796462;
  wire [7:0] sel_796463;
  wire [7:0] add_796466;
  wire [7:0] sel_796467;
  wire [7:0] add_796470;
  wire [7:0] sel_796471;
  wire [7:0] add_796474;
  wire [7:0] sel_796475;
  wire [7:0] add_796478;
  wire [7:0] sel_796479;
  wire [7:0] add_796482;
  wire [7:0] sel_796483;
  wire [7:0] add_796486;
  wire [7:0] sel_796487;
  wire [7:0] add_796490;
  wire [7:0] sel_796491;
  wire [7:0] add_796494;
  wire [7:0] sel_796495;
  wire [7:0] add_796498;
  wire [7:0] sel_796499;
  wire [7:0] add_796502;
  wire [7:0] sel_796503;
  wire [7:0] add_796506;
  wire [7:0] sel_796507;
  wire [7:0] add_796510;
  wire [7:0] sel_796511;
  wire [7:0] add_796514;
  wire [7:0] sel_796515;
  wire [7:0] add_796518;
  wire [7:0] sel_796519;
  wire [7:0] add_796522;
  wire [7:0] sel_796523;
  wire [7:0] add_796526;
  wire [7:0] sel_796527;
  wire [7:0] add_796530;
  wire [7:0] sel_796531;
  wire [7:0] add_796534;
  wire [7:0] sel_796535;
  wire [7:0] add_796538;
  wire [7:0] sel_796539;
  wire [7:0] add_796542;
  wire [7:0] sel_796543;
  wire [7:0] add_796546;
  wire [7:0] sel_796547;
  wire [7:0] add_796550;
  wire [7:0] sel_796551;
  wire [7:0] add_796554;
  wire [7:0] sel_796555;
  wire [7:0] add_796558;
  wire [7:0] sel_796559;
  wire [7:0] add_796562;
  wire [7:0] sel_796563;
  wire [7:0] add_796566;
  wire [7:0] sel_796567;
  wire [7:0] add_796570;
  wire [7:0] sel_796571;
  wire [7:0] add_796574;
  wire [7:0] sel_796575;
  wire [7:0] add_796578;
  wire [7:0] sel_796579;
  wire [7:0] add_796582;
  wire [7:0] sel_796583;
  wire [7:0] add_796586;
  wire [7:0] sel_796587;
  wire [7:0] add_796590;
  wire [7:0] sel_796591;
  wire [7:0] add_796594;
  wire [7:0] sel_796595;
  wire [7:0] add_796598;
  wire [7:0] sel_796599;
  wire [7:0] add_796602;
  wire [7:0] sel_796603;
  wire [7:0] add_796606;
  wire [7:0] sel_796607;
  wire [7:0] add_796610;
  wire [7:0] sel_796611;
  wire [7:0] add_796614;
  wire [7:0] sel_796615;
  wire [7:0] add_796618;
  wire [7:0] sel_796619;
  wire [7:0] add_796622;
  wire [7:0] sel_796623;
  wire [7:0] add_796626;
  wire [7:0] sel_796627;
  wire [7:0] add_796630;
  wire [7:0] sel_796631;
  wire [7:0] add_796634;
  wire [7:0] sel_796635;
  wire [7:0] add_796638;
  wire [7:0] sel_796639;
  wire [7:0] add_796642;
  wire [7:0] sel_796643;
  wire [7:0] add_796646;
  wire [7:0] sel_796647;
  wire [7:0] add_796650;
  wire [7:0] sel_796651;
  wire [7:0] add_796654;
  wire [7:0] sel_796655;
  wire [7:0] add_796658;
  wire [7:0] sel_796659;
  wire [7:0] add_796662;
  wire [7:0] sel_796663;
  wire [7:0] add_796666;
  wire [7:0] sel_796667;
  wire [7:0] add_796670;
  wire [7:0] sel_796671;
  wire [7:0] add_796674;
  wire [7:0] sel_796675;
  wire [7:0] add_796678;
  wire [7:0] sel_796679;
  wire [7:0] add_796682;
  wire [7:0] sel_796683;
  wire [7:0] add_796686;
  wire [7:0] sel_796687;
  wire [7:0] add_796690;
  wire [7:0] sel_796691;
  wire [7:0] add_796694;
  wire [7:0] sel_796695;
  wire [7:0] add_796698;
  wire [7:0] sel_796699;
  wire [7:0] add_796702;
  wire [7:0] sel_796703;
  wire [7:0] add_796706;
  wire [7:0] sel_796707;
  wire [7:0] add_796711;
  wire [15:0] array_index_796712;
  wire [7:0] sel_796713;
  wire [7:0] add_796716;
  wire [7:0] sel_796717;
  wire [7:0] add_796720;
  wire [7:0] sel_796721;
  wire [7:0] add_796724;
  wire [7:0] sel_796725;
  wire [7:0] add_796728;
  wire [7:0] sel_796729;
  wire [7:0] add_796732;
  wire [7:0] sel_796733;
  wire [7:0] add_796736;
  wire [7:0] sel_796737;
  wire [7:0] add_796740;
  wire [7:0] sel_796741;
  wire [7:0] add_796744;
  wire [7:0] sel_796745;
  wire [7:0] add_796748;
  wire [7:0] sel_796749;
  wire [7:0] add_796752;
  wire [7:0] sel_796753;
  wire [7:0] add_796756;
  wire [7:0] sel_796757;
  wire [7:0] add_796760;
  wire [7:0] sel_796761;
  wire [7:0] add_796764;
  wire [7:0] sel_796765;
  wire [7:0] add_796768;
  wire [7:0] sel_796769;
  wire [7:0] add_796772;
  wire [7:0] sel_796773;
  wire [7:0] add_796776;
  wire [7:0] sel_796777;
  wire [7:0] add_796780;
  wire [7:0] sel_796781;
  wire [7:0] add_796784;
  wire [7:0] sel_796785;
  wire [7:0] add_796788;
  wire [7:0] sel_796789;
  wire [7:0] add_796792;
  wire [7:0] sel_796793;
  wire [7:0] add_796796;
  wire [7:0] sel_796797;
  wire [7:0] add_796800;
  wire [7:0] sel_796801;
  wire [7:0] add_796804;
  wire [7:0] sel_796805;
  wire [7:0] add_796808;
  wire [7:0] sel_796809;
  wire [7:0] add_796812;
  wire [7:0] sel_796813;
  wire [7:0] add_796816;
  wire [7:0] sel_796817;
  wire [7:0] add_796820;
  wire [7:0] sel_796821;
  wire [7:0] add_796824;
  wire [7:0] sel_796825;
  wire [7:0] add_796828;
  wire [7:0] sel_796829;
  wire [7:0] add_796832;
  wire [7:0] sel_796833;
  wire [7:0] add_796836;
  wire [7:0] sel_796837;
  wire [7:0] add_796840;
  wire [7:0] sel_796841;
  wire [7:0] add_796844;
  wire [7:0] sel_796845;
  wire [7:0] add_796848;
  wire [7:0] sel_796849;
  wire [7:0] add_796852;
  wire [7:0] sel_796853;
  wire [7:0] add_796856;
  wire [7:0] sel_796857;
  wire [7:0] add_796860;
  wire [7:0] sel_796861;
  wire [7:0] add_796864;
  wire [7:0] sel_796865;
  wire [7:0] add_796868;
  wire [7:0] sel_796869;
  wire [7:0] add_796872;
  wire [7:0] sel_796873;
  wire [7:0] add_796876;
  wire [7:0] sel_796877;
  wire [7:0] add_796880;
  wire [7:0] sel_796881;
  wire [7:0] add_796884;
  wire [7:0] sel_796885;
  wire [7:0] add_796888;
  wire [7:0] sel_796889;
  wire [7:0] add_796892;
  wire [7:0] sel_796893;
  wire [7:0] add_796896;
  wire [7:0] sel_796897;
  wire [7:0] add_796900;
  wire [7:0] sel_796901;
  wire [7:0] add_796904;
  wire [7:0] sel_796905;
  wire [7:0] add_796908;
  wire [7:0] sel_796909;
  wire [7:0] add_796912;
  wire [7:0] sel_796913;
  wire [7:0] add_796916;
  wire [7:0] sel_796917;
  wire [7:0] add_796920;
  wire [7:0] sel_796921;
  wire [7:0] add_796924;
  wire [7:0] sel_796925;
  wire [7:0] add_796928;
  wire [7:0] sel_796929;
  wire [7:0] add_796932;
  wire [7:0] sel_796933;
  wire [7:0] add_796936;
  wire [7:0] sel_796937;
  wire [7:0] add_796940;
  wire [7:0] sel_796941;
  wire [7:0] add_796944;
  wire [7:0] sel_796945;
  wire [7:0] add_796948;
  wire [7:0] sel_796949;
  wire [7:0] add_796952;
  wire [7:0] sel_796953;
  wire [7:0] add_796956;
  wire [7:0] sel_796957;
  wire [7:0] add_796960;
  wire [7:0] sel_796961;
  wire [7:0] add_796964;
  wire [7:0] sel_796965;
  wire [7:0] add_796968;
  wire [7:0] sel_796969;
  wire [7:0] add_796972;
  wire [7:0] sel_796973;
  wire [7:0] add_796976;
  wire [7:0] sel_796977;
  wire [7:0] add_796980;
  wire [7:0] sel_796981;
  wire [7:0] add_796984;
  wire [7:0] sel_796985;
  wire [7:0] add_796988;
  wire [7:0] sel_796989;
  wire [7:0] add_796992;
  wire [7:0] sel_796993;
  wire [7:0] add_796996;
  wire [7:0] sel_796997;
  wire [7:0] add_797000;
  wire [7:0] sel_797001;
  wire [7:0] add_797004;
  wire [7:0] sel_797005;
  wire [7:0] add_797008;
  wire [7:0] sel_797009;
  wire [7:0] add_797012;
  wire [7:0] sel_797013;
  wire [7:0] add_797016;
  wire [7:0] sel_797017;
  wire [7:0] add_797020;
  wire [7:0] sel_797021;
  wire [7:0] add_797024;
  wire [7:0] sel_797025;
  wire [7:0] add_797028;
  wire [7:0] sel_797029;
  wire [7:0] add_797032;
  wire [7:0] sel_797033;
  wire [7:0] add_797036;
  wire [7:0] sel_797037;
  wire [7:0] add_797040;
  wire [7:0] sel_797041;
  wire [7:0] add_797044;
  wire [7:0] sel_797045;
  wire [7:0] add_797048;
  wire [7:0] sel_797049;
  wire [7:0] add_797052;
  wire [7:0] sel_797053;
  wire [7:0] add_797056;
  wire [7:0] sel_797057;
  wire [7:0] add_797060;
  wire [7:0] sel_797061;
  wire [7:0] add_797064;
  wire [7:0] sel_797065;
  wire [7:0] add_797068;
  wire [7:0] sel_797069;
  wire [7:0] add_797073;
  wire [15:0] array_index_797074;
  wire [7:0] sel_797075;
  wire [7:0] add_797078;
  wire [7:0] sel_797079;
  wire [7:0] add_797082;
  wire [7:0] sel_797083;
  wire [7:0] add_797086;
  wire [7:0] sel_797087;
  wire [7:0] add_797090;
  wire [7:0] sel_797091;
  wire [7:0] add_797094;
  wire [7:0] sel_797095;
  wire [7:0] add_797098;
  wire [7:0] sel_797099;
  wire [7:0] add_797102;
  wire [7:0] sel_797103;
  wire [7:0] add_797106;
  wire [7:0] sel_797107;
  wire [7:0] add_797110;
  wire [7:0] sel_797111;
  wire [7:0] add_797114;
  wire [7:0] sel_797115;
  wire [7:0] add_797118;
  wire [7:0] sel_797119;
  wire [7:0] add_797122;
  wire [7:0] sel_797123;
  wire [7:0] add_797126;
  wire [7:0] sel_797127;
  wire [7:0] add_797130;
  wire [7:0] sel_797131;
  wire [7:0] add_797134;
  wire [7:0] sel_797135;
  wire [7:0] add_797138;
  wire [7:0] sel_797139;
  wire [7:0] add_797142;
  wire [7:0] sel_797143;
  wire [7:0] add_797146;
  wire [7:0] sel_797147;
  wire [7:0] add_797150;
  wire [7:0] sel_797151;
  wire [7:0] add_797154;
  wire [7:0] sel_797155;
  wire [7:0] add_797158;
  wire [7:0] sel_797159;
  wire [7:0] add_797162;
  wire [7:0] sel_797163;
  wire [7:0] add_797166;
  wire [7:0] sel_797167;
  wire [7:0] add_797170;
  wire [7:0] sel_797171;
  wire [7:0] add_797174;
  wire [7:0] sel_797175;
  wire [7:0] add_797178;
  wire [7:0] sel_797179;
  wire [7:0] add_797182;
  wire [7:0] sel_797183;
  wire [7:0] add_797186;
  wire [7:0] sel_797187;
  wire [7:0] add_797190;
  wire [7:0] sel_797191;
  wire [7:0] add_797194;
  wire [7:0] sel_797195;
  wire [7:0] add_797198;
  wire [7:0] sel_797199;
  wire [7:0] add_797202;
  wire [7:0] sel_797203;
  wire [7:0] add_797206;
  wire [7:0] sel_797207;
  wire [7:0] add_797210;
  wire [7:0] sel_797211;
  wire [7:0] add_797214;
  wire [7:0] sel_797215;
  wire [7:0] add_797218;
  wire [7:0] sel_797219;
  wire [7:0] add_797222;
  wire [7:0] sel_797223;
  wire [7:0] add_797226;
  wire [7:0] sel_797227;
  wire [7:0] add_797230;
  wire [7:0] sel_797231;
  wire [7:0] add_797234;
  wire [7:0] sel_797235;
  wire [7:0] add_797238;
  wire [7:0] sel_797239;
  wire [7:0] add_797242;
  wire [7:0] sel_797243;
  wire [7:0] add_797246;
  wire [7:0] sel_797247;
  wire [7:0] add_797250;
  wire [7:0] sel_797251;
  wire [7:0] add_797254;
  wire [7:0] sel_797255;
  wire [7:0] add_797258;
  wire [7:0] sel_797259;
  wire [7:0] add_797262;
  wire [7:0] sel_797263;
  wire [7:0] add_797266;
  wire [7:0] sel_797267;
  wire [7:0] add_797270;
  wire [7:0] sel_797271;
  wire [7:0] add_797274;
  wire [7:0] sel_797275;
  wire [7:0] add_797278;
  wire [7:0] sel_797279;
  wire [7:0] add_797282;
  wire [7:0] sel_797283;
  wire [7:0] add_797286;
  wire [7:0] sel_797287;
  wire [7:0] add_797290;
  wire [7:0] sel_797291;
  wire [7:0] add_797294;
  wire [7:0] sel_797295;
  wire [7:0] add_797298;
  wire [7:0] sel_797299;
  wire [7:0] add_797302;
  wire [7:0] sel_797303;
  wire [7:0] add_797306;
  wire [7:0] sel_797307;
  wire [7:0] add_797310;
  wire [7:0] sel_797311;
  wire [7:0] add_797314;
  wire [7:0] sel_797315;
  wire [7:0] add_797318;
  wire [7:0] sel_797319;
  wire [7:0] add_797322;
  wire [7:0] sel_797323;
  wire [7:0] add_797326;
  wire [7:0] sel_797327;
  wire [7:0] add_797330;
  wire [7:0] sel_797331;
  wire [7:0] add_797334;
  wire [7:0] sel_797335;
  wire [7:0] add_797338;
  wire [7:0] sel_797339;
  wire [7:0] add_797342;
  wire [7:0] sel_797343;
  wire [7:0] add_797346;
  wire [7:0] sel_797347;
  wire [7:0] add_797350;
  wire [7:0] sel_797351;
  wire [7:0] add_797354;
  wire [7:0] sel_797355;
  wire [7:0] add_797358;
  wire [7:0] sel_797359;
  wire [7:0] add_797362;
  wire [7:0] sel_797363;
  wire [7:0] add_797366;
  wire [7:0] sel_797367;
  wire [7:0] add_797370;
  wire [7:0] sel_797371;
  wire [7:0] add_797374;
  wire [7:0] sel_797375;
  wire [7:0] add_797378;
  wire [7:0] sel_797379;
  wire [7:0] add_797382;
  wire [7:0] sel_797383;
  wire [7:0] add_797386;
  wire [7:0] sel_797387;
  wire [7:0] add_797390;
  wire [7:0] sel_797391;
  wire [7:0] add_797394;
  wire [7:0] sel_797395;
  wire [7:0] add_797398;
  wire [7:0] sel_797399;
  wire [7:0] add_797402;
  wire [7:0] sel_797403;
  wire [7:0] add_797406;
  wire [7:0] sel_797407;
  wire [7:0] add_797410;
  wire [7:0] sel_797411;
  wire [7:0] add_797414;
  wire [7:0] sel_797415;
  wire [7:0] add_797418;
  wire [7:0] sel_797419;
  wire [7:0] add_797422;
  wire [7:0] sel_797423;
  wire [7:0] add_797426;
  wire [7:0] sel_797427;
  wire [7:0] add_797430;
  wire [7:0] sel_797431;
  wire [7:0] add_797435;
  wire [15:0] array_index_797436;
  wire [7:0] sel_797437;
  wire [7:0] add_797440;
  wire [7:0] sel_797441;
  wire [7:0] add_797444;
  wire [7:0] sel_797445;
  wire [7:0] add_797448;
  wire [7:0] sel_797449;
  wire [7:0] add_797452;
  wire [7:0] sel_797453;
  wire [7:0] add_797456;
  wire [7:0] sel_797457;
  wire [7:0] add_797460;
  wire [7:0] sel_797461;
  wire [7:0] add_797464;
  wire [7:0] sel_797465;
  wire [7:0] add_797468;
  wire [7:0] sel_797469;
  wire [7:0] add_797472;
  wire [7:0] sel_797473;
  wire [7:0] add_797476;
  wire [7:0] sel_797477;
  wire [7:0] add_797480;
  wire [7:0] sel_797481;
  wire [7:0] add_797484;
  wire [7:0] sel_797485;
  wire [7:0] add_797488;
  wire [7:0] sel_797489;
  wire [7:0] add_797492;
  wire [7:0] sel_797493;
  wire [7:0] add_797496;
  wire [7:0] sel_797497;
  wire [7:0] add_797500;
  wire [7:0] sel_797501;
  wire [7:0] add_797504;
  wire [7:0] sel_797505;
  wire [7:0] add_797508;
  wire [7:0] sel_797509;
  wire [7:0] add_797512;
  wire [7:0] sel_797513;
  wire [7:0] add_797516;
  wire [7:0] sel_797517;
  wire [7:0] add_797520;
  wire [7:0] sel_797521;
  wire [7:0] add_797524;
  wire [7:0] sel_797525;
  wire [7:0] add_797528;
  wire [7:0] sel_797529;
  wire [7:0] add_797532;
  wire [7:0] sel_797533;
  wire [7:0] add_797536;
  wire [7:0] sel_797537;
  wire [7:0] add_797540;
  wire [7:0] sel_797541;
  wire [7:0] add_797544;
  wire [7:0] sel_797545;
  wire [7:0] add_797548;
  wire [7:0] sel_797549;
  wire [7:0] add_797552;
  wire [7:0] sel_797553;
  wire [7:0] add_797556;
  wire [7:0] sel_797557;
  wire [7:0] add_797560;
  wire [7:0] sel_797561;
  wire [7:0] add_797564;
  wire [7:0] sel_797565;
  wire [7:0] add_797568;
  wire [7:0] sel_797569;
  wire [7:0] add_797572;
  wire [7:0] sel_797573;
  wire [7:0] add_797576;
  wire [7:0] sel_797577;
  wire [7:0] add_797580;
  wire [7:0] sel_797581;
  wire [7:0] add_797584;
  wire [7:0] sel_797585;
  wire [7:0] add_797588;
  wire [7:0] sel_797589;
  wire [7:0] add_797592;
  wire [7:0] sel_797593;
  wire [7:0] add_797596;
  wire [7:0] sel_797597;
  wire [7:0] add_797600;
  wire [7:0] sel_797601;
  wire [7:0] add_797604;
  wire [7:0] sel_797605;
  wire [7:0] add_797608;
  wire [7:0] sel_797609;
  wire [7:0] add_797612;
  wire [7:0] sel_797613;
  wire [7:0] add_797616;
  wire [7:0] sel_797617;
  wire [7:0] add_797620;
  wire [7:0] sel_797621;
  wire [7:0] add_797624;
  wire [7:0] sel_797625;
  wire [7:0] add_797628;
  wire [7:0] sel_797629;
  wire [7:0] add_797632;
  wire [7:0] sel_797633;
  wire [7:0] add_797636;
  wire [7:0] sel_797637;
  wire [7:0] add_797640;
  wire [7:0] sel_797641;
  wire [7:0] add_797644;
  wire [7:0] sel_797645;
  wire [7:0] add_797648;
  wire [7:0] sel_797649;
  wire [7:0] add_797652;
  wire [7:0] sel_797653;
  wire [7:0] add_797656;
  wire [7:0] sel_797657;
  wire [7:0] add_797660;
  wire [7:0] sel_797661;
  wire [7:0] add_797664;
  wire [7:0] sel_797665;
  wire [7:0] add_797668;
  wire [7:0] sel_797669;
  wire [7:0] add_797672;
  wire [7:0] sel_797673;
  wire [7:0] add_797676;
  wire [7:0] sel_797677;
  wire [7:0] add_797680;
  wire [7:0] sel_797681;
  wire [7:0] add_797684;
  wire [7:0] sel_797685;
  wire [7:0] add_797688;
  wire [7:0] sel_797689;
  wire [7:0] add_797692;
  wire [7:0] sel_797693;
  wire [7:0] add_797696;
  wire [7:0] sel_797697;
  wire [7:0] add_797700;
  wire [7:0] sel_797701;
  wire [7:0] add_797704;
  wire [7:0] sel_797705;
  wire [7:0] add_797708;
  wire [7:0] sel_797709;
  wire [7:0] add_797712;
  wire [7:0] sel_797713;
  wire [7:0] add_797716;
  wire [7:0] sel_797717;
  wire [7:0] add_797720;
  wire [7:0] sel_797721;
  wire [7:0] add_797724;
  wire [7:0] sel_797725;
  wire [7:0] add_797728;
  wire [7:0] sel_797729;
  wire [7:0] add_797732;
  wire [7:0] sel_797733;
  wire [7:0] add_797736;
  wire [7:0] sel_797737;
  wire [7:0] add_797740;
  wire [7:0] sel_797741;
  wire [7:0] add_797744;
  wire [7:0] sel_797745;
  wire [7:0] add_797748;
  wire [7:0] sel_797749;
  wire [7:0] add_797752;
  wire [7:0] sel_797753;
  wire [7:0] add_797756;
  wire [7:0] sel_797757;
  wire [7:0] add_797760;
  wire [7:0] sel_797761;
  wire [7:0] add_797764;
  wire [7:0] sel_797765;
  wire [7:0] add_797768;
  wire [7:0] sel_797769;
  wire [7:0] add_797772;
  wire [7:0] sel_797773;
  wire [7:0] add_797776;
  wire [7:0] sel_797777;
  wire [7:0] add_797780;
  wire [7:0] sel_797781;
  wire [7:0] add_797784;
  wire [7:0] sel_797785;
  wire [7:0] add_797788;
  wire [7:0] sel_797789;
  wire [7:0] add_797792;
  wire [7:0] sel_797793;
  wire [7:0] add_797797;
  wire [15:0] array_index_797798;
  wire [7:0] sel_797799;
  wire [7:0] add_797802;
  wire [7:0] sel_797803;
  wire [7:0] add_797806;
  wire [7:0] sel_797807;
  wire [7:0] add_797810;
  wire [7:0] sel_797811;
  wire [7:0] add_797814;
  wire [7:0] sel_797815;
  wire [7:0] add_797818;
  wire [7:0] sel_797819;
  wire [7:0] add_797822;
  wire [7:0] sel_797823;
  wire [7:0] add_797826;
  wire [7:0] sel_797827;
  wire [7:0] add_797830;
  wire [7:0] sel_797831;
  wire [7:0] add_797834;
  wire [7:0] sel_797835;
  wire [7:0] add_797838;
  wire [7:0] sel_797839;
  wire [7:0] add_797842;
  wire [7:0] sel_797843;
  wire [7:0] add_797846;
  wire [7:0] sel_797847;
  wire [7:0] add_797850;
  wire [7:0] sel_797851;
  wire [7:0] add_797854;
  wire [7:0] sel_797855;
  wire [7:0] add_797858;
  wire [7:0] sel_797859;
  wire [7:0] add_797862;
  wire [7:0] sel_797863;
  wire [7:0] add_797866;
  wire [7:0] sel_797867;
  wire [7:0] add_797870;
  wire [7:0] sel_797871;
  wire [7:0] add_797874;
  wire [7:0] sel_797875;
  wire [7:0] add_797878;
  wire [7:0] sel_797879;
  wire [7:0] add_797882;
  wire [7:0] sel_797883;
  wire [7:0] add_797886;
  wire [7:0] sel_797887;
  wire [7:0] add_797890;
  wire [7:0] sel_797891;
  wire [7:0] add_797894;
  wire [7:0] sel_797895;
  wire [7:0] add_797898;
  wire [7:0] sel_797899;
  wire [7:0] add_797902;
  wire [7:0] sel_797903;
  wire [7:0] add_797906;
  wire [7:0] sel_797907;
  wire [7:0] add_797910;
  wire [7:0] sel_797911;
  wire [7:0] add_797914;
  wire [7:0] sel_797915;
  wire [7:0] add_797918;
  wire [7:0] sel_797919;
  wire [7:0] add_797922;
  wire [7:0] sel_797923;
  wire [7:0] add_797926;
  wire [7:0] sel_797927;
  wire [7:0] add_797930;
  wire [7:0] sel_797931;
  wire [7:0] add_797934;
  wire [7:0] sel_797935;
  wire [7:0] add_797938;
  wire [7:0] sel_797939;
  wire [7:0] add_797942;
  wire [7:0] sel_797943;
  wire [7:0] add_797946;
  wire [7:0] sel_797947;
  wire [7:0] add_797950;
  wire [7:0] sel_797951;
  wire [7:0] add_797954;
  wire [7:0] sel_797955;
  wire [7:0] add_797958;
  wire [7:0] sel_797959;
  wire [7:0] add_797962;
  wire [7:0] sel_797963;
  wire [7:0] add_797966;
  wire [7:0] sel_797967;
  wire [7:0] add_797970;
  wire [7:0] sel_797971;
  wire [7:0] add_797974;
  wire [7:0] sel_797975;
  wire [7:0] add_797978;
  wire [7:0] sel_797979;
  wire [7:0] add_797982;
  wire [7:0] sel_797983;
  wire [7:0] add_797986;
  wire [7:0] sel_797987;
  wire [7:0] add_797990;
  wire [7:0] sel_797991;
  wire [7:0] add_797994;
  wire [7:0] sel_797995;
  wire [7:0] add_797998;
  wire [7:0] sel_797999;
  wire [7:0] add_798002;
  wire [7:0] sel_798003;
  wire [7:0] add_798006;
  wire [7:0] sel_798007;
  wire [7:0] add_798010;
  wire [7:0] sel_798011;
  wire [7:0] add_798014;
  wire [7:0] sel_798015;
  wire [7:0] add_798018;
  wire [7:0] sel_798019;
  wire [7:0] add_798022;
  wire [7:0] sel_798023;
  wire [7:0] add_798026;
  wire [7:0] sel_798027;
  wire [7:0] add_798030;
  wire [7:0] sel_798031;
  wire [7:0] add_798034;
  wire [7:0] sel_798035;
  wire [7:0] add_798038;
  wire [7:0] sel_798039;
  wire [7:0] add_798042;
  wire [7:0] sel_798043;
  wire [7:0] add_798046;
  wire [7:0] sel_798047;
  wire [7:0] add_798050;
  wire [7:0] sel_798051;
  wire [7:0] add_798054;
  wire [7:0] sel_798055;
  wire [7:0] add_798058;
  wire [7:0] sel_798059;
  wire [7:0] add_798062;
  wire [7:0] sel_798063;
  wire [7:0] add_798066;
  wire [7:0] sel_798067;
  wire [7:0] add_798070;
  wire [7:0] sel_798071;
  wire [7:0] add_798074;
  wire [7:0] sel_798075;
  wire [7:0] add_798078;
  wire [7:0] sel_798079;
  wire [7:0] add_798082;
  wire [7:0] sel_798083;
  wire [7:0] add_798086;
  wire [7:0] sel_798087;
  wire [7:0] add_798090;
  wire [7:0] sel_798091;
  wire [7:0] add_798094;
  wire [7:0] sel_798095;
  wire [7:0] add_798098;
  wire [7:0] sel_798099;
  wire [7:0] add_798102;
  wire [7:0] sel_798103;
  wire [7:0] add_798106;
  wire [7:0] sel_798107;
  wire [7:0] add_798110;
  wire [7:0] sel_798111;
  wire [7:0] add_798114;
  wire [7:0] sel_798115;
  wire [7:0] add_798118;
  wire [7:0] sel_798119;
  wire [7:0] add_798122;
  wire [7:0] sel_798123;
  wire [7:0] add_798126;
  wire [7:0] sel_798127;
  wire [7:0] add_798130;
  wire [7:0] sel_798131;
  wire [7:0] add_798134;
  wire [7:0] sel_798135;
  wire [7:0] add_798138;
  wire [7:0] sel_798139;
  wire [7:0] add_798142;
  wire [7:0] sel_798143;
  wire [7:0] add_798146;
  wire [7:0] sel_798147;
  wire [7:0] add_798150;
  wire [7:0] sel_798151;
  wire [7:0] add_798154;
  wire [7:0] sel_798155;
  wire [7:0] add_798159;
  wire [15:0] array_index_798160;
  wire [7:0] sel_798161;
  wire [7:0] add_798164;
  wire [7:0] sel_798165;
  wire [7:0] add_798168;
  wire [7:0] sel_798169;
  wire [7:0] add_798172;
  wire [7:0] sel_798173;
  wire [7:0] add_798176;
  wire [7:0] sel_798177;
  wire [7:0] add_798180;
  wire [7:0] sel_798181;
  wire [7:0] add_798184;
  wire [7:0] sel_798185;
  wire [7:0] add_798188;
  wire [7:0] sel_798189;
  wire [7:0] add_798192;
  wire [7:0] sel_798193;
  wire [7:0] add_798196;
  wire [7:0] sel_798197;
  wire [7:0] add_798200;
  wire [7:0] sel_798201;
  wire [7:0] add_798204;
  wire [7:0] sel_798205;
  wire [7:0] add_798208;
  wire [7:0] sel_798209;
  wire [7:0] add_798212;
  wire [7:0] sel_798213;
  wire [7:0] add_798216;
  wire [7:0] sel_798217;
  wire [7:0] add_798220;
  wire [7:0] sel_798221;
  wire [7:0] add_798224;
  wire [7:0] sel_798225;
  wire [7:0] add_798228;
  wire [7:0] sel_798229;
  wire [7:0] add_798232;
  wire [7:0] sel_798233;
  wire [7:0] add_798236;
  wire [7:0] sel_798237;
  wire [7:0] add_798240;
  wire [7:0] sel_798241;
  wire [7:0] add_798244;
  wire [7:0] sel_798245;
  wire [7:0] add_798248;
  wire [7:0] sel_798249;
  wire [7:0] add_798252;
  wire [7:0] sel_798253;
  wire [7:0] add_798256;
  wire [7:0] sel_798257;
  wire [7:0] add_798260;
  wire [7:0] sel_798261;
  wire [7:0] add_798264;
  wire [7:0] sel_798265;
  wire [7:0] add_798268;
  wire [7:0] sel_798269;
  wire [7:0] add_798272;
  wire [7:0] sel_798273;
  wire [7:0] add_798276;
  wire [7:0] sel_798277;
  wire [7:0] add_798280;
  wire [7:0] sel_798281;
  wire [7:0] add_798284;
  wire [7:0] sel_798285;
  wire [7:0] add_798288;
  wire [7:0] sel_798289;
  wire [7:0] add_798292;
  wire [7:0] sel_798293;
  wire [7:0] add_798296;
  wire [7:0] sel_798297;
  wire [7:0] add_798300;
  wire [7:0] sel_798301;
  wire [7:0] add_798304;
  wire [7:0] sel_798305;
  wire [7:0] add_798308;
  wire [7:0] sel_798309;
  wire [7:0] add_798312;
  wire [7:0] sel_798313;
  wire [7:0] add_798316;
  wire [7:0] sel_798317;
  wire [7:0] add_798320;
  wire [7:0] sel_798321;
  wire [7:0] add_798324;
  wire [7:0] sel_798325;
  wire [7:0] add_798328;
  wire [7:0] sel_798329;
  wire [7:0] add_798332;
  wire [7:0] sel_798333;
  wire [7:0] add_798336;
  wire [7:0] sel_798337;
  wire [7:0] add_798340;
  wire [7:0] sel_798341;
  wire [7:0] add_798344;
  wire [7:0] sel_798345;
  wire [7:0] add_798348;
  wire [7:0] sel_798349;
  wire [7:0] add_798352;
  wire [7:0] sel_798353;
  wire [7:0] add_798356;
  wire [7:0] sel_798357;
  wire [7:0] add_798360;
  wire [7:0] sel_798361;
  wire [7:0] add_798364;
  wire [7:0] sel_798365;
  wire [7:0] add_798368;
  wire [7:0] sel_798369;
  wire [7:0] add_798372;
  wire [7:0] sel_798373;
  wire [7:0] add_798376;
  wire [7:0] sel_798377;
  wire [7:0] add_798380;
  wire [7:0] sel_798381;
  wire [7:0] add_798384;
  wire [7:0] sel_798385;
  wire [7:0] add_798388;
  wire [7:0] sel_798389;
  wire [7:0] add_798392;
  wire [7:0] sel_798393;
  wire [7:0] add_798396;
  wire [7:0] sel_798397;
  wire [7:0] add_798400;
  wire [7:0] sel_798401;
  wire [7:0] add_798404;
  wire [7:0] sel_798405;
  wire [7:0] add_798408;
  wire [7:0] sel_798409;
  wire [7:0] add_798412;
  wire [7:0] sel_798413;
  wire [7:0] add_798416;
  wire [7:0] sel_798417;
  wire [7:0] add_798420;
  wire [7:0] sel_798421;
  wire [7:0] add_798424;
  wire [7:0] sel_798425;
  wire [7:0] add_798428;
  wire [7:0] sel_798429;
  wire [7:0] add_798432;
  wire [7:0] sel_798433;
  wire [7:0] add_798436;
  wire [7:0] sel_798437;
  wire [7:0] add_798440;
  wire [7:0] sel_798441;
  wire [7:0] add_798444;
  wire [7:0] sel_798445;
  wire [7:0] add_798448;
  wire [7:0] sel_798449;
  wire [7:0] add_798452;
  wire [7:0] sel_798453;
  wire [7:0] add_798456;
  wire [7:0] sel_798457;
  wire [7:0] add_798460;
  wire [7:0] sel_798461;
  wire [7:0] add_798464;
  wire [7:0] sel_798465;
  wire [7:0] add_798468;
  wire [7:0] sel_798469;
  wire [7:0] add_798472;
  wire [7:0] sel_798473;
  wire [7:0] add_798476;
  wire [7:0] sel_798477;
  wire [7:0] add_798480;
  wire [7:0] sel_798481;
  wire [7:0] add_798484;
  wire [7:0] sel_798485;
  wire [7:0] add_798488;
  wire [7:0] sel_798489;
  wire [7:0] add_798492;
  wire [7:0] sel_798493;
  wire [7:0] add_798496;
  wire [7:0] sel_798497;
  wire [7:0] add_798500;
  wire [7:0] sel_798501;
  wire [7:0] add_798504;
  wire [7:0] sel_798505;
  wire [7:0] add_798508;
  wire [7:0] sel_798509;
  wire [7:0] add_798512;
  wire [7:0] sel_798513;
  wire [7:0] add_798516;
  wire [7:0] sel_798517;
  wire [7:0] add_798521;
  wire [15:0] array_index_798522;
  wire [7:0] sel_798523;
  wire [7:0] add_798526;
  wire [7:0] sel_798527;
  wire [7:0] add_798530;
  wire [7:0] sel_798531;
  wire [7:0] add_798534;
  wire [7:0] sel_798535;
  wire [7:0] add_798538;
  wire [7:0] sel_798539;
  wire [7:0] add_798542;
  wire [7:0] sel_798543;
  wire [7:0] add_798546;
  wire [7:0] sel_798547;
  wire [7:0] add_798550;
  wire [7:0] sel_798551;
  wire [7:0] add_798554;
  wire [7:0] sel_798555;
  wire [7:0] add_798558;
  wire [7:0] sel_798559;
  wire [7:0] add_798562;
  wire [7:0] sel_798563;
  wire [7:0] add_798566;
  wire [7:0] sel_798567;
  wire [7:0] add_798570;
  wire [7:0] sel_798571;
  wire [7:0] add_798574;
  wire [7:0] sel_798575;
  wire [7:0] add_798578;
  wire [7:0] sel_798579;
  wire [7:0] add_798582;
  wire [7:0] sel_798583;
  wire [7:0] add_798586;
  wire [7:0] sel_798587;
  wire [7:0] add_798590;
  wire [7:0] sel_798591;
  wire [7:0] add_798594;
  wire [7:0] sel_798595;
  wire [7:0] add_798598;
  wire [7:0] sel_798599;
  wire [7:0] add_798602;
  wire [7:0] sel_798603;
  wire [7:0] add_798606;
  wire [7:0] sel_798607;
  wire [7:0] add_798610;
  wire [7:0] sel_798611;
  wire [7:0] add_798614;
  wire [7:0] sel_798615;
  wire [7:0] add_798618;
  wire [7:0] sel_798619;
  wire [7:0] add_798622;
  wire [7:0] sel_798623;
  wire [7:0] add_798626;
  wire [7:0] sel_798627;
  wire [7:0] add_798630;
  wire [7:0] sel_798631;
  wire [7:0] add_798634;
  wire [7:0] sel_798635;
  wire [7:0] add_798638;
  wire [7:0] sel_798639;
  wire [7:0] add_798642;
  wire [7:0] sel_798643;
  wire [7:0] add_798646;
  wire [7:0] sel_798647;
  wire [7:0] add_798650;
  wire [7:0] sel_798651;
  wire [7:0] add_798654;
  wire [7:0] sel_798655;
  wire [7:0] add_798658;
  wire [7:0] sel_798659;
  wire [7:0] add_798662;
  wire [7:0] sel_798663;
  wire [7:0] add_798666;
  wire [7:0] sel_798667;
  wire [7:0] add_798670;
  wire [7:0] sel_798671;
  wire [7:0] add_798674;
  wire [7:0] sel_798675;
  wire [7:0] add_798678;
  wire [7:0] sel_798679;
  wire [7:0] add_798682;
  wire [7:0] sel_798683;
  wire [7:0] add_798686;
  wire [7:0] sel_798687;
  wire [7:0] add_798690;
  wire [7:0] sel_798691;
  wire [7:0] add_798694;
  wire [7:0] sel_798695;
  wire [7:0] add_798698;
  wire [7:0] sel_798699;
  wire [7:0] add_798702;
  wire [7:0] sel_798703;
  wire [7:0] add_798706;
  wire [7:0] sel_798707;
  wire [7:0] add_798710;
  wire [7:0] sel_798711;
  wire [7:0] add_798714;
  wire [7:0] sel_798715;
  wire [7:0] add_798718;
  wire [7:0] sel_798719;
  wire [7:0] add_798722;
  wire [7:0] sel_798723;
  wire [7:0] add_798726;
  wire [7:0] sel_798727;
  wire [7:0] add_798730;
  wire [7:0] sel_798731;
  wire [7:0] add_798734;
  wire [7:0] sel_798735;
  wire [7:0] add_798738;
  wire [7:0] sel_798739;
  wire [7:0] add_798742;
  wire [7:0] sel_798743;
  wire [7:0] add_798746;
  wire [7:0] sel_798747;
  wire [7:0] add_798750;
  wire [7:0] sel_798751;
  wire [7:0] add_798754;
  wire [7:0] sel_798755;
  wire [7:0] add_798758;
  wire [7:0] sel_798759;
  wire [7:0] add_798762;
  wire [7:0] sel_798763;
  wire [7:0] add_798766;
  wire [7:0] sel_798767;
  wire [7:0] add_798770;
  wire [7:0] sel_798771;
  wire [7:0] add_798774;
  wire [7:0] sel_798775;
  wire [7:0] add_798778;
  wire [7:0] sel_798779;
  wire [7:0] add_798782;
  wire [7:0] sel_798783;
  wire [7:0] add_798786;
  wire [7:0] sel_798787;
  wire [7:0] add_798790;
  wire [7:0] sel_798791;
  wire [7:0] add_798794;
  wire [7:0] sel_798795;
  wire [7:0] add_798798;
  wire [7:0] sel_798799;
  wire [7:0] add_798802;
  wire [7:0] sel_798803;
  wire [7:0] add_798806;
  wire [7:0] sel_798807;
  wire [7:0] add_798810;
  wire [7:0] sel_798811;
  wire [7:0] add_798814;
  wire [7:0] sel_798815;
  wire [7:0] add_798818;
  wire [7:0] sel_798819;
  wire [7:0] add_798822;
  wire [7:0] sel_798823;
  wire [7:0] add_798826;
  wire [7:0] sel_798827;
  wire [7:0] add_798830;
  wire [7:0] sel_798831;
  wire [7:0] add_798834;
  wire [7:0] sel_798835;
  wire [7:0] add_798838;
  wire [7:0] sel_798839;
  wire [7:0] add_798842;
  wire [7:0] sel_798843;
  wire [7:0] add_798846;
  wire [7:0] sel_798847;
  wire [7:0] add_798850;
  wire [7:0] sel_798851;
  wire [7:0] add_798854;
  wire [7:0] sel_798855;
  wire [7:0] add_798858;
  wire [7:0] sel_798859;
  wire [7:0] add_798862;
  wire [7:0] sel_798863;
  wire [7:0] add_798866;
  wire [7:0] sel_798867;
  wire [7:0] add_798870;
  wire [7:0] sel_798871;
  wire [7:0] add_798874;
  wire [7:0] sel_798875;
  wire [7:0] add_798878;
  wire [7:0] sel_798879;
  wire [7:0] add_798883;
  wire [15:0] array_index_798884;
  wire [7:0] sel_798885;
  wire [7:0] add_798888;
  wire [7:0] sel_798889;
  wire [7:0] add_798892;
  wire [7:0] sel_798893;
  wire [7:0] add_798896;
  wire [7:0] sel_798897;
  wire [7:0] add_798900;
  wire [7:0] sel_798901;
  wire [7:0] add_798904;
  wire [7:0] sel_798905;
  wire [7:0] add_798908;
  wire [7:0] sel_798909;
  wire [7:0] add_798912;
  wire [7:0] sel_798913;
  wire [7:0] add_798916;
  wire [7:0] sel_798917;
  wire [7:0] add_798920;
  wire [7:0] sel_798921;
  wire [7:0] add_798924;
  wire [7:0] sel_798925;
  wire [7:0] add_798928;
  wire [7:0] sel_798929;
  wire [7:0] add_798932;
  wire [7:0] sel_798933;
  wire [7:0] add_798936;
  wire [7:0] sel_798937;
  wire [7:0] add_798940;
  wire [7:0] sel_798941;
  wire [7:0] add_798944;
  wire [7:0] sel_798945;
  wire [7:0] add_798948;
  wire [7:0] sel_798949;
  wire [7:0] add_798952;
  wire [7:0] sel_798953;
  wire [7:0] add_798956;
  wire [7:0] sel_798957;
  wire [7:0] add_798960;
  wire [7:0] sel_798961;
  wire [7:0] add_798964;
  wire [7:0] sel_798965;
  wire [7:0] add_798968;
  wire [7:0] sel_798969;
  wire [7:0] add_798972;
  wire [7:0] sel_798973;
  wire [7:0] add_798976;
  wire [7:0] sel_798977;
  wire [7:0] add_798980;
  wire [7:0] sel_798981;
  wire [7:0] add_798984;
  wire [7:0] sel_798985;
  wire [7:0] add_798988;
  wire [7:0] sel_798989;
  wire [7:0] add_798992;
  wire [7:0] sel_798993;
  wire [7:0] add_798996;
  wire [7:0] sel_798997;
  wire [7:0] add_799000;
  wire [7:0] sel_799001;
  wire [7:0] add_799004;
  wire [7:0] sel_799005;
  wire [7:0] add_799008;
  wire [7:0] sel_799009;
  wire [7:0] add_799012;
  wire [7:0] sel_799013;
  wire [7:0] add_799016;
  wire [7:0] sel_799017;
  wire [7:0] add_799020;
  wire [7:0] sel_799021;
  wire [7:0] add_799024;
  wire [7:0] sel_799025;
  wire [7:0] add_799028;
  wire [7:0] sel_799029;
  wire [7:0] add_799032;
  wire [7:0] sel_799033;
  wire [7:0] add_799036;
  wire [7:0] sel_799037;
  wire [7:0] add_799040;
  wire [7:0] sel_799041;
  wire [7:0] add_799044;
  wire [7:0] sel_799045;
  wire [7:0] add_799048;
  wire [7:0] sel_799049;
  wire [7:0] add_799052;
  wire [7:0] sel_799053;
  wire [7:0] add_799056;
  wire [7:0] sel_799057;
  wire [7:0] add_799060;
  wire [7:0] sel_799061;
  wire [7:0] add_799064;
  wire [7:0] sel_799065;
  wire [7:0] add_799068;
  wire [7:0] sel_799069;
  wire [7:0] add_799072;
  wire [7:0] sel_799073;
  wire [7:0] add_799076;
  wire [7:0] sel_799077;
  wire [7:0] add_799080;
  wire [7:0] sel_799081;
  wire [7:0] add_799084;
  wire [7:0] sel_799085;
  wire [7:0] add_799088;
  wire [7:0] sel_799089;
  wire [7:0] add_799092;
  wire [7:0] sel_799093;
  wire [7:0] add_799096;
  wire [7:0] sel_799097;
  wire [7:0] add_799100;
  wire [7:0] sel_799101;
  wire [7:0] add_799104;
  wire [7:0] sel_799105;
  wire [7:0] add_799108;
  wire [7:0] sel_799109;
  wire [7:0] add_799112;
  wire [7:0] sel_799113;
  wire [7:0] add_799116;
  wire [7:0] sel_799117;
  wire [7:0] add_799120;
  wire [7:0] sel_799121;
  wire [7:0] add_799124;
  wire [7:0] sel_799125;
  wire [7:0] add_799128;
  wire [7:0] sel_799129;
  wire [7:0] add_799132;
  wire [7:0] sel_799133;
  wire [7:0] add_799136;
  wire [7:0] sel_799137;
  wire [7:0] add_799140;
  wire [7:0] sel_799141;
  wire [7:0] add_799144;
  wire [7:0] sel_799145;
  wire [7:0] add_799148;
  wire [7:0] sel_799149;
  wire [7:0] add_799152;
  wire [7:0] sel_799153;
  wire [7:0] add_799156;
  wire [7:0] sel_799157;
  wire [7:0] add_799160;
  wire [7:0] sel_799161;
  wire [7:0] add_799164;
  wire [7:0] sel_799165;
  wire [7:0] add_799168;
  wire [7:0] sel_799169;
  wire [7:0] add_799172;
  wire [7:0] sel_799173;
  wire [7:0] add_799176;
  wire [7:0] sel_799177;
  wire [7:0] add_799180;
  wire [7:0] sel_799181;
  wire [7:0] add_799184;
  wire [7:0] sel_799185;
  wire [7:0] add_799188;
  wire [7:0] sel_799189;
  wire [7:0] add_799192;
  wire [7:0] sel_799193;
  wire [7:0] add_799196;
  wire [7:0] sel_799197;
  wire [7:0] add_799200;
  wire [7:0] sel_799201;
  wire [7:0] add_799204;
  wire [7:0] sel_799205;
  wire [7:0] add_799208;
  wire [7:0] sel_799209;
  wire [7:0] add_799212;
  wire [7:0] sel_799213;
  wire [7:0] add_799216;
  wire [7:0] sel_799217;
  wire [7:0] add_799220;
  wire [7:0] sel_799221;
  wire [7:0] add_799224;
  wire [7:0] sel_799225;
  wire [7:0] add_799228;
  wire [7:0] sel_799229;
  wire [7:0] add_799232;
  wire [7:0] sel_799233;
  wire [7:0] add_799236;
  wire [7:0] sel_799237;
  wire [7:0] add_799240;
  wire [7:0] sel_799241;
  wire [7:0] add_799245;
  wire [15:0] array_index_799246;
  wire [7:0] sel_799247;
  wire [7:0] add_799250;
  wire [7:0] sel_799251;
  wire [7:0] add_799254;
  wire [7:0] sel_799255;
  wire [7:0] add_799258;
  wire [7:0] sel_799259;
  wire [7:0] add_799262;
  wire [7:0] sel_799263;
  wire [7:0] add_799266;
  wire [7:0] sel_799267;
  wire [7:0] add_799270;
  wire [7:0] sel_799271;
  wire [7:0] add_799274;
  wire [7:0] sel_799275;
  wire [7:0] add_799278;
  wire [7:0] sel_799279;
  wire [7:0] add_799282;
  wire [7:0] sel_799283;
  wire [7:0] add_799286;
  wire [7:0] sel_799287;
  wire [7:0] add_799290;
  wire [7:0] sel_799291;
  wire [7:0] add_799294;
  wire [7:0] sel_799295;
  wire [7:0] add_799298;
  wire [7:0] sel_799299;
  wire [7:0] add_799302;
  wire [7:0] sel_799303;
  wire [7:0] add_799306;
  wire [7:0] sel_799307;
  wire [7:0] add_799310;
  wire [7:0] sel_799311;
  wire [7:0] add_799314;
  wire [7:0] sel_799315;
  wire [7:0] add_799318;
  wire [7:0] sel_799319;
  wire [7:0] add_799322;
  wire [7:0] sel_799323;
  wire [7:0] add_799326;
  wire [7:0] sel_799327;
  wire [7:0] add_799330;
  wire [7:0] sel_799331;
  wire [7:0] add_799334;
  wire [7:0] sel_799335;
  wire [7:0] add_799338;
  wire [7:0] sel_799339;
  wire [7:0] add_799342;
  wire [7:0] sel_799343;
  wire [7:0] add_799346;
  wire [7:0] sel_799347;
  wire [7:0] add_799350;
  wire [7:0] sel_799351;
  wire [7:0] add_799354;
  wire [7:0] sel_799355;
  wire [7:0] add_799358;
  wire [7:0] sel_799359;
  wire [7:0] add_799362;
  wire [7:0] sel_799363;
  wire [7:0] add_799366;
  wire [7:0] sel_799367;
  wire [7:0] add_799370;
  wire [7:0] sel_799371;
  wire [7:0] add_799374;
  wire [7:0] sel_799375;
  wire [7:0] add_799378;
  wire [7:0] sel_799379;
  wire [7:0] add_799382;
  wire [7:0] sel_799383;
  wire [7:0] add_799386;
  wire [7:0] sel_799387;
  wire [7:0] add_799390;
  wire [7:0] sel_799391;
  wire [7:0] add_799394;
  wire [7:0] sel_799395;
  wire [7:0] add_799398;
  wire [7:0] sel_799399;
  wire [7:0] add_799402;
  wire [7:0] sel_799403;
  wire [7:0] add_799406;
  wire [7:0] sel_799407;
  wire [7:0] add_799410;
  wire [7:0] sel_799411;
  wire [7:0] add_799414;
  wire [7:0] sel_799415;
  wire [7:0] add_799418;
  wire [7:0] sel_799419;
  wire [7:0] add_799422;
  wire [7:0] sel_799423;
  wire [7:0] add_799426;
  wire [7:0] sel_799427;
  wire [7:0] add_799430;
  wire [7:0] sel_799431;
  wire [7:0] add_799434;
  wire [7:0] sel_799435;
  wire [7:0] add_799438;
  wire [7:0] sel_799439;
  wire [7:0] add_799442;
  wire [7:0] sel_799443;
  wire [7:0] add_799446;
  wire [7:0] sel_799447;
  wire [7:0] add_799450;
  wire [7:0] sel_799451;
  wire [7:0] add_799454;
  wire [7:0] sel_799455;
  wire [7:0] add_799458;
  wire [7:0] sel_799459;
  wire [7:0] add_799462;
  wire [7:0] sel_799463;
  wire [7:0] add_799466;
  wire [7:0] sel_799467;
  wire [7:0] add_799470;
  wire [7:0] sel_799471;
  wire [7:0] add_799474;
  wire [7:0] sel_799475;
  wire [7:0] add_799478;
  wire [7:0] sel_799479;
  wire [7:0] add_799482;
  wire [7:0] sel_799483;
  wire [7:0] add_799486;
  wire [7:0] sel_799487;
  wire [7:0] add_799490;
  wire [7:0] sel_799491;
  wire [7:0] add_799494;
  wire [7:0] sel_799495;
  wire [7:0] add_799498;
  wire [7:0] sel_799499;
  wire [7:0] add_799502;
  wire [7:0] sel_799503;
  wire [7:0] add_799506;
  wire [7:0] sel_799507;
  wire [7:0] add_799510;
  wire [7:0] sel_799511;
  wire [7:0] add_799514;
  wire [7:0] sel_799515;
  wire [7:0] add_799518;
  wire [7:0] sel_799519;
  wire [7:0] add_799522;
  wire [7:0] sel_799523;
  wire [7:0] add_799526;
  wire [7:0] sel_799527;
  wire [7:0] add_799530;
  wire [7:0] sel_799531;
  wire [7:0] add_799534;
  wire [7:0] sel_799535;
  wire [7:0] add_799538;
  wire [7:0] sel_799539;
  wire [7:0] add_799542;
  wire [7:0] sel_799543;
  wire [7:0] add_799546;
  wire [7:0] sel_799547;
  wire [7:0] add_799550;
  wire [7:0] sel_799551;
  wire [7:0] add_799554;
  wire [7:0] sel_799555;
  wire [7:0] add_799558;
  wire [7:0] sel_799559;
  wire [7:0] add_799562;
  wire [7:0] sel_799563;
  wire [7:0] add_799566;
  wire [7:0] sel_799567;
  wire [7:0] add_799570;
  wire [7:0] sel_799571;
  wire [7:0] add_799574;
  wire [7:0] sel_799575;
  wire [7:0] add_799578;
  wire [7:0] sel_799579;
  wire [7:0] add_799582;
  wire [7:0] sel_799583;
  wire [7:0] add_799586;
  wire [7:0] sel_799587;
  wire [7:0] add_799590;
  wire [7:0] sel_799591;
  wire [7:0] add_799594;
  wire [7:0] sel_799595;
  wire [7:0] add_799598;
  wire [7:0] sel_799599;
  wire [7:0] add_799602;
  wire [7:0] sel_799603;
  wire [7:0] add_799607;
  wire [15:0] array_index_799608;
  wire [7:0] sel_799609;
  wire [7:0] add_799612;
  wire [7:0] sel_799613;
  wire [7:0] add_799616;
  wire [7:0] sel_799617;
  wire [7:0] add_799620;
  wire [7:0] sel_799621;
  wire [7:0] add_799624;
  wire [7:0] sel_799625;
  wire [7:0] add_799628;
  wire [7:0] sel_799629;
  wire [7:0] add_799632;
  wire [7:0] sel_799633;
  wire [7:0] add_799636;
  wire [7:0] sel_799637;
  wire [7:0] add_799640;
  wire [7:0] sel_799641;
  wire [7:0] add_799644;
  wire [7:0] sel_799645;
  wire [7:0] add_799648;
  wire [7:0] sel_799649;
  wire [7:0] add_799652;
  wire [7:0] sel_799653;
  wire [7:0] add_799656;
  wire [7:0] sel_799657;
  wire [7:0] add_799660;
  wire [7:0] sel_799661;
  wire [7:0] add_799664;
  wire [7:0] sel_799665;
  wire [7:0] add_799668;
  wire [7:0] sel_799669;
  wire [7:0] add_799672;
  wire [7:0] sel_799673;
  wire [7:0] add_799676;
  wire [7:0] sel_799677;
  wire [7:0] add_799680;
  wire [7:0] sel_799681;
  wire [7:0] add_799684;
  wire [7:0] sel_799685;
  wire [7:0] add_799688;
  wire [7:0] sel_799689;
  wire [7:0] add_799692;
  wire [7:0] sel_799693;
  wire [7:0] add_799696;
  wire [7:0] sel_799697;
  wire [7:0] add_799700;
  wire [7:0] sel_799701;
  wire [7:0] add_799704;
  wire [7:0] sel_799705;
  wire [7:0] add_799708;
  wire [7:0] sel_799709;
  wire [7:0] add_799712;
  wire [7:0] sel_799713;
  wire [7:0] add_799716;
  wire [7:0] sel_799717;
  wire [7:0] add_799720;
  wire [7:0] sel_799721;
  wire [7:0] add_799724;
  wire [7:0] sel_799725;
  wire [7:0] add_799728;
  wire [7:0] sel_799729;
  wire [7:0] add_799732;
  wire [7:0] sel_799733;
  wire [7:0] add_799736;
  wire [7:0] sel_799737;
  wire [7:0] add_799740;
  wire [7:0] sel_799741;
  wire [7:0] add_799744;
  wire [7:0] sel_799745;
  wire [7:0] add_799748;
  wire [7:0] sel_799749;
  wire [7:0] add_799752;
  wire [7:0] sel_799753;
  wire [7:0] add_799756;
  wire [7:0] sel_799757;
  wire [7:0] add_799760;
  wire [7:0] sel_799761;
  wire [7:0] add_799764;
  wire [7:0] sel_799765;
  wire [7:0] add_799768;
  wire [7:0] sel_799769;
  wire [7:0] add_799772;
  wire [7:0] sel_799773;
  wire [7:0] add_799776;
  wire [7:0] sel_799777;
  wire [7:0] add_799780;
  wire [7:0] sel_799781;
  wire [7:0] add_799784;
  wire [7:0] sel_799785;
  wire [7:0] add_799788;
  wire [7:0] sel_799789;
  wire [7:0] add_799792;
  wire [7:0] sel_799793;
  wire [7:0] add_799796;
  wire [7:0] sel_799797;
  wire [7:0] add_799800;
  wire [7:0] sel_799801;
  wire [7:0] add_799804;
  wire [7:0] sel_799805;
  wire [7:0] add_799808;
  wire [7:0] sel_799809;
  wire [7:0] add_799812;
  wire [7:0] sel_799813;
  wire [7:0] add_799816;
  wire [7:0] sel_799817;
  wire [7:0] add_799820;
  wire [7:0] sel_799821;
  wire [7:0] add_799824;
  wire [7:0] sel_799825;
  wire [7:0] add_799828;
  wire [7:0] sel_799829;
  wire [7:0] add_799832;
  wire [7:0] sel_799833;
  wire [7:0] add_799836;
  wire [7:0] sel_799837;
  wire [7:0] add_799840;
  wire [7:0] sel_799841;
  wire [7:0] add_799844;
  wire [7:0] sel_799845;
  wire [7:0] add_799848;
  wire [7:0] sel_799849;
  wire [7:0] add_799852;
  wire [7:0] sel_799853;
  wire [7:0] add_799856;
  wire [7:0] sel_799857;
  wire [7:0] add_799860;
  wire [7:0] sel_799861;
  wire [7:0] add_799864;
  wire [7:0] sel_799865;
  wire [7:0] add_799868;
  wire [7:0] sel_799869;
  wire [7:0] add_799872;
  wire [7:0] sel_799873;
  wire [7:0] add_799876;
  wire [7:0] sel_799877;
  wire [7:0] add_799880;
  wire [7:0] sel_799881;
  wire [7:0] add_799884;
  wire [7:0] sel_799885;
  wire [7:0] add_799888;
  wire [7:0] sel_799889;
  wire [7:0] add_799892;
  wire [7:0] sel_799893;
  wire [7:0] add_799896;
  wire [7:0] sel_799897;
  wire [7:0] add_799900;
  wire [7:0] sel_799901;
  wire [7:0] add_799904;
  wire [7:0] sel_799905;
  wire [7:0] add_799908;
  wire [7:0] sel_799909;
  wire [7:0] add_799912;
  wire [7:0] sel_799913;
  wire [7:0] add_799916;
  wire [7:0] sel_799917;
  wire [7:0] add_799920;
  wire [7:0] sel_799921;
  wire [7:0] add_799924;
  wire [7:0] sel_799925;
  wire [7:0] add_799928;
  wire [7:0] sel_799929;
  wire [7:0] add_799932;
  wire [7:0] sel_799933;
  wire [7:0] add_799936;
  wire [7:0] sel_799937;
  wire [7:0] add_799940;
  wire [7:0] sel_799941;
  wire [7:0] add_799944;
  wire [7:0] sel_799945;
  wire [7:0] add_799948;
  wire [7:0] sel_799949;
  wire [7:0] add_799952;
  wire [7:0] sel_799953;
  wire [7:0] add_799956;
  wire [7:0] sel_799957;
  wire [7:0] add_799960;
  wire [7:0] sel_799961;
  wire [7:0] add_799964;
  wire [7:0] sel_799965;
  wire [7:0] add_799969;
  wire [15:0] array_index_799970;
  wire [7:0] sel_799971;
  wire [7:0] add_799974;
  wire [7:0] sel_799975;
  wire [7:0] add_799978;
  wire [7:0] sel_799979;
  wire [7:0] add_799982;
  wire [7:0] sel_799983;
  wire [7:0] add_799986;
  wire [7:0] sel_799987;
  wire [7:0] add_799990;
  wire [7:0] sel_799991;
  wire [7:0] add_799994;
  wire [7:0] sel_799995;
  wire [7:0] add_799998;
  wire [7:0] sel_799999;
  wire [7:0] add_800002;
  wire [7:0] sel_800003;
  wire [7:0] add_800006;
  wire [7:0] sel_800007;
  wire [7:0] add_800010;
  wire [7:0] sel_800011;
  wire [7:0] add_800014;
  wire [7:0] sel_800015;
  wire [7:0] add_800018;
  wire [7:0] sel_800019;
  wire [7:0] add_800022;
  wire [7:0] sel_800023;
  wire [7:0] add_800026;
  wire [7:0] sel_800027;
  wire [7:0] add_800030;
  wire [7:0] sel_800031;
  wire [7:0] add_800034;
  wire [7:0] sel_800035;
  wire [7:0] add_800038;
  wire [7:0] sel_800039;
  wire [7:0] add_800042;
  wire [7:0] sel_800043;
  wire [7:0] add_800046;
  wire [7:0] sel_800047;
  wire [7:0] add_800050;
  wire [7:0] sel_800051;
  wire [7:0] add_800054;
  wire [7:0] sel_800055;
  wire [7:0] add_800058;
  wire [7:0] sel_800059;
  wire [7:0] add_800062;
  wire [7:0] sel_800063;
  wire [7:0] add_800066;
  wire [7:0] sel_800067;
  wire [7:0] add_800070;
  wire [7:0] sel_800071;
  wire [7:0] add_800074;
  wire [7:0] sel_800075;
  wire [7:0] add_800078;
  wire [7:0] sel_800079;
  wire [7:0] add_800082;
  wire [7:0] sel_800083;
  wire [7:0] add_800086;
  wire [7:0] sel_800087;
  wire [7:0] add_800090;
  wire [7:0] sel_800091;
  wire [7:0] add_800094;
  wire [7:0] sel_800095;
  wire [7:0] add_800098;
  wire [7:0] sel_800099;
  wire [7:0] add_800102;
  wire [7:0] sel_800103;
  wire [7:0] add_800106;
  wire [7:0] sel_800107;
  wire [7:0] add_800110;
  wire [7:0] sel_800111;
  wire [7:0] add_800114;
  wire [7:0] sel_800115;
  wire [7:0] add_800118;
  wire [7:0] sel_800119;
  wire [7:0] add_800122;
  wire [7:0] sel_800123;
  wire [7:0] add_800126;
  wire [7:0] sel_800127;
  wire [7:0] add_800130;
  wire [7:0] sel_800131;
  wire [7:0] add_800134;
  wire [7:0] sel_800135;
  wire [7:0] add_800138;
  wire [7:0] sel_800139;
  wire [7:0] add_800142;
  wire [7:0] sel_800143;
  wire [7:0] add_800146;
  wire [7:0] sel_800147;
  wire [7:0] add_800150;
  wire [7:0] sel_800151;
  wire [7:0] add_800154;
  wire [7:0] sel_800155;
  wire [7:0] add_800158;
  wire [7:0] sel_800159;
  wire [7:0] add_800162;
  wire [7:0] sel_800163;
  wire [7:0] add_800166;
  wire [7:0] sel_800167;
  wire [7:0] add_800170;
  wire [7:0] sel_800171;
  wire [7:0] add_800174;
  wire [7:0] sel_800175;
  wire [7:0] add_800178;
  wire [7:0] sel_800179;
  wire [7:0] add_800182;
  wire [7:0] sel_800183;
  wire [7:0] add_800186;
  wire [7:0] sel_800187;
  wire [7:0] add_800190;
  wire [7:0] sel_800191;
  wire [7:0] add_800194;
  wire [7:0] sel_800195;
  wire [7:0] add_800198;
  wire [7:0] sel_800199;
  wire [7:0] add_800202;
  wire [7:0] sel_800203;
  wire [7:0] add_800206;
  wire [7:0] sel_800207;
  wire [7:0] add_800210;
  wire [7:0] sel_800211;
  wire [7:0] add_800214;
  wire [7:0] sel_800215;
  wire [7:0] add_800218;
  wire [7:0] sel_800219;
  wire [7:0] add_800222;
  wire [7:0] sel_800223;
  wire [7:0] add_800226;
  wire [7:0] sel_800227;
  wire [7:0] add_800230;
  wire [7:0] sel_800231;
  wire [7:0] add_800234;
  wire [7:0] sel_800235;
  wire [7:0] add_800238;
  wire [7:0] sel_800239;
  wire [7:0] add_800242;
  wire [7:0] sel_800243;
  wire [7:0] add_800246;
  wire [7:0] sel_800247;
  wire [7:0] add_800250;
  wire [7:0] sel_800251;
  wire [7:0] add_800254;
  wire [7:0] sel_800255;
  wire [7:0] add_800258;
  wire [7:0] sel_800259;
  wire [7:0] add_800262;
  wire [7:0] sel_800263;
  wire [7:0] add_800266;
  wire [7:0] sel_800267;
  wire [7:0] add_800270;
  wire [7:0] sel_800271;
  wire [7:0] add_800274;
  wire [7:0] sel_800275;
  wire [7:0] add_800278;
  wire [7:0] sel_800279;
  wire [7:0] add_800282;
  wire [7:0] sel_800283;
  wire [7:0] add_800286;
  wire [7:0] sel_800287;
  wire [7:0] add_800290;
  wire [7:0] sel_800291;
  wire [7:0] add_800294;
  wire [7:0] sel_800295;
  wire [7:0] add_800298;
  wire [7:0] sel_800299;
  wire [7:0] add_800302;
  wire [7:0] sel_800303;
  wire [7:0] add_800306;
  wire [7:0] sel_800307;
  wire [7:0] add_800310;
  wire [7:0] sel_800311;
  wire [7:0] add_800314;
  wire [7:0] sel_800315;
  wire [7:0] add_800318;
  wire [7:0] sel_800319;
  wire [7:0] add_800322;
  wire [7:0] sel_800323;
  wire [7:0] add_800326;
  wire [7:0] sel_800327;
  wire [7:0] add_800331;
  wire [15:0] array_index_800332;
  wire [7:0] sel_800333;
  wire [7:0] add_800336;
  wire [7:0] sel_800337;
  wire [7:0] add_800340;
  wire [7:0] sel_800341;
  wire [7:0] add_800344;
  wire [7:0] sel_800345;
  wire [7:0] add_800348;
  wire [7:0] sel_800349;
  wire [7:0] add_800352;
  wire [7:0] sel_800353;
  wire [7:0] add_800356;
  wire [7:0] sel_800357;
  wire [7:0] add_800360;
  wire [7:0] sel_800361;
  wire [7:0] add_800364;
  wire [7:0] sel_800365;
  wire [7:0] add_800368;
  wire [7:0] sel_800369;
  wire [7:0] add_800372;
  wire [7:0] sel_800373;
  wire [7:0] add_800376;
  wire [7:0] sel_800377;
  wire [7:0] add_800380;
  wire [7:0] sel_800381;
  wire [7:0] add_800384;
  wire [7:0] sel_800385;
  wire [7:0] add_800388;
  wire [7:0] sel_800389;
  wire [7:0] add_800392;
  wire [7:0] sel_800393;
  wire [7:0] add_800396;
  wire [7:0] sel_800397;
  wire [7:0] add_800400;
  wire [7:0] sel_800401;
  wire [7:0] add_800404;
  wire [7:0] sel_800405;
  wire [7:0] add_800408;
  wire [7:0] sel_800409;
  wire [7:0] add_800412;
  wire [7:0] sel_800413;
  wire [7:0] add_800416;
  wire [7:0] sel_800417;
  wire [7:0] add_800420;
  wire [7:0] sel_800421;
  wire [7:0] add_800424;
  wire [7:0] sel_800425;
  wire [7:0] add_800428;
  wire [7:0] sel_800429;
  wire [7:0] add_800432;
  wire [7:0] sel_800433;
  wire [7:0] add_800436;
  wire [7:0] sel_800437;
  wire [7:0] add_800440;
  wire [7:0] sel_800441;
  wire [7:0] add_800444;
  wire [7:0] sel_800445;
  wire [7:0] add_800448;
  wire [7:0] sel_800449;
  wire [7:0] add_800452;
  wire [7:0] sel_800453;
  wire [7:0] add_800456;
  wire [7:0] sel_800457;
  wire [7:0] add_800460;
  wire [7:0] sel_800461;
  wire [7:0] add_800464;
  wire [7:0] sel_800465;
  wire [7:0] add_800468;
  wire [7:0] sel_800469;
  wire [7:0] add_800472;
  wire [7:0] sel_800473;
  wire [7:0] add_800476;
  wire [7:0] sel_800477;
  wire [7:0] add_800480;
  wire [7:0] sel_800481;
  wire [7:0] add_800484;
  wire [7:0] sel_800485;
  wire [7:0] add_800488;
  wire [7:0] sel_800489;
  wire [7:0] add_800492;
  wire [7:0] sel_800493;
  wire [7:0] add_800496;
  wire [7:0] sel_800497;
  wire [7:0] add_800500;
  wire [7:0] sel_800501;
  wire [7:0] add_800504;
  wire [7:0] sel_800505;
  wire [7:0] add_800508;
  wire [7:0] sel_800509;
  wire [7:0] add_800512;
  wire [7:0] sel_800513;
  wire [7:0] add_800516;
  wire [7:0] sel_800517;
  wire [7:0] add_800520;
  wire [7:0] sel_800521;
  wire [7:0] add_800524;
  wire [7:0] sel_800525;
  wire [7:0] add_800528;
  wire [7:0] sel_800529;
  wire [7:0] add_800532;
  wire [7:0] sel_800533;
  wire [7:0] add_800536;
  wire [7:0] sel_800537;
  wire [7:0] add_800540;
  wire [7:0] sel_800541;
  wire [7:0] add_800544;
  wire [7:0] sel_800545;
  wire [7:0] add_800548;
  wire [7:0] sel_800549;
  wire [7:0] add_800552;
  wire [7:0] sel_800553;
  wire [7:0] add_800556;
  wire [7:0] sel_800557;
  wire [7:0] add_800560;
  wire [7:0] sel_800561;
  wire [7:0] add_800564;
  wire [7:0] sel_800565;
  wire [7:0] add_800568;
  wire [7:0] sel_800569;
  wire [7:0] add_800572;
  wire [7:0] sel_800573;
  wire [7:0] add_800576;
  wire [7:0] sel_800577;
  wire [7:0] add_800580;
  wire [7:0] sel_800581;
  wire [7:0] add_800584;
  wire [7:0] sel_800585;
  wire [7:0] add_800588;
  wire [7:0] sel_800589;
  wire [7:0] add_800592;
  wire [7:0] sel_800593;
  wire [7:0] add_800596;
  wire [7:0] sel_800597;
  wire [7:0] add_800600;
  wire [7:0] sel_800601;
  wire [7:0] add_800604;
  wire [7:0] sel_800605;
  wire [7:0] add_800608;
  wire [7:0] sel_800609;
  wire [7:0] add_800612;
  wire [7:0] sel_800613;
  wire [7:0] add_800616;
  wire [7:0] sel_800617;
  wire [7:0] add_800620;
  wire [7:0] sel_800621;
  wire [7:0] add_800624;
  wire [7:0] sel_800625;
  wire [7:0] add_800628;
  wire [7:0] sel_800629;
  wire [7:0] add_800632;
  wire [7:0] sel_800633;
  wire [7:0] add_800636;
  wire [7:0] sel_800637;
  wire [7:0] add_800640;
  wire [7:0] sel_800641;
  wire [7:0] add_800644;
  wire [7:0] sel_800645;
  wire [7:0] add_800648;
  wire [7:0] sel_800649;
  wire [7:0] add_800652;
  wire [7:0] sel_800653;
  wire [7:0] add_800656;
  wire [7:0] sel_800657;
  wire [7:0] add_800660;
  wire [7:0] sel_800661;
  wire [7:0] add_800664;
  wire [7:0] sel_800665;
  wire [7:0] add_800668;
  wire [7:0] sel_800669;
  wire [7:0] add_800672;
  wire [7:0] sel_800673;
  wire [7:0] add_800676;
  wire [7:0] sel_800677;
  wire [7:0] add_800680;
  wire [7:0] sel_800681;
  wire [7:0] add_800684;
  wire [7:0] sel_800685;
  wire [7:0] add_800688;
  wire [7:0] sel_800689;
  wire [7:0] add_800693;
  wire [15:0] array_index_800694;
  wire [7:0] sel_800695;
  wire [7:0] add_800698;
  wire [7:0] sel_800699;
  wire [7:0] add_800702;
  wire [7:0] sel_800703;
  wire [7:0] add_800706;
  wire [7:0] sel_800707;
  wire [7:0] add_800710;
  wire [7:0] sel_800711;
  wire [7:0] add_800714;
  wire [7:0] sel_800715;
  wire [7:0] add_800718;
  wire [7:0] sel_800719;
  wire [7:0] add_800722;
  wire [7:0] sel_800723;
  wire [7:0] add_800726;
  wire [7:0] sel_800727;
  wire [7:0] add_800730;
  wire [7:0] sel_800731;
  wire [7:0] add_800734;
  wire [7:0] sel_800735;
  wire [7:0] add_800738;
  wire [7:0] sel_800739;
  wire [7:0] add_800742;
  wire [7:0] sel_800743;
  wire [7:0] add_800746;
  wire [7:0] sel_800747;
  wire [7:0] add_800750;
  wire [7:0] sel_800751;
  wire [7:0] add_800754;
  wire [7:0] sel_800755;
  wire [7:0] add_800758;
  wire [7:0] sel_800759;
  wire [7:0] add_800762;
  wire [7:0] sel_800763;
  wire [7:0] add_800766;
  wire [7:0] sel_800767;
  wire [7:0] add_800770;
  wire [7:0] sel_800771;
  wire [7:0] add_800774;
  wire [7:0] sel_800775;
  wire [7:0] add_800778;
  wire [7:0] sel_800779;
  wire [7:0] add_800782;
  wire [7:0] sel_800783;
  wire [7:0] add_800786;
  wire [7:0] sel_800787;
  wire [7:0] add_800790;
  wire [7:0] sel_800791;
  wire [7:0] add_800794;
  wire [7:0] sel_800795;
  wire [7:0] add_800798;
  wire [7:0] sel_800799;
  wire [7:0] add_800802;
  wire [7:0] sel_800803;
  wire [7:0] add_800806;
  wire [7:0] sel_800807;
  wire [7:0] add_800810;
  wire [7:0] sel_800811;
  wire [7:0] add_800814;
  wire [7:0] sel_800815;
  wire [7:0] add_800818;
  wire [7:0] sel_800819;
  wire [7:0] add_800822;
  wire [7:0] sel_800823;
  wire [7:0] add_800826;
  wire [7:0] sel_800827;
  wire [7:0] add_800830;
  wire [7:0] sel_800831;
  wire [7:0] add_800834;
  wire [7:0] sel_800835;
  wire [7:0] add_800838;
  wire [7:0] sel_800839;
  wire [7:0] add_800842;
  wire [7:0] sel_800843;
  wire [7:0] add_800846;
  wire [7:0] sel_800847;
  wire [7:0] add_800850;
  wire [7:0] sel_800851;
  wire [7:0] add_800854;
  wire [7:0] sel_800855;
  wire [7:0] add_800858;
  wire [7:0] sel_800859;
  wire [7:0] add_800862;
  wire [7:0] sel_800863;
  wire [7:0] add_800866;
  wire [7:0] sel_800867;
  wire [7:0] add_800870;
  wire [7:0] sel_800871;
  wire [7:0] add_800874;
  wire [7:0] sel_800875;
  wire [7:0] add_800878;
  wire [7:0] sel_800879;
  wire [7:0] add_800882;
  wire [7:0] sel_800883;
  wire [7:0] add_800886;
  wire [7:0] sel_800887;
  wire [7:0] add_800890;
  wire [7:0] sel_800891;
  wire [7:0] add_800894;
  wire [7:0] sel_800895;
  wire [7:0] add_800898;
  wire [7:0] sel_800899;
  wire [7:0] add_800902;
  wire [7:0] sel_800903;
  wire [7:0] add_800906;
  wire [7:0] sel_800907;
  wire [7:0] add_800910;
  wire [7:0] sel_800911;
  wire [7:0] add_800914;
  wire [7:0] sel_800915;
  wire [7:0] add_800918;
  wire [7:0] sel_800919;
  wire [7:0] add_800922;
  wire [7:0] sel_800923;
  wire [7:0] add_800926;
  wire [7:0] sel_800927;
  wire [7:0] add_800930;
  wire [7:0] sel_800931;
  wire [7:0] add_800934;
  wire [7:0] sel_800935;
  wire [7:0] add_800938;
  wire [7:0] sel_800939;
  wire [7:0] add_800942;
  wire [7:0] sel_800943;
  wire [7:0] add_800946;
  wire [7:0] sel_800947;
  wire [7:0] add_800950;
  wire [7:0] sel_800951;
  wire [7:0] add_800954;
  wire [7:0] sel_800955;
  wire [7:0] add_800958;
  wire [7:0] sel_800959;
  wire [7:0] add_800962;
  wire [7:0] sel_800963;
  wire [7:0] add_800966;
  wire [7:0] sel_800967;
  wire [7:0] add_800970;
  wire [7:0] sel_800971;
  wire [7:0] add_800974;
  wire [7:0] sel_800975;
  wire [7:0] add_800978;
  wire [7:0] sel_800979;
  wire [7:0] add_800982;
  wire [7:0] sel_800983;
  wire [7:0] add_800986;
  wire [7:0] sel_800987;
  wire [7:0] add_800990;
  wire [7:0] sel_800991;
  wire [7:0] add_800994;
  wire [7:0] sel_800995;
  wire [7:0] add_800998;
  wire [7:0] sel_800999;
  wire [7:0] add_801002;
  wire [7:0] sel_801003;
  wire [7:0] add_801006;
  wire [7:0] sel_801007;
  wire [7:0] add_801010;
  wire [7:0] sel_801011;
  wire [7:0] add_801014;
  wire [7:0] sel_801015;
  wire [7:0] add_801018;
  wire [7:0] sel_801019;
  wire [7:0] add_801022;
  wire [7:0] sel_801023;
  wire [7:0] add_801026;
  wire [7:0] sel_801027;
  wire [7:0] add_801030;
  wire [7:0] sel_801031;
  wire [7:0] add_801034;
  wire [7:0] sel_801035;
  wire [7:0] add_801038;
  wire [7:0] sel_801039;
  wire [7:0] add_801042;
  wire [7:0] sel_801043;
  wire [7:0] add_801046;
  wire [7:0] sel_801047;
  wire [7:0] add_801050;
  wire [7:0] sel_801051;
  wire [7:0] add_801055;
  wire [15:0] array_index_801056;
  wire [7:0] sel_801057;
  wire [7:0] add_801060;
  wire [7:0] sel_801061;
  wire [7:0] add_801064;
  wire [7:0] sel_801065;
  wire [7:0] add_801068;
  wire [7:0] sel_801069;
  wire [7:0] add_801072;
  wire [7:0] sel_801073;
  wire [7:0] add_801076;
  wire [7:0] sel_801077;
  wire [7:0] add_801080;
  wire [7:0] sel_801081;
  wire [7:0] add_801084;
  wire [7:0] sel_801085;
  wire [7:0] add_801088;
  wire [7:0] sel_801089;
  wire [7:0] add_801092;
  wire [7:0] sel_801093;
  wire [7:0] add_801096;
  wire [7:0] sel_801097;
  wire [7:0] add_801100;
  wire [7:0] sel_801101;
  wire [7:0] add_801104;
  wire [7:0] sel_801105;
  wire [7:0] add_801108;
  wire [7:0] sel_801109;
  wire [7:0] add_801112;
  wire [7:0] sel_801113;
  wire [7:0] add_801116;
  wire [7:0] sel_801117;
  wire [7:0] add_801120;
  wire [7:0] sel_801121;
  wire [7:0] add_801124;
  wire [7:0] sel_801125;
  wire [7:0] add_801128;
  wire [7:0] sel_801129;
  wire [7:0] add_801132;
  wire [7:0] sel_801133;
  wire [7:0] add_801136;
  wire [7:0] sel_801137;
  wire [7:0] add_801140;
  wire [7:0] sel_801141;
  wire [7:0] add_801144;
  wire [7:0] sel_801145;
  wire [7:0] add_801148;
  wire [7:0] sel_801149;
  wire [7:0] add_801152;
  wire [7:0] sel_801153;
  wire [7:0] add_801156;
  wire [7:0] sel_801157;
  wire [7:0] add_801160;
  wire [7:0] sel_801161;
  wire [7:0] add_801164;
  wire [7:0] sel_801165;
  wire [7:0] add_801168;
  wire [7:0] sel_801169;
  wire [7:0] add_801172;
  wire [7:0] sel_801173;
  wire [7:0] add_801176;
  wire [7:0] sel_801177;
  wire [7:0] add_801180;
  wire [7:0] sel_801181;
  wire [7:0] add_801184;
  wire [7:0] sel_801185;
  wire [7:0] add_801188;
  wire [7:0] sel_801189;
  wire [7:0] add_801192;
  wire [7:0] sel_801193;
  wire [7:0] add_801196;
  wire [7:0] sel_801197;
  wire [7:0] add_801200;
  wire [7:0] sel_801201;
  wire [7:0] add_801204;
  wire [7:0] sel_801205;
  wire [7:0] add_801208;
  wire [7:0] sel_801209;
  wire [7:0] add_801212;
  wire [7:0] sel_801213;
  wire [7:0] add_801216;
  wire [7:0] sel_801217;
  wire [7:0] add_801220;
  wire [7:0] sel_801221;
  wire [7:0] add_801224;
  wire [7:0] sel_801225;
  wire [7:0] add_801228;
  wire [7:0] sel_801229;
  wire [7:0] add_801232;
  wire [7:0] sel_801233;
  wire [7:0] add_801236;
  wire [7:0] sel_801237;
  wire [7:0] add_801240;
  wire [7:0] sel_801241;
  wire [7:0] add_801244;
  wire [7:0] sel_801245;
  wire [7:0] add_801248;
  wire [7:0] sel_801249;
  wire [7:0] add_801252;
  wire [7:0] sel_801253;
  wire [7:0] add_801256;
  wire [7:0] sel_801257;
  wire [7:0] add_801260;
  wire [7:0] sel_801261;
  wire [7:0] add_801264;
  wire [7:0] sel_801265;
  wire [7:0] add_801268;
  wire [7:0] sel_801269;
  wire [7:0] add_801272;
  wire [7:0] sel_801273;
  wire [7:0] add_801276;
  wire [7:0] sel_801277;
  wire [7:0] add_801280;
  wire [7:0] sel_801281;
  wire [7:0] add_801284;
  wire [7:0] sel_801285;
  wire [7:0] add_801288;
  wire [7:0] sel_801289;
  wire [7:0] add_801292;
  wire [7:0] sel_801293;
  wire [7:0] add_801296;
  wire [7:0] sel_801297;
  wire [7:0] add_801300;
  wire [7:0] sel_801301;
  wire [7:0] add_801304;
  wire [7:0] sel_801305;
  wire [7:0] add_801308;
  wire [7:0] sel_801309;
  wire [7:0] add_801312;
  wire [7:0] sel_801313;
  wire [7:0] add_801316;
  wire [7:0] sel_801317;
  wire [7:0] add_801320;
  wire [7:0] sel_801321;
  wire [7:0] add_801324;
  wire [7:0] sel_801325;
  wire [7:0] add_801328;
  wire [7:0] sel_801329;
  wire [7:0] add_801332;
  wire [7:0] sel_801333;
  wire [7:0] add_801336;
  wire [7:0] sel_801337;
  wire [7:0] add_801340;
  wire [7:0] sel_801341;
  wire [7:0] add_801344;
  wire [7:0] sel_801345;
  wire [7:0] add_801348;
  wire [7:0] sel_801349;
  wire [7:0] add_801352;
  wire [7:0] sel_801353;
  wire [7:0] add_801356;
  wire [7:0] sel_801357;
  wire [7:0] add_801360;
  wire [7:0] sel_801361;
  wire [7:0] add_801364;
  wire [7:0] sel_801365;
  wire [7:0] add_801368;
  wire [7:0] sel_801369;
  wire [7:0] add_801372;
  wire [7:0] sel_801373;
  wire [7:0] add_801376;
  wire [7:0] sel_801377;
  wire [7:0] add_801380;
  wire [7:0] sel_801381;
  wire [7:0] add_801384;
  wire [7:0] sel_801385;
  wire [7:0] add_801388;
  wire [7:0] sel_801389;
  wire [7:0] add_801392;
  wire [7:0] sel_801393;
  wire [7:0] add_801396;
  wire [7:0] sel_801397;
  wire [7:0] add_801400;
  wire [7:0] sel_801401;
  wire [7:0] add_801404;
  wire [7:0] sel_801405;
  wire [7:0] add_801408;
  wire [7:0] sel_801409;
  wire [7:0] add_801412;
  wire [7:0] sel_801413;
  wire [7:0] add_801417;
  wire [15:0] array_index_801418;
  wire [7:0] sel_801419;
  wire [7:0] add_801422;
  wire [7:0] sel_801423;
  wire [7:0] add_801426;
  wire [7:0] sel_801427;
  wire [7:0] add_801430;
  wire [7:0] sel_801431;
  wire [7:0] add_801434;
  wire [7:0] sel_801435;
  wire [7:0] add_801438;
  wire [7:0] sel_801439;
  wire [7:0] add_801442;
  wire [7:0] sel_801443;
  wire [7:0] add_801446;
  wire [7:0] sel_801447;
  wire [7:0] add_801450;
  wire [7:0] sel_801451;
  wire [7:0] add_801454;
  wire [7:0] sel_801455;
  wire [7:0] add_801458;
  wire [7:0] sel_801459;
  wire [7:0] add_801462;
  wire [7:0] sel_801463;
  wire [7:0] add_801466;
  wire [7:0] sel_801467;
  wire [7:0] add_801470;
  wire [7:0] sel_801471;
  wire [7:0] add_801474;
  wire [7:0] sel_801475;
  wire [7:0] add_801478;
  wire [7:0] sel_801479;
  wire [7:0] add_801482;
  wire [7:0] sel_801483;
  wire [7:0] add_801486;
  wire [7:0] sel_801487;
  wire [7:0] add_801490;
  wire [7:0] sel_801491;
  wire [7:0] add_801494;
  wire [7:0] sel_801495;
  wire [7:0] add_801498;
  wire [7:0] sel_801499;
  wire [7:0] add_801502;
  wire [7:0] sel_801503;
  wire [7:0] add_801506;
  wire [7:0] sel_801507;
  wire [7:0] add_801510;
  wire [7:0] sel_801511;
  wire [7:0] add_801514;
  wire [7:0] sel_801515;
  wire [7:0] add_801518;
  wire [7:0] sel_801519;
  wire [7:0] add_801522;
  wire [7:0] sel_801523;
  wire [7:0] add_801526;
  wire [7:0] sel_801527;
  wire [7:0] add_801530;
  wire [7:0] sel_801531;
  wire [7:0] add_801534;
  wire [7:0] sel_801535;
  wire [7:0] add_801538;
  wire [7:0] sel_801539;
  wire [7:0] add_801542;
  wire [7:0] sel_801543;
  wire [7:0] add_801546;
  wire [7:0] sel_801547;
  wire [7:0] add_801550;
  wire [7:0] sel_801551;
  wire [7:0] add_801554;
  wire [7:0] sel_801555;
  wire [7:0] add_801558;
  wire [7:0] sel_801559;
  wire [7:0] add_801562;
  wire [7:0] sel_801563;
  wire [7:0] add_801566;
  wire [7:0] sel_801567;
  wire [7:0] add_801570;
  wire [7:0] sel_801571;
  wire [7:0] add_801574;
  wire [7:0] sel_801575;
  wire [7:0] add_801578;
  wire [7:0] sel_801579;
  wire [7:0] add_801582;
  wire [7:0] sel_801583;
  wire [7:0] add_801586;
  wire [7:0] sel_801587;
  wire [7:0] add_801590;
  wire [7:0] sel_801591;
  wire [7:0] add_801594;
  wire [7:0] sel_801595;
  wire [7:0] add_801598;
  wire [7:0] sel_801599;
  wire [7:0] add_801602;
  wire [7:0] sel_801603;
  wire [7:0] add_801606;
  wire [7:0] sel_801607;
  wire [7:0] add_801610;
  wire [7:0] sel_801611;
  wire [7:0] add_801614;
  wire [7:0] sel_801615;
  wire [7:0] add_801618;
  wire [7:0] sel_801619;
  wire [7:0] add_801622;
  wire [7:0] sel_801623;
  wire [7:0] add_801626;
  wire [7:0] sel_801627;
  wire [7:0] add_801630;
  wire [7:0] sel_801631;
  wire [7:0] add_801634;
  wire [7:0] sel_801635;
  wire [7:0] add_801638;
  wire [7:0] sel_801639;
  wire [7:0] add_801642;
  wire [7:0] sel_801643;
  wire [7:0] add_801646;
  wire [7:0] sel_801647;
  wire [7:0] add_801650;
  wire [7:0] sel_801651;
  wire [7:0] add_801654;
  wire [7:0] sel_801655;
  wire [7:0] add_801658;
  wire [7:0] sel_801659;
  wire [7:0] add_801662;
  wire [7:0] sel_801663;
  wire [7:0] add_801666;
  wire [7:0] sel_801667;
  wire [7:0] add_801670;
  wire [7:0] sel_801671;
  wire [7:0] add_801674;
  wire [7:0] sel_801675;
  wire [7:0] add_801678;
  wire [7:0] sel_801679;
  wire [7:0] add_801682;
  wire [7:0] sel_801683;
  wire [7:0] add_801686;
  wire [7:0] sel_801687;
  wire [7:0] add_801690;
  wire [7:0] sel_801691;
  wire [7:0] add_801694;
  wire [7:0] sel_801695;
  wire [7:0] add_801698;
  wire [7:0] sel_801699;
  wire [7:0] add_801702;
  wire [7:0] sel_801703;
  wire [7:0] add_801706;
  wire [7:0] sel_801707;
  wire [7:0] add_801710;
  wire [7:0] sel_801711;
  wire [7:0] add_801714;
  wire [7:0] sel_801715;
  wire [7:0] add_801718;
  wire [7:0] sel_801719;
  wire [7:0] add_801722;
  wire [7:0] sel_801723;
  wire [7:0] add_801726;
  wire [7:0] sel_801727;
  wire [7:0] add_801730;
  wire [7:0] sel_801731;
  wire [7:0] add_801734;
  wire [7:0] sel_801735;
  wire [7:0] add_801738;
  wire [7:0] sel_801739;
  wire [7:0] add_801742;
  wire [7:0] sel_801743;
  wire [7:0] add_801746;
  wire [7:0] sel_801747;
  wire [7:0] add_801750;
  wire [7:0] sel_801751;
  wire [7:0] add_801754;
  wire [7:0] sel_801755;
  wire [7:0] add_801758;
  wire [7:0] sel_801759;
  wire [7:0] add_801762;
  wire [7:0] sel_801763;
  wire [7:0] add_801766;
  wire [7:0] sel_801767;
  wire [7:0] add_801770;
  wire [7:0] sel_801771;
  wire [7:0] add_801774;
  wire [7:0] sel_801775;
  wire [7:0] add_801779;
  wire [15:0] array_index_801780;
  wire [7:0] sel_801781;
  wire [7:0] add_801784;
  wire [7:0] sel_801785;
  wire [7:0] add_801788;
  wire [7:0] sel_801789;
  wire [7:0] add_801792;
  wire [7:0] sel_801793;
  wire [7:0] add_801796;
  wire [7:0] sel_801797;
  wire [7:0] add_801800;
  wire [7:0] sel_801801;
  wire [7:0] add_801804;
  wire [7:0] sel_801805;
  wire [7:0] add_801808;
  wire [7:0] sel_801809;
  wire [7:0] add_801812;
  wire [7:0] sel_801813;
  wire [7:0] add_801816;
  wire [7:0] sel_801817;
  wire [7:0] add_801820;
  wire [7:0] sel_801821;
  wire [7:0] add_801824;
  wire [7:0] sel_801825;
  wire [7:0] add_801828;
  wire [7:0] sel_801829;
  wire [7:0] add_801832;
  wire [7:0] sel_801833;
  wire [7:0] add_801836;
  wire [7:0] sel_801837;
  wire [7:0] add_801840;
  wire [7:0] sel_801841;
  wire [7:0] add_801844;
  wire [7:0] sel_801845;
  wire [7:0] add_801848;
  wire [7:0] sel_801849;
  wire [7:0] add_801852;
  wire [7:0] sel_801853;
  wire [7:0] add_801856;
  wire [7:0] sel_801857;
  wire [7:0] add_801860;
  wire [7:0] sel_801861;
  wire [7:0] add_801864;
  wire [7:0] sel_801865;
  wire [7:0] add_801868;
  wire [7:0] sel_801869;
  wire [7:0] add_801872;
  wire [7:0] sel_801873;
  wire [7:0] add_801876;
  wire [7:0] sel_801877;
  wire [7:0] add_801880;
  wire [7:0] sel_801881;
  wire [7:0] add_801884;
  wire [7:0] sel_801885;
  wire [7:0] add_801888;
  wire [7:0] sel_801889;
  wire [7:0] add_801892;
  wire [7:0] sel_801893;
  wire [7:0] add_801896;
  wire [7:0] sel_801897;
  wire [7:0] add_801900;
  wire [7:0] sel_801901;
  wire [7:0] add_801904;
  wire [7:0] sel_801905;
  wire [7:0] add_801908;
  wire [7:0] sel_801909;
  wire [7:0] add_801912;
  wire [7:0] sel_801913;
  wire [7:0] add_801916;
  wire [7:0] sel_801917;
  wire [7:0] add_801920;
  wire [7:0] sel_801921;
  wire [7:0] add_801924;
  wire [7:0] sel_801925;
  wire [7:0] add_801928;
  wire [7:0] sel_801929;
  wire [7:0] add_801932;
  wire [7:0] sel_801933;
  wire [7:0] add_801936;
  wire [7:0] sel_801937;
  wire [7:0] add_801940;
  wire [7:0] sel_801941;
  wire [7:0] add_801944;
  wire [7:0] sel_801945;
  wire [7:0] add_801948;
  wire [7:0] sel_801949;
  wire [7:0] add_801952;
  wire [7:0] sel_801953;
  wire [7:0] add_801956;
  wire [7:0] sel_801957;
  wire [7:0] add_801960;
  wire [7:0] sel_801961;
  wire [7:0] add_801964;
  wire [7:0] sel_801965;
  wire [7:0] add_801968;
  wire [7:0] sel_801969;
  wire [7:0] add_801972;
  wire [7:0] sel_801973;
  wire [7:0] add_801976;
  wire [7:0] sel_801977;
  wire [7:0] add_801980;
  wire [7:0] sel_801981;
  wire [7:0] add_801984;
  wire [7:0] sel_801985;
  wire [7:0] add_801988;
  wire [7:0] sel_801989;
  wire [7:0] add_801992;
  wire [7:0] sel_801993;
  wire [7:0] add_801996;
  wire [7:0] sel_801997;
  wire [7:0] add_802000;
  wire [7:0] sel_802001;
  wire [7:0] add_802004;
  wire [7:0] sel_802005;
  wire [7:0] add_802008;
  wire [7:0] sel_802009;
  wire [7:0] add_802012;
  wire [7:0] sel_802013;
  wire [7:0] add_802016;
  wire [7:0] sel_802017;
  wire [7:0] add_802020;
  wire [7:0] sel_802021;
  wire [7:0] add_802024;
  wire [7:0] sel_802025;
  wire [7:0] add_802028;
  wire [7:0] sel_802029;
  wire [7:0] add_802032;
  wire [7:0] sel_802033;
  wire [7:0] add_802036;
  wire [7:0] sel_802037;
  wire [7:0] add_802040;
  wire [7:0] sel_802041;
  wire [7:0] add_802044;
  wire [7:0] sel_802045;
  wire [7:0] add_802048;
  wire [7:0] sel_802049;
  wire [7:0] add_802052;
  wire [7:0] sel_802053;
  wire [7:0] add_802056;
  wire [7:0] sel_802057;
  wire [7:0] add_802060;
  wire [7:0] sel_802061;
  wire [7:0] add_802064;
  wire [7:0] sel_802065;
  wire [7:0] add_802068;
  wire [7:0] sel_802069;
  wire [7:0] add_802072;
  wire [7:0] sel_802073;
  wire [7:0] add_802076;
  wire [7:0] sel_802077;
  wire [7:0] add_802080;
  wire [7:0] sel_802081;
  wire [7:0] add_802084;
  wire [7:0] sel_802085;
  wire [7:0] add_802088;
  wire [7:0] sel_802089;
  wire [7:0] add_802092;
  wire [7:0] sel_802093;
  wire [7:0] add_802096;
  wire [7:0] sel_802097;
  wire [7:0] add_802100;
  wire [7:0] sel_802101;
  wire [7:0] add_802104;
  wire [7:0] sel_802105;
  wire [7:0] add_802108;
  wire [7:0] sel_802109;
  wire [7:0] add_802112;
  wire [7:0] sel_802113;
  wire [7:0] add_802116;
  wire [7:0] sel_802117;
  wire [7:0] add_802120;
  wire [7:0] sel_802121;
  wire [7:0] add_802124;
  wire [7:0] sel_802125;
  wire [7:0] add_802128;
  wire [7:0] sel_802129;
  wire [7:0] add_802132;
  wire [7:0] sel_802133;
  wire [7:0] add_802136;
  wire [7:0] sel_802137;
  wire [7:0] add_802141;
  wire [15:0] array_index_802142;
  wire [7:0] sel_802143;
  wire [7:0] add_802146;
  wire [7:0] sel_802147;
  wire [7:0] add_802150;
  wire [7:0] sel_802151;
  wire [7:0] add_802154;
  wire [7:0] sel_802155;
  wire [7:0] add_802158;
  wire [7:0] sel_802159;
  wire [7:0] add_802162;
  wire [7:0] sel_802163;
  wire [7:0] add_802166;
  wire [7:0] sel_802167;
  wire [7:0] add_802170;
  wire [7:0] sel_802171;
  wire [7:0] add_802174;
  wire [7:0] sel_802175;
  wire [7:0] add_802178;
  wire [7:0] sel_802179;
  wire [7:0] add_802182;
  wire [7:0] sel_802183;
  wire [7:0] add_802186;
  wire [7:0] sel_802187;
  wire [7:0] add_802190;
  wire [7:0] sel_802191;
  wire [7:0] add_802194;
  wire [7:0] sel_802195;
  wire [7:0] add_802198;
  wire [7:0] sel_802199;
  wire [7:0] add_802202;
  wire [7:0] sel_802203;
  wire [7:0] add_802206;
  wire [7:0] sel_802207;
  wire [7:0] add_802210;
  wire [7:0] sel_802211;
  wire [7:0] add_802214;
  wire [7:0] sel_802215;
  wire [7:0] add_802218;
  wire [7:0] sel_802219;
  wire [7:0] add_802222;
  wire [7:0] sel_802223;
  wire [7:0] add_802226;
  wire [7:0] sel_802227;
  wire [7:0] add_802230;
  wire [7:0] sel_802231;
  wire [7:0] add_802234;
  wire [7:0] sel_802235;
  wire [7:0] add_802238;
  wire [7:0] sel_802239;
  wire [7:0] add_802242;
  wire [7:0] sel_802243;
  wire [7:0] add_802246;
  wire [7:0] sel_802247;
  wire [7:0] add_802250;
  wire [7:0] sel_802251;
  wire [7:0] add_802254;
  wire [7:0] sel_802255;
  wire [7:0] add_802258;
  wire [7:0] sel_802259;
  wire [7:0] add_802262;
  wire [7:0] sel_802263;
  wire [7:0] add_802266;
  wire [7:0] sel_802267;
  wire [7:0] add_802270;
  wire [7:0] sel_802271;
  wire [7:0] add_802274;
  wire [7:0] sel_802275;
  wire [7:0] add_802278;
  wire [7:0] sel_802279;
  wire [7:0] add_802282;
  wire [7:0] sel_802283;
  wire [7:0] add_802286;
  wire [7:0] sel_802287;
  wire [7:0] add_802290;
  wire [7:0] sel_802291;
  wire [7:0] add_802294;
  wire [7:0] sel_802295;
  wire [7:0] add_802298;
  wire [7:0] sel_802299;
  wire [7:0] add_802302;
  wire [7:0] sel_802303;
  wire [7:0] add_802306;
  wire [7:0] sel_802307;
  wire [7:0] add_802310;
  wire [7:0] sel_802311;
  wire [7:0] add_802314;
  wire [7:0] sel_802315;
  wire [7:0] add_802318;
  wire [7:0] sel_802319;
  wire [7:0] add_802322;
  wire [7:0] sel_802323;
  wire [7:0] add_802326;
  wire [7:0] sel_802327;
  wire [7:0] add_802330;
  wire [7:0] sel_802331;
  wire [7:0] add_802334;
  wire [7:0] sel_802335;
  wire [7:0] add_802338;
  wire [7:0] sel_802339;
  wire [7:0] add_802342;
  wire [7:0] sel_802343;
  wire [7:0] add_802346;
  wire [7:0] sel_802347;
  wire [7:0] add_802350;
  wire [7:0] sel_802351;
  wire [7:0] add_802354;
  wire [7:0] sel_802355;
  wire [7:0] add_802358;
  wire [7:0] sel_802359;
  wire [7:0] add_802362;
  wire [7:0] sel_802363;
  wire [7:0] add_802366;
  wire [7:0] sel_802367;
  wire [7:0] add_802370;
  wire [7:0] sel_802371;
  wire [7:0] add_802374;
  wire [7:0] sel_802375;
  wire [7:0] add_802378;
  wire [7:0] sel_802379;
  wire [7:0] add_802382;
  wire [7:0] sel_802383;
  wire [7:0] add_802386;
  wire [7:0] sel_802387;
  wire [7:0] add_802390;
  wire [7:0] sel_802391;
  wire [7:0] add_802394;
  wire [7:0] sel_802395;
  wire [7:0] add_802398;
  wire [7:0] sel_802399;
  wire [7:0] add_802402;
  wire [7:0] sel_802403;
  wire [7:0] add_802406;
  wire [7:0] sel_802407;
  wire [7:0] add_802410;
  wire [7:0] sel_802411;
  wire [7:0] add_802414;
  wire [7:0] sel_802415;
  wire [7:0] add_802418;
  wire [7:0] sel_802419;
  wire [7:0] add_802422;
  wire [7:0] sel_802423;
  wire [7:0] add_802426;
  wire [7:0] sel_802427;
  wire [7:0] add_802430;
  wire [7:0] sel_802431;
  wire [7:0] add_802434;
  wire [7:0] sel_802435;
  wire [7:0] add_802438;
  wire [7:0] sel_802439;
  wire [7:0] add_802442;
  wire [7:0] sel_802443;
  wire [7:0] add_802446;
  wire [7:0] sel_802447;
  wire [7:0] add_802450;
  wire [7:0] sel_802451;
  wire [7:0] add_802454;
  wire [7:0] sel_802455;
  wire [7:0] add_802458;
  wire [7:0] sel_802459;
  wire [7:0] add_802462;
  wire [7:0] sel_802463;
  wire [7:0] add_802466;
  wire [7:0] sel_802467;
  wire [7:0] add_802470;
  wire [7:0] sel_802471;
  wire [7:0] add_802474;
  wire [7:0] sel_802475;
  wire [7:0] add_802478;
  wire [7:0] sel_802479;
  wire [7:0] add_802482;
  wire [7:0] sel_802483;
  wire [7:0] add_802486;
  wire [7:0] sel_802487;
  wire [7:0] add_802490;
  wire [7:0] sel_802491;
  wire [7:0] add_802494;
  wire [7:0] sel_802495;
  wire [7:0] add_802498;
  wire [7:0] sel_802499;
  wire [7:0] add_802503;
  wire [15:0] array_index_802504;
  wire [7:0] sel_802505;
  wire [7:0] add_802508;
  wire [7:0] sel_802509;
  wire [7:0] add_802512;
  wire [7:0] sel_802513;
  wire [7:0] add_802516;
  wire [7:0] sel_802517;
  wire [7:0] add_802520;
  wire [7:0] sel_802521;
  wire [7:0] add_802524;
  wire [7:0] sel_802525;
  wire [7:0] add_802528;
  wire [7:0] sel_802529;
  wire [7:0] add_802532;
  wire [7:0] sel_802533;
  wire [7:0] add_802536;
  wire [7:0] sel_802537;
  wire [7:0] add_802540;
  wire [7:0] sel_802541;
  wire [7:0] add_802544;
  wire [7:0] sel_802545;
  wire [7:0] add_802548;
  wire [7:0] sel_802549;
  wire [7:0] add_802552;
  wire [7:0] sel_802553;
  wire [7:0] add_802556;
  wire [7:0] sel_802557;
  wire [7:0] add_802560;
  wire [7:0] sel_802561;
  wire [7:0] add_802564;
  wire [7:0] sel_802565;
  wire [7:0] add_802568;
  wire [7:0] sel_802569;
  wire [7:0] add_802572;
  wire [7:0] sel_802573;
  wire [7:0] add_802576;
  wire [7:0] sel_802577;
  wire [7:0] add_802580;
  wire [7:0] sel_802581;
  wire [7:0] add_802584;
  wire [7:0] sel_802585;
  wire [7:0] add_802588;
  wire [7:0] sel_802589;
  wire [7:0] add_802592;
  wire [7:0] sel_802593;
  wire [7:0] add_802596;
  wire [7:0] sel_802597;
  wire [7:0] add_802600;
  wire [7:0] sel_802601;
  wire [7:0] add_802604;
  wire [7:0] sel_802605;
  wire [7:0] add_802608;
  wire [7:0] sel_802609;
  wire [7:0] add_802612;
  wire [7:0] sel_802613;
  wire [7:0] add_802616;
  wire [7:0] sel_802617;
  wire [7:0] add_802620;
  wire [7:0] sel_802621;
  wire [7:0] add_802624;
  wire [7:0] sel_802625;
  wire [7:0] add_802628;
  wire [7:0] sel_802629;
  wire [7:0] add_802632;
  wire [7:0] sel_802633;
  wire [7:0] add_802636;
  wire [7:0] sel_802637;
  wire [7:0] add_802640;
  wire [7:0] sel_802641;
  wire [7:0] add_802644;
  wire [7:0] sel_802645;
  wire [7:0] add_802648;
  wire [7:0] sel_802649;
  wire [7:0] add_802652;
  wire [7:0] sel_802653;
  wire [7:0] add_802656;
  wire [7:0] sel_802657;
  wire [7:0] add_802660;
  wire [7:0] sel_802661;
  wire [7:0] add_802664;
  wire [7:0] sel_802665;
  wire [7:0] add_802668;
  wire [7:0] sel_802669;
  wire [7:0] add_802672;
  wire [7:0] sel_802673;
  wire [7:0] add_802676;
  wire [7:0] sel_802677;
  wire [7:0] add_802680;
  wire [7:0] sel_802681;
  wire [7:0] add_802684;
  wire [7:0] sel_802685;
  wire [7:0] add_802688;
  wire [7:0] sel_802689;
  wire [7:0] add_802692;
  wire [7:0] sel_802693;
  wire [7:0] add_802696;
  wire [7:0] sel_802697;
  wire [7:0] add_802700;
  wire [7:0] sel_802701;
  wire [7:0] add_802704;
  wire [7:0] sel_802705;
  wire [7:0] add_802708;
  wire [7:0] sel_802709;
  wire [7:0] add_802712;
  wire [7:0] sel_802713;
  wire [7:0] add_802716;
  wire [7:0] sel_802717;
  wire [7:0] add_802720;
  wire [7:0] sel_802721;
  wire [7:0] add_802724;
  wire [7:0] sel_802725;
  wire [7:0] add_802728;
  wire [7:0] sel_802729;
  wire [7:0] add_802732;
  wire [7:0] sel_802733;
  wire [7:0] add_802736;
  wire [7:0] sel_802737;
  wire [7:0] add_802740;
  wire [7:0] sel_802741;
  wire [7:0] add_802744;
  wire [7:0] sel_802745;
  wire [7:0] add_802748;
  wire [7:0] sel_802749;
  wire [7:0] add_802752;
  wire [7:0] sel_802753;
  wire [7:0] add_802756;
  wire [7:0] sel_802757;
  wire [7:0] add_802760;
  wire [7:0] sel_802761;
  wire [7:0] add_802764;
  wire [7:0] sel_802765;
  wire [7:0] add_802768;
  wire [7:0] sel_802769;
  wire [7:0] add_802772;
  wire [7:0] sel_802773;
  wire [7:0] add_802776;
  wire [7:0] sel_802777;
  wire [7:0] add_802780;
  wire [7:0] sel_802781;
  wire [7:0] add_802784;
  wire [7:0] sel_802785;
  wire [7:0] add_802788;
  wire [7:0] sel_802789;
  wire [7:0] add_802792;
  wire [7:0] sel_802793;
  wire [7:0] add_802796;
  wire [7:0] sel_802797;
  wire [7:0] add_802800;
  wire [7:0] sel_802801;
  wire [7:0] add_802804;
  wire [7:0] sel_802805;
  wire [7:0] add_802808;
  wire [7:0] sel_802809;
  wire [7:0] add_802812;
  wire [7:0] sel_802813;
  wire [7:0] add_802816;
  wire [7:0] sel_802817;
  wire [7:0] add_802820;
  wire [7:0] sel_802821;
  wire [7:0] add_802824;
  wire [7:0] sel_802825;
  wire [7:0] add_802828;
  wire [7:0] sel_802829;
  wire [7:0] add_802832;
  wire [7:0] sel_802833;
  wire [7:0] add_802836;
  wire [7:0] sel_802837;
  wire [7:0] add_802840;
  wire [7:0] sel_802841;
  wire [7:0] add_802844;
  wire [7:0] sel_802845;
  wire [7:0] add_802848;
  wire [7:0] sel_802849;
  wire [7:0] add_802852;
  wire [7:0] sel_802853;
  wire [7:0] add_802856;
  wire [7:0] sel_802857;
  wire [7:0] add_802860;
  wire [7:0] sel_802861;
  wire [7:0] add_802865;
  wire [15:0] array_index_802866;
  wire [7:0] sel_802867;
  wire [7:0] add_802870;
  wire [7:0] sel_802871;
  wire [7:0] add_802874;
  wire [7:0] sel_802875;
  wire [7:0] add_802878;
  wire [7:0] sel_802879;
  wire [7:0] add_802882;
  wire [7:0] sel_802883;
  wire [7:0] add_802886;
  wire [7:0] sel_802887;
  wire [7:0] add_802890;
  wire [7:0] sel_802891;
  wire [7:0] add_802894;
  wire [7:0] sel_802895;
  wire [7:0] add_802898;
  wire [7:0] sel_802899;
  wire [7:0] add_802902;
  wire [7:0] sel_802903;
  wire [7:0] add_802906;
  wire [7:0] sel_802907;
  wire [7:0] add_802910;
  wire [7:0] sel_802911;
  wire [7:0] add_802914;
  wire [7:0] sel_802915;
  wire [7:0] add_802918;
  wire [7:0] sel_802919;
  wire [7:0] add_802922;
  wire [7:0] sel_802923;
  wire [7:0] add_802926;
  wire [7:0] sel_802927;
  wire [7:0] add_802930;
  wire [7:0] sel_802931;
  wire [7:0] add_802934;
  wire [7:0] sel_802935;
  wire [7:0] add_802938;
  wire [7:0] sel_802939;
  wire [7:0] add_802942;
  wire [7:0] sel_802943;
  wire [7:0] add_802946;
  wire [7:0] sel_802947;
  wire [7:0] add_802950;
  wire [7:0] sel_802951;
  wire [7:0] add_802954;
  wire [7:0] sel_802955;
  wire [7:0] add_802958;
  wire [7:0] sel_802959;
  wire [7:0] add_802962;
  wire [7:0] sel_802963;
  wire [7:0] add_802966;
  wire [7:0] sel_802967;
  wire [7:0] add_802970;
  wire [7:0] sel_802971;
  wire [7:0] add_802974;
  wire [7:0] sel_802975;
  wire [7:0] add_802978;
  wire [7:0] sel_802979;
  wire [7:0] add_802982;
  wire [7:0] sel_802983;
  wire [7:0] add_802986;
  wire [7:0] sel_802987;
  wire [7:0] add_802990;
  wire [7:0] sel_802991;
  wire [7:0] add_802994;
  wire [7:0] sel_802995;
  wire [7:0] add_802998;
  wire [7:0] sel_802999;
  wire [7:0] add_803002;
  wire [7:0] sel_803003;
  wire [7:0] add_803006;
  wire [7:0] sel_803007;
  wire [7:0] add_803010;
  wire [7:0] sel_803011;
  wire [7:0] add_803014;
  wire [7:0] sel_803015;
  wire [7:0] add_803018;
  wire [7:0] sel_803019;
  wire [7:0] add_803022;
  wire [7:0] sel_803023;
  wire [7:0] add_803026;
  wire [7:0] sel_803027;
  wire [7:0] add_803030;
  wire [7:0] sel_803031;
  wire [7:0] add_803034;
  wire [7:0] sel_803035;
  wire [7:0] add_803038;
  wire [7:0] sel_803039;
  wire [7:0] add_803042;
  wire [7:0] sel_803043;
  wire [7:0] add_803046;
  wire [7:0] sel_803047;
  wire [7:0] add_803050;
  wire [7:0] sel_803051;
  wire [7:0] add_803054;
  wire [7:0] sel_803055;
  wire [7:0] add_803058;
  wire [7:0] sel_803059;
  wire [7:0] add_803062;
  wire [7:0] sel_803063;
  wire [7:0] add_803066;
  wire [7:0] sel_803067;
  wire [7:0] add_803070;
  wire [7:0] sel_803071;
  wire [7:0] add_803074;
  wire [7:0] sel_803075;
  wire [7:0] add_803078;
  wire [7:0] sel_803079;
  wire [7:0] add_803082;
  wire [7:0] sel_803083;
  wire [7:0] add_803086;
  wire [7:0] sel_803087;
  wire [7:0] add_803090;
  wire [7:0] sel_803091;
  wire [7:0] add_803094;
  wire [7:0] sel_803095;
  wire [7:0] add_803098;
  wire [7:0] sel_803099;
  wire [7:0] add_803102;
  wire [7:0] sel_803103;
  wire [7:0] add_803106;
  wire [7:0] sel_803107;
  wire [7:0] add_803110;
  wire [7:0] sel_803111;
  wire [7:0] add_803114;
  wire [7:0] sel_803115;
  wire [7:0] add_803118;
  wire [7:0] sel_803119;
  wire [7:0] add_803122;
  wire [7:0] sel_803123;
  wire [7:0] add_803126;
  wire [7:0] sel_803127;
  wire [7:0] add_803130;
  wire [7:0] sel_803131;
  wire [7:0] add_803134;
  wire [7:0] sel_803135;
  wire [7:0] add_803138;
  wire [7:0] sel_803139;
  wire [7:0] add_803142;
  wire [7:0] sel_803143;
  wire [7:0] add_803146;
  wire [7:0] sel_803147;
  wire [7:0] add_803150;
  wire [7:0] sel_803151;
  wire [7:0] add_803154;
  wire [7:0] sel_803155;
  wire [7:0] add_803158;
  wire [7:0] sel_803159;
  wire [7:0] add_803162;
  wire [7:0] sel_803163;
  wire [7:0] add_803166;
  wire [7:0] sel_803167;
  wire [7:0] add_803170;
  wire [7:0] sel_803171;
  wire [7:0] add_803174;
  wire [7:0] sel_803175;
  wire [7:0] add_803178;
  wire [7:0] sel_803179;
  wire [7:0] add_803182;
  wire [7:0] sel_803183;
  wire [7:0] add_803186;
  wire [7:0] sel_803187;
  wire [7:0] add_803190;
  wire [7:0] sel_803191;
  wire [7:0] add_803194;
  wire [7:0] sel_803195;
  wire [7:0] add_803198;
  wire [7:0] sel_803199;
  wire [7:0] add_803202;
  wire [7:0] sel_803203;
  wire [7:0] add_803206;
  wire [7:0] sel_803207;
  wire [7:0] add_803210;
  wire [7:0] sel_803211;
  wire [7:0] add_803214;
  wire [7:0] sel_803215;
  wire [7:0] add_803218;
  wire [7:0] sel_803219;
  wire [7:0] add_803222;
  wire [7:0] sel_803223;
  wire [7:0] add_803227;
  wire [15:0] array_index_803228;
  wire [7:0] sel_803229;
  wire [7:0] add_803232;
  wire [7:0] sel_803233;
  wire [7:0] add_803236;
  wire [7:0] sel_803237;
  wire [7:0] add_803240;
  wire [7:0] sel_803241;
  wire [7:0] add_803244;
  wire [7:0] sel_803245;
  wire [7:0] add_803248;
  wire [7:0] sel_803249;
  wire [7:0] add_803252;
  wire [7:0] sel_803253;
  wire [7:0] add_803256;
  wire [7:0] sel_803257;
  wire [7:0] add_803260;
  wire [7:0] sel_803261;
  wire [7:0] add_803264;
  wire [7:0] sel_803265;
  wire [7:0] add_803268;
  wire [7:0] sel_803269;
  wire [7:0] add_803272;
  wire [7:0] sel_803273;
  wire [7:0] add_803276;
  wire [7:0] sel_803277;
  wire [7:0] add_803280;
  wire [7:0] sel_803281;
  wire [7:0] add_803284;
  wire [7:0] sel_803285;
  wire [7:0] add_803288;
  wire [7:0] sel_803289;
  wire [7:0] add_803292;
  wire [7:0] sel_803293;
  wire [7:0] add_803296;
  wire [7:0] sel_803297;
  wire [7:0] add_803300;
  wire [7:0] sel_803301;
  wire [7:0] add_803304;
  wire [7:0] sel_803305;
  wire [7:0] add_803308;
  wire [7:0] sel_803309;
  wire [7:0] add_803312;
  wire [7:0] sel_803313;
  wire [7:0] add_803316;
  wire [7:0] sel_803317;
  wire [7:0] add_803320;
  wire [7:0] sel_803321;
  wire [7:0] add_803324;
  wire [7:0] sel_803325;
  wire [7:0] add_803328;
  wire [7:0] sel_803329;
  wire [7:0] add_803332;
  wire [7:0] sel_803333;
  wire [7:0] add_803336;
  wire [7:0] sel_803337;
  wire [7:0] add_803340;
  wire [7:0] sel_803341;
  wire [7:0] add_803344;
  wire [7:0] sel_803345;
  wire [7:0] add_803348;
  wire [7:0] sel_803349;
  wire [7:0] add_803352;
  wire [7:0] sel_803353;
  wire [7:0] add_803356;
  wire [7:0] sel_803357;
  wire [7:0] add_803360;
  wire [7:0] sel_803361;
  wire [7:0] add_803364;
  wire [7:0] sel_803365;
  wire [7:0] add_803368;
  wire [7:0] sel_803369;
  wire [7:0] add_803372;
  wire [7:0] sel_803373;
  wire [7:0] add_803376;
  wire [7:0] sel_803377;
  wire [7:0] add_803380;
  wire [7:0] sel_803381;
  wire [7:0] add_803384;
  wire [7:0] sel_803385;
  wire [7:0] add_803388;
  wire [7:0] sel_803389;
  wire [7:0] add_803392;
  wire [7:0] sel_803393;
  wire [7:0] add_803396;
  wire [7:0] sel_803397;
  wire [7:0] add_803400;
  wire [7:0] sel_803401;
  wire [7:0] add_803404;
  wire [7:0] sel_803405;
  wire [7:0] add_803408;
  wire [7:0] sel_803409;
  wire [7:0] add_803412;
  wire [7:0] sel_803413;
  wire [7:0] add_803416;
  wire [7:0] sel_803417;
  wire [7:0] add_803420;
  wire [7:0] sel_803421;
  wire [7:0] add_803424;
  wire [7:0] sel_803425;
  wire [7:0] add_803428;
  wire [7:0] sel_803429;
  wire [7:0] add_803432;
  wire [7:0] sel_803433;
  wire [7:0] add_803436;
  wire [7:0] sel_803437;
  wire [7:0] add_803440;
  wire [7:0] sel_803441;
  wire [7:0] add_803444;
  wire [7:0] sel_803445;
  wire [7:0] add_803448;
  wire [7:0] sel_803449;
  wire [7:0] add_803452;
  wire [7:0] sel_803453;
  wire [7:0] add_803456;
  wire [7:0] sel_803457;
  wire [7:0] add_803460;
  wire [7:0] sel_803461;
  wire [7:0] add_803464;
  wire [7:0] sel_803465;
  wire [7:0] add_803468;
  wire [7:0] sel_803469;
  wire [7:0] add_803472;
  wire [7:0] sel_803473;
  wire [7:0] add_803476;
  wire [7:0] sel_803477;
  wire [7:0] add_803480;
  wire [7:0] sel_803481;
  wire [7:0] add_803484;
  wire [7:0] sel_803485;
  wire [7:0] add_803488;
  wire [7:0] sel_803489;
  wire [7:0] add_803492;
  wire [7:0] sel_803493;
  wire [7:0] add_803496;
  wire [7:0] sel_803497;
  wire [7:0] add_803500;
  wire [7:0] sel_803501;
  wire [7:0] add_803504;
  wire [7:0] sel_803505;
  wire [7:0] add_803508;
  wire [7:0] sel_803509;
  wire [7:0] add_803512;
  wire [7:0] sel_803513;
  wire [7:0] add_803516;
  wire [7:0] sel_803517;
  wire [7:0] add_803520;
  wire [7:0] sel_803521;
  wire [7:0] add_803524;
  wire [7:0] sel_803525;
  wire [7:0] add_803528;
  wire [7:0] sel_803529;
  wire [7:0] add_803532;
  wire [7:0] sel_803533;
  wire [7:0] add_803536;
  wire [7:0] sel_803537;
  wire [7:0] add_803540;
  wire [7:0] sel_803541;
  wire [7:0] add_803544;
  wire [7:0] sel_803545;
  wire [7:0] add_803548;
  wire [7:0] sel_803549;
  wire [7:0] add_803552;
  wire [7:0] sel_803553;
  wire [7:0] add_803556;
  wire [7:0] sel_803557;
  wire [7:0] add_803560;
  wire [7:0] sel_803561;
  wire [7:0] add_803564;
  wire [7:0] sel_803565;
  wire [7:0] add_803568;
  wire [7:0] sel_803569;
  wire [7:0] add_803572;
  wire [7:0] sel_803573;
  wire [7:0] add_803576;
  wire [7:0] sel_803577;
  wire [7:0] add_803580;
  wire [7:0] sel_803581;
  wire [7:0] add_803584;
  wire [7:0] sel_803585;
  wire [7:0] add_803589;
  wire [15:0] array_index_803590;
  wire [7:0] sel_803591;
  wire [7:0] add_803594;
  wire [7:0] sel_803595;
  wire [7:0] add_803598;
  wire [7:0] sel_803599;
  wire [7:0] add_803602;
  wire [7:0] sel_803603;
  wire [7:0] add_803606;
  wire [7:0] sel_803607;
  wire [7:0] add_803610;
  wire [7:0] sel_803611;
  wire [7:0] add_803614;
  wire [7:0] sel_803615;
  wire [7:0] add_803618;
  wire [7:0] sel_803619;
  wire [7:0] add_803622;
  wire [7:0] sel_803623;
  wire [7:0] add_803626;
  wire [7:0] sel_803627;
  wire [7:0] add_803630;
  wire [7:0] sel_803631;
  wire [7:0] add_803634;
  wire [7:0] sel_803635;
  wire [7:0] add_803638;
  wire [7:0] sel_803639;
  wire [7:0] add_803642;
  wire [7:0] sel_803643;
  wire [7:0] add_803646;
  wire [7:0] sel_803647;
  wire [7:0] add_803650;
  wire [7:0] sel_803651;
  wire [7:0] add_803654;
  wire [7:0] sel_803655;
  wire [7:0] add_803658;
  wire [7:0] sel_803659;
  wire [7:0] add_803662;
  wire [7:0] sel_803663;
  wire [7:0] add_803666;
  wire [7:0] sel_803667;
  wire [7:0] add_803670;
  wire [7:0] sel_803671;
  wire [7:0] add_803674;
  wire [7:0] sel_803675;
  wire [7:0] add_803678;
  wire [7:0] sel_803679;
  wire [7:0] add_803682;
  wire [7:0] sel_803683;
  wire [7:0] add_803686;
  wire [7:0] sel_803687;
  wire [7:0] add_803690;
  wire [7:0] sel_803691;
  wire [7:0] add_803694;
  wire [7:0] sel_803695;
  wire [7:0] add_803698;
  wire [7:0] sel_803699;
  wire [7:0] add_803702;
  wire [7:0] sel_803703;
  wire [7:0] add_803706;
  wire [7:0] sel_803707;
  wire [7:0] add_803710;
  wire [7:0] sel_803711;
  wire [7:0] add_803714;
  wire [7:0] sel_803715;
  wire [7:0] add_803718;
  wire [7:0] sel_803719;
  wire [7:0] add_803722;
  wire [7:0] sel_803723;
  wire [7:0] add_803726;
  wire [7:0] sel_803727;
  wire [7:0] add_803730;
  wire [7:0] sel_803731;
  wire [7:0] add_803734;
  wire [7:0] sel_803735;
  wire [7:0] add_803738;
  wire [7:0] sel_803739;
  wire [7:0] add_803742;
  wire [7:0] sel_803743;
  wire [7:0] add_803746;
  wire [7:0] sel_803747;
  wire [7:0] add_803750;
  wire [7:0] sel_803751;
  wire [7:0] add_803754;
  wire [7:0] sel_803755;
  wire [7:0] add_803758;
  wire [7:0] sel_803759;
  wire [7:0] add_803762;
  wire [7:0] sel_803763;
  wire [7:0] add_803766;
  wire [7:0] sel_803767;
  wire [7:0] add_803770;
  wire [7:0] sel_803771;
  wire [7:0] add_803774;
  wire [7:0] sel_803775;
  wire [7:0] add_803778;
  wire [7:0] sel_803779;
  wire [7:0] add_803782;
  wire [7:0] sel_803783;
  wire [7:0] add_803786;
  wire [7:0] sel_803787;
  wire [7:0] add_803790;
  wire [7:0] sel_803791;
  wire [7:0] add_803794;
  wire [7:0] sel_803795;
  wire [7:0] add_803798;
  wire [7:0] sel_803799;
  wire [7:0] add_803802;
  wire [7:0] sel_803803;
  wire [7:0] add_803806;
  wire [7:0] sel_803807;
  wire [7:0] add_803810;
  wire [7:0] sel_803811;
  wire [7:0] add_803814;
  wire [7:0] sel_803815;
  wire [7:0] add_803818;
  wire [7:0] sel_803819;
  wire [7:0] add_803822;
  wire [7:0] sel_803823;
  wire [7:0] add_803826;
  wire [7:0] sel_803827;
  wire [7:0] add_803830;
  wire [7:0] sel_803831;
  wire [7:0] add_803834;
  wire [7:0] sel_803835;
  wire [7:0] add_803838;
  wire [7:0] sel_803839;
  wire [7:0] add_803842;
  wire [7:0] sel_803843;
  wire [7:0] add_803846;
  wire [7:0] sel_803847;
  wire [7:0] add_803850;
  wire [7:0] sel_803851;
  wire [7:0] add_803854;
  wire [7:0] sel_803855;
  wire [7:0] add_803858;
  wire [7:0] sel_803859;
  wire [7:0] add_803862;
  wire [7:0] sel_803863;
  wire [7:0] add_803866;
  wire [7:0] sel_803867;
  wire [7:0] add_803870;
  wire [7:0] sel_803871;
  wire [7:0] add_803874;
  wire [7:0] sel_803875;
  wire [7:0] add_803878;
  wire [7:0] sel_803879;
  wire [7:0] add_803882;
  wire [7:0] sel_803883;
  wire [7:0] add_803886;
  wire [7:0] sel_803887;
  wire [7:0] add_803890;
  wire [7:0] sel_803891;
  wire [7:0] add_803894;
  wire [7:0] sel_803895;
  wire [7:0] add_803898;
  wire [7:0] sel_803899;
  wire [7:0] add_803902;
  wire [7:0] sel_803903;
  wire [7:0] add_803906;
  wire [7:0] sel_803907;
  wire [7:0] add_803910;
  wire [7:0] sel_803911;
  wire [7:0] add_803914;
  wire [7:0] sel_803915;
  wire [7:0] add_803918;
  wire [7:0] sel_803919;
  wire [7:0] add_803922;
  wire [7:0] sel_803923;
  wire [7:0] add_803926;
  wire [7:0] sel_803927;
  wire [7:0] add_803930;
  wire [7:0] sel_803931;
  wire [7:0] add_803934;
  wire [7:0] sel_803935;
  wire [7:0] add_803938;
  wire [7:0] sel_803939;
  wire [7:0] add_803942;
  wire [7:0] sel_803943;
  wire [7:0] add_803946;
  wire [7:0] sel_803947;
  wire [7:0] add_803951;
  wire [15:0] array_index_803952;
  wire [7:0] sel_803953;
  wire [7:0] add_803956;
  wire [7:0] sel_803957;
  wire [7:0] add_803960;
  wire [7:0] sel_803961;
  wire [7:0] add_803964;
  wire [7:0] sel_803965;
  wire [7:0] add_803968;
  wire [7:0] sel_803969;
  wire [7:0] add_803972;
  wire [7:0] sel_803973;
  wire [7:0] add_803976;
  wire [7:0] sel_803977;
  wire [7:0] add_803980;
  wire [7:0] sel_803981;
  wire [7:0] add_803984;
  wire [7:0] sel_803985;
  wire [7:0] add_803988;
  wire [7:0] sel_803989;
  wire [7:0] add_803992;
  wire [7:0] sel_803993;
  wire [7:0] add_803996;
  wire [7:0] sel_803997;
  wire [7:0] add_804000;
  wire [7:0] sel_804001;
  wire [7:0] add_804004;
  wire [7:0] sel_804005;
  wire [7:0] add_804008;
  wire [7:0] sel_804009;
  wire [7:0] add_804012;
  wire [7:0] sel_804013;
  wire [7:0] add_804016;
  wire [7:0] sel_804017;
  wire [7:0] add_804020;
  wire [7:0] sel_804021;
  wire [7:0] add_804024;
  wire [7:0] sel_804025;
  wire [7:0] add_804028;
  wire [7:0] sel_804029;
  wire [7:0] add_804032;
  wire [7:0] sel_804033;
  wire [7:0] add_804036;
  wire [7:0] sel_804037;
  wire [7:0] add_804040;
  wire [7:0] sel_804041;
  wire [7:0] add_804044;
  wire [7:0] sel_804045;
  wire [7:0] add_804048;
  wire [7:0] sel_804049;
  wire [7:0] add_804052;
  wire [7:0] sel_804053;
  wire [7:0] add_804056;
  wire [7:0] sel_804057;
  wire [7:0] add_804060;
  wire [7:0] sel_804061;
  wire [7:0] add_804064;
  wire [7:0] sel_804065;
  wire [7:0] add_804068;
  wire [7:0] sel_804069;
  wire [7:0] add_804072;
  wire [7:0] sel_804073;
  wire [7:0] add_804076;
  wire [7:0] sel_804077;
  wire [7:0] add_804080;
  wire [7:0] sel_804081;
  wire [7:0] add_804084;
  wire [7:0] sel_804085;
  wire [7:0] add_804088;
  wire [7:0] sel_804089;
  wire [7:0] add_804092;
  wire [7:0] sel_804093;
  wire [7:0] add_804096;
  wire [7:0] sel_804097;
  wire [7:0] add_804100;
  wire [7:0] sel_804101;
  wire [7:0] add_804104;
  wire [7:0] sel_804105;
  wire [7:0] add_804108;
  wire [7:0] sel_804109;
  wire [7:0] add_804112;
  wire [7:0] sel_804113;
  wire [7:0] add_804116;
  wire [7:0] sel_804117;
  wire [7:0] add_804120;
  wire [7:0] sel_804121;
  wire [7:0] add_804124;
  wire [7:0] sel_804125;
  wire [7:0] add_804128;
  wire [7:0] sel_804129;
  wire [7:0] add_804132;
  wire [7:0] sel_804133;
  wire [7:0] add_804136;
  wire [7:0] sel_804137;
  wire [7:0] add_804140;
  wire [7:0] sel_804141;
  wire [7:0] add_804144;
  wire [7:0] sel_804145;
  wire [7:0] add_804148;
  wire [7:0] sel_804149;
  wire [7:0] add_804152;
  wire [7:0] sel_804153;
  wire [7:0] add_804156;
  wire [7:0] sel_804157;
  wire [7:0] add_804160;
  wire [7:0] sel_804161;
  wire [7:0] add_804164;
  wire [7:0] sel_804165;
  wire [7:0] add_804168;
  wire [7:0] sel_804169;
  wire [7:0] add_804172;
  wire [7:0] sel_804173;
  wire [7:0] add_804176;
  wire [7:0] sel_804177;
  wire [7:0] add_804180;
  wire [7:0] sel_804181;
  wire [7:0] add_804184;
  wire [7:0] sel_804185;
  wire [7:0] add_804188;
  wire [7:0] sel_804189;
  wire [7:0] add_804192;
  wire [7:0] sel_804193;
  wire [7:0] add_804196;
  wire [7:0] sel_804197;
  wire [7:0] add_804200;
  wire [7:0] sel_804201;
  wire [7:0] add_804204;
  wire [7:0] sel_804205;
  wire [7:0] add_804208;
  wire [7:0] sel_804209;
  wire [7:0] add_804212;
  wire [7:0] sel_804213;
  wire [7:0] add_804216;
  wire [7:0] sel_804217;
  wire [7:0] add_804220;
  wire [7:0] sel_804221;
  wire [7:0] add_804224;
  wire [7:0] sel_804225;
  wire [7:0] add_804228;
  wire [7:0] sel_804229;
  wire [7:0] add_804232;
  wire [7:0] sel_804233;
  wire [7:0] add_804236;
  wire [7:0] sel_804237;
  wire [7:0] add_804240;
  wire [7:0] sel_804241;
  wire [7:0] add_804244;
  wire [7:0] sel_804245;
  wire [7:0] add_804248;
  wire [7:0] sel_804249;
  wire [7:0] add_804252;
  wire [7:0] sel_804253;
  wire [7:0] add_804256;
  wire [7:0] sel_804257;
  wire [7:0] add_804260;
  wire [7:0] sel_804261;
  wire [7:0] add_804264;
  wire [7:0] sel_804265;
  wire [7:0] add_804268;
  wire [7:0] sel_804269;
  wire [7:0] add_804272;
  wire [7:0] sel_804273;
  wire [7:0] add_804276;
  wire [7:0] sel_804277;
  wire [7:0] add_804280;
  wire [7:0] sel_804281;
  wire [7:0] add_804284;
  wire [7:0] sel_804285;
  wire [7:0] add_804288;
  wire [7:0] sel_804289;
  wire [7:0] add_804292;
  wire [7:0] sel_804293;
  wire [7:0] add_804296;
  wire [7:0] sel_804297;
  wire [7:0] add_804300;
  wire [7:0] sel_804301;
  wire [7:0] add_804304;
  wire [7:0] sel_804305;
  wire [7:0] add_804308;
  wire [7:0] sel_804309;
  wire [7:0] add_804313;
  wire [15:0] array_index_804314;
  wire [7:0] sel_804315;
  wire [7:0] add_804318;
  wire [7:0] sel_804319;
  wire [7:0] add_804322;
  wire [7:0] sel_804323;
  wire [7:0] add_804326;
  wire [7:0] sel_804327;
  wire [7:0] add_804330;
  wire [7:0] sel_804331;
  wire [7:0] add_804334;
  wire [7:0] sel_804335;
  wire [7:0] add_804338;
  wire [7:0] sel_804339;
  wire [7:0] add_804342;
  wire [7:0] sel_804343;
  wire [7:0] add_804346;
  wire [7:0] sel_804347;
  wire [7:0] add_804350;
  wire [7:0] sel_804351;
  wire [7:0] add_804354;
  wire [7:0] sel_804355;
  wire [7:0] add_804358;
  wire [7:0] sel_804359;
  wire [7:0] add_804362;
  wire [7:0] sel_804363;
  wire [7:0] add_804366;
  wire [7:0] sel_804367;
  wire [7:0] add_804370;
  wire [7:0] sel_804371;
  wire [7:0] add_804374;
  wire [7:0] sel_804375;
  wire [7:0] add_804378;
  wire [7:0] sel_804379;
  wire [7:0] add_804382;
  wire [7:0] sel_804383;
  wire [7:0] add_804386;
  wire [7:0] sel_804387;
  wire [7:0] add_804390;
  wire [7:0] sel_804391;
  wire [7:0] add_804394;
  wire [7:0] sel_804395;
  wire [7:0] add_804398;
  wire [7:0] sel_804399;
  wire [7:0] add_804402;
  wire [7:0] sel_804403;
  wire [7:0] add_804406;
  wire [7:0] sel_804407;
  wire [7:0] add_804410;
  wire [7:0] sel_804411;
  wire [7:0] add_804414;
  wire [7:0] sel_804415;
  wire [7:0] add_804418;
  wire [7:0] sel_804419;
  wire [7:0] add_804422;
  wire [7:0] sel_804423;
  wire [7:0] add_804426;
  wire [7:0] sel_804427;
  wire [7:0] add_804430;
  wire [7:0] sel_804431;
  wire [7:0] add_804434;
  wire [7:0] sel_804435;
  wire [7:0] add_804438;
  wire [7:0] sel_804439;
  wire [7:0] add_804442;
  wire [7:0] sel_804443;
  wire [7:0] add_804446;
  wire [7:0] sel_804447;
  wire [7:0] add_804450;
  wire [7:0] sel_804451;
  wire [7:0] add_804454;
  wire [7:0] sel_804455;
  wire [7:0] add_804458;
  wire [7:0] sel_804459;
  wire [7:0] add_804462;
  wire [7:0] sel_804463;
  wire [7:0] add_804466;
  wire [7:0] sel_804467;
  wire [7:0] add_804470;
  wire [7:0] sel_804471;
  wire [7:0] add_804474;
  wire [7:0] sel_804475;
  wire [7:0] add_804478;
  wire [7:0] sel_804479;
  wire [7:0] add_804482;
  wire [7:0] sel_804483;
  wire [7:0] add_804486;
  wire [7:0] sel_804487;
  wire [7:0] add_804490;
  wire [7:0] sel_804491;
  wire [7:0] add_804494;
  wire [7:0] sel_804495;
  wire [7:0] add_804498;
  wire [7:0] sel_804499;
  wire [7:0] add_804502;
  wire [7:0] sel_804503;
  wire [7:0] add_804506;
  wire [7:0] sel_804507;
  wire [7:0] add_804510;
  wire [7:0] sel_804511;
  wire [7:0] add_804514;
  wire [7:0] sel_804515;
  wire [7:0] add_804518;
  wire [7:0] sel_804519;
  wire [7:0] add_804522;
  wire [7:0] sel_804523;
  wire [7:0] add_804526;
  wire [7:0] sel_804527;
  wire [7:0] add_804530;
  wire [7:0] sel_804531;
  wire [7:0] add_804534;
  wire [7:0] sel_804535;
  wire [7:0] add_804538;
  wire [7:0] sel_804539;
  wire [7:0] add_804542;
  wire [7:0] sel_804543;
  wire [7:0] add_804546;
  wire [7:0] sel_804547;
  wire [7:0] add_804550;
  wire [7:0] sel_804551;
  wire [7:0] add_804554;
  wire [7:0] sel_804555;
  wire [7:0] add_804558;
  wire [7:0] sel_804559;
  wire [7:0] add_804562;
  wire [7:0] sel_804563;
  wire [7:0] add_804566;
  wire [7:0] sel_804567;
  wire [7:0] add_804570;
  wire [7:0] sel_804571;
  wire [7:0] add_804574;
  wire [7:0] sel_804575;
  wire [7:0] add_804578;
  wire [7:0] sel_804579;
  wire [7:0] add_804582;
  wire [7:0] sel_804583;
  wire [7:0] add_804586;
  wire [7:0] sel_804587;
  wire [7:0] add_804590;
  wire [7:0] sel_804591;
  wire [7:0] add_804594;
  wire [7:0] sel_804595;
  wire [7:0] add_804598;
  wire [7:0] sel_804599;
  wire [7:0] add_804602;
  wire [7:0] sel_804603;
  wire [7:0] add_804606;
  wire [7:0] sel_804607;
  wire [7:0] add_804610;
  wire [7:0] sel_804611;
  wire [7:0] add_804614;
  wire [7:0] sel_804615;
  wire [7:0] add_804618;
  wire [7:0] sel_804619;
  wire [7:0] add_804622;
  wire [7:0] sel_804623;
  wire [7:0] add_804626;
  wire [7:0] sel_804627;
  wire [7:0] add_804630;
  wire [7:0] sel_804631;
  wire [7:0] add_804634;
  wire [7:0] sel_804635;
  wire [7:0] add_804638;
  wire [7:0] sel_804639;
  wire [7:0] add_804642;
  wire [7:0] sel_804643;
  wire [7:0] add_804646;
  wire [7:0] sel_804647;
  wire [7:0] add_804650;
  wire [7:0] sel_804651;
  wire [7:0] add_804654;
  wire [7:0] sel_804655;
  wire [7:0] add_804658;
  wire [7:0] sel_804659;
  wire [7:0] add_804662;
  wire [7:0] sel_804663;
  wire [7:0] add_804666;
  wire [7:0] sel_804667;
  wire [7:0] add_804670;
  wire [7:0] sel_804671;
  wire [7:0] add_804675;
  wire [15:0] array_index_804676;
  wire [7:0] sel_804677;
  wire [7:0] add_804680;
  wire [7:0] sel_804681;
  wire [7:0] add_804684;
  wire [7:0] sel_804685;
  wire [7:0] add_804688;
  wire [7:0] sel_804689;
  wire [7:0] add_804692;
  wire [7:0] sel_804693;
  wire [7:0] add_804696;
  wire [7:0] sel_804697;
  wire [7:0] add_804700;
  wire [7:0] sel_804701;
  wire [7:0] add_804704;
  wire [7:0] sel_804705;
  wire [7:0] add_804708;
  wire [7:0] sel_804709;
  wire [7:0] add_804712;
  wire [7:0] sel_804713;
  wire [7:0] add_804716;
  wire [7:0] sel_804717;
  wire [7:0] add_804720;
  wire [7:0] sel_804721;
  wire [7:0] add_804724;
  wire [7:0] sel_804725;
  wire [7:0] add_804728;
  wire [7:0] sel_804729;
  wire [7:0] add_804732;
  wire [7:0] sel_804733;
  wire [7:0] add_804736;
  wire [7:0] sel_804737;
  wire [7:0] add_804740;
  wire [7:0] sel_804741;
  wire [7:0] add_804744;
  wire [7:0] sel_804745;
  wire [7:0] add_804748;
  wire [7:0] sel_804749;
  wire [7:0] add_804752;
  wire [7:0] sel_804753;
  wire [7:0] add_804756;
  wire [7:0] sel_804757;
  wire [7:0] add_804760;
  wire [7:0] sel_804761;
  wire [7:0] add_804764;
  wire [7:0] sel_804765;
  wire [7:0] add_804768;
  wire [7:0] sel_804769;
  wire [7:0] add_804772;
  wire [7:0] sel_804773;
  wire [7:0] add_804776;
  wire [7:0] sel_804777;
  wire [7:0] add_804780;
  wire [7:0] sel_804781;
  wire [7:0] add_804784;
  wire [7:0] sel_804785;
  wire [7:0] add_804788;
  wire [7:0] sel_804789;
  wire [7:0] add_804792;
  wire [7:0] sel_804793;
  wire [7:0] add_804796;
  wire [7:0] sel_804797;
  wire [7:0] add_804800;
  wire [7:0] sel_804801;
  wire [7:0] add_804804;
  wire [7:0] sel_804805;
  wire [7:0] add_804808;
  wire [7:0] sel_804809;
  wire [7:0] add_804812;
  wire [7:0] sel_804813;
  wire [7:0] add_804816;
  wire [7:0] sel_804817;
  wire [7:0] add_804820;
  wire [7:0] sel_804821;
  wire [7:0] add_804824;
  wire [7:0] sel_804825;
  wire [7:0] add_804828;
  wire [7:0] sel_804829;
  wire [7:0] add_804832;
  wire [7:0] sel_804833;
  wire [7:0] add_804836;
  wire [7:0] sel_804837;
  wire [7:0] add_804840;
  wire [7:0] sel_804841;
  wire [7:0] add_804844;
  wire [7:0] sel_804845;
  wire [7:0] add_804848;
  wire [7:0] sel_804849;
  wire [7:0] add_804852;
  wire [7:0] sel_804853;
  wire [7:0] add_804856;
  wire [7:0] sel_804857;
  wire [7:0] add_804860;
  wire [7:0] sel_804861;
  wire [7:0] add_804864;
  wire [7:0] sel_804865;
  wire [7:0] add_804868;
  wire [7:0] sel_804869;
  wire [7:0] add_804872;
  wire [7:0] sel_804873;
  wire [7:0] add_804876;
  wire [7:0] sel_804877;
  wire [7:0] add_804880;
  wire [7:0] sel_804881;
  wire [7:0] add_804884;
  wire [7:0] sel_804885;
  wire [7:0] add_804888;
  wire [7:0] sel_804889;
  wire [7:0] add_804892;
  wire [7:0] sel_804893;
  wire [7:0] add_804896;
  wire [7:0] sel_804897;
  wire [7:0] add_804900;
  wire [7:0] sel_804901;
  wire [7:0] add_804904;
  wire [7:0] sel_804905;
  wire [7:0] add_804908;
  wire [7:0] sel_804909;
  wire [7:0] add_804912;
  wire [7:0] sel_804913;
  wire [7:0] add_804916;
  wire [7:0] sel_804917;
  wire [7:0] add_804920;
  wire [7:0] sel_804921;
  wire [7:0] add_804924;
  wire [7:0] sel_804925;
  wire [7:0] add_804928;
  wire [7:0] sel_804929;
  wire [7:0] add_804932;
  wire [7:0] sel_804933;
  wire [7:0] add_804936;
  wire [7:0] sel_804937;
  wire [7:0] add_804940;
  wire [7:0] sel_804941;
  wire [7:0] add_804944;
  wire [7:0] sel_804945;
  wire [7:0] add_804948;
  wire [7:0] sel_804949;
  wire [7:0] add_804952;
  wire [7:0] sel_804953;
  wire [7:0] add_804956;
  wire [7:0] sel_804957;
  wire [7:0] add_804960;
  wire [7:0] sel_804961;
  wire [7:0] add_804964;
  wire [7:0] sel_804965;
  wire [7:0] add_804968;
  wire [7:0] sel_804969;
  wire [7:0] add_804972;
  wire [7:0] sel_804973;
  wire [7:0] add_804976;
  wire [7:0] sel_804977;
  wire [7:0] add_804980;
  wire [7:0] sel_804981;
  wire [7:0] add_804984;
  wire [7:0] sel_804985;
  wire [7:0] add_804988;
  wire [7:0] sel_804989;
  wire [7:0] add_804992;
  wire [7:0] sel_804993;
  wire [7:0] add_804996;
  wire [7:0] sel_804997;
  wire [7:0] add_805000;
  wire [7:0] sel_805001;
  wire [7:0] add_805004;
  wire [7:0] sel_805005;
  wire [7:0] add_805008;
  wire [7:0] sel_805009;
  wire [7:0] add_805012;
  wire [7:0] sel_805013;
  wire [7:0] add_805016;
  wire [7:0] sel_805017;
  wire [7:0] add_805020;
  wire [7:0] sel_805021;
  wire [7:0] add_805024;
  wire [7:0] sel_805025;
  wire [7:0] add_805028;
  wire [7:0] sel_805029;
  wire [7:0] add_805032;
  wire [7:0] sel_805033;
  wire [7:0] add_805037;
  wire [15:0] array_index_805038;
  wire [7:0] sel_805039;
  wire [7:0] add_805042;
  wire [7:0] sel_805043;
  wire [7:0] add_805046;
  wire [7:0] sel_805047;
  wire [7:0] add_805050;
  wire [7:0] sel_805051;
  wire [7:0] add_805054;
  wire [7:0] sel_805055;
  wire [7:0] add_805058;
  wire [7:0] sel_805059;
  wire [7:0] add_805062;
  wire [7:0] sel_805063;
  wire [7:0] add_805066;
  wire [7:0] sel_805067;
  wire [7:0] add_805070;
  wire [7:0] sel_805071;
  wire [7:0] add_805074;
  wire [7:0] sel_805075;
  wire [7:0] add_805078;
  wire [7:0] sel_805079;
  wire [7:0] add_805082;
  wire [7:0] sel_805083;
  wire [7:0] add_805086;
  wire [7:0] sel_805087;
  wire [7:0] add_805090;
  wire [7:0] sel_805091;
  wire [7:0] add_805094;
  wire [7:0] sel_805095;
  wire [7:0] add_805098;
  wire [7:0] sel_805099;
  wire [7:0] add_805102;
  wire [7:0] sel_805103;
  wire [7:0] add_805106;
  wire [7:0] sel_805107;
  wire [7:0] add_805110;
  wire [7:0] sel_805111;
  wire [7:0] add_805114;
  wire [7:0] sel_805115;
  wire [7:0] add_805118;
  wire [7:0] sel_805119;
  wire [7:0] add_805122;
  wire [7:0] sel_805123;
  wire [7:0] add_805126;
  wire [7:0] sel_805127;
  wire [7:0] add_805130;
  wire [7:0] sel_805131;
  wire [7:0] add_805134;
  wire [7:0] sel_805135;
  wire [7:0] add_805138;
  wire [7:0] sel_805139;
  wire [7:0] add_805142;
  wire [7:0] sel_805143;
  wire [7:0] add_805146;
  wire [7:0] sel_805147;
  wire [7:0] add_805150;
  wire [7:0] sel_805151;
  wire [7:0] add_805154;
  wire [7:0] sel_805155;
  wire [7:0] add_805158;
  wire [7:0] sel_805159;
  wire [7:0] add_805162;
  wire [7:0] sel_805163;
  wire [7:0] add_805166;
  wire [7:0] sel_805167;
  wire [7:0] add_805170;
  wire [7:0] sel_805171;
  wire [7:0] add_805174;
  wire [7:0] sel_805175;
  wire [7:0] add_805178;
  wire [7:0] sel_805179;
  wire [7:0] add_805182;
  wire [7:0] sel_805183;
  wire [7:0] add_805186;
  wire [7:0] sel_805187;
  wire [7:0] add_805190;
  wire [7:0] sel_805191;
  wire [7:0] add_805194;
  wire [7:0] sel_805195;
  wire [7:0] add_805198;
  wire [7:0] sel_805199;
  wire [7:0] add_805202;
  wire [7:0] sel_805203;
  wire [7:0] add_805206;
  wire [7:0] sel_805207;
  wire [7:0] add_805210;
  wire [7:0] sel_805211;
  wire [7:0] add_805214;
  wire [7:0] sel_805215;
  wire [7:0] add_805218;
  wire [7:0] sel_805219;
  wire [7:0] add_805222;
  wire [7:0] sel_805223;
  wire [7:0] add_805226;
  wire [7:0] sel_805227;
  wire [7:0] add_805230;
  wire [7:0] sel_805231;
  wire [7:0] add_805234;
  wire [7:0] sel_805235;
  wire [7:0] add_805238;
  wire [7:0] sel_805239;
  wire [7:0] add_805242;
  wire [7:0] sel_805243;
  wire [7:0] add_805246;
  wire [7:0] sel_805247;
  wire [7:0] add_805250;
  wire [7:0] sel_805251;
  wire [7:0] add_805254;
  wire [7:0] sel_805255;
  wire [7:0] add_805258;
  wire [7:0] sel_805259;
  wire [7:0] add_805262;
  wire [7:0] sel_805263;
  wire [7:0] add_805266;
  wire [7:0] sel_805267;
  wire [7:0] add_805270;
  wire [7:0] sel_805271;
  wire [7:0] add_805274;
  wire [7:0] sel_805275;
  wire [7:0] add_805278;
  wire [7:0] sel_805279;
  wire [7:0] add_805282;
  wire [7:0] sel_805283;
  wire [7:0] add_805286;
  wire [7:0] sel_805287;
  wire [7:0] add_805290;
  wire [7:0] sel_805291;
  wire [7:0] add_805294;
  wire [7:0] sel_805295;
  wire [7:0] add_805298;
  wire [7:0] sel_805299;
  wire [7:0] add_805302;
  wire [7:0] sel_805303;
  wire [7:0] add_805306;
  wire [7:0] sel_805307;
  wire [7:0] add_805310;
  wire [7:0] sel_805311;
  wire [7:0] add_805314;
  wire [7:0] sel_805315;
  wire [7:0] add_805318;
  wire [7:0] sel_805319;
  wire [7:0] add_805322;
  wire [7:0] sel_805323;
  wire [7:0] add_805326;
  wire [7:0] sel_805327;
  wire [7:0] add_805330;
  wire [7:0] sel_805331;
  wire [7:0] add_805334;
  wire [7:0] sel_805335;
  wire [7:0] add_805338;
  wire [7:0] sel_805339;
  wire [7:0] add_805342;
  wire [7:0] sel_805343;
  wire [7:0] add_805346;
  wire [7:0] sel_805347;
  wire [7:0] add_805350;
  wire [7:0] sel_805351;
  wire [7:0] add_805354;
  wire [7:0] sel_805355;
  wire [7:0] add_805358;
  wire [7:0] sel_805359;
  wire [7:0] add_805362;
  wire [7:0] sel_805363;
  wire [7:0] add_805366;
  wire [7:0] sel_805367;
  wire [7:0] add_805370;
  wire [7:0] sel_805371;
  wire [7:0] add_805374;
  wire [7:0] sel_805375;
  wire [7:0] add_805378;
  wire [7:0] sel_805379;
  wire [7:0] add_805382;
  wire [7:0] sel_805383;
  wire [7:0] add_805386;
  wire [7:0] sel_805387;
  wire [7:0] add_805390;
  wire [7:0] sel_805391;
  wire [7:0] add_805394;
  wire [7:0] sel_805395;
  wire [7:0] add_805398;
  assign array_index_772631 = set1_unflattened[7'h00];
  assign array_index_772632 = set2_unflattened[7'h00];
  assign array_index_772636 = set2_unflattened[7'h01];
  assign concat_772637 = {1'h0, array_index_772631 == array_index_772632};
  assign add_772640 = concat_772637 + 2'h1;
  assign array_index_772644 = set2_unflattened[7'h02];
  assign concat_772645 = {1'h0, array_index_772631 == array_index_772636 ? add_772640 : concat_772637};
  assign add_772648 = concat_772645 + 3'h1;
  assign array_index_772652 = set2_unflattened[7'h03];
  assign concat_772653 = {1'h0, array_index_772631 == array_index_772644 ? add_772648 : concat_772645};
  assign add_772656 = concat_772653 + 4'h1;
  assign array_index_772660 = set2_unflattened[7'h04];
  assign concat_772661 = {1'h0, array_index_772631 == array_index_772652 ? add_772656 : concat_772653};
  assign add_772664 = concat_772661 + 5'h01;
  assign array_index_772668 = set2_unflattened[7'h05];
  assign concat_772669 = {1'h0, array_index_772631 == array_index_772660 ? add_772664 : concat_772661};
  assign add_772672 = concat_772669 + 6'h01;
  assign array_index_772676 = set2_unflattened[7'h06];
  assign concat_772677 = {1'h0, array_index_772631 == array_index_772668 ? add_772672 : concat_772669};
  assign add_772680 = concat_772677 + 7'h01;
  assign array_index_772684 = set2_unflattened[7'h07];
  assign concat_772685 = {1'h0, array_index_772631 == array_index_772676 ? add_772680 : concat_772677};
  assign add_772689 = concat_772685 + 8'h01;
  assign array_index_772690 = set2_unflattened[7'h08];
  assign sel_772691 = array_index_772631 == array_index_772684 ? add_772689 : concat_772685;
  assign add_772695 = sel_772691 + 8'h01;
  assign array_index_772696 = set2_unflattened[7'h09];
  assign sel_772697 = array_index_772631 == array_index_772690 ? add_772695 : sel_772691;
  assign add_772701 = sel_772697 + 8'h01;
  assign array_index_772702 = set2_unflattened[7'h0a];
  assign sel_772703 = array_index_772631 == array_index_772696 ? add_772701 : sel_772697;
  assign add_772707 = sel_772703 + 8'h01;
  assign array_index_772708 = set2_unflattened[7'h0b];
  assign sel_772709 = array_index_772631 == array_index_772702 ? add_772707 : sel_772703;
  assign add_772713 = sel_772709 + 8'h01;
  assign array_index_772714 = set2_unflattened[7'h0c];
  assign sel_772715 = array_index_772631 == array_index_772708 ? add_772713 : sel_772709;
  assign add_772719 = sel_772715 + 8'h01;
  assign array_index_772720 = set2_unflattened[7'h0d];
  assign sel_772721 = array_index_772631 == array_index_772714 ? add_772719 : sel_772715;
  assign add_772725 = sel_772721 + 8'h01;
  assign array_index_772726 = set2_unflattened[7'h0e];
  assign sel_772727 = array_index_772631 == array_index_772720 ? add_772725 : sel_772721;
  assign add_772731 = sel_772727 + 8'h01;
  assign array_index_772732 = set2_unflattened[7'h0f];
  assign sel_772733 = array_index_772631 == array_index_772726 ? add_772731 : sel_772727;
  assign add_772737 = sel_772733 + 8'h01;
  assign array_index_772738 = set2_unflattened[7'h10];
  assign sel_772739 = array_index_772631 == array_index_772732 ? add_772737 : sel_772733;
  assign add_772743 = sel_772739 + 8'h01;
  assign array_index_772744 = set2_unflattened[7'h11];
  assign sel_772745 = array_index_772631 == array_index_772738 ? add_772743 : sel_772739;
  assign add_772749 = sel_772745 + 8'h01;
  assign array_index_772750 = set2_unflattened[7'h12];
  assign sel_772751 = array_index_772631 == array_index_772744 ? add_772749 : sel_772745;
  assign add_772755 = sel_772751 + 8'h01;
  assign array_index_772756 = set2_unflattened[7'h13];
  assign sel_772757 = array_index_772631 == array_index_772750 ? add_772755 : sel_772751;
  assign add_772761 = sel_772757 + 8'h01;
  assign array_index_772762 = set2_unflattened[7'h14];
  assign sel_772763 = array_index_772631 == array_index_772756 ? add_772761 : sel_772757;
  assign add_772767 = sel_772763 + 8'h01;
  assign array_index_772768 = set2_unflattened[7'h15];
  assign sel_772769 = array_index_772631 == array_index_772762 ? add_772767 : sel_772763;
  assign add_772773 = sel_772769 + 8'h01;
  assign array_index_772774 = set2_unflattened[7'h16];
  assign sel_772775 = array_index_772631 == array_index_772768 ? add_772773 : sel_772769;
  assign add_772779 = sel_772775 + 8'h01;
  assign array_index_772780 = set2_unflattened[7'h17];
  assign sel_772781 = array_index_772631 == array_index_772774 ? add_772779 : sel_772775;
  assign add_772785 = sel_772781 + 8'h01;
  assign array_index_772786 = set2_unflattened[7'h18];
  assign sel_772787 = array_index_772631 == array_index_772780 ? add_772785 : sel_772781;
  assign add_772791 = sel_772787 + 8'h01;
  assign array_index_772792 = set2_unflattened[7'h19];
  assign sel_772793 = array_index_772631 == array_index_772786 ? add_772791 : sel_772787;
  assign add_772797 = sel_772793 + 8'h01;
  assign array_index_772798 = set2_unflattened[7'h1a];
  assign sel_772799 = array_index_772631 == array_index_772792 ? add_772797 : sel_772793;
  assign add_772803 = sel_772799 + 8'h01;
  assign array_index_772804 = set2_unflattened[7'h1b];
  assign sel_772805 = array_index_772631 == array_index_772798 ? add_772803 : sel_772799;
  assign add_772809 = sel_772805 + 8'h01;
  assign array_index_772810 = set2_unflattened[7'h1c];
  assign sel_772811 = array_index_772631 == array_index_772804 ? add_772809 : sel_772805;
  assign add_772815 = sel_772811 + 8'h01;
  assign array_index_772816 = set2_unflattened[7'h1d];
  assign sel_772817 = array_index_772631 == array_index_772810 ? add_772815 : sel_772811;
  assign add_772821 = sel_772817 + 8'h01;
  assign array_index_772822 = set2_unflattened[7'h1e];
  assign sel_772823 = array_index_772631 == array_index_772816 ? add_772821 : sel_772817;
  assign add_772827 = sel_772823 + 8'h01;
  assign array_index_772828 = set2_unflattened[7'h1f];
  assign sel_772829 = array_index_772631 == array_index_772822 ? add_772827 : sel_772823;
  assign add_772833 = sel_772829 + 8'h01;
  assign array_index_772834 = set2_unflattened[7'h20];
  assign sel_772835 = array_index_772631 == array_index_772828 ? add_772833 : sel_772829;
  assign add_772839 = sel_772835 + 8'h01;
  assign array_index_772840 = set2_unflattened[7'h21];
  assign sel_772841 = array_index_772631 == array_index_772834 ? add_772839 : sel_772835;
  assign add_772845 = sel_772841 + 8'h01;
  assign array_index_772846 = set2_unflattened[7'h22];
  assign sel_772847 = array_index_772631 == array_index_772840 ? add_772845 : sel_772841;
  assign add_772851 = sel_772847 + 8'h01;
  assign array_index_772852 = set2_unflattened[7'h23];
  assign sel_772853 = array_index_772631 == array_index_772846 ? add_772851 : sel_772847;
  assign add_772857 = sel_772853 + 8'h01;
  assign array_index_772858 = set2_unflattened[7'h24];
  assign sel_772859 = array_index_772631 == array_index_772852 ? add_772857 : sel_772853;
  assign add_772863 = sel_772859 + 8'h01;
  assign array_index_772864 = set2_unflattened[7'h25];
  assign sel_772865 = array_index_772631 == array_index_772858 ? add_772863 : sel_772859;
  assign add_772869 = sel_772865 + 8'h01;
  assign array_index_772870 = set2_unflattened[7'h26];
  assign sel_772871 = array_index_772631 == array_index_772864 ? add_772869 : sel_772865;
  assign add_772875 = sel_772871 + 8'h01;
  assign array_index_772876 = set2_unflattened[7'h27];
  assign sel_772877 = array_index_772631 == array_index_772870 ? add_772875 : sel_772871;
  assign add_772881 = sel_772877 + 8'h01;
  assign array_index_772882 = set2_unflattened[7'h28];
  assign sel_772883 = array_index_772631 == array_index_772876 ? add_772881 : sel_772877;
  assign add_772887 = sel_772883 + 8'h01;
  assign array_index_772888 = set2_unflattened[7'h29];
  assign sel_772889 = array_index_772631 == array_index_772882 ? add_772887 : sel_772883;
  assign add_772893 = sel_772889 + 8'h01;
  assign array_index_772894 = set2_unflattened[7'h2a];
  assign sel_772895 = array_index_772631 == array_index_772888 ? add_772893 : sel_772889;
  assign add_772899 = sel_772895 + 8'h01;
  assign array_index_772900 = set2_unflattened[7'h2b];
  assign sel_772901 = array_index_772631 == array_index_772894 ? add_772899 : sel_772895;
  assign add_772905 = sel_772901 + 8'h01;
  assign array_index_772906 = set2_unflattened[7'h2c];
  assign sel_772907 = array_index_772631 == array_index_772900 ? add_772905 : sel_772901;
  assign add_772911 = sel_772907 + 8'h01;
  assign array_index_772912 = set2_unflattened[7'h2d];
  assign sel_772913 = array_index_772631 == array_index_772906 ? add_772911 : sel_772907;
  assign add_772917 = sel_772913 + 8'h01;
  assign array_index_772918 = set2_unflattened[7'h2e];
  assign sel_772919 = array_index_772631 == array_index_772912 ? add_772917 : sel_772913;
  assign add_772923 = sel_772919 + 8'h01;
  assign array_index_772924 = set2_unflattened[7'h2f];
  assign sel_772925 = array_index_772631 == array_index_772918 ? add_772923 : sel_772919;
  assign add_772929 = sel_772925 + 8'h01;
  assign array_index_772930 = set2_unflattened[7'h30];
  assign sel_772931 = array_index_772631 == array_index_772924 ? add_772929 : sel_772925;
  assign add_772935 = sel_772931 + 8'h01;
  assign array_index_772936 = set2_unflattened[7'h31];
  assign sel_772937 = array_index_772631 == array_index_772930 ? add_772935 : sel_772931;
  assign add_772941 = sel_772937 + 8'h01;
  assign array_index_772942 = set2_unflattened[7'h32];
  assign sel_772943 = array_index_772631 == array_index_772936 ? add_772941 : sel_772937;
  assign add_772947 = sel_772943 + 8'h01;
  assign array_index_772948 = set2_unflattened[7'h33];
  assign sel_772949 = array_index_772631 == array_index_772942 ? add_772947 : sel_772943;
  assign add_772953 = sel_772949 + 8'h01;
  assign array_index_772954 = set2_unflattened[7'h34];
  assign sel_772955 = array_index_772631 == array_index_772948 ? add_772953 : sel_772949;
  assign add_772959 = sel_772955 + 8'h01;
  assign array_index_772960 = set2_unflattened[7'h35];
  assign sel_772961 = array_index_772631 == array_index_772954 ? add_772959 : sel_772955;
  assign add_772965 = sel_772961 + 8'h01;
  assign array_index_772966 = set2_unflattened[7'h36];
  assign sel_772967 = array_index_772631 == array_index_772960 ? add_772965 : sel_772961;
  assign add_772971 = sel_772967 + 8'h01;
  assign array_index_772972 = set2_unflattened[7'h37];
  assign sel_772973 = array_index_772631 == array_index_772966 ? add_772971 : sel_772967;
  assign add_772977 = sel_772973 + 8'h01;
  assign array_index_772978 = set2_unflattened[7'h38];
  assign sel_772979 = array_index_772631 == array_index_772972 ? add_772977 : sel_772973;
  assign add_772983 = sel_772979 + 8'h01;
  assign array_index_772984 = set2_unflattened[7'h39];
  assign sel_772985 = array_index_772631 == array_index_772978 ? add_772983 : sel_772979;
  assign add_772989 = sel_772985 + 8'h01;
  assign array_index_772990 = set2_unflattened[7'h3a];
  assign sel_772991 = array_index_772631 == array_index_772984 ? add_772989 : sel_772985;
  assign add_772995 = sel_772991 + 8'h01;
  assign array_index_772996 = set2_unflattened[7'h3b];
  assign sel_772997 = array_index_772631 == array_index_772990 ? add_772995 : sel_772991;
  assign add_773001 = sel_772997 + 8'h01;
  assign array_index_773002 = set2_unflattened[7'h3c];
  assign sel_773003 = array_index_772631 == array_index_772996 ? add_773001 : sel_772997;
  assign add_773007 = sel_773003 + 8'h01;
  assign array_index_773008 = set2_unflattened[7'h3d];
  assign sel_773009 = array_index_772631 == array_index_773002 ? add_773007 : sel_773003;
  assign add_773013 = sel_773009 + 8'h01;
  assign array_index_773014 = set2_unflattened[7'h3e];
  assign sel_773015 = array_index_772631 == array_index_773008 ? add_773013 : sel_773009;
  assign add_773019 = sel_773015 + 8'h01;
  assign array_index_773020 = set2_unflattened[7'h3f];
  assign sel_773021 = array_index_772631 == array_index_773014 ? add_773019 : sel_773015;
  assign add_773025 = sel_773021 + 8'h01;
  assign array_index_773026 = set2_unflattened[7'h40];
  assign sel_773027 = array_index_772631 == array_index_773020 ? add_773025 : sel_773021;
  assign add_773031 = sel_773027 + 8'h01;
  assign array_index_773032 = set2_unflattened[7'h41];
  assign sel_773033 = array_index_772631 == array_index_773026 ? add_773031 : sel_773027;
  assign add_773037 = sel_773033 + 8'h01;
  assign array_index_773038 = set2_unflattened[7'h42];
  assign sel_773039 = array_index_772631 == array_index_773032 ? add_773037 : sel_773033;
  assign add_773043 = sel_773039 + 8'h01;
  assign array_index_773044 = set2_unflattened[7'h43];
  assign sel_773045 = array_index_772631 == array_index_773038 ? add_773043 : sel_773039;
  assign add_773049 = sel_773045 + 8'h01;
  assign array_index_773050 = set2_unflattened[7'h44];
  assign sel_773051 = array_index_772631 == array_index_773044 ? add_773049 : sel_773045;
  assign add_773055 = sel_773051 + 8'h01;
  assign array_index_773056 = set2_unflattened[7'h45];
  assign sel_773057 = array_index_772631 == array_index_773050 ? add_773055 : sel_773051;
  assign add_773061 = sel_773057 + 8'h01;
  assign array_index_773062 = set2_unflattened[7'h46];
  assign sel_773063 = array_index_772631 == array_index_773056 ? add_773061 : sel_773057;
  assign add_773067 = sel_773063 + 8'h01;
  assign array_index_773068 = set2_unflattened[7'h47];
  assign sel_773069 = array_index_772631 == array_index_773062 ? add_773067 : sel_773063;
  assign add_773073 = sel_773069 + 8'h01;
  assign array_index_773074 = set2_unflattened[7'h48];
  assign sel_773075 = array_index_772631 == array_index_773068 ? add_773073 : sel_773069;
  assign add_773079 = sel_773075 + 8'h01;
  assign array_index_773080 = set2_unflattened[7'h49];
  assign sel_773081 = array_index_772631 == array_index_773074 ? add_773079 : sel_773075;
  assign add_773085 = sel_773081 + 8'h01;
  assign array_index_773086 = set2_unflattened[7'h4a];
  assign sel_773087 = array_index_772631 == array_index_773080 ? add_773085 : sel_773081;
  assign add_773091 = sel_773087 + 8'h01;
  assign array_index_773092 = set2_unflattened[7'h4b];
  assign sel_773093 = array_index_772631 == array_index_773086 ? add_773091 : sel_773087;
  assign add_773097 = sel_773093 + 8'h01;
  assign array_index_773098 = set2_unflattened[7'h4c];
  assign sel_773099 = array_index_772631 == array_index_773092 ? add_773097 : sel_773093;
  assign add_773103 = sel_773099 + 8'h01;
  assign array_index_773104 = set2_unflattened[7'h4d];
  assign sel_773105 = array_index_772631 == array_index_773098 ? add_773103 : sel_773099;
  assign add_773109 = sel_773105 + 8'h01;
  assign array_index_773110 = set2_unflattened[7'h4e];
  assign sel_773111 = array_index_772631 == array_index_773104 ? add_773109 : sel_773105;
  assign add_773115 = sel_773111 + 8'h01;
  assign array_index_773116 = set2_unflattened[7'h4f];
  assign sel_773117 = array_index_772631 == array_index_773110 ? add_773115 : sel_773111;
  assign add_773121 = sel_773117 + 8'h01;
  assign array_index_773122 = set2_unflattened[7'h50];
  assign sel_773123 = array_index_772631 == array_index_773116 ? add_773121 : sel_773117;
  assign add_773127 = sel_773123 + 8'h01;
  assign array_index_773128 = set2_unflattened[7'h51];
  assign sel_773129 = array_index_772631 == array_index_773122 ? add_773127 : sel_773123;
  assign add_773133 = sel_773129 + 8'h01;
  assign array_index_773134 = set2_unflattened[7'h52];
  assign sel_773135 = array_index_772631 == array_index_773128 ? add_773133 : sel_773129;
  assign add_773139 = sel_773135 + 8'h01;
  assign array_index_773140 = set2_unflattened[7'h53];
  assign sel_773141 = array_index_772631 == array_index_773134 ? add_773139 : sel_773135;
  assign add_773145 = sel_773141 + 8'h01;
  assign array_index_773146 = set2_unflattened[7'h54];
  assign sel_773147 = array_index_772631 == array_index_773140 ? add_773145 : sel_773141;
  assign add_773151 = sel_773147 + 8'h01;
  assign array_index_773152 = set2_unflattened[7'h55];
  assign sel_773153 = array_index_772631 == array_index_773146 ? add_773151 : sel_773147;
  assign add_773157 = sel_773153 + 8'h01;
  assign array_index_773158 = set2_unflattened[7'h56];
  assign sel_773159 = array_index_772631 == array_index_773152 ? add_773157 : sel_773153;
  assign add_773163 = sel_773159 + 8'h01;
  assign array_index_773164 = set2_unflattened[7'h57];
  assign sel_773165 = array_index_772631 == array_index_773158 ? add_773163 : sel_773159;
  assign add_773169 = sel_773165 + 8'h01;
  assign array_index_773170 = set2_unflattened[7'h58];
  assign sel_773171 = array_index_772631 == array_index_773164 ? add_773169 : sel_773165;
  assign add_773175 = sel_773171 + 8'h01;
  assign array_index_773176 = set2_unflattened[7'h59];
  assign sel_773177 = array_index_772631 == array_index_773170 ? add_773175 : sel_773171;
  assign add_773181 = sel_773177 + 8'h01;
  assign array_index_773182 = set1_unflattened[7'h01];
  assign sel_773183 = array_index_772631 == array_index_773176 ? add_773181 : sel_773177;
  assign add_773186 = sel_773183 + 8'h01;
  assign sel_773187 = array_index_773182 == array_index_772632 ? add_773186 : sel_773183;
  assign add_773190 = sel_773187 + 8'h01;
  assign sel_773191 = array_index_773182 == array_index_772636 ? add_773190 : sel_773187;
  assign add_773194 = sel_773191 + 8'h01;
  assign sel_773195 = array_index_773182 == array_index_772644 ? add_773194 : sel_773191;
  assign add_773198 = sel_773195 + 8'h01;
  assign sel_773199 = array_index_773182 == array_index_772652 ? add_773198 : sel_773195;
  assign add_773202 = sel_773199 + 8'h01;
  assign sel_773203 = array_index_773182 == array_index_772660 ? add_773202 : sel_773199;
  assign add_773206 = sel_773203 + 8'h01;
  assign sel_773207 = array_index_773182 == array_index_772668 ? add_773206 : sel_773203;
  assign add_773210 = sel_773207 + 8'h01;
  assign sel_773211 = array_index_773182 == array_index_772676 ? add_773210 : sel_773207;
  assign add_773214 = sel_773211 + 8'h01;
  assign sel_773215 = array_index_773182 == array_index_772684 ? add_773214 : sel_773211;
  assign add_773218 = sel_773215 + 8'h01;
  assign sel_773219 = array_index_773182 == array_index_772690 ? add_773218 : sel_773215;
  assign add_773222 = sel_773219 + 8'h01;
  assign sel_773223 = array_index_773182 == array_index_772696 ? add_773222 : sel_773219;
  assign add_773226 = sel_773223 + 8'h01;
  assign sel_773227 = array_index_773182 == array_index_772702 ? add_773226 : sel_773223;
  assign add_773230 = sel_773227 + 8'h01;
  assign sel_773231 = array_index_773182 == array_index_772708 ? add_773230 : sel_773227;
  assign add_773234 = sel_773231 + 8'h01;
  assign sel_773235 = array_index_773182 == array_index_772714 ? add_773234 : sel_773231;
  assign add_773238 = sel_773235 + 8'h01;
  assign sel_773239 = array_index_773182 == array_index_772720 ? add_773238 : sel_773235;
  assign add_773242 = sel_773239 + 8'h01;
  assign sel_773243 = array_index_773182 == array_index_772726 ? add_773242 : sel_773239;
  assign add_773246 = sel_773243 + 8'h01;
  assign sel_773247 = array_index_773182 == array_index_772732 ? add_773246 : sel_773243;
  assign add_773250 = sel_773247 + 8'h01;
  assign sel_773251 = array_index_773182 == array_index_772738 ? add_773250 : sel_773247;
  assign add_773254 = sel_773251 + 8'h01;
  assign sel_773255 = array_index_773182 == array_index_772744 ? add_773254 : sel_773251;
  assign add_773258 = sel_773255 + 8'h01;
  assign sel_773259 = array_index_773182 == array_index_772750 ? add_773258 : sel_773255;
  assign add_773262 = sel_773259 + 8'h01;
  assign sel_773263 = array_index_773182 == array_index_772756 ? add_773262 : sel_773259;
  assign add_773266 = sel_773263 + 8'h01;
  assign sel_773267 = array_index_773182 == array_index_772762 ? add_773266 : sel_773263;
  assign add_773270 = sel_773267 + 8'h01;
  assign sel_773271 = array_index_773182 == array_index_772768 ? add_773270 : sel_773267;
  assign add_773274 = sel_773271 + 8'h01;
  assign sel_773275 = array_index_773182 == array_index_772774 ? add_773274 : sel_773271;
  assign add_773278 = sel_773275 + 8'h01;
  assign sel_773279 = array_index_773182 == array_index_772780 ? add_773278 : sel_773275;
  assign add_773282 = sel_773279 + 8'h01;
  assign sel_773283 = array_index_773182 == array_index_772786 ? add_773282 : sel_773279;
  assign add_773286 = sel_773283 + 8'h01;
  assign sel_773287 = array_index_773182 == array_index_772792 ? add_773286 : sel_773283;
  assign add_773290 = sel_773287 + 8'h01;
  assign sel_773291 = array_index_773182 == array_index_772798 ? add_773290 : sel_773287;
  assign add_773294 = sel_773291 + 8'h01;
  assign sel_773295 = array_index_773182 == array_index_772804 ? add_773294 : sel_773291;
  assign add_773298 = sel_773295 + 8'h01;
  assign sel_773299 = array_index_773182 == array_index_772810 ? add_773298 : sel_773295;
  assign add_773302 = sel_773299 + 8'h01;
  assign sel_773303 = array_index_773182 == array_index_772816 ? add_773302 : sel_773299;
  assign add_773306 = sel_773303 + 8'h01;
  assign sel_773307 = array_index_773182 == array_index_772822 ? add_773306 : sel_773303;
  assign add_773310 = sel_773307 + 8'h01;
  assign sel_773311 = array_index_773182 == array_index_772828 ? add_773310 : sel_773307;
  assign add_773314 = sel_773311 + 8'h01;
  assign sel_773315 = array_index_773182 == array_index_772834 ? add_773314 : sel_773311;
  assign add_773318 = sel_773315 + 8'h01;
  assign sel_773319 = array_index_773182 == array_index_772840 ? add_773318 : sel_773315;
  assign add_773322 = sel_773319 + 8'h01;
  assign sel_773323 = array_index_773182 == array_index_772846 ? add_773322 : sel_773319;
  assign add_773326 = sel_773323 + 8'h01;
  assign sel_773327 = array_index_773182 == array_index_772852 ? add_773326 : sel_773323;
  assign add_773330 = sel_773327 + 8'h01;
  assign sel_773331 = array_index_773182 == array_index_772858 ? add_773330 : sel_773327;
  assign add_773334 = sel_773331 + 8'h01;
  assign sel_773335 = array_index_773182 == array_index_772864 ? add_773334 : sel_773331;
  assign add_773338 = sel_773335 + 8'h01;
  assign sel_773339 = array_index_773182 == array_index_772870 ? add_773338 : sel_773335;
  assign add_773342 = sel_773339 + 8'h01;
  assign sel_773343 = array_index_773182 == array_index_772876 ? add_773342 : sel_773339;
  assign add_773346 = sel_773343 + 8'h01;
  assign sel_773347 = array_index_773182 == array_index_772882 ? add_773346 : sel_773343;
  assign add_773350 = sel_773347 + 8'h01;
  assign sel_773351 = array_index_773182 == array_index_772888 ? add_773350 : sel_773347;
  assign add_773354 = sel_773351 + 8'h01;
  assign sel_773355 = array_index_773182 == array_index_772894 ? add_773354 : sel_773351;
  assign add_773358 = sel_773355 + 8'h01;
  assign sel_773359 = array_index_773182 == array_index_772900 ? add_773358 : sel_773355;
  assign add_773362 = sel_773359 + 8'h01;
  assign sel_773363 = array_index_773182 == array_index_772906 ? add_773362 : sel_773359;
  assign add_773366 = sel_773363 + 8'h01;
  assign sel_773367 = array_index_773182 == array_index_772912 ? add_773366 : sel_773363;
  assign add_773370 = sel_773367 + 8'h01;
  assign sel_773371 = array_index_773182 == array_index_772918 ? add_773370 : sel_773367;
  assign add_773374 = sel_773371 + 8'h01;
  assign sel_773375 = array_index_773182 == array_index_772924 ? add_773374 : sel_773371;
  assign add_773378 = sel_773375 + 8'h01;
  assign sel_773379 = array_index_773182 == array_index_772930 ? add_773378 : sel_773375;
  assign add_773382 = sel_773379 + 8'h01;
  assign sel_773383 = array_index_773182 == array_index_772936 ? add_773382 : sel_773379;
  assign add_773386 = sel_773383 + 8'h01;
  assign sel_773387 = array_index_773182 == array_index_772942 ? add_773386 : sel_773383;
  assign add_773390 = sel_773387 + 8'h01;
  assign sel_773391 = array_index_773182 == array_index_772948 ? add_773390 : sel_773387;
  assign add_773394 = sel_773391 + 8'h01;
  assign sel_773395 = array_index_773182 == array_index_772954 ? add_773394 : sel_773391;
  assign add_773398 = sel_773395 + 8'h01;
  assign sel_773399 = array_index_773182 == array_index_772960 ? add_773398 : sel_773395;
  assign add_773402 = sel_773399 + 8'h01;
  assign sel_773403 = array_index_773182 == array_index_772966 ? add_773402 : sel_773399;
  assign add_773406 = sel_773403 + 8'h01;
  assign sel_773407 = array_index_773182 == array_index_772972 ? add_773406 : sel_773403;
  assign add_773410 = sel_773407 + 8'h01;
  assign sel_773411 = array_index_773182 == array_index_772978 ? add_773410 : sel_773407;
  assign add_773414 = sel_773411 + 8'h01;
  assign sel_773415 = array_index_773182 == array_index_772984 ? add_773414 : sel_773411;
  assign add_773418 = sel_773415 + 8'h01;
  assign sel_773419 = array_index_773182 == array_index_772990 ? add_773418 : sel_773415;
  assign add_773422 = sel_773419 + 8'h01;
  assign sel_773423 = array_index_773182 == array_index_772996 ? add_773422 : sel_773419;
  assign add_773426 = sel_773423 + 8'h01;
  assign sel_773427 = array_index_773182 == array_index_773002 ? add_773426 : sel_773423;
  assign add_773430 = sel_773427 + 8'h01;
  assign sel_773431 = array_index_773182 == array_index_773008 ? add_773430 : sel_773427;
  assign add_773434 = sel_773431 + 8'h01;
  assign sel_773435 = array_index_773182 == array_index_773014 ? add_773434 : sel_773431;
  assign add_773438 = sel_773435 + 8'h01;
  assign sel_773439 = array_index_773182 == array_index_773020 ? add_773438 : sel_773435;
  assign add_773442 = sel_773439 + 8'h01;
  assign sel_773443 = array_index_773182 == array_index_773026 ? add_773442 : sel_773439;
  assign add_773446 = sel_773443 + 8'h01;
  assign sel_773447 = array_index_773182 == array_index_773032 ? add_773446 : sel_773443;
  assign add_773450 = sel_773447 + 8'h01;
  assign sel_773451 = array_index_773182 == array_index_773038 ? add_773450 : sel_773447;
  assign add_773454 = sel_773451 + 8'h01;
  assign sel_773455 = array_index_773182 == array_index_773044 ? add_773454 : sel_773451;
  assign add_773458 = sel_773455 + 8'h01;
  assign sel_773459 = array_index_773182 == array_index_773050 ? add_773458 : sel_773455;
  assign add_773462 = sel_773459 + 8'h01;
  assign sel_773463 = array_index_773182 == array_index_773056 ? add_773462 : sel_773459;
  assign add_773466 = sel_773463 + 8'h01;
  assign sel_773467 = array_index_773182 == array_index_773062 ? add_773466 : sel_773463;
  assign add_773470 = sel_773467 + 8'h01;
  assign sel_773471 = array_index_773182 == array_index_773068 ? add_773470 : sel_773467;
  assign add_773474 = sel_773471 + 8'h01;
  assign sel_773475 = array_index_773182 == array_index_773074 ? add_773474 : sel_773471;
  assign add_773478 = sel_773475 + 8'h01;
  assign sel_773479 = array_index_773182 == array_index_773080 ? add_773478 : sel_773475;
  assign add_773482 = sel_773479 + 8'h01;
  assign sel_773483 = array_index_773182 == array_index_773086 ? add_773482 : sel_773479;
  assign add_773486 = sel_773483 + 8'h01;
  assign sel_773487 = array_index_773182 == array_index_773092 ? add_773486 : sel_773483;
  assign add_773490 = sel_773487 + 8'h01;
  assign sel_773491 = array_index_773182 == array_index_773098 ? add_773490 : sel_773487;
  assign add_773494 = sel_773491 + 8'h01;
  assign sel_773495 = array_index_773182 == array_index_773104 ? add_773494 : sel_773491;
  assign add_773498 = sel_773495 + 8'h01;
  assign sel_773499 = array_index_773182 == array_index_773110 ? add_773498 : sel_773495;
  assign add_773502 = sel_773499 + 8'h01;
  assign sel_773503 = array_index_773182 == array_index_773116 ? add_773502 : sel_773499;
  assign add_773506 = sel_773503 + 8'h01;
  assign sel_773507 = array_index_773182 == array_index_773122 ? add_773506 : sel_773503;
  assign add_773510 = sel_773507 + 8'h01;
  assign sel_773511 = array_index_773182 == array_index_773128 ? add_773510 : sel_773507;
  assign add_773514 = sel_773511 + 8'h01;
  assign sel_773515 = array_index_773182 == array_index_773134 ? add_773514 : sel_773511;
  assign add_773518 = sel_773515 + 8'h01;
  assign sel_773519 = array_index_773182 == array_index_773140 ? add_773518 : sel_773515;
  assign add_773522 = sel_773519 + 8'h01;
  assign sel_773523 = array_index_773182 == array_index_773146 ? add_773522 : sel_773519;
  assign add_773526 = sel_773523 + 8'h01;
  assign sel_773527 = array_index_773182 == array_index_773152 ? add_773526 : sel_773523;
  assign add_773530 = sel_773527 + 8'h01;
  assign sel_773531 = array_index_773182 == array_index_773158 ? add_773530 : sel_773527;
  assign add_773534 = sel_773531 + 8'h01;
  assign sel_773535 = array_index_773182 == array_index_773164 ? add_773534 : sel_773531;
  assign add_773538 = sel_773535 + 8'h01;
  assign sel_773539 = array_index_773182 == array_index_773170 ? add_773538 : sel_773535;
  assign add_773543 = sel_773539 + 8'h01;
  assign array_index_773544 = set1_unflattened[7'h02];
  assign sel_773545 = array_index_773182 == array_index_773176 ? add_773543 : sel_773539;
  assign add_773548 = sel_773545 + 8'h01;
  assign sel_773549 = array_index_773544 == array_index_772632 ? add_773548 : sel_773545;
  assign add_773552 = sel_773549 + 8'h01;
  assign sel_773553 = array_index_773544 == array_index_772636 ? add_773552 : sel_773549;
  assign add_773556 = sel_773553 + 8'h01;
  assign sel_773557 = array_index_773544 == array_index_772644 ? add_773556 : sel_773553;
  assign add_773560 = sel_773557 + 8'h01;
  assign sel_773561 = array_index_773544 == array_index_772652 ? add_773560 : sel_773557;
  assign add_773564 = sel_773561 + 8'h01;
  assign sel_773565 = array_index_773544 == array_index_772660 ? add_773564 : sel_773561;
  assign add_773568 = sel_773565 + 8'h01;
  assign sel_773569 = array_index_773544 == array_index_772668 ? add_773568 : sel_773565;
  assign add_773572 = sel_773569 + 8'h01;
  assign sel_773573 = array_index_773544 == array_index_772676 ? add_773572 : sel_773569;
  assign add_773576 = sel_773573 + 8'h01;
  assign sel_773577 = array_index_773544 == array_index_772684 ? add_773576 : sel_773573;
  assign add_773580 = sel_773577 + 8'h01;
  assign sel_773581 = array_index_773544 == array_index_772690 ? add_773580 : sel_773577;
  assign add_773584 = sel_773581 + 8'h01;
  assign sel_773585 = array_index_773544 == array_index_772696 ? add_773584 : sel_773581;
  assign add_773588 = sel_773585 + 8'h01;
  assign sel_773589 = array_index_773544 == array_index_772702 ? add_773588 : sel_773585;
  assign add_773592 = sel_773589 + 8'h01;
  assign sel_773593 = array_index_773544 == array_index_772708 ? add_773592 : sel_773589;
  assign add_773596 = sel_773593 + 8'h01;
  assign sel_773597 = array_index_773544 == array_index_772714 ? add_773596 : sel_773593;
  assign add_773600 = sel_773597 + 8'h01;
  assign sel_773601 = array_index_773544 == array_index_772720 ? add_773600 : sel_773597;
  assign add_773604 = sel_773601 + 8'h01;
  assign sel_773605 = array_index_773544 == array_index_772726 ? add_773604 : sel_773601;
  assign add_773608 = sel_773605 + 8'h01;
  assign sel_773609 = array_index_773544 == array_index_772732 ? add_773608 : sel_773605;
  assign add_773612 = sel_773609 + 8'h01;
  assign sel_773613 = array_index_773544 == array_index_772738 ? add_773612 : sel_773609;
  assign add_773616 = sel_773613 + 8'h01;
  assign sel_773617 = array_index_773544 == array_index_772744 ? add_773616 : sel_773613;
  assign add_773620 = sel_773617 + 8'h01;
  assign sel_773621 = array_index_773544 == array_index_772750 ? add_773620 : sel_773617;
  assign add_773624 = sel_773621 + 8'h01;
  assign sel_773625 = array_index_773544 == array_index_772756 ? add_773624 : sel_773621;
  assign add_773628 = sel_773625 + 8'h01;
  assign sel_773629 = array_index_773544 == array_index_772762 ? add_773628 : sel_773625;
  assign add_773632 = sel_773629 + 8'h01;
  assign sel_773633 = array_index_773544 == array_index_772768 ? add_773632 : sel_773629;
  assign add_773636 = sel_773633 + 8'h01;
  assign sel_773637 = array_index_773544 == array_index_772774 ? add_773636 : sel_773633;
  assign add_773640 = sel_773637 + 8'h01;
  assign sel_773641 = array_index_773544 == array_index_772780 ? add_773640 : sel_773637;
  assign add_773644 = sel_773641 + 8'h01;
  assign sel_773645 = array_index_773544 == array_index_772786 ? add_773644 : sel_773641;
  assign add_773648 = sel_773645 + 8'h01;
  assign sel_773649 = array_index_773544 == array_index_772792 ? add_773648 : sel_773645;
  assign add_773652 = sel_773649 + 8'h01;
  assign sel_773653 = array_index_773544 == array_index_772798 ? add_773652 : sel_773649;
  assign add_773656 = sel_773653 + 8'h01;
  assign sel_773657 = array_index_773544 == array_index_772804 ? add_773656 : sel_773653;
  assign add_773660 = sel_773657 + 8'h01;
  assign sel_773661 = array_index_773544 == array_index_772810 ? add_773660 : sel_773657;
  assign add_773664 = sel_773661 + 8'h01;
  assign sel_773665 = array_index_773544 == array_index_772816 ? add_773664 : sel_773661;
  assign add_773668 = sel_773665 + 8'h01;
  assign sel_773669 = array_index_773544 == array_index_772822 ? add_773668 : sel_773665;
  assign add_773672 = sel_773669 + 8'h01;
  assign sel_773673 = array_index_773544 == array_index_772828 ? add_773672 : sel_773669;
  assign add_773676 = sel_773673 + 8'h01;
  assign sel_773677 = array_index_773544 == array_index_772834 ? add_773676 : sel_773673;
  assign add_773680 = sel_773677 + 8'h01;
  assign sel_773681 = array_index_773544 == array_index_772840 ? add_773680 : sel_773677;
  assign add_773684 = sel_773681 + 8'h01;
  assign sel_773685 = array_index_773544 == array_index_772846 ? add_773684 : sel_773681;
  assign add_773688 = sel_773685 + 8'h01;
  assign sel_773689 = array_index_773544 == array_index_772852 ? add_773688 : sel_773685;
  assign add_773692 = sel_773689 + 8'h01;
  assign sel_773693 = array_index_773544 == array_index_772858 ? add_773692 : sel_773689;
  assign add_773696 = sel_773693 + 8'h01;
  assign sel_773697 = array_index_773544 == array_index_772864 ? add_773696 : sel_773693;
  assign add_773700 = sel_773697 + 8'h01;
  assign sel_773701 = array_index_773544 == array_index_772870 ? add_773700 : sel_773697;
  assign add_773704 = sel_773701 + 8'h01;
  assign sel_773705 = array_index_773544 == array_index_772876 ? add_773704 : sel_773701;
  assign add_773708 = sel_773705 + 8'h01;
  assign sel_773709 = array_index_773544 == array_index_772882 ? add_773708 : sel_773705;
  assign add_773712 = sel_773709 + 8'h01;
  assign sel_773713 = array_index_773544 == array_index_772888 ? add_773712 : sel_773709;
  assign add_773716 = sel_773713 + 8'h01;
  assign sel_773717 = array_index_773544 == array_index_772894 ? add_773716 : sel_773713;
  assign add_773720 = sel_773717 + 8'h01;
  assign sel_773721 = array_index_773544 == array_index_772900 ? add_773720 : sel_773717;
  assign add_773724 = sel_773721 + 8'h01;
  assign sel_773725 = array_index_773544 == array_index_772906 ? add_773724 : sel_773721;
  assign add_773728 = sel_773725 + 8'h01;
  assign sel_773729 = array_index_773544 == array_index_772912 ? add_773728 : sel_773725;
  assign add_773732 = sel_773729 + 8'h01;
  assign sel_773733 = array_index_773544 == array_index_772918 ? add_773732 : sel_773729;
  assign add_773736 = sel_773733 + 8'h01;
  assign sel_773737 = array_index_773544 == array_index_772924 ? add_773736 : sel_773733;
  assign add_773740 = sel_773737 + 8'h01;
  assign sel_773741 = array_index_773544 == array_index_772930 ? add_773740 : sel_773737;
  assign add_773744 = sel_773741 + 8'h01;
  assign sel_773745 = array_index_773544 == array_index_772936 ? add_773744 : sel_773741;
  assign add_773748 = sel_773745 + 8'h01;
  assign sel_773749 = array_index_773544 == array_index_772942 ? add_773748 : sel_773745;
  assign add_773752 = sel_773749 + 8'h01;
  assign sel_773753 = array_index_773544 == array_index_772948 ? add_773752 : sel_773749;
  assign add_773756 = sel_773753 + 8'h01;
  assign sel_773757 = array_index_773544 == array_index_772954 ? add_773756 : sel_773753;
  assign add_773760 = sel_773757 + 8'h01;
  assign sel_773761 = array_index_773544 == array_index_772960 ? add_773760 : sel_773757;
  assign add_773764 = sel_773761 + 8'h01;
  assign sel_773765 = array_index_773544 == array_index_772966 ? add_773764 : sel_773761;
  assign add_773768 = sel_773765 + 8'h01;
  assign sel_773769 = array_index_773544 == array_index_772972 ? add_773768 : sel_773765;
  assign add_773772 = sel_773769 + 8'h01;
  assign sel_773773 = array_index_773544 == array_index_772978 ? add_773772 : sel_773769;
  assign add_773776 = sel_773773 + 8'h01;
  assign sel_773777 = array_index_773544 == array_index_772984 ? add_773776 : sel_773773;
  assign add_773780 = sel_773777 + 8'h01;
  assign sel_773781 = array_index_773544 == array_index_772990 ? add_773780 : sel_773777;
  assign add_773784 = sel_773781 + 8'h01;
  assign sel_773785 = array_index_773544 == array_index_772996 ? add_773784 : sel_773781;
  assign add_773788 = sel_773785 + 8'h01;
  assign sel_773789 = array_index_773544 == array_index_773002 ? add_773788 : sel_773785;
  assign add_773792 = sel_773789 + 8'h01;
  assign sel_773793 = array_index_773544 == array_index_773008 ? add_773792 : sel_773789;
  assign add_773796 = sel_773793 + 8'h01;
  assign sel_773797 = array_index_773544 == array_index_773014 ? add_773796 : sel_773793;
  assign add_773800 = sel_773797 + 8'h01;
  assign sel_773801 = array_index_773544 == array_index_773020 ? add_773800 : sel_773797;
  assign add_773804 = sel_773801 + 8'h01;
  assign sel_773805 = array_index_773544 == array_index_773026 ? add_773804 : sel_773801;
  assign add_773808 = sel_773805 + 8'h01;
  assign sel_773809 = array_index_773544 == array_index_773032 ? add_773808 : sel_773805;
  assign add_773812 = sel_773809 + 8'h01;
  assign sel_773813 = array_index_773544 == array_index_773038 ? add_773812 : sel_773809;
  assign add_773816 = sel_773813 + 8'h01;
  assign sel_773817 = array_index_773544 == array_index_773044 ? add_773816 : sel_773813;
  assign add_773820 = sel_773817 + 8'h01;
  assign sel_773821 = array_index_773544 == array_index_773050 ? add_773820 : sel_773817;
  assign add_773824 = sel_773821 + 8'h01;
  assign sel_773825 = array_index_773544 == array_index_773056 ? add_773824 : sel_773821;
  assign add_773828 = sel_773825 + 8'h01;
  assign sel_773829 = array_index_773544 == array_index_773062 ? add_773828 : sel_773825;
  assign add_773832 = sel_773829 + 8'h01;
  assign sel_773833 = array_index_773544 == array_index_773068 ? add_773832 : sel_773829;
  assign add_773836 = sel_773833 + 8'h01;
  assign sel_773837 = array_index_773544 == array_index_773074 ? add_773836 : sel_773833;
  assign add_773840 = sel_773837 + 8'h01;
  assign sel_773841 = array_index_773544 == array_index_773080 ? add_773840 : sel_773837;
  assign add_773844 = sel_773841 + 8'h01;
  assign sel_773845 = array_index_773544 == array_index_773086 ? add_773844 : sel_773841;
  assign add_773848 = sel_773845 + 8'h01;
  assign sel_773849 = array_index_773544 == array_index_773092 ? add_773848 : sel_773845;
  assign add_773852 = sel_773849 + 8'h01;
  assign sel_773853 = array_index_773544 == array_index_773098 ? add_773852 : sel_773849;
  assign add_773856 = sel_773853 + 8'h01;
  assign sel_773857 = array_index_773544 == array_index_773104 ? add_773856 : sel_773853;
  assign add_773860 = sel_773857 + 8'h01;
  assign sel_773861 = array_index_773544 == array_index_773110 ? add_773860 : sel_773857;
  assign add_773864 = sel_773861 + 8'h01;
  assign sel_773865 = array_index_773544 == array_index_773116 ? add_773864 : sel_773861;
  assign add_773868 = sel_773865 + 8'h01;
  assign sel_773869 = array_index_773544 == array_index_773122 ? add_773868 : sel_773865;
  assign add_773872 = sel_773869 + 8'h01;
  assign sel_773873 = array_index_773544 == array_index_773128 ? add_773872 : sel_773869;
  assign add_773876 = sel_773873 + 8'h01;
  assign sel_773877 = array_index_773544 == array_index_773134 ? add_773876 : sel_773873;
  assign add_773880 = sel_773877 + 8'h01;
  assign sel_773881 = array_index_773544 == array_index_773140 ? add_773880 : sel_773877;
  assign add_773884 = sel_773881 + 8'h01;
  assign sel_773885 = array_index_773544 == array_index_773146 ? add_773884 : sel_773881;
  assign add_773888 = sel_773885 + 8'h01;
  assign sel_773889 = array_index_773544 == array_index_773152 ? add_773888 : sel_773885;
  assign add_773892 = sel_773889 + 8'h01;
  assign sel_773893 = array_index_773544 == array_index_773158 ? add_773892 : sel_773889;
  assign add_773896 = sel_773893 + 8'h01;
  assign sel_773897 = array_index_773544 == array_index_773164 ? add_773896 : sel_773893;
  assign add_773900 = sel_773897 + 8'h01;
  assign sel_773901 = array_index_773544 == array_index_773170 ? add_773900 : sel_773897;
  assign add_773905 = sel_773901 + 8'h01;
  assign array_index_773906 = set1_unflattened[7'h03];
  assign sel_773907 = array_index_773544 == array_index_773176 ? add_773905 : sel_773901;
  assign add_773910 = sel_773907 + 8'h01;
  assign sel_773911 = array_index_773906 == array_index_772632 ? add_773910 : sel_773907;
  assign add_773914 = sel_773911 + 8'h01;
  assign sel_773915 = array_index_773906 == array_index_772636 ? add_773914 : sel_773911;
  assign add_773918 = sel_773915 + 8'h01;
  assign sel_773919 = array_index_773906 == array_index_772644 ? add_773918 : sel_773915;
  assign add_773922 = sel_773919 + 8'h01;
  assign sel_773923 = array_index_773906 == array_index_772652 ? add_773922 : sel_773919;
  assign add_773926 = sel_773923 + 8'h01;
  assign sel_773927 = array_index_773906 == array_index_772660 ? add_773926 : sel_773923;
  assign add_773930 = sel_773927 + 8'h01;
  assign sel_773931 = array_index_773906 == array_index_772668 ? add_773930 : sel_773927;
  assign add_773934 = sel_773931 + 8'h01;
  assign sel_773935 = array_index_773906 == array_index_772676 ? add_773934 : sel_773931;
  assign add_773938 = sel_773935 + 8'h01;
  assign sel_773939 = array_index_773906 == array_index_772684 ? add_773938 : sel_773935;
  assign add_773942 = sel_773939 + 8'h01;
  assign sel_773943 = array_index_773906 == array_index_772690 ? add_773942 : sel_773939;
  assign add_773946 = sel_773943 + 8'h01;
  assign sel_773947 = array_index_773906 == array_index_772696 ? add_773946 : sel_773943;
  assign add_773950 = sel_773947 + 8'h01;
  assign sel_773951 = array_index_773906 == array_index_772702 ? add_773950 : sel_773947;
  assign add_773954 = sel_773951 + 8'h01;
  assign sel_773955 = array_index_773906 == array_index_772708 ? add_773954 : sel_773951;
  assign add_773958 = sel_773955 + 8'h01;
  assign sel_773959 = array_index_773906 == array_index_772714 ? add_773958 : sel_773955;
  assign add_773962 = sel_773959 + 8'h01;
  assign sel_773963 = array_index_773906 == array_index_772720 ? add_773962 : sel_773959;
  assign add_773966 = sel_773963 + 8'h01;
  assign sel_773967 = array_index_773906 == array_index_772726 ? add_773966 : sel_773963;
  assign add_773970 = sel_773967 + 8'h01;
  assign sel_773971 = array_index_773906 == array_index_772732 ? add_773970 : sel_773967;
  assign add_773974 = sel_773971 + 8'h01;
  assign sel_773975 = array_index_773906 == array_index_772738 ? add_773974 : sel_773971;
  assign add_773978 = sel_773975 + 8'h01;
  assign sel_773979 = array_index_773906 == array_index_772744 ? add_773978 : sel_773975;
  assign add_773982 = sel_773979 + 8'h01;
  assign sel_773983 = array_index_773906 == array_index_772750 ? add_773982 : sel_773979;
  assign add_773986 = sel_773983 + 8'h01;
  assign sel_773987 = array_index_773906 == array_index_772756 ? add_773986 : sel_773983;
  assign add_773990 = sel_773987 + 8'h01;
  assign sel_773991 = array_index_773906 == array_index_772762 ? add_773990 : sel_773987;
  assign add_773994 = sel_773991 + 8'h01;
  assign sel_773995 = array_index_773906 == array_index_772768 ? add_773994 : sel_773991;
  assign add_773998 = sel_773995 + 8'h01;
  assign sel_773999 = array_index_773906 == array_index_772774 ? add_773998 : sel_773995;
  assign add_774002 = sel_773999 + 8'h01;
  assign sel_774003 = array_index_773906 == array_index_772780 ? add_774002 : sel_773999;
  assign add_774006 = sel_774003 + 8'h01;
  assign sel_774007 = array_index_773906 == array_index_772786 ? add_774006 : sel_774003;
  assign add_774010 = sel_774007 + 8'h01;
  assign sel_774011 = array_index_773906 == array_index_772792 ? add_774010 : sel_774007;
  assign add_774014 = sel_774011 + 8'h01;
  assign sel_774015 = array_index_773906 == array_index_772798 ? add_774014 : sel_774011;
  assign add_774018 = sel_774015 + 8'h01;
  assign sel_774019 = array_index_773906 == array_index_772804 ? add_774018 : sel_774015;
  assign add_774022 = sel_774019 + 8'h01;
  assign sel_774023 = array_index_773906 == array_index_772810 ? add_774022 : sel_774019;
  assign add_774026 = sel_774023 + 8'h01;
  assign sel_774027 = array_index_773906 == array_index_772816 ? add_774026 : sel_774023;
  assign add_774030 = sel_774027 + 8'h01;
  assign sel_774031 = array_index_773906 == array_index_772822 ? add_774030 : sel_774027;
  assign add_774034 = sel_774031 + 8'h01;
  assign sel_774035 = array_index_773906 == array_index_772828 ? add_774034 : sel_774031;
  assign add_774038 = sel_774035 + 8'h01;
  assign sel_774039 = array_index_773906 == array_index_772834 ? add_774038 : sel_774035;
  assign add_774042 = sel_774039 + 8'h01;
  assign sel_774043 = array_index_773906 == array_index_772840 ? add_774042 : sel_774039;
  assign add_774046 = sel_774043 + 8'h01;
  assign sel_774047 = array_index_773906 == array_index_772846 ? add_774046 : sel_774043;
  assign add_774050 = sel_774047 + 8'h01;
  assign sel_774051 = array_index_773906 == array_index_772852 ? add_774050 : sel_774047;
  assign add_774054 = sel_774051 + 8'h01;
  assign sel_774055 = array_index_773906 == array_index_772858 ? add_774054 : sel_774051;
  assign add_774058 = sel_774055 + 8'h01;
  assign sel_774059 = array_index_773906 == array_index_772864 ? add_774058 : sel_774055;
  assign add_774062 = sel_774059 + 8'h01;
  assign sel_774063 = array_index_773906 == array_index_772870 ? add_774062 : sel_774059;
  assign add_774066 = sel_774063 + 8'h01;
  assign sel_774067 = array_index_773906 == array_index_772876 ? add_774066 : sel_774063;
  assign add_774070 = sel_774067 + 8'h01;
  assign sel_774071 = array_index_773906 == array_index_772882 ? add_774070 : sel_774067;
  assign add_774074 = sel_774071 + 8'h01;
  assign sel_774075 = array_index_773906 == array_index_772888 ? add_774074 : sel_774071;
  assign add_774078 = sel_774075 + 8'h01;
  assign sel_774079 = array_index_773906 == array_index_772894 ? add_774078 : sel_774075;
  assign add_774082 = sel_774079 + 8'h01;
  assign sel_774083 = array_index_773906 == array_index_772900 ? add_774082 : sel_774079;
  assign add_774086 = sel_774083 + 8'h01;
  assign sel_774087 = array_index_773906 == array_index_772906 ? add_774086 : sel_774083;
  assign add_774090 = sel_774087 + 8'h01;
  assign sel_774091 = array_index_773906 == array_index_772912 ? add_774090 : sel_774087;
  assign add_774094 = sel_774091 + 8'h01;
  assign sel_774095 = array_index_773906 == array_index_772918 ? add_774094 : sel_774091;
  assign add_774098 = sel_774095 + 8'h01;
  assign sel_774099 = array_index_773906 == array_index_772924 ? add_774098 : sel_774095;
  assign add_774102 = sel_774099 + 8'h01;
  assign sel_774103 = array_index_773906 == array_index_772930 ? add_774102 : sel_774099;
  assign add_774106 = sel_774103 + 8'h01;
  assign sel_774107 = array_index_773906 == array_index_772936 ? add_774106 : sel_774103;
  assign add_774110 = sel_774107 + 8'h01;
  assign sel_774111 = array_index_773906 == array_index_772942 ? add_774110 : sel_774107;
  assign add_774114 = sel_774111 + 8'h01;
  assign sel_774115 = array_index_773906 == array_index_772948 ? add_774114 : sel_774111;
  assign add_774118 = sel_774115 + 8'h01;
  assign sel_774119 = array_index_773906 == array_index_772954 ? add_774118 : sel_774115;
  assign add_774122 = sel_774119 + 8'h01;
  assign sel_774123 = array_index_773906 == array_index_772960 ? add_774122 : sel_774119;
  assign add_774126 = sel_774123 + 8'h01;
  assign sel_774127 = array_index_773906 == array_index_772966 ? add_774126 : sel_774123;
  assign add_774130 = sel_774127 + 8'h01;
  assign sel_774131 = array_index_773906 == array_index_772972 ? add_774130 : sel_774127;
  assign add_774134 = sel_774131 + 8'h01;
  assign sel_774135 = array_index_773906 == array_index_772978 ? add_774134 : sel_774131;
  assign add_774138 = sel_774135 + 8'h01;
  assign sel_774139 = array_index_773906 == array_index_772984 ? add_774138 : sel_774135;
  assign add_774142 = sel_774139 + 8'h01;
  assign sel_774143 = array_index_773906 == array_index_772990 ? add_774142 : sel_774139;
  assign add_774146 = sel_774143 + 8'h01;
  assign sel_774147 = array_index_773906 == array_index_772996 ? add_774146 : sel_774143;
  assign add_774150 = sel_774147 + 8'h01;
  assign sel_774151 = array_index_773906 == array_index_773002 ? add_774150 : sel_774147;
  assign add_774154 = sel_774151 + 8'h01;
  assign sel_774155 = array_index_773906 == array_index_773008 ? add_774154 : sel_774151;
  assign add_774158 = sel_774155 + 8'h01;
  assign sel_774159 = array_index_773906 == array_index_773014 ? add_774158 : sel_774155;
  assign add_774162 = sel_774159 + 8'h01;
  assign sel_774163 = array_index_773906 == array_index_773020 ? add_774162 : sel_774159;
  assign add_774166 = sel_774163 + 8'h01;
  assign sel_774167 = array_index_773906 == array_index_773026 ? add_774166 : sel_774163;
  assign add_774170 = sel_774167 + 8'h01;
  assign sel_774171 = array_index_773906 == array_index_773032 ? add_774170 : sel_774167;
  assign add_774174 = sel_774171 + 8'h01;
  assign sel_774175 = array_index_773906 == array_index_773038 ? add_774174 : sel_774171;
  assign add_774178 = sel_774175 + 8'h01;
  assign sel_774179 = array_index_773906 == array_index_773044 ? add_774178 : sel_774175;
  assign add_774182 = sel_774179 + 8'h01;
  assign sel_774183 = array_index_773906 == array_index_773050 ? add_774182 : sel_774179;
  assign add_774186 = sel_774183 + 8'h01;
  assign sel_774187 = array_index_773906 == array_index_773056 ? add_774186 : sel_774183;
  assign add_774190 = sel_774187 + 8'h01;
  assign sel_774191 = array_index_773906 == array_index_773062 ? add_774190 : sel_774187;
  assign add_774194 = sel_774191 + 8'h01;
  assign sel_774195 = array_index_773906 == array_index_773068 ? add_774194 : sel_774191;
  assign add_774198 = sel_774195 + 8'h01;
  assign sel_774199 = array_index_773906 == array_index_773074 ? add_774198 : sel_774195;
  assign add_774202 = sel_774199 + 8'h01;
  assign sel_774203 = array_index_773906 == array_index_773080 ? add_774202 : sel_774199;
  assign add_774206 = sel_774203 + 8'h01;
  assign sel_774207 = array_index_773906 == array_index_773086 ? add_774206 : sel_774203;
  assign add_774210 = sel_774207 + 8'h01;
  assign sel_774211 = array_index_773906 == array_index_773092 ? add_774210 : sel_774207;
  assign add_774214 = sel_774211 + 8'h01;
  assign sel_774215 = array_index_773906 == array_index_773098 ? add_774214 : sel_774211;
  assign add_774218 = sel_774215 + 8'h01;
  assign sel_774219 = array_index_773906 == array_index_773104 ? add_774218 : sel_774215;
  assign add_774222 = sel_774219 + 8'h01;
  assign sel_774223 = array_index_773906 == array_index_773110 ? add_774222 : sel_774219;
  assign add_774226 = sel_774223 + 8'h01;
  assign sel_774227 = array_index_773906 == array_index_773116 ? add_774226 : sel_774223;
  assign add_774230 = sel_774227 + 8'h01;
  assign sel_774231 = array_index_773906 == array_index_773122 ? add_774230 : sel_774227;
  assign add_774234 = sel_774231 + 8'h01;
  assign sel_774235 = array_index_773906 == array_index_773128 ? add_774234 : sel_774231;
  assign add_774238 = sel_774235 + 8'h01;
  assign sel_774239 = array_index_773906 == array_index_773134 ? add_774238 : sel_774235;
  assign add_774242 = sel_774239 + 8'h01;
  assign sel_774243 = array_index_773906 == array_index_773140 ? add_774242 : sel_774239;
  assign add_774246 = sel_774243 + 8'h01;
  assign sel_774247 = array_index_773906 == array_index_773146 ? add_774246 : sel_774243;
  assign add_774250 = sel_774247 + 8'h01;
  assign sel_774251 = array_index_773906 == array_index_773152 ? add_774250 : sel_774247;
  assign add_774254 = sel_774251 + 8'h01;
  assign sel_774255 = array_index_773906 == array_index_773158 ? add_774254 : sel_774251;
  assign add_774258 = sel_774255 + 8'h01;
  assign sel_774259 = array_index_773906 == array_index_773164 ? add_774258 : sel_774255;
  assign add_774262 = sel_774259 + 8'h01;
  assign sel_774263 = array_index_773906 == array_index_773170 ? add_774262 : sel_774259;
  assign add_774267 = sel_774263 + 8'h01;
  assign array_index_774268 = set1_unflattened[7'h04];
  assign sel_774269 = array_index_773906 == array_index_773176 ? add_774267 : sel_774263;
  assign add_774272 = sel_774269 + 8'h01;
  assign sel_774273 = array_index_774268 == array_index_772632 ? add_774272 : sel_774269;
  assign add_774276 = sel_774273 + 8'h01;
  assign sel_774277 = array_index_774268 == array_index_772636 ? add_774276 : sel_774273;
  assign add_774280 = sel_774277 + 8'h01;
  assign sel_774281 = array_index_774268 == array_index_772644 ? add_774280 : sel_774277;
  assign add_774284 = sel_774281 + 8'h01;
  assign sel_774285 = array_index_774268 == array_index_772652 ? add_774284 : sel_774281;
  assign add_774288 = sel_774285 + 8'h01;
  assign sel_774289 = array_index_774268 == array_index_772660 ? add_774288 : sel_774285;
  assign add_774292 = sel_774289 + 8'h01;
  assign sel_774293 = array_index_774268 == array_index_772668 ? add_774292 : sel_774289;
  assign add_774296 = sel_774293 + 8'h01;
  assign sel_774297 = array_index_774268 == array_index_772676 ? add_774296 : sel_774293;
  assign add_774300 = sel_774297 + 8'h01;
  assign sel_774301 = array_index_774268 == array_index_772684 ? add_774300 : sel_774297;
  assign add_774304 = sel_774301 + 8'h01;
  assign sel_774305 = array_index_774268 == array_index_772690 ? add_774304 : sel_774301;
  assign add_774308 = sel_774305 + 8'h01;
  assign sel_774309 = array_index_774268 == array_index_772696 ? add_774308 : sel_774305;
  assign add_774312 = sel_774309 + 8'h01;
  assign sel_774313 = array_index_774268 == array_index_772702 ? add_774312 : sel_774309;
  assign add_774316 = sel_774313 + 8'h01;
  assign sel_774317 = array_index_774268 == array_index_772708 ? add_774316 : sel_774313;
  assign add_774320 = sel_774317 + 8'h01;
  assign sel_774321 = array_index_774268 == array_index_772714 ? add_774320 : sel_774317;
  assign add_774324 = sel_774321 + 8'h01;
  assign sel_774325 = array_index_774268 == array_index_772720 ? add_774324 : sel_774321;
  assign add_774328 = sel_774325 + 8'h01;
  assign sel_774329 = array_index_774268 == array_index_772726 ? add_774328 : sel_774325;
  assign add_774332 = sel_774329 + 8'h01;
  assign sel_774333 = array_index_774268 == array_index_772732 ? add_774332 : sel_774329;
  assign add_774336 = sel_774333 + 8'h01;
  assign sel_774337 = array_index_774268 == array_index_772738 ? add_774336 : sel_774333;
  assign add_774340 = sel_774337 + 8'h01;
  assign sel_774341 = array_index_774268 == array_index_772744 ? add_774340 : sel_774337;
  assign add_774344 = sel_774341 + 8'h01;
  assign sel_774345 = array_index_774268 == array_index_772750 ? add_774344 : sel_774341;
  assign add_774348 = sel_774345 + 8'h01;
  assign sel_774349 = array_index_774268 == array_index_772756 ? add_774348 : sel_774345;
  assign add_774352 = sel_774349 + 8'h01;
  assign sel_774353 = array_index_774268 == array_index_772762 ? add_774352 : sel_774349;
  assign add_774356 = sel_774353 + 8'h01;
  assign sel_774357 = array_index_774268 == array_index_772768 ? add_774356 : sel_774353;
  assign add_774360 = sel_774357 + 8'h01;
  assign sel_774361 = array_index_774268 == array_index_772774 ? add_774360 : sel_774357;
  assign add_774364 = sel_774361 + 8'h01;
  assign sel_774365 = array_index_774268 == array_index_772780 ? add_774364 : sel_774361;
  assign add_774368 = sel_774365 + 8'h01;
  assign sel_774369 = array_index_774268 == array_index_772786 ? add_774368 : sel_774365;
  assign add_774372 = sel_774369 + 8'h01;
  assign sel_774373 = array_index_774268 == array_index_772792 ? add_774372 : sel_774369;
  assign add_774376 = sel_774373 + 8'h01;
  assign sel_774377 = array_index_774268 == array_index_772798 ? add_774376 : sel_774373;
  assign add_774380 = sel_774377 + 8'h01;
  assign sel_774381 = array_index_774268 == array_index_772804 ? add_774380 : sel_774377;
  assign add_774384 = sel_774381 + 8'h01;
  assign sel_774385 = array_index_774268 == array_index_772810 ? add_774384 : sel_774381;
  assign add_774388 = sel_774385 + 8'h01;
  assign sel_774389 = array_index_774268 == array_index_772816 ? add_774388 : sel_774385;
  assign add_774392 = sel_774389 + 8'h01;
  assign sel_774393 = array_index_774268 == array_index_772822 ? add_774392 : sel_774389;
  assign add_774396 = sel_774393 + 8'h01;
  assign sel_774397 = array_index_774268 == array_index_772828 ? add_774396 : sel_774393;
  assign add_774400 = sel_774397 + 8'h01;
  assign sel_774401 = array_index_774268 == array_index_772834 ? add_774400 : sel_774397;
  assign add_774404 = sel_774401 + 8'h01;
  assign sel_774405 = array_index_774268 == array_index_772840 ? add_774404 : sel_774401;
  assign add_774408 = sel_774405 + 8'h01;
  assign sel_774409 = array_index_774268 == array_index_772846 ? add_774408 : sel_774405;
  assign add_774412 = sel_774409 + 8'h01;
  assign sel_774413 = array_index_774268 == array_index_772852 ? add_774412 : sel_774409;
  assign add_774416 = sel_774413 + 8'h01;
  assign sel_774417 = array_index_774268 == array_index_772858 ? add_774416 : sel_774413;
  assign add_774420 = sel_774417 + 8'h01;
  assign sel_774421 = array_index_774268 == array_index_772864 ? add_774420 : sel_774417;
  assign add_774424 = sel_774421 + 8'h01;
  assign sel_774425 = array_index_774268 == array_index_772870 ? add_774424 : sel_774421;
  assign add_774428 = sel_774425 + 8'h01;
  assign sel_774429 = array_index_774268 == array_index_772876 ? add_774428 : sel_774425;
  assign add_774432 = sel_774429 + 8'h01;
  assign sel_774433 = array_index_774268 == array_index_772882 ? add_774432 : sel_774429;
  assign add_774436 = sel_774433 + 8'h01;
  assign sel_774437 = array_index_774268 == array_index_772888 ? add_774436 : sel_774433;
  assign add_774440 = sel_774437 + 8'h01;
  assign sel_774441 = array_index_774268 == array_index_772894 ? add_774440 : sel_774437;
  assign add_774444 = sel_774441 + 8'h01;
  assign sel_774445 = array_index_774268 == array_index_772900 ? add_774444 : sel_774441;
  assign add_774448 = sel_774445 + 8'h01;
  assign sel_774449 = array_index_774268 == array_index_772906 ? add_774448 : sel_774445;
  assign add_774452 = sel_774449 + 8'h01;
  assign sel_774453 = array_index_774268 == array_index_772912 ? add_774452 : sel_774449;
  assign add_774456 = sel_774453 + 8'h01;
  assign sel_774457 = array_index_774268 == array_index_772918 ? add_774456 : sel_774453;
  assign add_774460 = sel_774457 + 8'h01;
  assign sel_774461 = array_index_774268 == array_index_772924 ? add_774460 : sel_774457;
  assign add_774464 = sel_774461 + 8'h01;
  assign sel_774465 = array_index_774268 == array_index_772930 ? add_774464 : sel_774461;
  assign add_774468 = sel_774465 + 8'h01;
  assign sel_774469 = array_index_774268 == array_index_772936 ? add_774468 : sel_774465;
  assign add_774472 = sel_774469 + 8'h01;
  assign sel_774473 = array_index_774268 == array_index_772942 ? add_774472 : sel_774469;
  assign add_774476 = sel_774473 + 8'h01;
  assign sel_774477 = array_index_774268 == array_index_772948 ? add_774476 : sel_774473;
  assign add_774480 = sel_774477 + 8'h01;
  assign sel_774481 = array_index_774268 == array_index_772954 ? add_774480 : sel_774477;
  assign add_774484 = sel_774481 + 8'h01;
  assign sel_774485 = array_index_774268 == array_index_772960 ? add_774484 : sel_774481;
  assign add_774488 = sel_774485 + 8'h01;
  assign sel_774489 = array_index_774268 == array_index_772966 ? add_774488 : sel_774485;
  assign add_774492 = sel_774489 + 8'h01;
  assign sel_774493 = array_index_774268 == array_index_772972 ? add_774492 : sel_774489;
  assign add_774496 = sel_774493 + 8'h01;
  assign sel_774497 = array_index_774268 == array_index_772978 ? add_774496 : sel_774493;
  assign add_774500 = sel_774497 + 8'h01;
  assign sel_774501 = array_index_774268 == array_index_772984 ? add_774500 : sel_774497;
  assign add_774504 = sel_774501 + 8'h01;
  assign sel_774505 = array_index_774268 == array_index_772990 ? add_774504 : sel_774501;
  assign add_774508 = sel_774505 + 8'h01;
  assign sel_774509 = array_index_774268 == array_index_772996 ? add_774508 : sel_774505;
  assign add_774512 = sel_774509 + 8'h01;
  assign sel_774513 = array_index_774268 == array_index_773002 ? add_774512 : sel_774509;
  assign add_774516 = sel_774513 + 8'h01;
  assign sel_774517 = array_index_774268 == array_index_773008 ? add_774516 : sel_774513;
  assign add_774520 = sel_774517 + 8'h01;
  assign sel_774521 = array_index_774268 == array_index_773014 ? add_774520 : sel_774517;
  assign add_774524 = sel_774521 + 8'h01;
  assign sel_774525 = array_index_774268 == array_index_773020 ? add_774524 : sel_774521;
  assign add_774528 = sel_774525 + 8'h01;
  assign sel_774529 = array_index_774268 == array_index_773026 ? add_774528 : sel_774525;
  assign add_774532 = sel_774529 + 8'h01;
  assign sel_774533 = array_index_774268 == array_index_773032 ? add_774532 : sel_774529;
  assign add_774536 = sel_774533 + 8'h01;
  assign sel_774537 = array_index_774268 == array_index_773038 ? add_774536 : sel_774533;
  assign add_774540 = sel_774537 + 8'h01;
  assign sel_774541 = array_index_774268 == array_index_773044 ? add_774540 : sel_774537;
  assign add_774544 = sel_774541 + 8'h01;
  assign sel_774545 = array_index_774268 == array_index_773050 ? add_774544 : sel_774541;
  assign add_774548 = sel_774545 + 8'h01;
  assign sel_774549 = array_index_774268 == array_index_773056 ? add_774548 : sel_774545;
  assign add_774552 = sel_774549 + 8'h01;
  assign sel_774553 = array_index_774268 == array_index_773062 ? add_774552 : sel_774549;
  assign add_774556 = sel_774553 + 8'h01;
  assign sel_774557 = array_index_774268 == array_index_773068 ? add_774556 : sel_774553;
  assign add_774560 = sel_774557 + 8'h01;
  assign sel_774561 = array_index_774268 == array_index_773074 ? add_774560 : sel_774557;
  assign add_774564 = sel_774561 + 8'h01;
  assign sel_774565 = array_index_774268 == array_index_773080 ? add_774564 : sel_774561;
  assign add_774568 = sel_774565 + 8'h01;
  assign sel_774569 = array_index_774268 == array_index_773086 ? add_774568 : sel_774565;
  assign add_774572 = sel_774569 + 8'h01;
  assign sel_774573 = array_index_774268 == array_index_773092 ? add_774572 : sel_774569;
  assign add_774576 = sel_774573 + 8'h01;
  assign sel_774577 = array_index_774268 == array_index_773098 ? add_774576 : sel_774573;
  assign add_774580 = sel_774577 + 8'h01;
  assign sel_774581 = array_index_774268 == array_index_773104 ? add_774580 : sel_774577;
  assign add_774584 = sel_774581 + 8'h01;
  assign sel_774585 = array_index_774268 == array_index_773110 ? add_774584 : sel_774581;
  assign add_774588 = sel_774585 + 8'h01;
  assign sel_774589 = array_index_774268 == array_index_773116 ? add_774588 : sel_774585;
  assign add_774592 = sel_774589 + 8'h01;
  assign sel_774593 = array_index_774268 == array_index_773122 ? add_774592 : sel_774589;
  assign add_774596 = sel_774593 + 8'h01;
  assign sel_774597 = array_index_774268 == array_index_773128 ? add_774596 : sel_774593;
  assign add_774600 = sel_774597 + 8'h01;
  assign sel_774601 = array_index_774268 == array_index_773134 ? add_774600 : sel_774597;
  assign add_774604 = sel_774601 + 8'h01;
  assign sel_774605 = array_index_774268 == array_index_773140 ? add_774604 : sel_774601;
  assign add_774608 = sel_774605 + 8'h01;
  assign sel_774609 = array_index_774268 == array_index_773146 ? add_774608 : sel_774605;
  assign add_774612 = sel_774609 + 8'h01;
  assign sel_774613 = array_index_774268 == array_index_773152 ? add_774612 : sel_774609;
  assign add_774616 = sel_774613 + 8'h01;
  assign sel_774617 = array_index_774268 == array_index_773158 ? add_774616 : sel_774613;
  assign add_774620 = sel_774617 + 8'h01;
  assign sel_774621 = array_index_774268 == array_index_773164 ? add_774620 : sel_774617;
  assign add_774624 = sel_774621 + 8'h01;
  assign sel_774625 = array_index_774268 == array_index_773170 ? add_774624 : sel_774621;
  assign add_774629 = sel_774625 + 8'h01;
  assign array_index_774630 = set1_unflattened[7'h05];
  assign sel_774631 = array_index_774268 == array_index_773176 ? add_774629 : sel_774625;
  assign add_774634 = sel_774631 + 8'h01;
  assign sel_774635 = array_index_774630 == array_index_772632 ? add_774634 : sel_774631;
  assign add_774638 = sel_774635 + 8'h01;
  assign sel_774639 = array_index_774630 == array_index_772636 ? add_774638 : sel_774635;
  assign add_774642 = sel_774639 + 8'h01;
  assign sel_774643 = array_index_774630 == array_index_772644 ? add_774642 : sel_774639;
  assign add_774646 = sel_774643 + 8'h01;
  assign sel_774647 = array_index_774630 == array_index_772652 ? add_774646 : sel_774643;
  assign add_774650 = sel_774647 + 8'h01;
  assign sel_774651 = array_index_774630 == array_index_772660 ? add_774650 : sel_774647;
  assign add_774654 = sel_774651 + 8'h01;
  assign sel_774655 = array_index_774630 == array_index_772668 ? add_774654 : sel_774651;
  assign add_774658 = sel_774655 + 8'h01;
  assign sel_774659 = array_index_774630 == array_index_772676 ? add_774658 : sel_774655;
  assign add_774662 = sel_774659 + 8'h01;
  assign sel_774663 = array_index_774630 == array_index_772684 ? add_774662 : sel_774659;
  assign add_774666 = sel_774663 + 8'h01;
  assign sel_774667 = array_index_774630 == array_index_772690 ? add_774666 : sel_774663;
  assign add_774670 = sel_774667 + 8'h01;
  assign sel_774671 = array_index_774630 == array_index_772696 ? add_774670 : sel_774667;
  assign add_774674 = sel_774671 + 8'h01;
  assign sel_774675 = array_index_774630 == array_index_772702 ? add_774674 : sel_774671;
  assign add_774678 = sel_774675 + 8'h01;
  assign sel_774679 = array_index_774630 == array_index_772708 ? add_774678 : sel_774675;
  assign add_774682 = sel_774679 + 8'h01;
  assign sel_774683 = array_index_774630 == array_index_772714 ? add_774682 : sel_774679;
  assign add_774686 = sel_774683 + 8'h01;
  assign sel_774687 = array_index_774630 == array_index_772720 ? add_774686 : sel_774683;
  assign add_774690 = sel_774687 + 8'h01;
  assign sel_774691 = array_index_774630 == array_index_772726 ? add_774690 : sel_774687;
  assign add_774694 = sel_774691 + 8'h01;
  assign sel_774695 = array_index_774630 == array_index_772732 ? add_774694 : sel_774691;
  assign add_774698 = sel_774695 + 8'h01;
  assign sel_774699 = array_index_774630 == array_index_772738 ? add_774698 : sel_774695;
  assign add_774702 = sel_774699 + 8'h01;
  assign sel_774703 = array_index_774630 == array_index_772744 ? add_774702 : sel_774699;
  assign add_774706 = sel_774703 + 8'h01;
  assign sel_774707 = array_index_774630 == array_index_772750 ? add_774706 : sel_774703;
  assign add_774710 = sel_774707 + 8'h01;
  assign sel_774711 = array_index_774630 == array_index_772756 ? add_774710 : sel_774707;
  assign add_774714 = sel_774711 + 8'h01;
  assign sel_774715 = array_index_774630 == array_index_772762 ? add_774714 : sel_774711;
  assign add_774718 = sel_774715 + 8'h01;
  assign sel_774719 = array_index_774630 == array_index_772768 ? add_774718 : sel_774715;
  assign add_774722 = sel_774719 + 8'h01;
  assign sel_774723 = array_index_774630 == array_index_772774 ? add_774722 : sel_774719;
  assign add_774726 = sel_774723 + 8'h01;
  assign sel_774727 = array_index_774630 == array_index_772780 ? add_774726 : sel_774723;
  assign add_774730 = sel_774727 + 8'h01;
  assign sel_774731 = array_index_774630 == array_index_772786 ? add_774730 : sel_774727;
  assign add_774734 = sel_774731 + 8'h01;
  assign sel_774735 = array_index_774630 == array_index_772792 ? add_774734 : sel_774731;
  assign add_774738 = sel_774735 + 8'h01;
  assign sel_774739 = array_index_774630 == array_index_772798 ? add_774738 : sel_774735;
  assign add_774742 = sel_774739 + 8'h01;
  assign sel_774743 = array_index_774630 == array_index_772804 ? add_774742 : sel_774739;
  assign add_774746 = sel_774743 + 8'h01;
  assign sel_774747 = array_index_774630 == array_index_772810 ? add_774746 : sel_774743;
  assign add_774750 = sel_774747 + 8'h01;
  assign sel_774751 = array_index_774630 == array_index_772816 ? add_774750 : sel_774747;
  assign add_774754 = sel_774751 + 8'h01;
  assign sel_774755 = array_index_774630 == array_index_772822 ? add_774754 : sel_774751;
  assign add_774758 = sel_774755 + 8'h01;
  assign sel_774759 = array_index_774630 == array_index_772828 ? add_774758 : sel_774755;
  assign add_774762 = sel_774759 + 8'h01;
  assign sel_774763 = array_index_774630 == array_index_772834 ? add_774762 : sel_774759;
  assign add_774766 = sel_774763 + 8'h01;
  assign sel_774767 = array_index_774630 == array_index_772840 ? add_774766 : sel_774763;
  assign add_774770 = sel_774767 + 8'h01;
  assign sel_774771 = array_index_774630 == array_index_772846 ? add_774770 : sel_774767;
  assign add_774774 = sel_774771 + 8'h01;
  assign sel_774775 = array_index_774630 == array_index_772852 ? add_774774 : sel_774771;
  assign add_774778 = sel_774775 + 8'h01;
  assign sel_774779 = array_index_774630 == array_index_772858 ? add_774778 : sel_774775;
  assign add_774782 = sel_774779 + 8'h01;
  assign sel_774783 = array_index_774630 == array_index_772864 ? add_774782 : sel_774779;
  assign add_774786 = sel_774783 + 8'h01;
  assign sel_774787 = array_index_774630 == array_index_772870 ? add_774786 : sel_774783;
  assign add_774790 = sel_774787 + 8'h01;
  assign sel_774791 = array_index_774630 == array_index_772876 ? add_774790 : sel_774787;
  assign add_774794 = sel_774791 + 8'h01;
  assign sel_774795 = array_index_774630 == array_index_772882 ? add_774794 : sel_774791;
  assign add_774798 = sel_774795 + 8'h01;
  assign sel_774799 = array_index_774630 == array_index_772888 ? add_774798 : sel_774795;
  assign add_774802 = sel_774799 + 8'h01;
  assign sel_774803 = array_index_774630 == array_index_772894 ? add_774802 : sel_774799;
  assign add_774806 = sel_774803 + 8'h01;
  assign sel_774807 = array_index_774630 == array_index_772900 ? add_774806 : sel_774803;
  assign add_774810 = sel_774807 + 8'h01;
  assign sel_774811 = array_index_774630 == array_index_772906 ? add_774810 : sel_774807;
  assign add_774814 = sel_774811 + 8'h01;
  assign sel_774815 = array_index_774630 == array_index_772912 ? add_774814 : sel_774811;
  assign add_774818 = sel_774815 + 8'h01;
  assign sel_774819 = array_index_774630 == array_index_772918 ? add_774818 : sel_774815;
  assign add_774822 = sel_774819 + 8'h01;
  assign sel_774823 = array_index_774630 == array_index_772924 ? add_774822 : sel_774819;
  assign add_774826 = sel_774823 + 8'h01;
  assign sel_774827 = array_index_774630 == array_index_772930 ? add_774826 : sel_774823;
  assign add_774830 = sel_774827 + 8'h01;
  assign sel_774831 = array_index_774630 == array_index_772936 ? add_774830 : sel_774827;
  assign add_774834 = sel_774831 + 8'h01;
  assign sel_774835 = array_index_774630 == array_index_772942 ? add_774834 : sel_774831;
  assign add_774838 = sel_774835 + 8'h01;
  assign sel_774839 = array_index_774630 == array_index_772948 ? add_774838 : sel_774835;
  assign add_774842 = sel_774839 + 8'h01;
  assign sel_774843 = array_index_774630 == array_index_772954 ? add_774842 : sel_774839;
  assign add_774846 = sel_774843 + 8'h01;
  assign sel_774847 = array_index_774630 == array_index_772960 ? add_774846 : sel_774843;
  assign add_774850 = sel_774847 + 8'h01;
  assign sel_774851 = array_index_774630 == array_index_772966 ? add_774850 : sel_774847;
  assign add_774854 = sel_774851 + 8'h01;
  assign sel_774855 = array_index_774630 == array_index_772972 ? add_774854 : sel_774851;
  assign add_774858 = sel_774855 + 8'h01;
  assign sel_774859 = array_index_774630 == array_index_772978 ? add_774858 : sel_774855;
  assign add_774862 = sel_774859 + 8'h01;
  assign sel_774863 = array_index_774630 == array_index_772984 ? add_774862 : sel_774859;
  assign add_774866 = sel_774863 + 8'h01;
  assign sel_774867 = array_index_774630 == array_index_772990 ? add_774866 : sel_774863;
  assign add_774870 = sel_774867 + 8'h01;
  assign sel_774871 = array_index_774630 == array_index_772996 ? add_774870 : sel_774867;
  assign add_774874 = sel_774871 + 8'h01;
  assign sel_774875 = array_index_774630 == array_index_773002 ? add_774874 : sel_774871;
  assign add_774878 = sel_774875 + 8'h01;
  assign sel_774879 = array_index_774630 == array_index_773008 ? add_774878 : sel_774875;
  assign add_774882 = sel_774879 + 8'h01;
  assign sel_774883 = array_index_774630 == array_index_773014 ? add_774882 : sel_774879;
  assign add_774886 = sel_774883 + 8'h01;
  assign sel_774887 = array_index_774630 == array_index_773020 ? add_774886 : sel_774883;
  assign add_774890 = sel_774887 + 8'h01;
  assign sel_774891 = array_index_774630 == array_index_773026 ? add_774890 : sel_774887;
  assign add_774894 = sel_774891 + 8'h01;
  assign sel_774895 = array_index_774630 == array_index_773032 ? add_774894 : sel_774891;
  assign add_774898 = sel_774895 + 8'h01;
  assign sel_774899 = array_index_774630 == array_index_773038 ? add_774898 : sel_774895;
  assign add_774902 = sel_774899 + 8'h01;
  assign sel_774903 = array_index_774630 == array_index_773044 ? add_774902 : sel_774899;
  assign add_774906 = sel_774903 + 8'h01;
  assign sel_774907 = array_index_774630 == array_index_773050 ? add_774906 : sel_774903;
  assign add_774910 = sel_774907 + 8'h01;
  assign sel_774911 = array_index_774630 == array_index_773056 ? add_774910 : sel_774907;
  assign add_774914 = sel_774911 + 8'h01;
  assign sel_774915 = array_index_774630 == array_index_773062 ? add_774914 : sel_774911;
  assign add_774918 = sel_774915 + 8'h01;
  assign sel_774919 = array_index_774630 == array_index_773068 ? add_774918 : sel_774915;
  assign add_774922 = sel_774919 + 8'h01;
  assign sel_774923 = array_index_774630 == array_index_773074 ? add_774922 : sel_774919;
  assign add_774926 = sel_774923 + 8'h01;
  assign sel_774927 = array_index_774630 == array_index_773080 ? add_774926 : sel_774923;
  assign add_774930 = sel_774927 + 8'h01;
  assign sel_774931 = array_index_774630 == array_index_773086 ? add_774930 : sel_774927;
  assign add_774934 = sel_774931 + 8'h01;
  assign sel_774935 = array_index_774630 == array_index_773092 ? add_774934 : sel_774931;
  assign add_774938 = sel_774935 + 8'h01;
  assign sel_774939 = array_index_774630 == array_index_773098 ? add_774938 : sel_774935;
  assign add_774942 = sel_774939 + 8'h01;
  assign sel_774943 = array_index_774630 == array_index_773104 ? add_774942 : sel_774939;
  assign add_774946 = sel_774943 + 8'h01;
  assign sel_774947 = array_index_774630 == array_index_773110 ? add_774946 : sel_774943;
  assign add_774950 = sel_774947 + 8'h01;
  assign sel_774951 = array_index_774630 == array_index_773116 ? add_774950 : sel_774947;
  assign add_774954 = sel_774951 + 8'h01;
  assign sel_774955 = array_index_774630 == array_index_773122 ? add_774954 : sel_774951;
  assign add_774958 = sel_774955 + 8'h01;
  assign sel_774959 = array_index_774630 == array_index_773128 ? add_774958 : sel_774955;
  assign add_774962 = sel_774959 + 8'h01;
  assign sel_774963 = array_index_774630 == array_index_773134 ? add_774962 : sel_774959;
  assign add_774966 = sel_774963 + 8'h01;
  assign sel_774967 = array_index_774630 == array_index_773140 ? add_774966 : sel_774963;
  assign add_774970 = sel_774967 + 8'h01;
  assign sel_774971 = array_index_774630 == array_index_773146 ? add_774970 : sel_774967;
  assign add_774974 = sel_774971 + 8'h01;
  assign sel_774975 = array_index_774630 == array_index_773152 ? add_774974 : sel_774971;
  assign add_774978 = sel_774975 + 8'h01;
  assign sel_774979 = array_index_774630 == array_index_773158 ? add_774978 : sel_774975;
  assign add_774982 = sel_774979 + 8'h01;
  assign sel_774983 = array_index_774630 == array_index_773164 ? add_774982 : sel_774979;
  assign add_774986 = sel_774983 + 8'h01;
  assign sel_774987 = array_index_774630 == array_index_773170 ? add_774986 : sel_774983;
  assign add_774991 = sel_774987 + 8'h01;
  assign array_index_774992 = set1_unflattened[7'h06];
  assign sel_774993 = array_index_774630 == array_index_773176 ? add_774991 : sel_774987;
  assign add_774996 = sel_774993 + 8'h01;
  assign sel_774997 = array_index_774992 == array_index_772632 ? add_774996 : sel_774993;
  assign add_775000 = sel_774997 + 8'h01;
  assign sel_775001 = array_index_774992 == array_index_772636 ? add_775000 : sel_774997;
  assign add_775004 = sel_775001 + 8'h01;
  assign sel_775005 = array_index_774992 == array_index_772644 ? add_775004 : sel_775001;
  assign add_775008 = sel_775005 + 8'h01;
  assign sel_775009 = array_index_774992 == array_index_772652 ? add_775008 : sel_775005;
  assign add_775012 = sel_775009 + 8'h01;
  assign sel_775013 = array_index_774992 == array_index_772660 ? add_775012 : sel_775009;
  assign add_775016 = sel_775013 + 8'h01;
  assign sel_775017 = array_index_774992 == array_index_772668 ? add_775016 : sel_775013;
  assign add_775020 = sel_775017 + 8'h01;
  assign sel_775021 = array_index_774992 == array_index_772676 ? add_775020 : sel_775017;
  assign add_775024 = sel_775021 + 8'h01;
  assign sel_775025 = array_index_774992 == array_index_772684 ? add_775024 : sel_775021;
  assign add_775028 = sel_775025 + 8'h01;
  assign sel_775029 = array_index_774992 == array_index_772690 ? add_775028 : sel_775025;
  assign add_775032 = sel_775029 + 8'h01;
  assign sel_775033 = array_index_774992 == array_index_772696 ? add_775032 : sel_775029;
  assign add_775036 = sel_775033 + 8'h01;
  assign sel_775037 = array_index_774992 == array_index_772702 ? add_775036 : sel_775033;
  assign add_775040 = sel_775037 + 8'h01;
  assign sel_775041 = array_index_774992 == array_index_772708 ? add_775040 : sel_775037;
  assign add_775044 = sel_775041 + 8'h01;
  assign sel_775045 = array_index_774992 == array_index_772714 ? add_775044 : sel_775041;
  assign add_775048 = sel_775045 + 8'h01;
  assign sel_775049 = array_index_774992 == array_index_772720 ? add_775048 : sel_775045;
  assign add_775052 = sel_775049 + 8'h01;
  assign sel_775053 = array_index_774992 == array_index_772726 ? add_775052 : sel_775049;
  assign add_775056 = sel_775053 + 8'h01;
  assign sel_775057 = array_index_774992 == array_index_772732 ? add_775056 : sel_775053;
  assign add_775060 = sel_775057 + 8'h01;
  assign sel_775061 = array_index_774992 == array_index_772738 ? add_775060 : sel_775057;
  assign add_775064 = sel_775061 + 8'h01;
  assign sel_775065 = array_index_774992 == array_index_772744 ? add_775064 : sel_775061;
  assign add_775068 = sel_775065 + 8'h01;
  assign sel_775069 = array_index_774992 == array_index_772750 ? add_775068 : sel_775065;
  assign add_775072 = sel_775069 + 8'h01;
  assign sel_775073 = array_index_774992 == array_index_772756 ? add_775072 : sel_775069;
  assign add_775076 = sel_775073 + 8'h01;
  assign sel_775077 = array_index_774992 == array_index_772762 ? add_775076 : sel_775073;
  assign add_775080 = sel_775077 + 8'h01;
  assign sel_775081 = array_index_774992 == array_index_772768 ? add_775080 : sel_775077;
  assign add_775084 = sel_775081 + 8'h01;
  assign sel_775085 = array_index_774992 == array_index_772774 ? add_775084 : sel_775081;
  assign add_775088 = sel_775085 + 8'h01;
  assign sel_775089 = array_index_774992 == array_index_772780 ? add_775088 : sel_775085;
  assign add_775092 = sel_775089 + 8'h01;
  assign sel_775093 = array_index_774992 == array_index_772786 ? add_775092 : sel_775089;
  assign add_775096 = sel_775093 + 8'h01;
  assign sel_775097 = array_index_774992 == array_index_772792 ? add_775096 : sel_775093;
  assign add_775100 = sel_775097 + 8'h01;
  assign sel_775101 = array_index_774992 == array_index_772798 ? add_775100 : sel_775097;
  assign add_775104 = sel_775101 + 8'h01;
  assign sel_775105 = array_index_774992 == array_index_772804 ? add_775104 : sel_775101;
  assign add_775108 = sel_775105 + 8'h01;
  assign sel_775109 = array_index_774992 == array_index_772810 ? add_775108 : sel_775105;
  assign add_775112 = sel_775109 + 8'h01;
  assign sel_775113 = array_index_774992 == array_index_772816 ? add_775112 : sel_775109;
  assign add_775116 = sel_775113 + 8'h01;
  assign sel_775117 = array_index_774992 == array_index_772822 ? add_775116 : sel_775113;
  assign add_775120 = sel_775117 + 8'h01;
  assign sel_775121 = array_index_774992 == array_index_772828 ? add_775120 : sel_775117;
  assign add_775124 = sel_775121 + 8'h01;
  assign sel_775125 = array_index_774992 == array_index_772834 ? add_775124 : sel_775121;
  assign add_775128 = sel_775125 + 8'h01;
  assign sel_775129 = array_index_774992 == array_index_772840 ? add_775128 : sel_775125;
  assign add_775132 = sel_775129 + 8'h01;
  assign sel_775133 = array_index_774992 == array_index_772846 ? add_775132 : sel_775129;
  assign add_775136 = sel_775133 + 8'h01;
  assign sel_775137 = array_index_774992 == array_index_772852 ? add_775136 : sel_775133;
  assign add_775140 = sel_775137 + 8'h01;
  assign sel_775141 = array_index_774992 == array_index_772858 ? add_775140 : sel_775137;
  assign add_775144 = sel_775141 + 8'h01;
  assign sel_775145 = array_index_774992 == array_index_772864 ? add_775144 : sel_775141;
  assign add_775148 = sel_775145 + 8'h01;
  assign sel_775149 = array_index_774992 == array_index_772870 ? add_775148 : sel_775145;
  assign add_775152 = sel_775149 + 8'h01;
  assign sel_775153 = array_index_774992 == array_index_772876 ? add_775152 : sel_775149;
  assign add_775156 = sel_775153 + 8'h01;
  assign sel_775157 = array_index_774992 == array_index_772882 ? add_775156 : sel_775153;
  assign add_775160 = sel_775157 + 8'h01;
  assign sel_775161 = array_index_774992 == array_index_772888 ? add_775160 : sel_775157;
  assign add_775164 = sel_775161 + 8'h01;
  assign sel_775165 = array_index_774992 == array_index_772894 ? add_775164 : sel_775161;
  assign add_775168 = sel_775165 + 8'h01;
  assign sel_775169 = array_index_774992 == array_index_772900 ? add_775168 : sel_775165;
  assign add_775172 = sel_775169 + 8'h01;
  assign sel_775173 = array_index_774992 == array_index_772906 ? add_775172 : sel_775169;
  assign add_775176 = sel_775173 + 8'h01;
  assign sel_775177 = array_index_774992 == array_index_772912 ? add_775176 : sel_775173;
  assign add_775180 = sel_775177 + 8'h01;
  assign sel_775181 = array_index_774992 == array_index_772918 ? add_775180 : sel_775177;
  assign add_775184 = sel_775181 + 8'h01;
  assign sel_775185 = array_index_774992 == array_index_772924 ? add_775184 : sel_775181;
  assign add_775188 = sel_775185 + 8'h01;
  assign sel_775189 = array_index_774992 == array_index_772930 ? add_775188 : sel_775185;
  assign add_775192 = sel_775189 + 8'h01;
  assign sel_775193 = array_index_774992 == array_index_772936 ? add_775192 : sel_775189;
  assign add_775196 = sel_775193 + 8'h01;
  assign sel_775197 = array_index_774992 == array_index_772942 ? add_775196 : sel_775193;
  assign add_775200 = sel_775197 + 8'h01;
  assign sel_775201 = array_index_774992 == array_index_772948 ? add_775200 : sel_775197;
  assign add_775204 = sel_775201 + 8'h01;
  assign sel_775205 = array_index_774992 == array_index_772954 ? add_775204 : sel_775201;
  assign add_775208 = sel_775205 + 8'h01;
  assign sel_775209 = array_index_774992 == array_index_772960 ? add_775208 : sel_775205;
  assign add_775212 = sel_775209 + 8'h01;
  assign sel_775213 = array_index_774992 == array_index_772966 ? add_775212 : sel_775209;
  assign add_775216 = sel_775213 + 8'h01;
  assign sel_775217 = array_index_774992 == array_index_772972 ? add_775216 : sel_775213;
  assign add_775220 = sel_775217 + 8'h01;
  assign sel_775221 = array_index_774992 == array_index_772978 ? add_775220 : sel_775217;
  assign add_775224 = sel_775221 + 8'h01;
  assign sel_775225 = array_index_774992 == array_index_772984 ? add_775224 : sel_775221;
  assign add_775228 = sel_775225 + 8'h01;
  assign sel_775229 = array_index_774992 == array_index_772990 ? add_775228 : sel_775225;
  assign add_775232 = sel_775229 + 8'h01;
  assign sel_775233 = array_index_774992 == array_index_772996 ? add_775232 : sel_775229;
  assign add_775236 = sel_775233 + 8'h01;
  assign sel_775237 = array_index_774992 == array_index_773002 ? add_775236 : sel_775233;
  assign add_775240 = sel_775237 + 8'h01;
  assign sel_775241 = array_index_774992 == array_index_773008 ? add_775240 : sel_775237;
  assign add_775244 = sel_775241 + 8'h01;
  assign sel_775245 = array_index_774992 == array_index_773014 ? add_775244 : sel_775241;
  assign add_775248 = sel_775245 + 8'h01;
  assign sel_775249 = array_index_774992 == array_index_773020 ? add_775248 : sel_775245;
  assign add_775252 = sel_775249 + 8'h01;
  assign sel_775253 = array_index_774992 == array_index_773026 ? add_775252 : sel_775249;
  assign add_775256 = sel_775253 + 8'h01;
  assign sel_775257 = array_index_774992 == array_index_773032 ? add_775256 : sel_775253;
  assign add_775260 = sel_775257 + 8'h01;
  assign sel_775261 = array_index_774992 == array_index_773038 ? add_775260 : sel_775257;
  assign add_775264 = sel_775261 + 8'h01;
  assign sel_775265 = array_index_774992 == array_index_773044 ? add_775264 : sel_775261;
  assign add_775268 = sel_775265 + 8'h01;
  assign sel_775269 = array_index_774992 == array_index_773050 ? add_775268 : sel_775265;
  assign add_775272 = sel_775269 + 8'h01;
  assign sel_775273 = array_index_774992 == array_index_773056 ? add_775272 : sel_775269;
  assign add_775276 = sel_775273 + 8'h01;
  assign sel_775277 = array_index_774992 == array_index_773062 ? add_775276 : sel_775273;
  assign add_775280 = sel_775277 + 8'h01;
  assign sel_775281 = array_index_774992 == array_index_773068 ? add_775280 : sel_775277;
  assign add_775284 = sel_775281 + 8'h01;
  assign sel_775285 = array_index_774992 == array_index_773074 ? add_775284 : sel_775281;
  assign add_775288 = sel_775285 + 8'h01;
  assign sel_775289 = array_index_774992 == array_index_773080 ? add_775288 : sel_775285;
  assign add_775292 = sel_775289 + 8'h01;
  assign sel_775293 = array_index_774992 == array_index_773086 ? add_775292 : sel_775289;
  assign add_775296 = sel_775293 + 8'h01;
  assign sel_775297 = array_index_774992 == array_index_773092 ? add_775296 : sel_775293;
  assign add_775300 = sel_775297 + 8'h01;
  assign sel_775301 = array_index_774992 == array_index_773098 ? add_775300 : sel_775297;
  assign add_775304 = sel_775301 + 8'h01;
  assign sel_775305 = array_index_774992 == array_index_773104 ? add_775304 : sel_775301;
  assign add_775308 = sel_775305 + 8'h01;
  assign sel_775309 = array_index_774992 == array_index_773110 ? add_775308 : sel_775305;
  assign add_775312 = sel_775309 + 8'h01;
  assign sel_775313 = array_index_774992 == array_index_773116 ? add_775312 : sel_775309;
  assign add_775316 = sel_775313 + 8'h01;
  assign sel_775317 = array_index_774992 == array_index_773122 ? add_775316 : sel_775313;
  assign add_775320 = sel_775317 + 8'h01;
  assign sel_775321 = array_index_774992 == array_index_773128 ? add_775320 : sel_775317;
  assign add_775324 = sel_775321 + 8'h01;
  assign sel_775325 = array_index_774992 == array_index_773134 ? add_775324 : sel_775321;
  assign add_775328 = sel_775325 + 8'h01;
  assign sel_775329 = array_index_774992 == array_index_773140 ? add_775328 : sel_775325;
  assign add_775332 = sel_775329 + 8'h01;
  assign sel_775333 = array_index_774992 == array_index_773146 ? add_775332 : sel_775329;
  assign add_775336 = sel_775333 + 8'h01;
  assign sel_775337 = array_index_774992 == array_index_773152 ? add_775336 : sel_775333;
  assign add_775340 = sel_775337 + 8'h01;
  assign sel_775341 = array_index_774992 == array_index_773158 ? add_775340 : sel_775337;
  assign add_775344 = sel_775341 + 8'h01;
  assign sel_775345 = array_index_774992 == array_index_773164 ? add_775344 : sel_775341;
  assign add_775348 = sel_775345 + 8'h01;
  assign sel_775349 = array_index_774992 == array_index_773170 ? add_775348 : sel_775345;
  assign add_775353 = sel_775349 + 8'h01;
  assign array_index_775354 = set1_unflattened[7'h07];
  assign sel_775355 = array_index_774992 == array_index_773176 ? add_775353 : sel_775349;
  assign add_775358 = sel_775355 + 8'h01;
  assign sel_775359 = array_index_775354 == array_index_772632 ? add_775358 : sel_775355;
  assign add_775362 = sel_775359 + 8'h01;
  assign sel_775363 = array_index_775354 == array_index_772636 ? add_775362 : sel_775359;
  assign add_775366 = sel_775363 + 8'h01;
  assign sel_775367 = array_index_775354 == array_index_772644 ? add_775366 : sel_775363;
  assign add_775370 = sel_775367 + 8'h01;
  assign sel_775371 = array_index_775354 == array_index_772652 ? add_775370 : sel_775367;
  assign add_775374 = sel_775371 + 8'h01;
  assign sel_775375 = array_index_775354 == array_index_772660 ? add_775374 : sel_775371;
  assign add_775378 = sel_775375 + 8'h01;
  assign sel_775379 = array_index_775354 == array_index_772668 ? add_775378 : sel_775375;
  assign add_775382 = sel_775379 + 8'h01;
  assign sel_775383 = array_index_775354 == array_index_772676 ? add_775382 : sel_775379;
  assign add_775386 = sel_775383 + 8'h01;
  assign sel_775387 = array_index_775354 == array_index_772684 ? add_775386 : sel_775383;
  assign add_775390 = sel_775387 + 8'h01;
  assign sel_775391 = array_index_775354 == array_index_772690 ? add_775390 : sel_775387;
  assign add_775394 = sel_775391 + 8'h01;
  assign sel_775395 = array_index_775354 == array_index_772696 ? add_775394 : sel_775391;
  assign add_775398 = sel_775395 + 8'h01;
  assign sel_775399 = array_index_775354 == array_index_772702 ? add_775398 : sel_775395;
  assign add_775402 = sel_775399 + 8'h01;
  assign sel_775403 = array_index_775354 == array_index_772708 ? add_775402 : sel_775399;
  assign add_775406 = sel_775403 + 8'h01;
  assign sel_775407 = array_index_775354 == array_index_772714 ? add_775406 : sel_775403;
  assign add_775410 = sel_775407 + 8'h01;
  assign sel_775411 = array_index_775354 == array_index_772720 ? add_775410 : sel_775407;
  assign add_775414 = sel_775411 + 8'h01;
  assign sel_775415 = array_index_775354 == array_index_772726 ? add_775414 : sel_775411;
  assign add_775418 = sel_775415 + 8'h01;
  assign sel_775419 = array_index_775354 == array_index_772732 ? add_775418 : sel_775415;
  assign add_775422 = sel_775419 + 8'h01;
  assign sel_775423 = array_index_775354 == array_index_772738 ? add_775422 : sel_775419;
  assign add_775426 = sel_775423 + 8'h01;
  assign sel_775427 = array_index_775354 == array_index_772744 ? add_775426 : sel_775423;
  assign add_775430 = sel_775427 + 8'h01;
  assign sel_775431 = array_index_775354 == array_index_772750 ? add_775430 : sel_775427;
  assign add_775434 = sel_775431 + 8'h01;
  assign sel_775435 = array_index_775354 == array_index_772756 ? add_775434 : sel_775431;
  assign add_775438 = sel_775435 + 8'h01;
  assign sel_775439 = array_index_775354 == array_index_772762 ? add_775438 : sel_775435;
  assign add_775442 = sel_775439 + 8'h01;
  assign sel_775443 = array_index_775354 == array_index_772768 ? add_775442 : sel_775439;
  assign add_775446 = sel_775443 + 8'h01;
  assign sel_775447 = array_index_775354 == array_index_772774 ? add_775446 : sel_775443;
  assign add_775450 = sel_775447 + 8'h01;
  assign sel_775451 = array_index_775354 == array_index_772780 ? add_775450 : sel_775447;
  assign add_775454 = sel_775451 + 8'h01;
  assign sel_775455 = array_index_775354 == array_index_772786 ? add_775454 : sel_775451;
  assign add_775458 = sel_775455 + 8'h01;
  assign sel_775459 = array_index_775354 == array_index_772792 ? add_775458 : sel_775455;
  assign add_775462 = sel_775459 + 8'h01;
  assign sel_775463 = array_index_775354 == array_index_772798 ? add_775462 : sel_775459;
  assign add_775466 = sel_775463 + 8'h01;
  assign sel_775467 = array_index_775354 == array_index_772804 ? add_775466 : sel_775463;
  assign add_775470 = sel_775467 + 8'h01;
  assign sel_775471 = array_index_775354 == array_index_772810 ? add_775470 : sel_775467;
  assign add_775474 = sel_775471 + 8'h01;
  assign sel_775475 = array_index_775354 == array_index_772816 ? add_775474 : sel_775471;
  assign add_775478 = sel_775475 + 8'h01;
  assign sel_775479 = array_index_775354 == array_index_772822 ? add_775478 : sel_775475;
  assign add_775482 = sel_775479 + 8'h01;
  assign sel_775483 = array_index_775354 == array_index_772828 ? add_775482 : sel_775479;
  assign add_775486 = sel_775483 + 8'h01;
  assign sel_775487 = array_index_775354 == array_index_772834 ? add_775486 : sel_775483;
  assign add_775490 = sel_775487 + 8'h01;
  assign sel_775491 = array_index_775354 == array_index_772840 ? add_775490 : sel_775487;
  assign add_775494 = sel_775491 + 8'h01;
  assign sel_775495 = array_index_775354 == array_index_772846 ? add_775494 : sel_775491;
  assign add_775498 = sel_775495 + 8'h01;
  assign sel_775499 = array_index_775354 == array_index_772852 ? add_775498 : sel_775495;
  assign add_775502 = sel_775499 + 8'h01;
  assign sel_775503 = array_index_775354 == array_index_772858 ? add_775502 : sel_775499;
  assign add_775506 = sel_775503 + 8'h01;
  assign sel_775507 = array_index_775354 == array_index_772864 ? add_775506 : sel_775503;
  assign add_775510 = sel_775507 + 8'h01;
  assign sel_775511 = array_index_775354 == array_index_772870 ? add_775510 : sel_775507;
  assign add_775514 = sel_775511 + 8'h01;
  assign sel_775515 = array_index_775354 == array_index_772876 ? add_775514 : sel_775511;
  assign add_775518 = sel_775515 + 8'h01;
  assign sel_775519 = array_index_775354 == array_index_772882 ? add_775518 : sel_775515;
  assign add_775522 = sel_775519 + 8'h01;
  assign sel_775523 = array_index_775354 == array_index_772888 ? add_775522 : sel_775519;
  assign add_775526 = sel_775523 + 8'h01;
  assign sel_775527 = array_index_775354 == array_index_772894 ? add_775526 : sel_775523;
  assign add_775530 = sel_775527 + 8'h01;
  assign sel_775531 = array_index_775354 == array_index_772900 ? add_775530 : sel_775527;
  assign add_775534 = sel_775531 + 8'h01;
  assign sel_775535 = array_index_775354 == array_index_772906 ? add_775534 : sel_775531;
  assign add_775538 = sel_775535 + 8'h01;
  assign sel_775539 = array_index_775354 == array_index_772912 ? add_775538 : sel_775535;
  assign add_775542 = sel_775539 + 8'h01;
  assign sel_775543 = array_index_775354 == array_index_772918 ? add_775542 : sel_775539;
  assign add_775546 = sel_775543 + 8'h01;
  assign sel_775547 = array_index_775354 == array_index_772924 ? add_775546 : sel_775543;
  assign add_775550 = sel_775547 + 8'h01;
  assign sel_775551 = array_index_775354 == array_index_772930 ? add_775550 : sel_775547;
  assign add_775554 = sel_775551 + 8'h01;
  assign sel_775555 = array_index_775354 == array_index_772936 ? add_775554 : sel_775551;
  assign add_775558 = sel_775555 + 8'h01;
  assign sel_775559 = array_index_775354 == array_index_772942 ? add_775558 : sel_775555;
  assign add_775562 = sel_775559 + 8'h01;
  assign sel_775563 = array_index_775354 == array_index_772948 ? add_775562 : sel_775559;
  assign add_775566 = sel_775563 + 8'h01;
  assign sel_775567 = array_index_775354 == array_index_772954 ? add_775566 : sel_775563;
  assign add_775570 = sel_775567 + 8'h01;
  assign sel_775571 = array_index_775354 == array_index_772960 ? add_775570 : sel_775567;
  assign add_775574 = sel_775571 + 8'h01;
  assign sel_775575 = array_index_775354 == array_index_772966 ? add_775574 : sel_775571;
  assign add_775578 = sel_775575 + 8'h01;
  assign sel_775579 = array_index_775354 == array_index_772972 ? add_775578 : sel_775575;
  assign add_775582 = sel_775579 + 8'h01;
  assign sel_775583 = array_index_775354 == array_index_772978 ? add_775582 : sel_775579;
  assign add_775586 = sel_775583 + 8'h01;
  assign sel_775587 = array_index_775354 == array_index_772984 ? add_775586 : sel_775583;
  assign add_775590 = sel_775587 + 8'h01;
  assign sel_775591 = array_index_775354 == array_index_772990 ? add_775590 : sel_775587;
  assign add_775594 = sel_775591 + 8'h01;
  assign sel_775595 = array_index_775354 == array_index_772996 ? add_775594 : sel_775591;
  assign add_775598 = sel_775595 + 8'h01;
  assign sel_775599 = array_index_775354 == array_index_773002 ? add_775598 : sel_775595;
  assign add_775602 = sel_775599 + 8'h01;
  assign sel_775603 = array_index_775354 == array_index_773008 ? add_775602 : sel_775599;
  assign add_775606 = sel_775603 + 8'h01;
  assign sel_775607 = array_index_775354 == array_index_773014 ? add_775606 : sel_775603;
  assign add_775610 = sel_775607 + 8'h01;
  assign sel_775611 = array_index_775354 == array_index_773020 ? add_775610 : sel_775607;
  assign add_775614 = sel_775611 + 8'h01;
  assign sel_775615 = array_index_775354 == array_index_773026 ? add_775614 : sel_775611;
  assign add_775618 = sel_775615 + 8'h01;
  assign sel_775619 = array_index_775354 == array_index_773032 ? add_775618 : sel_775615;
  assign add_775622 = sel_775619 + 8'h01;
  assign sel_775623 = array_index_775354 == array_index_773038 ? add_775622 : sel_775619;
  assign add_775626 = sel_775623 + 8'h01;
  assign sel_775627 = array_index_775354 == array_index_773044 ? add_775626 : sel_775623;
  assign add_775630 = sel_775627 + 8'h01;
  assign sel_775631 = array_index_775354 == array_index_773050 ? add_775630 : sel_775627;
  assign add_775634 = sel_775631 + 8'h01;
  assign sel_775635 = array_index_775354 == array_index_773056 ? add_775634 : sel_775631;
  assign add_775638 = sel_775635 + 8'h01;
  assign sel_775639 = array_index_775354 == array_index_773062 ? add_775638 : sel_775635;
  assign add_775642 = sel_775639 + 8'h01;
  assign sel_775643 = array_index_775354 == array_index_773068 ? add_775642 : sel_775639;
  assign add_775646 = sel_775643 + 8'h01;
  assign sel_775647 = array_index_775354 == array_index_773074 ? add_775646 : sel_775643;
  assign add_775650 = sel_775647 + 8'h01;
  assign sel_775651 = array_index_775354 == array_index_773080 ? add_775650 : sel_775647;
  assign add_775654 = sel_775651 + 8'h01;
  assign sel_775655 = array_index_775354 == array_index_773086 ? add_775654 : sel_775651;
  assign add_775658 = sel_775655 + 8'h01;
  assign sel_775659 = array_index_775354 == array_index_773092 ? add_775658 : sel_775655;
  assign add_775662 = sel_775659 + 8'h01;
  assign sel_775663 = array_index_775354 == array_index_773098 ? add_775662 : sel_775659;
  assign add_775666 = sel_775663 + 8'h01;
  assign sel_775667 = array_index_775354 == array_index_773104 ? add_775666 : sel_775663;
  assign add_775670 = sel_775667 + 8'h01;
  assign sel_775671 = array_index_775354 == array_index_773110 ? add_775670 : sel_775667;
  assign add_775674 = sel_775671 + 8'h01;
  assign sel_775675 = array_index_775354 == array_index_773116 ? add_775674 : sel_775671;
  assign add_775678 = sel_775675 + 8'h01;
  assign sel_775679 = array_index_775354 == array_index_773122 ? add_775678 : sel_775675;
  assign add_775682 = sel_775679 + 8'h01;
  assign sel_775683 = array_index_775354 == array_index_773128 ? add_775682 : sel_775679;
  assign add_775686 = sel_775683 + 8'h01;
  assign sel_775687 = array_index_775354 == array_index_773134 ? add_775686 : sel_775683;
  assign add_775690 = sel_775687 + 8'h01;
  assign sel_775691 = array_index_775354 == array_index_773140 ? add_775690 : sel_775687;
  assign add_775694 = sel_775691 + 8'h01;
  assign sel_775695 = array_index_775354 == array_index_773146 ? add_775694 : sel_775691;
  assign add_775698 = sel_775695 + 8'h01;
  assign sel_775699 = array_index_775354 == array_index_773152 ? add_775698 : sel_775695;
  assign add_775702 = sel_775699 + 8'h01;
  assign sel_775703 = array_index_775354 == array_index_773158 ? add_775702 : sel_775699;
  assign add_775706 = sel_775703 + 8'h01;
  assign sel_775707 = array_index_775354 == array_index_773164 ? add_775706 : sel_775703;
  assign add_775710 = sel_775707 + 8'h01;
  assign sel_775711 = array_index_775354 == array_index_773170 ? add_775710 : sel_775707;
  assign add_775715 = sel_775711 + 8'h01;
  assign array_index_775716 = set1_unflattened[7'h08];
  assign sel_775717 = array_index_775354 == array_index_773176 ? add_775715 : sel_775711;
  assign add_775720 = sel_775717 + 8'h01;
  assign sel_775721 = array_index_775716 == array_index_772632 ? add_775720 : sel_775717;
  assign add_775724 = sel_775721 + 8'h01;
  assign sel_775725 = array_index_775716 == array_index_772636 ? add_775724 : sel_775721;
  assign add_775728 = sel_775725 + 8'h01;
  assign sel_775729 = array_index_775716 == array_index_772644 ? add_775728 : sel_775725;
  assign add_775732 = sel_775729 + 8'h01;
  assign sel_775733 = array_index_775716 == array_index_772652 ? add_775732 : sel_775729;
  assign add_775736 = sel_775733 + 8'h01;
  assign sel_775737 = array_index_775716 == array_index_772660 ? add_775736 : sel_775733;
  assign add_775740 = sel_775737 + 8'h01;
  assign sel_775741 = array_index_775716 == array_index_772668 ? add_775740 : sel_775737;
  assign add_775744 = sel_775741 + 8'h01;
  assign sel_775745 = array_index_775716 == array_index_772676 ? add_775744 : sel_775741;
  assign add_775748 = sel_775745 + 8'h01;
  assign sel_775749 = array_index_775716 == array_index_772684 ? add_775748 : sel_775745;
  assign add_775752 = sel_775749 + 8'h01;
  assign sel_775753 = array_index_775716 == array_index_772690 ? add_775752 : sel_775749;
  assign add_775756 = sel_775753 + 8'h01;
  assign sel_775757 = array_index_775716 == array_index_772696 ? add_775756 : sel_775753;
  assign add_775760 = sel_775757 + 8'h01;
  assign sel_775761 = array_index_775716 == array_index_772702 ? add_775760 : sel_775757;
  assign add_775764 = sel_775761 + 8'h01;
  assign sel_775765 = array_index_775716 == array_index_772708 ? add_775764 : sel_775761;
  assign add_775768 = sel_775765 + 8'h01;
  assign sel_775769 = array_index_775716 == array_index_772714 ? add_775768 : sel_775765;
  assign add_775772 = sel_775769 + 8'h01;
  assign sel_775773 = array_index_775716 == array_index_772720 ? add_775772 : sel_775769;
  assign add_775776 = sel_775773 + 8'h01;
  assign sel_775777 = array_index_775716 == array_index_772726 ? add_775776 : sel_775773;
  assign add_775780 = sel_775777 + 8'h01;
  assign sel_775781 = array_index_775716 == array_index_772732 ? add_775780 : sel_775777;
  assign add_775784 = sel_775781 + 8'h01;
  assign sel_775785 = array_index_775716 == array_index_772738 ? add_775784 : sel_775781;
  assign add_775788 = sel_775785 + 8'h01;
  assign sel_775789 = array_index_775716 == array_index_772744 ? add_775788 : sel_775785;
  assign add_775792 = sel_775789 + 8'h01;
  assign sel_775793 = array_index_775716 == array_index_772750 ? add_775792 : sel_775789;
  assign add_775796 = sel_775793 + 8'h01;
  assign sel_775797 = array_index_775716 == array_index_772756 ? add_775796 : sel_775793;
  assign add_775800 = sel_775797 + 8'h01;
  assign sel_775801 = array_index_775716 == array_index_772762 ? add_775800 : sel_775797;
  assign add_775804 = sel_775801 + 8'h01;
  assign sel_775805 = array_index_775716 == array_index_772768 ? add_775804 : sel_775801;
  assign add_775808 = sel_775805 + 8'h01;
  assign sel_775809 = array_index_775716 == array_index_772774 ? add_775808 : sel_775805;
  assign add_775812 = sel_775809 + 8'h01;
  assign sel_775813 = array_index_775716 == array_index_772780 ? add_775812 : sel_775809;
  assign add_775816 = sel_775813 + 8'h01;
  assign sel_775817 = array_index_775716 == array_index_772786 ? add_775816 : sel_775813;
  assign add_775820 = sel_775817 + 8'h01;
  assign sel_775821 = array_index_775716 == array_index_772792 ? add_775820 : sel_775817;
  assign add_775824 = sel_775821 + 8'h01;
  assign sel_775825 = array_index_775716 == array_index_772798 ? add_775824 : sel_775821;
  assign add_775828 = sel_775825 + 8'h01;
  assign sel_775829 = array_index_775716 == array_index_772804 ? add_775828 : sel_775825;
  assign add_775832 = sel_775829 + 8'h01;
  assign sel_775833 = array_index_775716 == array_index_772810 ? add_775832 : sel_775829;
  assign add_775836 = sel_775833 + 8'h01;
  assign sel_775837 = array_index_775716 == array_index_772816 ? add_775836 : sel_775833;
  assign add_775840 = sel_775837 + 8'h01;
  assign sel_775841 = array_index_775716 == array_index_772822 ? add_775840 : sel_775837;
  assign add_775844 = sel_775841 + 8'h01;
  assign sel_775845 = array_index_775716 == array_index_772828 ? add_775844 : sel_775841;
  assign add_775848 = sel_775845 + 8'h01;
  assign sel_775849 = array_index_775716 == array_index_772834 ? add_775848 : sel_775845;
  assign add_775852 = sel_775849 + 8'h01;
  assign sel_775853 = array_index_775716 == array_index_772840 ? add_775852 : sel_775849;
  assign add_775856 = sel_775853 + 8'h01;
  assign sel_775857 = array_index_775716 == array_index_772846 ? add_775856 : sel_775853;
  assign add_775860 = sel_775857 + 8'h01;
  assign sel_775861 = array_index_775716 == array_index_772852 ? add_775860 : sel_775857;
  assign add_775864 = sel_775861 + 8'h01;
  assign sel_775865 = array_index_775716 == array_index_772858 ? add_775864 : sel_775861;
  assign add_775868 = sel_775865 + 8'h01;
  assign sel_775869 = array_index_775716 == array_index_772864 ? add_775868 : sel_775865;
  assign add_775872 = sel_775869 + 8'h01;
  assign sel_775873 = array_index_775716 == array_index_772870 ? add_775872 : sel_775869;
  assign add_775876 = sel_775873 + 8'h01;
  assign sel_775877 = array_index_775716 == array_index_772876 ? add_775876 : sel_775873;
  assign add_775880 = sel_775877 + 8'h01;
  assign sel_775881 = array_index_775716 == array_index_772882 ? add_775880 : sel_775877;
  assign add_775884 = sel_775881 + 8'h01;
  assign sel_775885 = array_index_775716 == array_index_772888 ? add_775884 : sel_775881;
  assign add_775888 = sel_775885 + 8'h01;
  assign sel_775889 = array_index_775716 == array_index_772894 ? add_775888 : sel_775885;
  assign add_775892 = sel_775889 + 8'h01;
  assign sel_775893 = array_index_775716 == array_index_772900 ? add_775892 : sel_775889;
  assign add_775896 = sel_775893 + 8'h01;
  assign sel_775897 = array_index_775716 == array_index_772906 ? add_775896 : sel_775893;
  assign add_775900 = sel_775897 + 8'h01;
  assign sel_775901 = array_index_775716 == array_index_772912 ? add_775900 : sel_775897;
  assign add_775904 = sel_775901 + 8'h01;
  assign sel_775905 = array_index_775716 == array_index_772918 ? add_775904 : sel_775901;
  assign add_775908 = sel_775905 + 8'h01;
  assign sel_775909 = array_index_775716 == array_index_772924 ? add_775908 : sel_775905;
  assign add_775912 = sel_775909 + 8'h01;
  assign sel_775913 = array_index_775716 == array_index_772930 ? add_775912 : sel_775909;
  assign add_775916 = sel_775913 + 8'h01;
  assign sel_775917 = array_index_775716 == array_index_772936 ? add_775916 : sel_775913;
  assign add_775920 = sel_775917 + 8'h01;
  assign sel_775921 = array_index_775716 == array_index_772942 ? add_775920 : sel_775917;
  assign add_775924 = sel_775921 + 8'h01;
  assign sel_775925 = array_index_775716 == array_index_772948 ? add_775924 : sel_775921;
  assign add_775928 = sel_775925 + 8'h01;
  assign sel_775929 = array_index_775716 == array_index_772954 ? add_775928 : sel_775925;
  assign add_775932 = sel_775929 + 8'h01;
  assign sel_775933 = array_index_775716 == array_index_772960 ? add_775932 : sel_775929;
  assign add_775936 = sel_775933 + 8'h01;
  assign sel_775937 = array_index_775716 == array_index_772966 ? add_775936 : sel_775933;
  assign add_775940 = sel_775937 + 8'h01;
  assign sel_775941 = array_index_775716 == array_index_772972 ? add_775940 : sel_775937;
  assign add_775944 = sel_775941 + 8'h01;
  assign sel_775945 = array_index_775716 == array_index_772978 ? add_775944 : sel_775941;
  assign add_775948 = sel_775945 + 8'h01;
  assign sel_775949 = array_index_775716 == array_index_772984 ? add_775948 : sel_775945;
  assign add_775952 = sel_775949 + 8'h01;
  assign sel_775953 = array_index_775716 == array_index_772990 ? add_775952 : sel_775949;
  assign add_775956 = sel_775953 + 8'h01;
  assign sel_775957 = array_index_775716 == array_index_772996 ? add_775956 : sel_775953;
  assign add_775960 = sel_775957 + 8'h01;
  assign sel_775961 = array_index_775716 == array_index_773002 ? add_775960 : sel_775957;
  assign add_775964 = sel_775961 + 8'h01;
  assign sel_775965 = array_index_775716 == array_index_773008 ? add_775964 : sel_775961;
  assign add_775968 = sel_775965 + 8'h01;
  assign sel_775969 = array_index_775716 == array_index_773014 ? add_775968 : sel_775965;
  assign add_775972 = sel_775969 + 8'h01;
  assign sel_775973 = array_index_775716 == array_index_773020 ? add_775972 : sel_775969;
  assign add_775976 = sel_775973 + 8'h01;
  assign sel_775977 = array_index_775716 == array_index_773026 ? add_775976 : sel_775973;
  assign add_775980 = sel_775977 + 8'h01;
  assign sel_775981 = array_index_775716 == array_index_773032 ? add_775980 : sel_775977;
  assign add_775984 = sel_775981 + 8'h01;
  assign sel_775985 = array_index_775716 == array_index_773038 ? add_775984 : sel_775981;
  assign add_775988 = sel_775985 + 8'h01;
  assign sel_775989 = array_index_775716 == array_index_773044 ? add_775988 : sel_775985;
  assign add_775992 = sel_775989 + 8'h01;
  assign sel_775993 = array_index_775716 == array_index_773050 ? add_775992 : sel_775989;
  assign add_775996 = sel_775993 + 8'h01;
  assign sel_775997 = array_index_775716 == array_index_773056 ? add_775996 : sel_775993;
  assign add_776000 = sel_775997 + 8'h01;
  assign sel_776001 = array_index_775716 == array_index_773062 ? add_776000 : sel_775997;
  assign add_776004 = sel_776001 + 8'h01;
  assign sel_776005 = array_index_775716 == array_index_773068 ? add_776004 : sel_776001;
  assign add_776008 = sel_776005 + 8'h01;
  assign sel_776009 = array_index_775716 == array_index_773074 ? add_776008 : sel_776005;
  assign add_776012 = sel_776009 + 8'h01;
  assign sel_776013 = array_index_775716 == array_index_773080 ? add_776012 : sel_776009;
  assign add_776016 = sel_776013 + 8'h01;
  assign sel_776017 = array_index_775716 == array_index_773086 ? add_776016 : sel_776013;
  assign add_776020 = sel_776017 + 8'h01;
  assign sel_776021 = array_index_775716 == array_index_773092 ? add_776020 : sel_776017;
  assign add_776024 = sel_776021 + 8'h01;
  assign sel_776025 = array_index_775716 == array_index_773098 ? add_776024 : sel_776021;
  assign add_776028 = sel_776025 + 8'h01;
  assign sel_776029 = array_index_775716 == array_index_773104 ? add_776028 : sel_776025;
  assign add_776032 = sel_776029 + 8'h01;
  assign sel_776033 = array_index_775716 == array_index_773110 ? add_776032 : sel_776029;
  assign add_776036 = sel_776033 + 8'h01;
  assign sel_776037 = array_index_775716 == array_index_773116 ? add_776036 : sel_776033;
  assign add_776040 = sel_776037 + 8'h01;
  assign sel_776041 = array_index_775716 == array_index_773122 ? add_776040 : sel_776037;
  assign add_776044 = sel_776041 + 8'h01;
  assign sel_776045 = array_index_775716 == array_index_773128 ? add_776044 : sel_776041;
  assign add_776048 = sel_776045 + 8'h01;
  assign sel_776049 = array_index_775716 == array_index_773134 ? add_776048 : sel_776045;
  assign add_776052 = sel_776049 + 8'h01;
  assign sel_776053 = array_index_775716 == array_index_773140 ? add_776052 : sel_776049;
  assign add_776056 = sel_776053 + 8'h01;
  assign sel_776057 = array_index_775716 == array_index_773146 ? add_776056 : sel_776053;
  assign add_776060 = sel_776057 + 8'h01;
  assign sel_776061 = array_index_775716 == array_index_773152 ? add_776060 : sel_776057;
  assign add_776064 = sel_776061 + 8'h01;
  assign sel_776065 = array_index_775716 == array_index_773158 ? add_776064 : sel_776061;
  assign add_776068 = sel_776065 + 8'h01;
  assign sel_776069 = array_index_775716 == array_index_773164 ? add_776068 : sel_776065;
  assign add_776072 = sel_776069 + 8'h01;
  assign sel_776073 = array_index_775716 == array_index_773170 ? add_776072 : sel_776069;
  assign add_776077 = sel_776073 + 8'h01;
  assign array_index_776078 = set1_unflattened[7'h09];
  assign sel_776079 = array_index_775716 == array_index_773176 ? add_776077 : sel_776073;
  assign add_776082 = sel_776079 + 8'h01;
  assign sel_776083 = array_index_776078 == array_index_772632 ? add_776082 : sel_776079;
  assign add_776086 = sel_776083 + 8'h01;
  assign sel_776087 = array_index_776078 == array_index_772636 ? add_776086 : sel_776083;
  assign add_776090 = sel_776087 + 8'h01;
  assign sel_776091 = array_index_776078 == array_index_772644 ? add_776090 : sel_776087;
  assign add_776094 = sel_776091 + 8'h01;
  assign sel_776095 = array_index_776078 == array_index_772652 ? add_776094 : sel_776091;
  assign add_776098 = sel_776095 + 8'h01;
  assign sel_776099 = array_index_776078 == array_index_772660 ? add_776098 : sel_776095;
  assign add_776102 = sel_776099 + 8'h01;
  assign sel_776103 = array_index_776078 == array_index_772668 ? add_776102 : sel_776099;
  assign add_776106 = sel_776103 + 8'h01;
  assign sel_776107 = array_index_776078 == array_index_772676 ? add_776106 : sel_776103;
  assign add_776110 = sel_776107 + 8'h01;
  assign sel_776111 = array_index_776078 == array_index_772684 ? add_776110 : sel_776107;
  assign add_776114 = sel_776111 + 8'h01;
  assign sel_776115 = array_index_776078 == array_index_772690 ? add_776114 : sel_776111;
  assign add_776118 = sel_776115 + 8'h01;
  assign sel_776119 = array_index_776078 == array_index_772696 ? add_776118 : sel_776115;
  assign add_776122 = sel_776119 + 8'h01;
  assign sel_776123 = array_index_776078 == array_index_772702 ? add_776122 : sel_776119;
  assign add_776126 = sel_776123 + 8'h01;
  assign sel_776127 = array_index_776078 == array_index_772708 ? add_776126 : sel_776123;
  assign add_776130 = sel_776127 + 8'h01;
  assign sel_776131 = array_index_776078 == array_index_772714 ? add_776130 : sel_776127;
  assign add_776134 = sel_776131 + 8'h01;
  assign sel_776135 = array_index_776078 == array_index_772720 ? add_776134 : sel_776131;
  assign add_776138 = sel_776135 + 8'h01;
  assign sel_776139 = array_index_776078 == array_index_772726 ? add_776138 : sel_776135;
  assign add_776142 = sel_776139 + 8'h01;
  assign sel_776143 = array_index_776078 == array_index_772732 ? add_776142 : sel_776139;
  assign add_776146 = sel_776143 + 8'h01;
  assign sel_776147 = array_index_776078 == array_index_772738 ? add_776146 : sel_776143;
  assign add_776150 = sel_776147 + 8'h01;
  assign sel_776151 = array_index_776078 == array_index_772744 ? add_776150 : sel_776147;
  assign add_776154 = sel_776151 + 8'h01;
  assign sel_776155 = array_index_776078 == array_index_772750 ? add_776154 : sel_776151;
  assign add_776158 = sel_776155 + 8'h01;
  assign sel_776159 = array_index_776078 == array_index_772756 ? add_776158 : sel_776155;
  assign add_776162 = sel_776159 + 8'h01;
  assign sel_776163 = array_index_776078 == array_index_772762 ? add_776162 : sel_776159;
  assign add_776166 = sel_776163 + 8'h01;
  assign sel_776167 = array_index_776078 == array_index_772768 ? add_776166 : sel_776163;
  assign add_776170 = sel_776167 + 8'h01;
  assign sel_776171 = array_index_776078 == array_index_772774 ? add_776170 : sel_776167;
  assign add_776174 = sel_776171 + 8'h01;
  assign sel_776175 = array_index_776078 == array_index_772780 ? add_776174 : sel_776171;
  assign add_776178 = sel_776175 + 8'h01;
  assign sel_776179 = array_index_776078 == array_index_772786 ? add_776178 : sel_776175;
  assign add_776182 = sel_776179 + 8'h01;
  assign sel_776183 = array_index_776078 == array_index_772792 ? add_776182 : sel_776179;
  assign add_776186 = sel_776183 + 8'h01;
  assign sel_776187 = array_index_776078 == array_index_772798 ? add_776186 : sel_776183;
  assign add_776190 = sel_776187 + 8'h01;
  assign sel_776191 = array_index_776078 == array_index_772804 ? add_776190 : sel_776187;
  assign add_776194 = sel_776191 + 8'h01;
  assign sel_776195 = array_index_776078 == array_index_772810 ? add_776194 : sel_776191;
  assign add_776198 = sel_776195 + 8'h01;
  assign sel_776199 = array_index_776078 == array_index_772816 ? add_776198 : sel_776195;
  assign add_776202 = sel_776199 + 8'h01;
  assign sel_776203 = array_index_776078 == array_index_772822 ? add_776202 : sel_776199;
  assign add_776206 = sel_776203 + 8'h01;
  assign sel_776207 = array_index_776078 == array_index_772828 ? add_776206 : sel_776203;
  assign add_776210 = sel_776207 + 8'h01;
  assign sel_776211 = array_index_776078 == array_index_772834 ? add_776210 : sel_776207;
  assign add_776214 = sel_776211 + 8'h01;
  assign sel_776215 = array_index_776078 == array_index_772840 ? add_776214 : sel_776211;
  assign add_776218 = sel_776215 + 8'h01;
  assign sel_776219 = array_index_776078 == array_index_772846 ? add_776218 : sel_776215;
  assign add_776222 = sel_776219 + 8'h01;
  assign sel_776223 = array_index_776078 == array_index_772852 ? add_776222 : sel_776219;
  assign add_776226 = sel_776223 + 8'h01;
  assign sel_776227 = array_index_776078 == array_index_772858 ? add_776226 : sel_776223;
  assign add_776230 = sel_776227 + 8'h01;
  assign sel_776231 = array_index_776078 == array_index_772864 ? add_776230 : sel_776227;
  assign add_776234 = sel_776231 + 8'h01;
  assign sel_776235 = array_index_776078 == array_index_772870 ? add_776234 : sel_776231;
  assign add_776238 = sel_776235 + 8'h01;
  assign sel_776239 = array_index_776078 == array_index_772876 ? add_776238 : sel_776235;
  assign add_776242 = sel_776239 + 8'h01;
  assign sel_776243 = array_index_776078 == array_index_772882 ? add_776242 : sel_776239;
  assign add_776246 = sel_776243 + 8'h01;
  assign sel_776247 = array_index_776078 == array_index_772888 ? add_776246 : sel_776243;
  assign add_776250 = sel_776247 + 8'h01;
  assign sel_776251 = array_index_776078 == array_index_772894 ? add_776250 : sel_776247;
  assign add_776254 = sel_776251 + 8'h01;
  assign sel_776255 = array_index_776078 == array_index_772900 ? add_776254 : sel_776251;
  assign add_776258 = sel_776255 + 8'h01;
  assign sel_776259 = array_index_776078 == array_index_772906 ? add_776258 : sel_776255;
  assign add_776262 = sel_776259 + 8'h01;
  assign sel_776263 = array_index_776078 == array_index_772912 ? add_776262 : sel_776259;
  assign add_776266 = sel_776263 + 8'h01;
  assign sel_776267 = array_index_776078 == array_index_772918 ? add_776266 : sel_776263;
  assign add_776270 = sel_776267 + 8'h01;
  assign sel_776271 = array_index_776078 == array_index_772924 ? add_776270 : sel_776267;
  assign add_776274 = sel_776271 + 8'h01;
  assign sel_776275 = array_index_776078 == array_index_772930 ? add_776274 : sel_776271;
  assign add_776278 = sel_776275 + 8'h01;
  assign sel_776279 = array_index_776078 == array_index_772936 ? add_776278 : sel_776275;
  assign add_776282 = sel_776279 + 8'h01;
  assign sel_776283 = array_index_776078 == array_index_772942 ? add_776282 : sel_776279;
  assign add_776286 = sel_776283 + 8'h01;
  assign sel_776287 = array_index_776078 == array_index_772948 ? add_776286 : sel_776283;
  assign add_776290 = sel_776287 + 8'h01;
  assign sel_776291 = array_index_776078 == array_index_772954 ? add_776290 : sel_776287;
  assign add_776294 = sel_776291 + 8'h01;
  assign sel_776295 = array_index_776078 == array_index_772960 ? add_776294 : sel_776291;
  assign add_776298 = sel_776295 + 8'h01;
  assign sel_776299 = array_index_776078 == array_index_772966 ? add_776298 : sel_776295;
  assign add_776302 = sel_776299 + 8'h01;
  assign sel_776303 = array_index_776078 == array_index_772972 ? add_776302 : sel_776299;
  assign add_776306 = sel_776303 + 8'h01;
  assign sel_776307 = array_index_776078 == array_index_772978 ? add_776306 : sel_776303;
  assign add_776310 = sel_776307 + 8'h01;
  assign sel_776311 = array_index_776078 == array_index_772984 ? add_776310 : sel_776307;
  assign add_776314 = sel_776311 + 8'h01;
  assign sel_776315 = array_index_776078 == array_index_772990 ? add_776314 : sel_776311;
  assign add_776318 = sel_776315 + 8'h01;
  assign sel_776319 = array_index_776078 == array_index_772996 ? add_776318 : sel_776315;
  assign add_776322 = sel_776319 + 8'h01;
  assign sel_776323 = array_index_776078 == array_index_773002 ? add_776322 : sel_776319;
  assign add_776326 = sel_776323 + 8'h01;
  assign sel_776327 = array_index_776078 == array_index_773008 ? add_776326 : sel_776323;
  assign add_776330 = sel_776327 + 8'h01;
  assign sel_776331 = array_index_776078 == array_index_773014 ? add_776330 : sel_776327;
  assign add_776334 = sel_776331 + 8'h01;
  assign sel_776335 = array_index_776078 == array_index_773020 ? add_776334 : sel_776331;
  assign add_776338 = sel_776335 + 8'h01;
  assign sel_776339 = array_index_776078 == array_index_773026 ? add_776338 : sel_776335;
  assign add_776342 = sel_776339 + 8'h01;
  assign sel_776343 = array_index_776078 == array_index_773032 ? add_776342 : sel_776339;
  assign add_776346 = sel_776343 + 8'h01;
  assign sel_776347 = array_index_776078 == array_index_773038 ? add_776346 : sel_776343;
  assign add_776350 = sel_776347 + 8'h01;
  assign sel_776351 = array_index_776078 == array_index_773044 ? add_776350 : sel_776347;
  assign add_776354 = sel_776351 + 8'h01;
  assign sel_776355 = array_index_776078 == array_index_773050 ? add_776354 : sel_776351;
  assign add_776358 = sel_776355 + 8'h01;
  assign sel_776359 = array_index_776078 == array_index_773056 ? add_776358 : sel_776355;
  assign add_776362 = sel_776359 + 8'h01;
  assign sel_776363 = array_index_776078 == array_index_773062 ? add_776362 : sel_776359;
  assign add_776366 = sel_776363 + 8'h01;
  assign sel_776367 = array_index_776078 == array_index_773068 ? add_776366 : sel_776363;
  assign add_776370 = sel_776367 + 8'h01;
  assign sel_776371 = array_index_776078 == array_index_773074 ? add_776370 : sel_776367;
  assign add_776374 = sel_776371 + 8'h01;
  assign sel_776375 = array_index_776078 == array_index_773080 ? add_776374 : sel_776371;
  assign add_776378 = sel_776375 + 8'h01;
  assign sel_776379 = array_index_776078 == array_index_773086 ? add_776378 : sel_776375;
  assign add_776382 = sel_776379 + 8'h01;
  assign sel_776383 = array_index_776078 == array_index_773092 ? add_776382 : sel_776379;
  assign add_776386 = sel_776383 + 8'h01;
  assign sel_776387 = array_index_776078 == array_index_773098 ? add_776386 : sel_776383;
  assign add_776390 = sel_776387 + 8'h01;
  assign sel_776391 = array_index_776078 == array_index_773104 ? add_776390 : sel_776387;
  assign add_776394 = sel_776391 + 8'h01;
  assign sel_776395 = array_index_776078 == array_index_773110 ? add_776394 : sel_776391;
  assign add_776398 = sel_776395 + 8'h01;
  assign sel_776399 = array_index_776078 == array_index_773116 ? add_776398 : sel_776395;
  assign add_776402 = sel_776399 + 8'h01;
  assign sel_776403 = array_index_776078 == array_index_773122 ? add_776402 : sel_776399;
  assign add_776406 = sel_776403 + 8'h01;
  assign sel_776407 = array_index_776078 == array_index_773128 ? add_776406 : sel_776403;
  assign add_776410 = sel_776407 + 8'h01;
  assign sel_776411 = array_index_776078 == array_index_773134 ? add_776410 : sel_776407;
  assign add_776414 = sel_776411 + 8'h01;
  assign sel_776415 = array_index_776078 == array_index_773140 ? add_776414 : sel_776411;
  assign add_776418 = sel_776415 + 8'h01;
  assign sel_776419 = array_index_776078 == array_index_773146 ? add_776418 : sel_776415;
  assign add_776422 = sel_776419 + 8'h01;
  assign sel_776423 = array_index_776078 == array_index_773152 ? add_776422 : sel_776419;
  assign add_776426 = sel_776423 + 8'h01;
  assign sel_776427 = array_index_776078 == array_index_773158 ? add_776426 : sel_776423;
  assign add_776430 = sel_776427 + 8'h01;
  assign sel_776431 = array_index_776078 == array_index_773164 ? add_776430 : sel_776427;
  assign add_776434 = sel_776431 + 8'h01;
  assign sel_776435 = array_index_776078 == array_index_773170 ? add_776434 : sel_776431;
  assign add_776439 = sel_776435 + 8'h01;
  assign array_index_776440 = set1_unflattened[7'h0a];
  assign sel_776441 = array_index_776078 == array_index_773176 ? add_776439 : sel_776435;
  assign add_776444 = sel_776441 + 8'h01;
  assign sel_776445 = array_index_776440 == array_index_772632 ? add_776444 : sel_776441;
  assign add_776448 = sel_776445 + 8'h01;
  assign sel_776449 = array_index_776440 == array_index_772636 ? add_776448 : sel_776445;
  assign add_776452 = sel_776449 + 8'h01;
  assign sel_776453 = array_index_776440 == array_index_772644 ? add_776452 : sel_776449;
  assign add_776456 = sel_776453 + 8'h01;
  assign sel_776457 = array_index_776440 == array_index_772652 ? add_776456 : sel_776453;
  assign add_776460 = sel_776457 + 8'h01;
  assign sel_776461 = array_index_776440 == array_index_772660 ? add_776460 : sel_776457;
  assign add_776464 = sel_776461 + 8'h01;
  assign sel_776465 = array_index_776440 == array_index_772668 ? add_776464 : sel_776461;
  assign add_776468 = sel_776465 + 8'h01;
  assign sel_776469 = array_index_776440 == array_index_772676 ? add_776468 : sel_776465;
  assign add_776472 = sel_776469 + 8'h01;
  assign sel_776473 = array_index_776440 == array_index_772684 ? add_776472 : sel_776469;
  assign add_776476 = sel_776473 + 8'h01;
  assign sel_776477 = array_index_776440 == array_index_772690 ? add_776476 : sel_776473;
  assign add_776480 = sel_776477 + 8'h01;
  assign sel_776481 = array_index_776440 == array_index_772696 ? add_776480 : sel_776477;
  assign add_776484 = sel_776481 + 8'h01;
  assign sel_776485 = array_index_776440 == array_index_772702 ? add_776484 : sel_776481;
  assign add_776488 = sel_776485 + 8'h01;
  assign sel_776489 = array_index_776440 == array_index_772708 ? add_776488 : sel_776485;
  assign add_776492 = sel_776489 + 8'h01;
  assign sel_776493 = array_index_776440 == array_index_772714 ? add_776492 : sel_776489;
  assign add_776496 = sel_776493 + 8'h01;
  assign sel_776497 = array_index_776440 == array_index_772720 ? add_776496 : sel_776493;
  assign add_776500 = sel_776497 + 8'h01;
  assign sel_776501 = array_index_776440 == array_index_772726 ? add_776500 : sel_776497;
  assign add_776504 = sel_776501 + 8'h01;
  assign sel_776505 = array_index_776440 == array_index_772732 ? add_776504 : sel_776501;
  assign add_776508 = sel_776505 + 8'h01;
  assign sel_776509 = array_index_776440 == array_index_772738 ? add_776508 : sel_776505;
  assign add_776512 = sel_776509 + 8'h01;
  assign sel_776513 = array_index_776440 == array_index_772744 ? add_776512 : sel_776509;
  assign add_776516 = sel_776513 + 8'h01;
  assign sel_776517 = array_index_776440 == array_index_772750 ? add_776516 : sel_776513;
  assign add_776520 = sel_776517 + 8'h01;
  assign sel_776521 = array_index_776440 == array_index_772756 ? add_776520 : sel_776517;
  assign add_776524 = sel_776521 + 8'h01;
  assign sel_776525 = array_index_776440 == array_index_772762 ? add_776524 : sel_776521;
  assign add_776528 = sel_776525 + 8'h01;
  assign sel_776529 = array_index_776440 == array_index_772768 ? add_776528 : sel_776525;
  assign add_776532 = sel_776529 + 8'h01;
  assign sel_776533 = array_index_776440 == array_index_772774 ? add_776532 : sel_776529;
  assign add_776536 = sel_776533 + 8'h01;
  assign sel_776537 = array_index_776440 == array_index_772780 ? add_776536 : sel_776533;
  assign add_776540 = sel_776537 + 8'h01;
  assign sel_776541 = array_index_776440 == array_index_772786 ? add_776540 : sel_776537;
  assign add_776544 = sel_776541 + 8'h01;
  assign sel_776545 = array_index_776440 == array_index_772792 ? add_776544 : sel_776541;
  assign add_776548 = sel_776545 + 8'h01;
  assign sel_776549 = array_index_776440 == array_index_772798 ? add_776548 : sel_776545;
  assign add_776552 = sel_776549 + 8'h01;
  assign sel_776553 = array_index_776440 == array_index_772804 ? add_776552 : sel_776549;
  assign add_776556 = sel_776553 + 8'h01;
  assign sel_776557 = array_index_776440 == array_index_772810 ? add_776556 : sel_776553;
  assign add_776560 = sel_776557 + 8'h01;
  assign sel_776561 = array_index_776440 == array_index_772816 ? add_776560 : sel_776557;
  assign add_776564 = sel_776561 + 8'h01;
  assign sel_776565 = array_index_776440 == array_index_772822 ? add_776564 : sel_776561;
  assign add_776568 = sel_776565 + 8'h01;
  assign sel_776569 = array_index_776440 == array_index_772828 ? add_776568 : sel_776565;
  assign add_776572 = sel_776569 + 8'h01;
  assign sel_776573 = array_index_776440 == array_index_772834 ? add_776572 : sel_776569;
  assign add_776576 = sel_776573 + 8'h01;
  assign sel_776577 = array_index_776440 == array_index_772840 ? add_776576 : sel_776573;
  assign add_776580 = sel_776577 + 8'h01;
  assign sel_776581 = array_index_776440 == array_index_772846 ? add_776580 : sel_776577;
  assign add_776584 = sel_776581 + 8'h01;
  assign sel_776585 = array_index_776440 == array_index_772852 ? add_776584 : sel_776581;
  assign add_776588 = sel_776585 + 8'h01;
  assign sel_776589 = array_index_776440 == array_index_772858 ? add_776588 : sel_776585;
  assign add_776592 = sel_776589 + 8'h01;
  assign sel_776593 = array_index_776440 == array_index_772864 ? add_776592 : sel_776589;
  assign add_776596 = sel_776593 + 8'h01;
  assign sel_776597 = array_index_776440 == array_index_772870 ? add_776596 : sel_776593;
  assign add_776600 = sel_776597 + 8'h01;
  assign sel_776601 = array_index_776440 == array_index_772876 ? add_776600 : sel_776597;
  assign add_776604 = sel_776601 + 8'h01;
  assign sel_776605 = array_index_776440 == array_index_772882 ? add_776604 : sel_776601;
  assign add_776608 = sel_776605 + 8'h01;
  assign sel_776609 = array_index_776440 == array_index_772888 ? add_776608 : sel_776605;
  assign add_776612 = sel_776609 + 8'h01;
  assign sel_776613 = array_index_776440 == array_index_772894 ? add_776612 : sel_776609;
  assign add_776616 = sel_776613 + 8'h01;
  assign sel_776617 = array_index_776440 == array_index_772900 ? add_776616 : sel_776613;
  assign add_776620 = sel_776617 + 8'h01;
  assign sel_776621 = array_index_776440 == array_index_772906 ? add_776620 : sel_776617;
  assign add_776624 = sel_776621 + 8'h01;
  assign sel_776625 = array_index_776440 == array_index_772912 ? add_776624 : sel_776621;
  assign add_776628 = sel_776625 + 8'h01;
  assign sel_776629 = array_index_776440 == array_index_772918 ? add_776628 : sel_776625;
  assign add_776632 = sel_776629 + 8'h01;
  assign sel_776633 = array_index_776440 == array_index_772924 ? add_776632 : sel_776629;
  assign add_776636 = sel_776633 + 8'h01;
  assign sel_776637 = array_index_776440 == array_index_772930 ? add_776636 : sel_776633;
  assign add_776640 = sel_776637 + 8'h01;
  assign sel_776641 = array_index_776440 == array_index_772936 ? add_776640 : sel_776637;
  assign add_776644 = sel_776641 + 8'h01;
  assign sel_776645 = array_index_776440 == array_index_772942 ? add_776644 : sel_776641;
  assign add_776648 = sel_776645 + 8'h01;
  assign sel_776649 = array_index_776440 == array_index_772948 ? add_776648 : sel_776645;
  assign add_776652 = sel_776649 + 8'h01;
  assign sel_776653 = array_index_776440 == array_index_772954 ? add_776652 : sel_776649;
  assign add_776656 = sel_776653 + 8'h01;
  assign sel_776657 = array_index_776440 == array_index_772960 ? add_776656 : sel_776653;
  assign add_776660 = sel_776657 + 8'h01;
  assign sel_776661 = array_index_776440 == array_index_772966 ? add_776660 : sel_776657;
  assign add_776664 = sel_776661 + 8'h01;
  assign sel_776665 = array_index_776440 == array_index_772972 ? add_776664 : sel_776661;
  assign add_776668 = sel_776665 + 8'h01;
  assign sel_776669 = array_index_776440 == array_index_772978 ? add_776668 : sel_776665;
  assign add_776672 = sel_776669 + 8'h01;
  assign sel_776673 = array_index_776440 == array_index_772984 ? add_776672 : sel_776669;
  assign add_776676 = sel_776673 + 8'h01;
  assign sel_776677 = array_index_776440 == array_index_772990 ? add_776676 : sel_776673;
  assign add_776680 = sel_776677 + 8'h01;
  assign sel_776681 = array_index_776440 == array_index_772996 ? add_776680 : sel_776677;
  assign add_776684 = sel_776681 + 8'h01;
  assign sel_776685 = array_index_776440 == array_index_773002 ? add_776684 : sel_776681;
  assign add_776688 = sel_776685 + 8'h01;
  assign sel_776689 = array_index_776440 == array_index_773008 ? add_776688 : sel_776685;
  assign add_776692 = sel_776689 + 8'h01;
  assign sel_776693 = array_index_776440 == array_index_773014 ? add_776692 : sel_776689;
  assign add_776696 = sel_776693 + 8'h01;
  assign sel_776697 = array_index_776440 == array_index_773020 ? add_776696 : sel_776693;
  assign add_776700 = sel_776697 + 8'h01;
  assign sel_776701 = array_index_776440 == array_index_773026 ? add_776700 : sel_776697;
  assign add_776704 = sel_776701 + 8'h01;
  assign sel_776705 = array_index_776440 == array_index_773032 ? add_776704 : sel_776701;
  assign add_776708 = sel_776705 + 8'h01;
  assign sel_776709 = array_index_776440 == array_index_773038 ? add_776708 : sel_776705;
  assign add_776712 = sel_776709 + 8'h01;
  assign sel_776713 = array_index_776440 == array_index_773044 ? add_776712 : sel_776709;
  assign add_776716 = sel_776713 + 8'h01;
  assign sel_776717 = array_index_776440 == array_index_773050 ? add_776716 : sel_776713;
  assign add_776720 = sel_776717 + 8'h01;
  assign sel_776721 = array_index_776440 == array_index_773056 ? add_776720 : sel_776717;
  assign add_776724 = sel_776721 + 8'h01;
  assign sel_776725 = array_index_776440 == array_index_773062 ? add_776724 : sel_776721;
  assign add_776728 = sel_776725 + 8'h01;
  assign sel_776729 = array_index_776440 == array_index_773068 ? add_776728 : sel_776725;
  assign add_776732 = sel_776729 + 8'h01;
  assign sel_776733 = array_index_776440 == array_index_773074 ? add_776732 : sel_776729;
  assign add_776736 = sel_776733 + 8'h01;
  assign sel_776737 = array_index_776440 == array_index_773080 ? add_776736 : sel_776733;
  assign add_776740 = sel_776737 + 8'h01;
  assign sel_776741 = array_index_776440 == array_index_773086 ? add_776740 : sel_776737;
  assign add_776744 = sel_776741 + 8'h01;
  assign sel_776745 = array_index_776440 == array_index_773092 ? add_776744 : sel_776741;
  assign add_776748 = sel_776745 + 8'h01;
  assign sel_776749 = array_index_776440 == array_index_773098 ? add_776748 : sel_776745;
  assign add_776752 = sel_776749 + 8'h01;
  assign sel_776753 = array_index_776440 == array_index_773104 ? add_776752 : sel_776749;
  assign add_776756 = sel_776753 + 8'h01;
  assign sel_776757 = array_index_776440 == array_index_773110 ? add_776756 : sel_776753;
  assign add_776760 = sel_776757 + 8'h01;
  assign sel_776761 = array_index_776440 == array_index_773116 ? add_776760 : sel_776757;
  assign add_776764 = sel_776761 + 8'h01;
  assign sel_776765 = array_index_776440 == array_index_773122 ? add_776764 : sel_776761;
  assign add_776768 = sel_776765 + 8'h01;
  assign sel_776769 = array_index_776440 == array_index_773128 ? add_776768 : sel_776765;
  assign add_776772 = sel_776769 + 8'h01;
  assign sel_776773 = array_index_776440 == array_index_773134 ? add_776772 : sel_776769;
  assign add_776776 = sel_776773 + 8'h01;
  assign sel_776777 = array_index_776440 == array_index_773140 ? add_776776 : sel_776773;
  assign add_776780 = sel_776777 + 8'h01;
  assign sel_776781 = array_index_776440 == array_index_773146 ? add_776780 : sel_776777;
  assign add_776784 = sel_776781 + 8'h01;
  assign sel_776785 = array_index_776440 == array_index_773152 ? add_776784 : sel_776781;
  assign add_776788 = sel_776785 + 8'h01;
  assign sel_776789 = array_index_776440 == array_index_773158 ? add_776788 : sel_776785;
  assign add_776792 = sel_776789 + 8'h01;
  assign sel_776793 = array_index_776440 == array_index_773164 ? add_776792 : sel_776789;
  assign add_776796 = sel_776793 + 8'h01;
  assign sel_776797 = array_index_776440 == array_index_773170 ? add_776796 : sel_776793;
  assign add_776801 = sel_776797 + 8'h01;
  assign array_index_776802 = set1_unflattened[7'h0b];
  assign sel_776803 = array_index_776440 == array_index_773176 ? add_776801 : sel_776797;
  assign add_776806 = sel_776803 + 8'h01;
  assign sel_776807 = array_index_776802 == array_index_772632 ? add_776806 : sel_776803;
  assign add_776810 = sel_776807 + 8'h01;
  assign sel_776811 = array_index_776802 == array_index_772636 ? add_776810 : sel_776807;
  assign add_776814 = sel_776811 + 8'h01;
  assign sel_776815 = array_index_776802 == array_index_772644 ? add_776814 : sel_776811;
  assign add_776818 = sel_776815 + 8'h01;
  assign sel_776819 = array_index_776802 == array_index_772652 ? add_776818 : sel_776815;
  assign add_776822 = sel_776819 + 8'h01;
  assign sel_776823 = array_index_776802 == array_index_772660 ? add_776822 : sel_776819;
  assign add_776826 = sel_776823 + 8'h01;
  assign sel_776827 = array_index_776802 == array_index_772668 ? add_776826 : sel_776823;
  assign add_776830 = sel_776827 + 8'h01;
  assign sel_776831 = array_index_776802 == array_index_772676 ? add_776830 : sel_776827;
  assign add_776834 = sel_776831 + 8'h01;
  assign sel_776835 = array_index_776802 == array_index_772684 ? add_776834 : sel_776831;
  assign add_776838 = sel_776835 + 8'h01;
  assign sel_776839 = array_index_776802 == array_index_772690 ? add_776838 : sel_776835;
  assign add_776842 = sel_776839 + 8'h01;
  assign sel_776843 = array_index_776802 == array_index_772696 ? add_776842 : sel_776839;
  assign add_776846 = sel_776843 + 8'h01;
  assign sel_776847 = array_index_776802 == array_index_772702 ? add_776846 : sel_776843;
  assign add_776850 = sel_776847 + 8'h01;
  assign sel_776851 = array_index_776802 == array_index_772708 ? add_776850 : sel_776847;
  assign add_776854 = sel_776851 + 8'h01;
  assign sel_776855 = array_index_776802 == array_index_772714 ? add_776854 : sel_776851;
  assign add_776858 = sel_776855 + 8'h01;
  assign sel_776859 = array_index_776802 == array_index_772720 ? add_776858 : sel_776855;
  assign add_776862 = sel_776859 + 8'h01;
  assign sel_776863 = array_index_776802 == array_index_772726 ? add_776862 : sel_776859;
  assign add_776866 = sel_776863 + 8'h01;
  assign sel_776867 = array_index_776802 == array_index_772732 ? add_776866 : sel_776863;
  assign add_776870 = sel_776867 + 8'h01;
  assign sel_776871 = array_index_776802 == array_index_772738 ? add_776870 : sel_776867;
  assign add_776874 = sel_776871 + 8'h01;
  assign sel_776875 = array_index_776802 == array_index_772744 ? add_776874 : sel_776871;
  assign add_776878 = sel_776875 + 8'h01;
  assign sel_776879 = array_index_776802 == array_index_772750 ? add_776878 : sel_776875;
  assign add_776882 = sel_776879 + 8'h01;
  assign sel_776883 = array_index_776802 == array_index_772756 ? add_776882 : sel_776879;
  assign add_776886 = sel_776883 + 8'h01;
  assign sel_776887 = array_index_776802 == array_index_772762 ? add_776886 : sel_776883;
  assign add_776890 = sel_776887 + 8'h01;
  assign sel_776891 = array_index_776802 == array_index_772768 ? add_776890 : sel_776887;
  assign add_776894 = sel_776891 + 8'h01;
  assign sel_776895 = array_index_776802 == array_index_772774 ? add_776894 : sel_776891;
  assign add_776898 = sel_776895 + 8'h01;
  assign sel_776899 = array_index_776802 == array_index_772780 ? add_776898 : sel_776895;
  assign add_776902 = sel_776899 + 8'h01;
  assign sel_776903 = array_index_776802 == array_index_772786 ? add_776902 : sel_776899;
  assign add_776906 = sel_776903 + 8'h01;
  assign sel_776907 = array_index_776802 == array_index_772792 ? add_776906 : sel_776903;
  assign add_776910 = sel_776907 + 8'h01;
  assign sel_776911 = array_index_776802 == array_index_772798 ? add_776910 : sel_776907;
  assign add_776914 = sel_776911 + 8'h01;
  assign sel_776915 = array_index_776802 == array_index_772804 ? add_776914 : sel_776911;
  assign add_776918 = sel_776915 + 8'h01;
  assign sel_776919 = array_index_776802 == array_index_772810 ? add_776918 : sel_776915;
  assign add_776922 = sel_776919 + 8'h01;
  assign sel_776923 = array_index_776802 == array_index_772816 ? add_776922 : sel_776919;
  assign add_776926 = sel_776923 + 8'h01;
  assign sel_776927 = array_index_776802 == array_index_772822 ? add_776926 : sel_776923;
  assign add_776930 = sel_776927 + 8'h01;
  assign sel_776931 = array_index_776802 == array_index_772828 ? add_776930 : sel_776927;
  assign add_776934 = sel_776931 + 8'h01;
  assign sel_776935 = array_index_776802 == array_index_772834 ? add_776934 : sel_776931;
  assign add_776938 = sel_776935 + 8'h01;
  assign sel_776939 = array_index_776802 == array_index_772840 ? add_776938 : sel_776935;
  assign add_776942 = sel_776939 + 8'h01;
  assign sel_776943 = array_index_776802 == array_index_772846 ? add_776942 : sel_776939;
  assign add_776946 = sel_776943 + 8'h01;
  assign sel_776947 = array_index_776802 == array_index_772852 ? add_776946 : sel_776943;
  assign add_776950 = sel_776947 + 8'h01;
  assign sel_776951 = array_index_776802 == array_index_772858 ? add_776950 : sel_776947;
  assign add_776954 = sel_776951 + 8'h01;
  assign sel_776955 = array_index_776802 == array_index_772864 ? add_776954 : sel_776951;
  assign add_776958 = sel_776955 + 8'h01;
  assign sel_776959 = array_index_776802 == array_index_772870 ? add_776958 : sel_776955;
  assign add_776962 = sel_776959 + 8'h01;
  assign sel_776963 = array_index_776802 == array_index_772876 ? add_776962 : sel_776959;
  assign add_776966 = sel_776963 + 8'h01;
  assign sel_776967 = array_index_776802 == array_index_772882 ? add_776966 : sel_776963;
  assign add_776970 = sel_776967 + 8'h01;
  assign sel_776971 = array_index_776802 == array_index_772888 ? add_776970 : sel_776967;
  assign add_776974 = sel_776971 + 8'h01;
  assign sel_776975 = array_index_776802 == array_index_772894 ? add_776974 : sel_776971;
  assign add_776978 = sel_776975 + 8'h01;
  assign sel_776979 = array_index_776802 == array_index_772900 ? add_776978 : sel_776975;
  assign add_776982 = sel_776979 + 8'h01;
  assign sel_776983 = array_index_776802 == array_index_772906 ? add_776982 : sel_776979;
  assign add_776986 = sel_776983 + 8'h01;
  assign sel_776987 = array_index_776802 == array_index_772912 ? add_776986 : sel_776983;
  assign add_776990 = sel_776987 + 8'h01;
  assign sel_776991 = array_index_776802 == array_index_772918 ? add_776990 : sel_776987;
  assign add_776994 = sel_776991 + 8'h01;
  assign sel_776995 = array_index_776802 == array_index_772924 ? add_776994 : sel_776991;
  assign add_776998 = sel_776995 + 8'h01;
  assign sel_776999 = array_index_776802 == array_index_772930 ? add_776998 : sel_776995;
  assign add_777002 = sel_776999 + 8'h01;
  assign sel_777003 = array_index_776802 == array_index_772936 ? add_777002 : sel_776999;
  assign add_777006 = sel_777003 + 8'h01;
  assign sel_777007 = array_index_776802 == array_index_772942 ? add_777006 : sel_777003;
  assign add_777010 = sel_777007 + 8'h01;
  assign sel_777011 = array_index_776802 == array_index_772948 ? add_777010 : sel_777007;
  assign add_777014 = sel_777011 + 8'h01;
  assign sel_777015 = array_index_776802 == array_index_772954 ? add_777014 : sel_777011;
  assign add_777018 = sel_777015 + 8'h01;
  assign sel_777019 = array_index_776802 == array_index_772960 ? add_777018 : sel_777015;
  assign add_777022 = sel_777019 + 8'h01;
  assign sel_777023 = array_index_776802 == array_index_772966 ? add_777022 : sel_777019;
  assign add_777026 = sel_777023 + 8'h01;
  assign sel_777027 = array_index_776802 == array_index_772972 ? add_777026 : sel_777023;
  assign add_777030 = sel_777027 + 8'h01;
  assign sel_777031 = array_index_776802 == array_index_772978 ? add_777030 : sel_777027;
  assign add_777034 = sel_777031 + 8'h01;
  assign sel_777035 = array_index_776802 == array_index_772984 ? add_777034 : sel_777031;
  assign add_777038 = sel_777035 + 8'h01;
  assign sel_777039 = array_index_776802 == array_index_772990 ? add_777038 : sel_777035;
  assign add_777042 = sel_777039 + 8'h01;
  assign sel_777043 = array_index_776802 == array_index_772996 ? add_777042 : sel_777039;
  assign add_777046 = sel_777043 + 8'h01;
  assign sel_777047 = array_index_776802 == array_index_773002 ? add_777046 : sel_777043;
  assign add_777050 = sel_777047 + 8'h01;
  assign sel_777051 = array_index_776802 == array_index_773008 ? add_777050 : sel_777047;
  assign add_777054 = sel_777051 + 8'h01;
  assign sel_777055 = array_index_776802 == array_index_773014 ? add_777054 : sel_777051;
  assign add_777058 = sel_777055 + 8'h01;
  assign sel_777059 = array_index_776802 == array_index_773020 ? add_777058 : sel_777055;
  assign add_777062 = sel_777059 + 8'h01;
  assign sel_777063 = array_index_776802 == array_index_773026 ? add_777062 : sel_777059;
  assign add_777066 = sel_777063 + 8'h01;
  assign sel_777067 = array_index_776802 == array_index_773032 ? add_777066 : sel_777063;
  assign add_777070 = sel_777067 + 8'h01;
  assign sel_777071 = array_index_776802 == array_index_773038 ? add_777070 : sel_777067;
  assign add_777074 = sel_777071 + 8'h01;
  assign sel_777075 = array_index_776802 == array_index_773044 ? add_777074 : sel_777071;
  assign add_777078 = sel_777075 + 8'h01;
  assign sel_777079 = array_index_776802 == array_index_773050 ? add_777078 : sel_777075;
  assign add_777082 = sel_777079 + 8'h01;
  assign sel_777083 = array_index_776802 == array_index_773056 ? add_777082 : sel_777079;
  assign add_777086 = sel_777083 + 8'h01;
  assign sel_777087 = array_index_776802 == array_index_773062 ? add_777086 : sel_777083;
  assign add_777090 = sel_777087 + 8'h01;
  assign sel_777091 = array_index_776802 == array_index_773068 ? add_777090 : sel_777087;
  assign add_777094 = sel_777091 + 8'h01;
  assign sel_777095 = array_index_776802 == array_index_773074 ? add_777094 : sel_777091;
  assign add_777098 = sel_777095 + 8'h01;
  assign sel_777099 = array_index_776802 == array_index_773080 ? add_777098 : sel_777095;
  assign add_777102 = sel_777099 + 8'h01;
  assign sel_777103 = array_index_776802 == array_index_773086 ? add_777102 : sel_777099;
  assign add_777106 = sel_777103 + 8'h01;
  assign sel_777107 = array_index_776802 == array_index_773092 ? add_777106 : sel_777103;
  assign add_777110 = sel_777107 + 8'h01;
  assign sel_777111 = array_index_776802 == array_index_773098 ? add_777110 : sel_777107;
  assign add_777114 = sel_777111 + 8'h01;
  assign sel_777115 = array_index_776802 == array_index_773104 ? add_777114 : sel_777111;
  assign add_777118 = sel_777115 + 8'h01;
  assign sel_777119 = array_index_776802 == array_index_773110 ? add_777118 : sel_777115;
  assign add_777122 = sel_777119 + 8'h01;
  assign sel_777123 = array_index_776802 == array_index_773116 ? add_777122 : sel_777119;
  assign add_777126 = sel_777123 + 8'h01;
  assign sel_777127 = array_index_776802 == array_index_773122 ? add_777126 : sel_777123;
  assign add_777130 = sel_777127 + 8'h01;
  assign sel_777131 = array_index_776802 == array_index_773128 ? add_777130 : sel_777127;
  assign add_777134 = sel_777131 + 8'h01;
  assign sel_777135 = array_index_776802 == array_index_773134 ? add_777134 : sel_777131;
  assign add_777138 = sel_777135 + 8'h01;
  assign sel_777139 = array_index_776802 == array_index_773140 ? add_777138 : sel_777135;
  assign add_777142 = sel_777139 + 8'h01;
  assign sel_777143 = array_index_776802 == array_index_773146 ? add_777142 : sel_777139;
  assign add_777146 = sel_777143 + 8'h01;
  assign sel_777147 = array_index_776802 == array_index_773152 ? add_777146 : sel_777143;
  assign add_777150 = sel_777147 + 8'h01;
  assign sel_777151 = array_index_776802 == array_index_773158 ? add_777150 : sel_777147;
  assign add_777154 = sel_777151 + 8'h01;
  assign sel_777155 = array_index_776802 == array_index_773164 ? add_777154 : sel_777151;
  assign add_777158 = sel_777155 + 8'h01;
  assign sel_777159 = array_index_776802 == array_index_773170 ? add_777158 : sel_777155;
  assign add_777163 = sel_777159 + 8'h01;
  assign array_index_777164 = set1_unflattened[7'h0c];
  assign sel_777165 = array_index_776802 == array_index_773176 ? add_777163 : sel_777159;
  assign add_777168 = sel_777165 + 8'h01;
  assign sel_777169 = array_index_777164 == array_index_772632 ? add_777168 : sel_777165;
  assign add_777172 = sel_777169 + 8'h01;
  assign sel_777173 = array_index_777164 == array_index_772636 ? add_777172 : sel_777169;
  assign add_777176 = sel_777173 + 8'h01;
  assign sel_777177 = array_index_777164 == array_index_772644 ? add_777176 : sel_777173;
  assign add_777180 = sel_777177 + 8'h01;
  assign sel_777181 = array_index_777164 == array_index_772652 ? add_777180 : sel_777177;
  assign add_777184 = sel_777181 + 8'h01;
  assign sel_777185 = array_index_777164 == array_index_772660 ? add_777184 : sel_777181;
  assign add_777188 = sel_777185 + 8'h01;
  assign sel_777189 = array_index_777164 == array_index_772668 ? add_777188 : sel_777185;
  assign add_777192 = sel_777189 + 8'h01;
  assign sel_777193 = array_index_777164 == array_index_772676 ? add_777192 : sel_777189;
  assign add_777196 = sel_777193 + 8'h01;
  assign sel_777197 = array_index_777164 == array_index_772684 ? add_777196 : sel_777193;
  assign add_777200 = sel_777197 + 8'h01;
  assign sel_777201 = array_index_777164 == array_index_772690 ? add_777200 : sel_777197;
  assign add_777204 = sel_777201 + 8'h01;
  assign sel_777205 = array_index_777164 == array_index_772696 ? add_777204 : sel_777201;
  assign add_777208 = sel_777205 + 8'h01;
  assign sel_777209 = array_index_777164 == array_index_772702 ? add_777208 : sel_777205;
  assign add_777212 = sel_777209 + 8'h01;
  assign sel_777213 = array_index_777164 == array_index_772708 ? add_777212 : sel_777209;
  assign add_777216 = sel_777213 + 8'h01;
  assign sel_777217 = array_index_777164 == array_index_772714 ? add_777216 : sel_777213;
  assign add_777220 = sel_777217 + 8'h01;
  assign sel_777221 = array_index_777164 == array_index_772720 ? add_777220 : sel_777217;
  assign add_777224 = sel_777221 + 8'h01;
  assign sel_777225 = array_index_777164 == array_index_772726 ? add_777224 : sel_777221;
  assign add_777228 = sel_777225 + 8'h01;
  assign sel_777229 = array_index_777164 == array_index_772732 ? add_777228 : sel_777225;
  assign add_777232 = sel_777229 + 8'h01;
  assign sel_777233 = array_index_777164 == array_index_772738 ? add_777232 : sel_777229;
  assign add_777236 = sel_777233 + 8'h01;
  assign sel_777237 = array_index_777164 == array_index_772744 ? add_777236 : sel_777233;
  assign add_777240 = sel_777237 + 8'h01;
  assign sel_777241 = array_index_777164 == array_index_772750 ? add_777240 : sel_777237;
  assign add_777244 = sel_777241 + 8'h01;
  assign sel_777245 = array_index_777164 == array_index_772756 ? add_777244 : sel_777241;
  assign add_777248 = sel_777245 + 8'h01;
  assign sel_777249 = array_index_777164 == array_index_772762 ? add_777248 : sel_777245;
  assign add_777252 = sel_777249 + 8'h01;
  assign sel_777253 = array_index_777164 == array_index_772768 ? add_777252 : sel_777249;
  assign add_777256 = sel_777253 + 8'h01;
  assign sel_777257 = array_index_777164 == array_index_772774 ? add_777256 : sel_777253;
  assign add_777260 = sel_777257 + 8'h01;
  assign sel_777261 = array_index_777164 == array_index_772780 ? add_777260 : sel_777257;
  assign add_777264 = sel_777261 + 8'h01;
  assign sel_777265 = array_index_777164 == array_index_772786 ? add_777264 : sel_777261;
  assign add_777268 = sel_777265 + 8'h01;
  assign sel_777269 = array_index_777164 == array_index_772792 ? add_777268 : sel_777265;
  assign add_777272 = sel_777269 + 8'h01;
  assign sel_777273 = array_index_777164 == array_index_772798 ? add_777272 : sel_777269;
  assign add_777276 = sel_777273 + 8'h01;
  assign sel_777277 = array_index_777164 == array_index_772804 ? add_777276 : sel_777273;
  assign add_777280 = sel_777277 + 8'h01;
  assign sel_777281 = array_index_777164 == array_index_772810 ? add_777280 : sel_777277;
  assign add_777284 = sel_777281 + 8'h01;
  assign sel_777285 = array_index_777164 == array_index_772816 ? add_777284 : sel_777281;
  assign add_777288 = sel_777285 + 8'h01;
  assign sel_777289 = array_index_777164 == array_index_772822 ? add_777288 : sel_777285;
  assign add_777292 = sel_777289 + 8'h01;
  assign sel_777293 = array_index_777164 == array_index_772828 ? add_777292 : sel_777289;
  assign add_777296 = sel_777293 + 8'h01;
  assign sel_777297 = array_index_777164 == array_index_772834 ? add_777296 : sel_777293;
  assign add_777300 = sel_777297 + 8'h01;
  assign sel_777301 = array_index_777164 == array_index_772840 ? add_777300 : sel_777297;
  assign add_777304 = sel_777301 + 8'h01;
  assign sel_777305 = array_index_777164 == array_index_772846 ? add_777304 : sel_777301;
  assign add_777308 = sel_777305 + 8'h01;
  assign sel_777309 = array_index_777164 == array_index_772852 ? add_777308 : sel_777305;
  assign add_777312 = sel_777309 + 8'h01;
  assign sel_777313 = array_index_777164 == array_index_772858 ? add_777312 : sel_777309;
  assign add_777316 = sel_777313 + 8'h01;
  assign sel_777317 = array_index_777164 == array_index_772864 ? add_777316 : sel_777313;
  assign add_777320 = sel_777317 + 8'h01;
  assign sel_777321 = array_index_777164 == array_index_772870 ? add_777320 : sel_777317;
  assign add_777324 = sel_777321 + 8'h01;
  assign sel_777325 = array_index_777164 == array_index_772876 ? add_777324 : sel_777321;
  assign add_777328 = sel_777325 + 8'h01;
  assign sel_777329 = array_index_777164 == array_index_772882 ? add_777328 : sel_777325;
  assign add_777332 = sel_777329 + 8'h01;
  assign sel_777333 = array_index_777164 == array_index_772888 ? add_777332 : sel_777329;
  assign add_777336 = sel_777333 + 8'h01;
  assign sel_777337 = array_index_777164 == array_index_772894 ? add_777336 : sel_777333;
  assign add_777340 = sel_777337 + 8'h01;
  assign sel_777341 = array_index_777164 == array_index_772900 ? add_777340 : sel_777337;
  assign add_777344 = sel_777341 + 8'h01;
  assign sel_777345 = array_index_777164 == array_index_772906 ? add_777344 : sel_777341;
  assign add_777348 = sel_777345 + 8'h01;
  assign sel_777349 = array_index_777164 == array_index_772912 ? add_777348 : sel_777345;
  assign add_777352 = sel_777349 + 8'h01;
  assign sel_777353 = array_index_777164 == array_index_772918 ? add_777352 : sel_777349;
  assign add_777356 = sel_777353 + 8'h01;
  assign sel_777357 = array_index_777164 == array_index_772924 ? add_777356 : sel_777353;
  assign add_777360 = sel_777357 + 8'h01;
  assign sel_777361 = array_index_777164 == array_index_772930 ? add_777360 : sel_777357;
  assign add_777364 = sel_777361 + 8'h01;
  assign sel_777365 = array_index_777164 == array_index_772936 ? add_777364 : sel_777361;
  assign add_777368 = sel_777365 + 8'h01;
  assign sel_777369 = array_index_777164 == array_index_772942 ? add_777368 : sel_777365;
  assign add_777372 = sel_777369 + 8'h01;
  assign sel_777373 = array_index_777164 == array_index_772948 ? add_777372 : sel_777369;
  assign add_777376 = sel_777373 + 8'h01;
  assign sel_777377 = array_index_777164 == array_index_772954 ? add_777376 : sel_777373;
  assign add_777380 = sel_777377 + 8'h01;
  assign sel_777381 = array_index_777164 == array_index_772960 ? add_777380 : sel_777377;
  assign add_777384 = sel_777381 + 8'h01;
  assign sel_777385 = array_index_777164 == array_index_772966 ? add_777384 : sel_777381;
  assign add_777388 = sel_777385 + 8'h01;
  assign sel_777389 = array_index_777164 == array_index_772972 ? add_777388 : sel_777385;
  assign add_777392 = sel_777389 + 8'h01;
  assign sel_777393 = array_index_777164 == array_index_772978 ? add_777392 : sel_777389;
  assign add_777396 = sel_777393 + 8'h01;
  assign sel_777397 = array_index_777164 == array_index_772984 ? add_777396 : sel_777393;
  assign add_777400 = sel_777397 + 8'h01;
  assign sel_777401 = array_index_777164 == array_index_772990 ? add_777400 : sel_777397;
  assign add_777404 = sel_777401 + 8'h01;
  assign sel_777405 = array_index_777164 == array_index_772996 ? add_777404 : sel_777401;
  assign add_777408 = sel_777405 + 8'h01;
  assign sel_777409 = array_index_777164 == array_index_773002 ? add_777408 : sel_777405;
  assign add_777412 = sel_777409 + 8'h01;
  assign sel_777413 = array_index_777164 == array_index_773008 ? add_777412 : sel_777409;
  assign add_777416 = sel_777413 + 8'h01;
  assign sel_777417 = array_index_777164 == array_index_773014 ? add_777416 : sel_777413;
  assign add_777420 = sel_777417 + 8'h01;
  assign sel_777421 = array_index_777164 == array_index_773020 ? add_777420 : sel_777417;
  assign add_777424 = sel_777421 + 8'h01;
  assign sel_777425 = array_index_777164 == array_index_773026 ? add_777424 : sel_777421;
  assign add_777428 = sel_777425 + 8'h01;
  assign sel_777429 = array_index_777164 == array_index_773032 ? add_777428 : sel_777425;
  assign add_777432 = sel_777429 + 8'h01;
  assign sel_777433 = array_index_777164 == array_index_773038 ? add_777432 : sel_777429;
  assign add_777436 = sel_777433 + 8'h01;
  assign sel_777437 = array_index_777164 == array_index_773044 ? add_777436 : sel_777433;
  assign add_777440 = sel_777437 + 8'h01;
  assign sel_777441 = array_index_777164 == array_index_773050 ? add_777440 : sel_777437;
  assign add_777444 = sel_777441 + 8'h01;
  assign sel_777445 = array_index_777164 == array_index_773056 ? add_777444 : sel_777441;
  assign add_777448 = sel_777445 + 8'h01;
  assign sel_777449 = array_index_777164 == array_index_773062 ? add_777448 : sel_777445;
  assign add_777452 = sel_777449 + 8'h01;
  assign sel_777453 = array_index_777164 == array_index_773068 ? add_777452 : sel_777449;
  assign add_777456 = sel_777453 + 8'h01;
  assign sel_777457 = array_index_777164 == array_index_773074 ? add_777456 : sel_777453;
  assign add_777460 = sel_777457 + 8'h01;
  assign sel_777461 = array_index_777164 == array_index_773080 ? add_777460 : sel_777457;
  assign add_777464 = sel_777461 + 8'h01;
  assign sel_777465 = array_index_777164 == array_index_773086 ? add_777464 : sel_777461;
  assign add_777468 = sel_777465 + 8'h01;
  assign sel_777469 = array_index_777164 == array_index_773092 ? add_777468 : sel_777465;
  assign add_777472 = sel_777469 + 8'h01;
  assign sel_777473 = array_index_777164 == array_index_773098 ? add_777472 : sel_777469;
  assign add_777476 = sel_777473 + 8'h01;
  assign sel_777477 = array_index_777164 == array_index_773104 ? add_777476 : sel_777473;
  assign add_777480 = sel_777477 + 8'h01;
  assign sel_777481 = array_index_777164 == array_index_773110 ? add_777480 : sel_777477;
  assign add_777484 = sel_777481 + 8'h01;
  assign sel_777485 = array_index_777164 == array_index_773116 ? add_777484 : sel_777481;
  assign add_777488 = sel_777485 + 8'h01;
  assign sel_777489 = array_index_777164 == array_index_773122 ? add_777488 : sel_777485;
  assign add_777492 = sel_777489 + 8'h01;
  assign sel_777493 = array_index_777164 == array_index_773128 ? add_777492 : sel_777489;
  assign add_777496 = sel_777493 + 8'h01;
  assign sel_777497 = array_index_777164 == array_index_773134 ? add_777496 : sel_777493;
  assign add_777500 = sel_777497 + 8'h01;
  assign sel_777501 = array_index_777164 == array_index_773140 ? add_777500 : sel_777497;
  assign add_777504 = sel_777501 + 8'h01;
  assign sel_777505 = array_index_777164 == array_index_773146 ? add_777504 : sel_777501;
  assign add_777508 = sel_777505 + 8'h01;
  assign sel_777509 = array_index_777164 == array_index_773152 ? add_777508 : sel_777505;
  assign add_777512 = sel_777509 + 8'h01;
  assign sel_777513 = array_index_777164 == array_index_773158 ? add_777512 : sel_777509;
  assign add_777516 = sel_777513 + 8'h01;
  assign sel_777517 = array_index_777164 == array_index_773164 ? add_777516 : sel_777513;
  assign add_777520 = sel_777517 + 8'h01;
  assign sel_777521 = array_index_777164 == array_index_773170 ? add_777520 : sel_777517;
  assign add_777525 = sel_777521 + 8'h01;
  assign array_index_777526 = set1_unflattened[7'h0d];
  assign sel_777527 = array_index_777164 == array_index_773176 ? add_777525 : sel_777521;
  assign add_777530 = sel_777527 + 8'h01;
  assign sel_777531 = array_index_777526 == array_index_772632 ? add_777530 : sel_777527;
  assign add_777534 = sel_777531 + 8'h01;
  assign sel_777535 = array_index_777526 == array_index_772636 ? add_777534 : sel_777531;
  assign add_777538 = sel_777535 + 8'h01;
  assign sel_777539 = array_index_777526 == array_index_772644 ? add_777538 : sel_777535;
  assign add_777542 = sel_777539 + 8'h01;
  assign sel_777543 = array_index_777526 == array_index_772652 ? add_777542 : sel_777539;
  assign add_777546 = sel_777543 + 8'h01;
  assign sel_777547 = array_index_777526 == array_index_772660 ? add_777546 : sel_777543;
  assign add_777550 = sel_777547 + 8'h01;
  assign sel_777551 = array_index_777526 == array_index_772668 ? add_777550 : sel_777547;
  assign add_777554 = sel_777551 + 8'h01;
  assign sel_777555 = array_index_777526 == array_index_772676 ? add_777554 : sel_777551;
  assign add_777558 = sel_777555 + 8'h01;
  assign sel_777559 = array_index_777526 == array_index_772684 ? add_777558 : sel_777555;
  assign add_777562 = sel_777559 + 8'h01;
  assign sel_777563 = array_index_777526 == array_index_772690 ? add_777562 : sel_777559;
  assign add_777566 = sel_777563 + 8'h01;
  assign sel_777567 = array_index_777526 == array_index_772696 ? add_777566 : sel_777563;
  assign add_777570 = sel_777567 + 8'h01;
  assign sel_777571 = array_index_777526 == array_index_772702 ? add_777570 : sel_777567;
  assign add_777574 = sel_777571 + 8'h01;
  assign sel_777575 = array_index_777526 == array_index_772708 ? add_777574 : sel_777571;
  assign add_777578 = sel_777575 + 8'h01;
  assign sel_777579 = array_index_777526 == array_index_772714 ? add_777578 : sel_777575;
  assign add_777582 = sel_777579 + 8'h01;
  assign sel_777583 = array_index_777526 == array_index_772720 ? add_777582 : sel_777579;
  assign add_777586 = sel_777583 + 8'h01;
  assign sel_777587 = array_index_777526 == array_index_772726 ? add_777586 : sel_777583;
  assign add_777590 = sel_777587 + 8'h01;
  assign sel_777591 = array_index_777526 == array_index_772732 ? add_777590 : sel_777587;
  assign add_777594 = sel_777591 + 8'h01;
  assign sel_777595 = array_index_777526 == array_index_772738 ? add_777594 : sel_777591;
  assign add_777598 = sel_777595 + 8'h01;
  assign sel_777599 = array_index_777526 == array_index_772744 ? add_777598 : sel_777595;
  assign add_777602 = sel_777599 + 8'h01;
  assign sel_777603 = array_index_777526 == array_index_772750 ? add_777602 : sel_777599;
  assign add_777606 = sel_777603 + 8'h01;
  assign sel_777607 = array_index_777526 == array_index_772756 ? add_777606 : sel_777603;
  assign add_777610 = sel_777607 + 8'h01;
  assign sel_777611 = array_index_777526 == array_index_772762 ? add_777610 : sel_777607;
  assign add_777614 = sel_777611 + 8'h01;
  assign sel_777615 = array_index_777526 == array_index_772768 ? add_777614 : sel_777611;
  assign add_777618 = sel_777615 + 8'h01;
  assign sel_777619 = array_index_777526 == array_index_772774 ? add_777618 : sel_777615;
  assign add_777622 = sel_777619 + 8'h01;
  assign sel_777623 = array_index_777526 == array_index_772780 ? add_777622 : sel_777619;
  assign add_777626 = sel_777623 + 8'h01;
  assign sel_777627 = array_index_777526 == array_index_772786 ? add_777626 : sel_777623;
  assign add_777630 = sel_777627 + 8'h01;
  assign sel_777631 = array_index_777526 == array_index_772792 ? add_777630 : sel_777627;
  assign add_777634 = sel_777631 + 8'h01;
  assign sel_777635 = array_index_777526 == array_index_772798 ? add_777634 : sel_777631;
  assign add_777638 = sel_777635 + 8'h01;
  assign sel_777639 = array_index_777526 == array_index_772804 ? add_777638 : sel_777635;
  assign add_777642 = sel_777639 + 8'h01;
  assign sel_777643 = array_index_777526 == array_index_772810 ? add_777642 : sel_777639;
  assign add_777646 = sel_777643 + 8'h01;
  assign sel_777647 = array_index_777526 == array_index_772816 ? add_777646 : sel_777643;
  assign add_777650 = sel_777647 + 8'h01;
  assign sel_777651 = array_index_777526 == array_index_772822 ? add_777650 : sel_777647;
  assign add_777654 = sel_777651 + 8'h01;
  assign sel_777655 = array_index_777526 == array_index_772828 ? add_777654 : sel_777651;
  assign add_777658 = sel_777655 + 8'h01;
  assign sel_777659 = array_index_777526 == array_index_772834 ? add_777658 : sel_777655;
  assign add_777662 = sel_777659 + 8'h01;
  assign sel_777663 = array_index_777526 == array_index_772840 ? add_777662 : sel_777659;
  assign add_777666 = sel_777663 + 8'h01;
  assign sel_777667 = array_index_777526 == array_index_772846 ? add_777666 : sel_777663;
  assign add_777670 = sel_777667 + 8'h01;
  assign sel_777671 = array_index_777526 == array_index_772852 ? add_777670 : sel_777667;
  assign add_777674 = sel_777671 + 8'h01;
  assign sel_777675 = array_index_777526 == array_index_772858 ? add_777674 : sel_777671;
  assign add_777678 = sel_777675 + 8'h01;
  assign sel_777679 = array_index_777526 == array_index_772864 ? add_777678 : sel_777675;
  assign add_777682 = sel_777679 + 8'h01;
  assign sel_777683 = array_index_777526 == array_index_772870 ? add_777682 : sel_777679;
  assign add_777686 = sel_777683 + 8'h01;
  assign sel_777687 = array_index_777526 == array_index_772876 ? add_777686 : sel_777683;
  assign add_777690 = sel_777687 + 8'h01;
  assign sel_777691 = array_index_777526 == array_index_772882 ? add_777690 : sel_777687;
  assign add_777694 = sel_777691 + 8'h01;
  assign sel_777695 = array_index_777526 == array_index_772888 ? add_777694 : sel_777691;
  assign add_777698 = sel_777695 + 8'h01;
  assign sel_777699 = array_index_777526 == array_index_772894 ? add_777698 : sel_777695;
  assign add_777702 = sel_777699 + 8'h01;
  assign sel_777703 = array_index_777526 == array_index_772900 ? add_777702 : sel_777699;
  assign add_777706 = sel_777703 + 8'h01;
  assign sel_777707 = array_index_777526 == array_index_772906 ? add_777706 : sel_777703;
  assign add_777710 = sel_777707 + 8'h01;
  assign sel_777711 = array_index_777526 == array_index_772912 ? add_777710 : sel_777707;
  assign add_777714 = sel_777711 + 8'h01;
  assign sel_777715 = array_index_777526 == array_index_772918 ? add_777714 : sel_777711;
  assign add_777718 = sel_777715 + 8'h01;
  assign sel_777719 = array_index_777526 == array_index_772924 ? add_777718 : sel_777715;
  assign add_777722 = sel_777719 + 8'h01;
  assign sel_777723 = array_index_777526 == array_index_772930 ? add_777722 : sel_777719;
  assign add_777726 = sel_777723 + 8'h01;
  assign sel_777727 = array_index_777526 == array_index_772936 ? add_777726 : sel_777723;
  assign add_777730 = sel_777727 + 8'h01;
  assign sel_777731 = array_index_777526 == array_index_772942 ? add_777730 : sel_777727;
  assign add_777734 = sel_777731 + 8'h01;
  assign sel_777735 = array_index_777526 == array_index_772948 ? add_777734 : sel_777731;
  assign add_777738 = sel_777735 + 8'h01;
  assign sel_777739 = array_index_777526 == array_index_772954 ? add_777738 : sel_777735;
  assign add_777742 = sel_777739 + 8'h01;
  assign sel_777743 = array_index_777526 == array_index_772960 ? add_777742 : sel_777739;
  assign add_777746 = sel_777743 + 8'h01;
  assign sel_777747 = array_index_777526 == array_index_772966 ? add_777746 : sel_777743;
  assign add_777750 = sel_777747 + 8'h01;
  assign sel_777751 = array_index_777526 == array_index_772972 ? add_777750 : sel_777747;
  assign add_777754 = sel_777751 + 8'h01;
  assign sel_777755 = array_index_777526 == array_index_772978 ? add_777754 : sel_777751;
  assign add_777758 = sel_777755 + 8'h01;
  assign sel_777759 = array_index_777526 == array_index_772984 ? add_777758 : sel_777755;
  assign add_777762 = sel_777759 + 8'h01;
  assign sel_777763 = array_index_777526 == array_index_772990 ? add_777762 : sel_777759;
  assign add_777766 = sel_777763 + 8'h01;
  assign sel_777767 = array_index_777526 == array_index_772996 ? add_777766 : sel_777763;
  assign add_777770 = sel_777767 + 8'h01;
  assign sel_777771 = array_index_777526 == array_index_773002 ? add_777770 : sel_777767;
  assign add_777774 = sel_777771 + 8'h01;
  assign sel_777775 = array_index_777526 == array_index_773008 ? add_777774 : sel_777771;
  assign add_777778 = sel_777775 + 8'h01;
  assign sel_777779 = array_index_777526 == array_index_773014 ? add_777778 : sel_777775;
  assign add_777782 = sel_777779 + 8'h01;
  assign sel_777783 = array_index_777526 == array_index_773020 ? add_777782 : sel_777779;
  assign add_777786 = sel_777783 + 8'h01;
  assign sel_777787 = array_index_777526 == array_index_773026 ? add_777786 : sel_777783;
  assign add_777790 = sel_777787 + 8'h01;
  assign sel_777791 = array_index_777526 == array_index_773032 ? add_777790 : sel_777787;
  assign add_777794 = sel_777791 + 8'h01;
  assign sel_777795 = array_index_777526 == array_index_773038 ? add_777794 : sel_777791;
  assign add_777798 = sel_777795 + 8'h01;
  assign sel_777799 = array_index_777526 == array_index_773044 ? add_777798 : sel_777795;
  assign add_777802 = sel_777799 + 8'h01;
  assign sel_777803 = array_index_777526 == array_index_773050 ? add_777802 : sel_777799;
  assign add_777806 = sel_777803 + 8'h01;
  assign sel_777807 = array_index_777526 == array_index_773056 ? add_777806 : sel_777803;
  assign add_777810 = sel_777807 + 8'h01;
  assign sel_777811 = array_index_777526 == array_index_773062 ? add_777810 : sel_777807;
  assign add_777814 = sel_777811 + 8'h01;
  assign sel_777815 = array_index_777526 == array_index_773068 ? add_777814 : sel_777811;
  assign add_777818 = sel_777815 + 8'h01;
  assign sel_777819 = array_index_777526 == array_index_773074 ? add_777818 : sel_777815;
  assign add_777822 = sel_777819 + 8'h01;
  assign sel_777823 = array_index_777526 == array_index_773080 ? add_777822 : sel_777819;
  assign add_777826 = sel_777823 + 8'h01;
  assign sel_777827 = array_index_777526 == array_index_773086 ? add_777826 : sel_777823;
  assign add_777830 = sel_777827 + 8'h01;
  assign sel_777831 = array_index_777526 == array_index_773092 ? add_777830 : sel_777827;
  assign add_777834 = sel_777831 + 8'h01;
  assign sel_777835 = array_index_777526 == array_index_773098 ? add_777834 : sel_777831;
  assign add_777838 = sel_777835 + 8'h01;
  assign sel_777839 = array_index_777526 == array_index_773104 ? add_777838 : sel_777835;
  assign add_777842 = sel_777839 + 8'h01;
  assign sel_777843 = array_index_777526 == array_index_773110 ? add_777842 : sel_777839;
  assign add_777846 = sel_777843 + 8'h01;
  assign sel_777847 = array_index_777526 == array_index_773116 ? add_777846 : sel_777843;
  assign add_777850 = sel_777847 + 8'h01;
  assign sel_777851 = array_index_777526 == array_index_773122 ? add_777850 : sel_777847;
  assign add_777854 = sel_777851 + 8'h01;
  assign sel_777855 = array_index_777526 == array_index_773128 ? add_777854 : sel_777851;
  assign add_777858 = sel_777855 + 8'h01;
  assign sel_777859 = array_index_777526 == array_index_773134 ? add_777858 : sel_777855;
  assign add_777862 = sel_777859 + 8'h01;
  assign sel_777863 = array_index_777526 == array_index_773140 ? add_777862 : sel_777859;
  assign add_777866 = sel_777863 + 8'h01;
  assign sel_777867 = array_index_777526 == array_index_773146 ? add_777866 : sel_777863;
  assign add_777870 = sel_777867 + 8'h01;
  assign sel_777871 = array_index_777526 == array_index_773152 ? add_777870 : sel_777867;
  assign add_777874 = sel_777871 + 8'h01;
  assign sel_777875 = array_index_777526 == array_index_773158 ? add_777874 : sel_777871;
  assign add_777878 = sel_777875 + 8'h01;
  assign sel_777879 = array_index_777526 == array_index_773164 ? add_777878 : sel_777875;
  assign add_777882 = sel_777879 + 8'h01;
  assign sel_777883 = array_index_777526 == array_index_773170 ? add_777882 : sel_777879;
  assign add_777887 = sel_777883 + 8'h01;
  assign array_index_777888 = set1_unflattened[7'h0e];
  assign sel_777889 = array_index_777526 == array_index_773176 ? add_777887 : sel_777883;
  assign add_777892 = sel_777889 + 8'h01;
  assign sel_777893 = array_index_777888 == array_index_772632 ? add_777892 : sel_777889;
  assign add_777896 = sel_777893 + 8'h01;
  assign sel_777897 = array_index_777888 == array_index_772636 ? add_777896 : sel_777893;
  assign add_777900 = sel_777897 + 8'h01;
  assign sel_777901 = array_index_777888 == array_index_772644 ? add_777900 : sel_777897;
  assign add_777904 = sel_777901 + 8'h01;
  assign sel_777905 = array_index_777888 == array_index_772652 ? add_777904 : sel_777901;
  assign add_777908 = sel_777905 + 8'h01;
  assign sel_777909 = array_index_777888 == array_index_772660 ? add_777908 : sel_777905;
  assign add_777912 = sel_777909 + 8'h01;
  assign sel_777913 = array_index_777888 == array_index_772668 ? add_777912 : sel_777909;
  assign add_777916 = sel_777913 + 8'h01;
  assign sel_777917 = array_index_777888 == array_index_772676 ? add_777916 : sel_777913;
  assign add_777920 = sel_777917 + 8'h01;
  assign sel_777921 = array_index_777888 == array_index_772684 ? add_777920 : sel_777917;
  assign add_777924 = sel_777921 + 8'h01;
  assign sel_777925 = array_index_777888 == array_index_772690 ? add_777924 : sel_777921;
  assign add_777928 = sel_777925 + 8'h01;
  assign sel_777929 = array_index_777888 == array_index_772696 ? add_777928 : sel_777925;
  assign add_777932 = sel_777929 + 8'h01;
  assign sel_777933 = array_index_777888 == array_index_772702 ? add_777932 : sel_777929;
  assign add_777936 = sel_777933 + 8'h01;
  assign sel_777937 = array_index_777888 == array_index_772708 ? add_777936 : sel_777933;
  assign add_777940 = sel_777937 + 8'h01;
  assign sel_777941 = array_index_777888 == array_index_772714 ? add_777940 : sel_777937;
  assign add_777944 = sel_777941 + 8'h01;
  assign sel_777945 = array_index_777888 == array_index_772720 ? add_777944 : sel_777941;
  assign add_777948 = sel_777945 + 8'h01;
  assign sel_777949 = array_index_777888 == array_index_772726 ? add_777948 : sel_777945;
  assign add_777952 = sel_777949 + 8'h01;
  assign sel_777953 = array_index_777888 == array_index_772732 ? add_777952 : sel_777949;
  assign add_777956 = sel_777953 + 8'h01;
  assign sel_777957 = array_index_777888 == array_index_772738 ? add_777956 : sel_777953;
  assign add_777960 = sel_777957 + 8'h01;
  assign sel_777961 = array_index_777888 == array_index_772744 ? add_777960 : sel_777957;
  assign add_777964 = sel_777961 + 8'h01;
  assign sel_777965 = array_index_777888 == array_index_772750 ? add_777964 : sel_777961;
  assign add_777968 = sel_777965 + 8'h01;
  assign sel_777969 = array_index_777888 == array_index_772756 ? add_777968 : sel_777965;
  assign add_777972 = sel_777969 + 8'h01;
  assign sel_777973 = array_index_777888 == array_index_772762 ? add_777972 : sel_777969;
  assign add_777976 = sel_777973 + 8'h01;
  assign sel_777977 = array_index_777888 == array_index_772768 ? add_777976 : sel_777973;
  assign add_777980 = sel_777977 + 8'h01;
  assign sel_777981 = array_index_777888 == array_index_772774 ? add_777980 : sel_777977;
  assign add_777984 = sel_777981 + 8'h01;
  assign sel_777985 = array_index_777888 == array_index_772780 ? add_777984 : sel_777981;
  assign add_777988 = sel_777985 + 8'h01;
  assign sel_777989 = array_index_777888 == array_index_772786 ? add_777988 : sel_777985;
  assign add_777992 = sel_777989 + 8'h01;
  assign sel_777993 = array_index_777888 == array_index_772792 ? add_777992 : sel_777989;
  assign add_777996 = sel_777993 + 8'h01;
  assign sel_777997 = array_index_777888 == array_index_772798 ? add_777996 : sel_777993;
  assign add_778000 = sel_777997 + 8'h01;
  assign sel_778001 = array_index_777888 == array_index_772804 ? add_778000 : sel_777997;
  assign add_778004 = sel_778001 + 8'h01;
  assign sel_778005 = array_index_777888 == array_index_772810 ? add_778004 : sel_778001;
  assign add_778008 = sel_778005 + 8'h01;
  assign sel_778009 = array_index_777888 == array_index_772816 ? add_778008 : sel_778005;
  assign add_778012 = sel_778009 + 8'h01;
  assign sel_778013 = array_index_777888 == array_index_772822 ? add_778012 : sel_778009;
  assign add_778016 = sel_778013 + 8'h01;
  assign sel_778017 = array_index_777888 == array_index_772828 ? add_778016 : sel_778013;
  assign add_778020 = sel_778017 + 8'h01;
  assign sel_778021 = array_index_777888 == array_index_772834 ? add_778020 : sel_778017;
  assign add_778024 = sel_778021 + 8'h01;
  assign sel_778025 = array_index_777888 == array_index_772840 ? add_778024 : sel_778021;
  assign add_778028 = sel_778025 + 8'h01;
  assign sel_778029 = array_index_777888 == array_index_772846 ? add_778028 : sel_778025;
  assign add_778032 = sel_778029 + 8'h01;
  assign sel_778033 = array_index_777888 == array_index_772852 ? add_778032 : sel_778029;
  assign add_778036 = sel_778033 + 8'h01;
  assign sel_778037 = array_index_777888 == array_index_772858 ? add_778036 : sel_778033;
  assign add_778040 = sel_778037 + 8'h01;
  assign sel_778041 = array_index_777888 == array_index_772864 ? add_778040 : sel_778037;
  assign add_778044 = sel_778041 + 8'h01;
  assign sel_778045 = array_index_777888 == array_index_772870 ? add_778044 : sel_778041;
  assign add_778048 = sel_778045 + 8'h01;
  assign sel_778049 = array_index_777888 == array_index_772876 ? add_778048 : sel_778045;
  assign add_778052 = sel_778049 + 8'h01;
  assign sel_778053 = array_index_777888 == array_index_772882 ? add_778052 : sel_778049;
  assign add_778056 = sel_778053 + 8'h01;
  assign sel_778057 = array_index_777888 == array_index_772888 ? add_778056 : sel_778053;
  assign add_778060 = sel_778057 + 8'h01;
  assign sel_778061 = array_index_777888 == array_index_772894 ? add_778060 : sel_778057;
  assign add_778064 = sel_778061 + 8'h01;
  assign sel_778065 = array_index_777888 == array_index_772900 ? add_778064 : sel_778061;
  assign add_778068 = sel_778065 + 8'h01;
  assign sel_778069 = array_index_777888 == array_index_772906 ? add_778068 : sel_778065;
  assign add_778072 = sel_778069 + 8'h01;
  assign sel_778073 = array_index_777888 == array_index_772912 ? add_778072 : sel_778069;
  assign add_778076 = sel_778073 + 8'h01;
  assign sel_778077 = array_index_777888 == array_index_772918 ? add_778076 : sel_778073;
  assign add_778080 = sel_778077 + 8'h01;
  assign sel_778081 = array_index_777888 == array_index_772924 ? add_778080 : sel_778077;
  assign add_778084 = sel_778081 + 8'h01;
  assign sel_778085 = array_index_777888 == array_index_772930 ? add_778084 : sel_778081;
  assign add_778088 = sel_778085 + 8'h01;
  assign sel_778089 = array_index_777888 == array_index_772936 ? add_778088 : sel_778085;
  assign add_778092 = sel_778089 + 8'h01;
  assign sel_778093 = array_index_777888 == array_index_772942 ? add_778092 : sel_778089;
  assign add_778096 = sel_778093 + 8'h01;
  assign sel_778097 = array_index_777888 == array_index_772948 ? add_778096 : sel_778093;
  assign add_778100 = sel_778097 + 8'h01;
  assign sel_778101 = array_index_777888 == array_index_772954 ? add_778100 : sel_778097;
  assign add_778104 = sel_778101 + 8'h01;
  assign sel_778105 = array_index_777888 == array_index_772960 ? add_778104 : sel_778101;
  assign add_778108 = sel_778105 + 8'h01;
  assign sel_778109 = array_index_777888 == array_index_772966 ? add_778108 : sel_778105;
  assign add_778112 = sel_778109 + 8'h01;
  assign sel_778113 = array_index_777888 == array_index_772972 ? add_778112 : sel_778109;
  assign add_778116 = sel_778113 + 8'h01;
  assign sel_778117 = array_index_777888 == array_index_772978 ? add_778116 : sel_778113;
  assign add_778120 = sel_778117 + 8'h01;
  assign sel_778121 = array_index_777888 == array_index_772984 ? add_778120 : sel_778117;
  assign add_778124 = sel_778121 + 8'h01;
  assign sel_778125 = array_index_777888 == array_index_772990 ? add_778124 : sel_778121;
  assign add_778128 = sel_778125 + 8'h01;
  assign sel_778129 = array_index_777888 == array_index_772996 ? add_778128 : sel_778125;
  assign add_778132 = sel_778129 + 8'h01;
  assign sel_778133 = array_index_777888 == array_index_773002 ? add_778132 : sel_778129;
  assign add_778136 = sel_778133 + 8'h01;
  assign sel_778137 = array_index_777888 == array_index_773008 ? add_778136 : sel_778133;
  assign add_778140 = sel_778137 + 8'h01;
  assign sel_778141 = array_index_777888 == array_index_773014 ? add_778140 : sel_778137;
  assign add_778144 = sel_778141 + 8'h01;
  assign sel_778145 = array_index_777888 == array_index_773020 ? add_778144 : sel_778141;
  assign add_778148 = sel_778145 + 8'h01;
  assign sel_778149 = array_index_777888 == array_index_773026 ? add_778148 : sel_778145;
  assign add_778152 = sel_778149 + 8'h01;
  assign sel_778153 = array_index_777888 == array_index_773032 ? add_778152 : sel_778149;
  assign add_778156 = sel_778153 + 8'h01;
  assign sel_778157 = array_index_777888 == array_index_773038 ? add_778156 : sel_778153;
  assign add_778160 = sel_778157 + 8'h01;
  assign sel_778161 = array_index_777888 == array_index_773044 ? add_778160 : sel_778157;
  assign add_778164 = sel_778161 + 8'h01;
  assign sel_778165 = array_index_777888 == array_index_773050 ? add_778164 : sel_778161;
  assign add_778168 = sel_778165 + 8'h01;
  assign sel_778169 = array_index_777888 == array_index_773056 ? add_778168 : sel_778165;
  assign add_778172 = sel_778169 + 8'h01;
  assign sel_778173 = array_index_777888 == array_index_773062 ? add_778172 : sel_778169;
  assign add_778176 = sel_778173 + 8'h01;
  assign sel_778177 = array_index_777888 == array_index_773068 ? add_778176 : sel_778173;
  assign add_778180 = sel_778177 + 8'h01;
  assign sel_778181 = array_index_777888 == array_index_773074 ? add_778180 : sel_778177;
  assign add_778184 = sel_778181 + 8'h01;
  assign sel_778185 = array_index_777888 == array_index_773080 ? add_778184 : sel_778181;
  assign add_778188 = sel_778185 + 8'h01;
  assign sel_778189 = array_index_777888 == array_index_773086 ? add_778188 : sel_778185;
  assign add_778192 = sel_778189 + 8'h01;
  assign sel_778193 = array_index_777888 == array_index_773092 ? add_778192 : sel_778189;
  assign add_778196 = sel_778193 + 8'h01;
  assign sel_778197 = array_index_777888 == array_index_773098 ? add_778196 : sel_778193;
  assign add_778200 = sel_778197 + 8'h01;
  assign sel_778201 = array_index_777888 == array_index_773104 ? add_778200 : sel_778197;
  assign add_778204 = sel_778201 + 8'h01;
  assign sel_778205 = array_index_777888 == array_index_773110 ? add_778204 : sel_778201;
  assign add_778208 = sel_778205 + 8'h01;
  assign sel_778209 = array_index_777888 == array_index_773116 ? add_778208 : sel_778205;
  assign add_778212 = sel_778209 + 8'h01;
  assign sel_778213 = array_index_777888 == array_index_773122 ? add_778212 : sel_778209;
  assign add_778216 = sel_778213 + 8'h01;
  assign sel_778217 = array_index_777888 == array_index_773128 ? add_778216 : sel_778213;
  assign add_778220 = sel_778217 + 8'h01;
  assign sel_778221 = array_index_777888 == array_index_773134 ? add_778220 : sel_778217;
  assign add_778224 = sel_778221 + 8'h01;
  assign sel_778225 = array_index_777888 == array_index_773140 ? add_778224 : sel_778221;
  assign add_778228 = sel_778225 + 8'h01;
  assign sel_778229 = array_index_777888 == array_index_773146 ? add_778228 : sel_778225;
  assign add_778232 = sel_778229 + 8'h01;
  assign sel_778233 = array_index_777888 == array_index_773152 ? add_778232 : sel_778229;
  assign add_778236 = sel_778233 + 8'h01;
  assign sel_778237 = array_index_777888 == array_index_773158 ? add_778236 : sel_778233;
  assign add_778240 = sel_778237 + 8'h01;
  assign sel_778241 = array_index_777888 == array_index_773164 ? add_778240 : sel_778237;
  assign add_778244 = sel_778241 + 8'h01;
  assign sel_778245 = array_index_777888 == array_index_773170 ? add_778244 : sel_778241;
  assign add_778249 = sel_778245 + 8'h01;
  assign array_index_778250 = set1_unflattened[7'h0f];
  assign sel_778251 = array_index_777888 == array_index_773176 ? add_778249 : sel_778245;
  assign add_778254 = sel_778251 + 8'h01;
  assign sel_778255 = array_index_778250 == array_index_772632 ? add_778254 : sel_778251;
  assign add_778258 = sel_778255 + 8'h01;
  assign sel_778259 = array_index_778250 == array_index_772636 ? add_778258 : sel_778255;
  assign add_778262 = sel_778259 + 8'h01;
  assign sel_778263 = array_index_778250 == array_index_772644 ? add_778262 : sel_778259;
  assign add_778266 = sel_778263 + 8'h01;
  assign sel_778267 = array_index_778250 == array_index_772652 ? add_778266 : sel_778263;
  assign add_778270 = sel_778267 + 8'h01;
  assign sel_778271 = array_index_778250 == array_index_772660 ? add_778270 : sel_778267;
  assign add_778274 = sel_778271 + 8'h01;
  assign sel_778275 = array_index_778250 == array_index_772668 ? add_778274 : sel_778271;
  assign add_778278 = sel_778275 + 8'h01;
  assign sel_778279 = array_index_778250 == array_index_772676 ? add_778278 : sel_778275;
  assign add_778282 = sel_778279 + 8'h01;
  assign sel_778283 = array_index_778250 == array_index_772684 ? add_778282 : sel_778279;
  assign add_778286 = sel_778283 + 8'h01;
  assign sel_778287 = array_index_778250 == array_index_772690 ? add_778286 : sel_778283;
  assign add_778290 = sel_778287 + 8'h01;
  assign sel_778291 = array_index_778250 == array_index_772696 ? add_778290 : sel_778287;
  assign add_778294 = sel_778291 + 8'h01;
  assign sel_778295 = array_index_778250 == array_index_772702 ? add_778294 : sel_778291;
  assign add_778298 = sel_778295 + 8'h01;
  assign sel_778299 = array_index_778250 == array_index_772708 ? add_778298 : sel_778295;
  assign add_778302 = sel_778299 + 8'h01;
  assign sel_778303 = array_index_778250 == array_index_772714 ? add_778302 : sel_778299;
  assign add_778306 = sel_778303 + 8'h01;
  assign sel_778307 = array_index_778250 == array_index_772720 ? add_778306 : sel_778303;
  assign add_778310 = sel_778307 + 8'h01;
  assign sel_778311 = array_index_778250 == array_index_772726 ? add_778310 : sel_778307;
  assign add_778314 = sel_778311 + 8'h01;
  assign sel_778315 = array_index_778250 == array_index_772732 ? add_778314 : sel_778311;
  assign add_778318 = sel_778315 + 8'h01;
  assign sel_778319 = array_index_778250 == array_index_772738 ? add_778318 : sel_778315;
  assign add_778322 = sel_778319 + 8'h01;
  assign sel_778323 = array_index_778250 == array_index_772744 ? add_778322 : sel_778319;
  assign add_778326 = sel_778323 + 8'h01;
  assign sel_778327 = array_index_778250 == array_index_772750 ? add_778326 : sel_778323;
  assign add_778330 = sel_778327 + 8'h01;
  assign sel_778331 = array_index_778250 == array_index_772756 ? add_778330 : sel_778327;
  assign add_778334 = sel_778331 + 8'h01;
  assign sel_778335 = array_index_778250 == array_index_772762 ? add_778334 : sel_778331;
  assign add_778338 = sel_778335 + 8'h01;
  assign sel_778339 = array_index_778250 == array_index_772768 ? add_778338 : sel_778335;
  assign add_778342 = sel_778339 + 8'h01;
  assign sel_778343 = array_index_778250 == array_index_772774 ? add_778342 : sel_778339;
  assign add_778346 = sel_778343 + 8'h01;
  assign sel_778347 = array_index_778250 == array_index_772780 ? add_778346 : sel_778343;
  assign add_778350 = sel_778347 + 8'h01;
  assign sel_778351 = array_index_778250 == array_index_772786 ? add_778350 : sel_778347;
  assign add_778354 = sel_778351 + 8'h01;
  assign sel_778355 = array_index_778250 == array_index_772792 ? add_778354 : sel_778351;
  assign add_778358 = sel_778355 + 8'h01;
  assign sel_778359 = array_index_778250 == array_index_772798 ? add_778358 : sel_778355;
  assign add_778362 = sel_778359 + 8'h01;
  assign sel_778363 = array_index_778250 == array_index_772804 ? add_778362 : sel_778359;
  assign add_778366 = sel_778363 + 8'h01;
  assign sel_778367 = array_index_778250 == array_index_772810 ? add_778366 : sel_778363;
  assign add_778370 = sel_778367 + 8'h01;
  assign sel_778371 = array_index_778250 == array_index_772816 ? add_778370 : sel_778367;
  assign add_778374 = sel_778371 + 8'h01;
  assign sel_778375 = array_index_778250 == array_index_772822 ? add_778374 : sel_778371;
  assign add_778378 = sel_778375 + 8'h01;
  assign sel_778379 = array_index_778250 == array_index_772828 ? add_778378 : sel_778375;
  assign add_778382 = sel_778379 + 8'h01;
  assign sel_778383 = array_index_778250 == array_index_772834 ? add_778382 : sel_778379;
  assign add_778386 = sel_778383 + 8'h01;
  assign sel_778387 = array_index_778250 == array_index_772840 ? add_778386 : sel_778383;
  assign add_778390 = sel_778387 + 8'h01;
  assign sel_778391 = array_index_778250 == array_index_772846 ? add_778390 : sel_778387;
  assign add_778394 = sel_778391 + 8'h01;
  assign sel_778395 = array_index_778250 == array_index_772852 ? add_778394 : sel_778391;
  assign add_778398 = sel_778395 + 8'h01;
  assign sel_778399 = array_index_778250 == array_index_772858 ? add_778398 : sel_778395;
  assign add_778402 = sel_778399 + 8'h01;
  assign sel_778403 = array_index_778250 == array_index_772864 ? add_778402 : sel_778399;
  assign add_778406 = sel_778403 + 8'h01;
  assign sel_778407 = array_index_778250 == array_index_772870 ? add_778406 : sel_778403;
  assign add_778410 = sel_778407 + 8'h01;
  assign sel_778411 = array_index_778250 == array_index_772876 ? add_778410 : sel_778407;
  assign add_778414 = sel_778411 + 8'h01;
  assign sel_778415 = array_index_778250 == array_index_772882 ? add_778414 : sel_778411;
  assign add_778418 = sel_778415 + 8'h01;
  assign sel_778419 = array_index_778250 == array_index_772888 ? add_778418 : sel_778415;
  assign add_778422 = sel_778419 + 8'h01;
  assign sel_778423 = array_index_778250 == array_index_772894 ? add_778422 : sel_778419;
  assign add_778426 = sel_778423 + 8'h01;
  assign sel_778427 = array_index_778250 == array_index_772900 ? add_778426 : sel_778423;
  assign add_778430 = sel_778427 + 8'h01;
  assign sel_778431 = array_index_778250 == array_index_772906 ? add_778430 : sel_778427;
  assign add_778434 = sel_778431 + 8'h01;
  assign sel_778435 = array_index_778250 == array_index_772912 ? add_778434 : sel_778431;
  assign add_778438 = sel_778435 + 8'h01;
  assign sel_778439 = array_index_778250 == array_index_772918 ? add_778438 : sel_778435;
  assign add_778442 = sel_778439 + 8'h01;
  assign sel_778443 = array_index_778250 == array_index_772924 ? add_778442 : sel_778439;
  assign add_778446 = sel_778443 + 8'h01;
  assign sel_778447 = array_index_778250 == array_index_772930 ? add_778446 : sel_778443;
  assign add_778450 = sel_778447 + 8'h01;
  assign sel_778451 = array_index_778250 == array_index_772936 ? add_778450 : sel_778447;
  assign add_778454 = sel_778451 + 8'h01;
  assign sel_778455 = array_index_778250 == array_index_772942 ? add_778454 : sel_778451;
  assign add_778458 = sel_778455 + 8'h01;
  assign sel_778459 = array_index_778250 == array_index_772948 ? add_778458 : sel_778455;
  assign add_778462 = sel_778459 + 8'h01;
  assign sel_778463 = array_index_778250 == array_index_772954 ? add_778462 : sel_778459;
  assign add_778466 = sel_778463 + 8'h01;
  assign sel_778467 = array_index_778250 == array_index_772960 ? add_778466 : sel_778463;
  assign add_778470 = sel_778467 + 8'h01;
  assign sel_778471 = array_index_778250 == array_index_772966 ? add_778470 : sel_778467;
  assign add_778474 = sel_778471 + 8'h01;
  assign sel_778475 = array_index_778250 == array_index_772972 ? add_778474 : sel_778471;
  assign add_778478 = sel_778475 + 8'h01;
  assign sel_778479 = array_index_778250 == array_index_772978 ? add_778478 : sel_778475;
  assign add_778482 = sel_778479 + 8'h01;
  assign sel_778483 = array_index_778250 == array_index_772984 ? add_778482 : sel_778479;
  assign add_778486 = sel_778483 + 8'h01;
  assign sel_778487 = array_index_778250 == array_index_772990 ? add_778486 : sel_778483;
  assign add_778490 = sel_778487 + 8'h01;
  assign sel_778491 = array_index_778250 == array_index_772996 ? add_778490 : sel_778487;
  assign add_778494 = sel_778491 + 8'h01;
  assign sel_778495 = array_index_778250 == array_index_773002 ? add_778494 : sel_778491;
  assign add_778498 = sel_778495 + 8'h01;
  assign sel_778499 = array_index_778250 == array_index_773008 ? add_778498 : sel_778495;
  assign add_778502 = sel_778499 + 8'h01;
  assign sel_778503 = array_index_778250 == array_index_773014 ? add_778502 : sel_778499;
  assign add_778506 = sel_778503 + 8'h01;
  assign sel_778507 = array_index_778250 == array_index_773020 ? add_778506 : sel_778503;
  assign add_778510 = sel_778507 + 8'h01;
  assign sel_778511 = array_index_778250 == array_index_773026 ? add_778510 : sel_778507;
  assign add_778514 = sel_778511 + 8'h01;
  assign sel_778515 = array_index_778250 == array_index_773032 ? add_778514 : sel_778511;
  assign add_778518 = sel_778515 + 8'h01;
  assign sel_778519 = array_index_778250 == array_index_773038 ? add_778518 : sel_778515;
  assign add_778522 = sel_778519 + 8'h01;
  assign sel_778523 = array_index_778250 == array_index_773044 ? add_778522 : sel_778519;
  assign add_778526 = sel_778523 + 8'h01;
  assign sel_778527 = array_index_778250 == array_index_773050 ? add_778526 : sel_778523;
  assign add_778530 = sel_778527 + 8'h01;
  assign sel_778531 = array_index_778250 == array_index_773056 ? add_778530 : sel_778527;
  assign add_778534 = sel_778531 + 8'h01;
  assign sel_778535 = array_index_778250 == array_index_773062 ? add_778534 : sel_778531;
  assign add_778538 = sel_778535 + 8'h01;
  assign sel_778539 = array_index_778250 == array_index_773068 ? add_778538 : sel_778535;
  assign add_778542 = sel_778539 + 8'h01;
  assign sel_778543 = array_index_778250 == array_index_773074 ? add_778542 : sel_778539;
  assign add_778546 = sel_778543 + 8'h01;
  assign sel_778547 = array_index_778250 == array_index_773080 ? add_778546 : sel_778543;
  assign add_778550 = sel_778547 + 8'h01;
  assign sel_778551 = array_index_778250 == array_index_773086 ? add_778550 : sel_778547;
  assign add_778554 = sel_778551 + 8'h01;
  assign sel_778555 = array_index_778250 == array_index_773092 ? add_778554 : sel_778551;
  assign add_778558 = sel_778555 + 8'h01;
  assign sel_778559 = array_index_778250 == array_index_773098 ? add_778558 : sel_778555;
  assign add_778562 = sel_778559 + 8'h01;
  assign sel_778563 = array_index_778250 == array_index_773104 ? add_778562 : sel_778559;
  assign add_778566 = sel_778563 + 8'h01;
  assign sel_778567 = array_index_778250 == array_index_773110 ? add_778566 : sel_778563;
  assign add_778570 = sel_778567 + 8'h01;
  assign sel_778571 = array_index_778250 == array_index_773116 ? add_778570 : sel_778567;
  assign add_778574 = sel_778571 + 8'h01;
  assign sel_778575 = array_index_778250 == array_index_773122 ? add_778574 : sel_778571;
  assign add_778578 = sel_778575 + 8'h01;
  assign sel_778579 = array_index_778250 == array_index_773128 ? add_778578 : sel_778575;
  assign add_778582 = sel_778579 + 8'h01;
  assign sel_778583 = array_index_778250 == array_index_773134 ? add_778582 : sel_778579;
  assign add_778586 = sel_778583 + 8'h01;
  assign sel_778587 = array_index_778250 == array_index_773140 ? add_778586 : sel_778583;
  assign add_778590 = sel_778587 + 8'h01;
  assign sel_778591 = array_index_778250 == array_index_773146 ? add_778590 : sel_778587;
  assign add_778594 = sel_778591 + 8'h01;
  assign sel_778595 = array_index_778250 == array_index_773152 ? add_778594 : sel_778591;
  assign add_778598 = sel_778595 + 8'h01;
  assign sel_778599 = array_index_778250 == array_index_773158 ? add_778598 : sel_778595;
  assign add_778602 = sel_778599 + 8'h01;
  assign sel_778603 = array_index_778250 == array_index_773164 ? add_778602 : sel_778599;
  assign add_778606 = sel_778603 + 8'h01;
  assign sel_778607 = array_index_778250 == array_index_773170 ? add_778606 : sel_778603;
  assign add_778611 = sel_778607 + 8'h01;
  assign array_index_778612 = set1_unflattened[7'h10];
  assign sel_778613 = array_index_778250 == array_index_773176 ? add_778611 : sel_778607;
  assign add_778616 = sel_778613 + 8'h01;
  assign sel_778617 = array_index_778612 == array_index_772632 ? add_778616 : sel_778613;
  assign add_778620 = sel_778617 + 8'h01;
  assign sel_778621 = array_index_778612 == array_index_772636 ? add_778620 : sel_778617;
  assign add_778624 = sel_778621 + 8'h01;
  assign sel_778625 = array_index_778612 == array_index_772644 ? add_778624 : sel_778621;
  assign add_778628 = sel_778625 + 8'h01;
  assign sel_778629 = array_index_778612 == array_index_772652 ? add_778628 : sel_778625;
  assign add_778632 = sel_778629 + 8'h01;
  assign sel_778633 = array_index_778612 == array_index_772660 ? add_778632 : sel_778629;
  assign add_778636 = sel_778633 + 8'h01;
  assign sel_778637 = array_index_778612 == array_index_772668 ? add_778636 : sel_778633;
  assign add_778640 = sel_778637 + 8'h01;
  assign sel_778641 = array_index_778612 == array_index_772676 ? add_778640 : sel_778637;
  assign add_778644 = sel_778641 + 8'h01;
  assign sel_778645 = array_index_778612 == array_index_772684 ? add_778644 : sel_778641;
  assign add_778648 = sel_778645 + 8'h01;
  assign sel_778649 = array_index_778612 == array_index_772690 ? add_778648 : sel_778645;
  assign add_778652 = sel_778649 + 8'h01;
  assign sel_778653 = array_index_778612 == array_index_772696 ? add_778652 : sel_778649;
  assign add_778656 = sel_778653 + 8'h01;
  assign sel_778657 = array_index_778612 == array_index_772702 ? add_778656 : sel_778653;
  assign add_778660 = sel_778657 + 8'h01;
  assign sel_778661 = array_index_778612 == array_index_772708 ? add_778660 : sel_778657;
  assign add_778664 = sel_778661 + 8'h01;
  assign sel_778665 = array_index_778612 == array_index_772714 ? add_778664 : sel_778661;
  assign add_778668 = sel_778665 + 8'h01;
  assign sel_778669 = array_index_778612 == array_index_772720 ? add_778668 : sel_778665;
  assign add_778672 = sel_778669 + 8'h01;
  assign sel_778673 = array_index_778612 == array_index_772726 ? add_778672 : sel_778669;
  assign add_778676 = sel_778673 + 8'h01;
  assign sel_778677 = array_index_778612 == array_index_772732 ? add_778676 : sel_778673;
  assign add_778680 = sel_778677 + 8'h01;
  assign sel_778681 = array_index_778612 == array_index_772738 ? add_778680 : sel_778677;
  assign add_778684 = sel_778681 + 8'h01;
  assign sel_778685 = array_index_778612 == array_index_772744 ? add_778684 : sel_778681;
  assign add_778688 = sel_778685 + 8'h01;
  assign sel_778689 = array_index_778612 == array_index_772750 ? add_778688 : sel_778685;
  assign add_778692 = sel_778689 + 8'h01;
  assign sel_778693 = array_index_778612 == array_index_772756 ? add_778692 : sel_778689;
  assign add_778696 = sel_778693 + 8'h01;
  assign sel_778697 = array_index_778612 == array_index_772762 ? add_778696 : sel_778693;
  assign add_778700 = sel_778697 + 8'h01;
  assign sel_778701 = array_index_778612 == array_index_772768 ? add_778700 : sel_778697;
  assign add_778704 = sel_778701 + 8'h01;
  assign sel_778705 = array_index_778612 == array_index_772774 ? add_778704 : sel_778701;
  assign add_778708 = sel_778705 + 8'h01;
  assign sel_778709 = array_index_778612 == array_index_772780 ? add_778708 : sel_778705;
  assign add_778712 = sel_778709 + 8'h01;
  assign sel_778713 = array_index_778612 == array_index_772786 ? add_778712 : sel_778709;
  assign add_778716 = sel_778713 + 8'h01;
  assign sel_778717 = array_index_778612 == array_index_772792 ? add_778716 : sel_778713;
  assign add_778720 = sel_778717 + 8'h01;
  assign sel_778721 = array_index_778612 == array_index_772798 ? add_778720 : sel_778717;
  assign add_778724 = sel_778721 + 8'h01;
  assign sel_778725 = array_index_778612 == array_index_772804 ? add_778724 : sel_778721;
  assign add_778728 = sel_778725 + 8'h01;
  assign sel_778729 = array_index_778612 == array_index_772810 ? add_778728 : sel_778725;
  assign add_778732 = sel_778729 + 8'h01;
  assign sel_778733 = array_index_778612 == array_index_772816 ? add_778732 : sel_778729;
  assign add_778736 = sel_778733 + 8'h01;
  assign sel_778737 = array_index_778612 == array_index_772822 ? add_778736 : sel_778733;
  assign add_778740 = sel_778737 + 8'h01;
  assign sel_778741 = array_index_778612 == array_index_772828 ? add_778740 : sel_778737;
  assign add_778744 = sel_778741 + 8'h01;
  assign sel_778745 = array_index_778612 == array_index_772834 ? add_778744 : sel_778741;
  assign add_778748 = sel_778745 + 8'h01;
  assign sel_778749 = array_index_778612 == array_index_772840 ? add_778748 : sel_778745;
  assign add_778752 = sel_778749 + 8'h01;
  assign sel_778753 = array_index_778612 == array_index_772846 ? add_778752 : sel_778749;
  assign add_778756 = sel_778753 + 8'h01;
  assign sel_778757 = array_index_778612 == array_index_772852 ? add_778756 : sel_778753;
  assign add_778760 = sel_778757 + 8'h01;
  assign sel_778761 = array_index_778612 == array_index_772858 ? add_778760 : sel_778757;
  assign add_778764 = sel_778761 + 8'h01;
  assign sel_778765 = array_index_778612 == array_index_772864 ? add_778764 : sel_778761;
  assign add_778768 = sel_778765 + 8'h01;
  assign sel_778769 = array_index_778612 == array_index_772870 ? add_778768 : sel_778765;
  assign add_778772 = sel_778769 + 8'h01;
  assign sel_778773 = array_index_778612 == array_index_772876 ? add_778772 : sel_778769;
  assign add_778776 = sel_778773 + 8'h01;
  assign sel_778777 = array_index_778612 == array_index_772882 ? add_778776 : sel_778773;
  assign add_778780 = sel_778777 + 8'h01;
  assign sel_778781 = array_index_778612 == array_index_772888 ? add_778780 : sel_778777;
  assign add_778784 = sel_778781 + 8'h01;
  assign sel_778785 = array_index_778612 == array_index_772894 ? add_778784 : sel_778781;
  assign add_778788 = sel_778785 + 8'h01;
  assign sel_778789 = array_index_778612 == array_index_772900 ? add_778788 : sel_778785;
  assign add_778792 = sel_778789 + 8'h01;
  assign sel_778793 = array_index_778612 == array_index_772906 ? add_778792 : sel_778789;
  assign add_778796 = sel_778793 + 8'h01;
  assign sel_778797 = array_index_778612 == array_index_772912 ? add_778796 : sel_778793;
  assign add_778800 = sel_778797 + 8'h01;
  assign sel_778801 = array_index_778612 == array_index_772918 ? add_778800 : sel_778797;
  assign add_778804 = sel_778801 + 8'h01;
  assign sel_778805 = array_index_778612 == array_index_772924 ? add_778804 : sel_778801;
  assign add_778808 = sel_778805 + 8'h01;
  assign sel_778809 = array_index_778612 == array_index_772930 ? add_778808 : sel_778805;
  assign add_778812 = sel_778809 + 8'h01;
  assign sel_778813 = array_index_778612 == array_index_772936 ? add_778812 : sel_778809;
  assign add_778816 = sel_778813 + 8'h01;
  assign sel_778817 = array_index_778612 == array_index_772942 ? add_778816 : sel_778813;
  assign add_778820 = sel_778817 + 8'h01;
  assign sel_778821 = array_index_778612 == array_index_772948 ? add_778820 : sel_778817;
  assign add_778824 = sel_778821 + 8'h01;
  assign sel_778825 = array_index_778612 == array_index_772954 ? add_778824 : sel_778821;
  assign add_778828 = sel_778825 + 8'h01;
  assign sel_778829 = array_index_778612 == array_index_772960 ? add_778828 : sel_778825;
  assign add_778832 = sel_778829 + 8'h01;
  assign sel_778833 = array_index_778612 == array_index_772966 ? add_778832 : sel_778829;
  assign add_778836 = sel_778833 + 8'h01;
  assign sel_778837 = array_index_778612 == array_index_772972 ? add_778836 : sel_778833;
  assign add_778840 = sel_778837 + 8'h01;
  assign sel_778841 = array_index_778612 == array_index_772978 ? add_778840 : sel_778837;
  assign add_778844 = sel_778841 + 8'h01;
  assign sel_778845 = array_index_778612 == array_index_772984 ? add_778844 : sel_778841;
  assign add_778848 = sel_778845 + 8'h01;
  assign sel_778849 = array_index_778612 == array_index_772990 ? add_778848 : sel_778845;
  assign add_778852 = sel_778849 + 8'h01;
  assign sel_778853 = array_index_778612 == array_index_772996 ? add_778852 : sel_778849;
  assign add_778856 = sel_778853 + 8'h01;
  assign sel_778857 = array_index_778612 == array_index_773002 ? add_778856 : sel_778853;
  assign add_778860 = sel_778857 + 8'h01;
  assign sel_778861 = array_index_778612 == array_index_773008 ? add_778860 : sel_778857;
  assign add_778864 = sel_778861 + 8'h01;
  assign sel_778865 = array_index_778612 == array_index_773014 ? add_778864 : sel_778861;
  assign add_778868 = sel_778865 + 8'h01;
  assign sel_778869 = array_index_778612 == array_index_773020 ? add_778868 : sel_778865;
  assign add_778872 = sel_778869 + 8'h01;
  assign sel_778873 = array_index_778612 == array_index_773026 ? add_778872 : sel_778869;
  assign add_778876 = sel_778873 + 8'h01;
  assign sel_778877 = array_index_778612 == array_index_773032 ? add_778876 : sel_778873;
  assign add_778880 = sel_778877 + 8'h01;
  assign sel_778881 = array_index_778612 == array_index_773038 ? add_778880 : sel_778877;
  assign add_778884 = sel_778881 + 8'h01;
  assign sel_778885 = array_index_778612 == array_index_773044 ? add_778884 : sel_778881;
  assign add_778888 = sel_778885 + 8'h01;
  assign sel_778889 = array_index_778612 == array_index_773050 ? add_778888 : sel_778885;
  assign add_778892 = sel_778889 + 8'h01;
  assign sel_778893 = array_index_778612 == array_index_773056 ? add_778892 : sel_778889;
  assign add_778896 = sel_778893 + 8'h01;
  assign sel_778897 = array_index_778612 == array_index_773062 ? add_778896 : sel_778893;
  assign add_778900 = sel_778897 + 8'h01;
  assign sel_778901 = array_index_778612 == array_index_773068 ? add_778900 : sel_778897;
  assign add_778904 = sel_778901 + 8'h01;
  assign sel_778905 = array_index_778612 == array_index_773074 ? add_778904 : sel_778901;
  assign add_778908 = sel_778905 + 8'h01;
  assign sel_778909 = array_index_778612 == array_index_773080 ? add_778908 : sel_778905;
  assign add_778912 = sel_778909 + 8'h01;
  assign sel_778913 = array_index_778612 == array_index_773086 ? add_778912 : sel_778909;
  assign add_778916 = sel_778913 + 8'h01;
  assign sel_778917 = array_index_778612 == array_index_773092 ? add_778916 : sel_778913;
  assign add_778920 = sel_778917 + 8'h01;
  assign sel_778921 = array_index_778612 == array_index_773098 ? add_778920 : sel_778917;
  assign add_778924 = sel_778921 + 8'h01;
  assign sel_778925 = array_index_778612 == array_index_773104 ? add_778924 : sel_778921;
  assign add_778928 = sel_778925 + 8'h01;
  assign sel_778929 = array_index_778612 == array_index_773110 ? add_778928 : sel_778925;
  assign add_778932 = sel_778929 + 8'h01;
  assign sel_778933 = array_index_778612 == array_index_773116 ? add_778932 : sel_778929;
  assign add_778936 = sel_778933 + 8'h01;
  assign sel_778937 = array_index_778612 == array_index_773122 ? add_778936 : sel_778933;
  assign add_778940 = sel_778937 + 8'h01;
  assign sel_778941 = array_index_778612 == array_index_773128 ? add_778940 : sel_778937;
  assign add_778944 = sel_778941 + 8'h01;
  assign sel_778945 = array_index_778612 == array_index_773134 ? add_778944 : sel_778941;
  assign add_778948 = sel_778945 + 8'h01;
  assign sel_778949 = array_index_778612 == array_index_773140 ? add_778948 : sel_778945;
  assign add_778952 = sel_778949 + 8'h01;
  assign sel_778953 = array_index_778612 == array_index_773146 ? add_778952 : sel_778949;
  assign add_778956 = sel_778953 + 8'h01;
  assign sel_778957 = array_index_778612 == array_index_773152 ? add_778956 : sel_778953;
  assign add_778960 = sel_778957 + 8'h01;
  assign sel_778961 = array_index_778612 == array_index_773158 ? add_778960 : sel_778957;
  assign add_778964 = sel_778961 + 8'h01;
  assign sel_778965 = array_index_778612 == array_index_773164 ? add_778964 : sel_778961;
  assign add_778968 = sel_778965 + 8'h01;
  assign sel_778969 = array_index_778612 == array_index_773170 ? add_778968 : sel_778965;
  assign add_778973 = sel_778969 + 8'h01;
  assign array_index_778974 = set1_unflattened[7'h11];
  assign sel_778975 = array_index_778612 == array_index_773176 ? add_778973 : sel_778969;
  assign add_778978 = sel_778975 + 8'h01;
  assign sel_778979 = array_index_778974 == array_index_772632 ? add_778978 : sel_778975;
  assign add_778982 = sel_778979 + 8'h01;
  assign sel_778983 = array_index_778974 == array_index_772636 ? add_778982 : sel_778979;
  assign add_778986 = sel_778983 + 8'h01;
  assign sel_778987 = array_index_778974 == array_index_772644 ? add_778986 : sel_778983;
  assign add_778990 = sel_778987 + 8'h01;
  assign sel_778991 = array_index_778974 == array_index_772652 ? add_778990 : sel_778987;
  assign add_778994 = sel_778991 + 8'h01;
  assign sel_778995 = array_index_778974 == array_index_772660 ? add_778994 : sel_778991;
  assign add_778998 = sel_778995 + 8'h01;
  assign sel_778999 = array_index_778974 == array_index_772668 ? add_778998 : sel_778995;
  assign add_779002 = sel_778999 + 8'h01;
  assign sel_779003 = array_index_778974 == array_index_772676 ? add_779002 : sel_778999;
  assign add_779006 = sel_779003 + 8'h01;
  assign sel_779007 = array_index_778974 == array_index_772684 ? add_779006 : sel_779003;
  assign add_779010 = sel_779007 + 8'h01;
  assign sel_779011 = array_index_778974 == array_index_772690 ? add_779010 : sel_779007;
  assign add_779014 = sel_779011 + 8'h01;
  assign sel_779015 = array_index_778974 == array_index_772696 ? add_779014 : sel_779011;
  assign add_779018 = sel_779015 + 8'h01;
  assign sel_779019 = array_index_778974 == array_index_772702 ? add_779018 : sel_779015;
  assign add_779022 = sel_779019 + 8'h01;
  assign sel_779023 = array_index_778974 == array_index_772708 ? add_779022 : sel_779019;
  assign add_779026 = sel_779023 + 8'h01;
  assign sel_779027 = array_index_778974 == array_index_772714 ? add_779026 : sel_779023;
  assign add_779030 = sel_779027 + 8'h01;
  assign sel_779031 = array_index_778974 == array_index_772720 ? add_779030 : sel_779027;
  assign add_779034 = sel_779031 + 8'h01;
  assign sel_779035 = array_index_778974 == array_index_772726 ? add_779034 : sel_779031;
  assign add_779038 = sel_779035 + 8'h01;
  assign sel_779039 = array_index_778974 == array_index_772732 ? add_779038 : sel_779035;
  assign add_779042 = sel_779039 + 8'h01;
  assign sel_779043 = array_index_778974 == array_index_772738 ? add_779042 : sel_779039;
  assign add_779046 = sel_779043 + 8'h01;
  assign sel_779047 = array_index_778974 == array_index_772744 ? add_779046 : sel_779043;
  assign add_779050 = sel_779047 + 8'h01;
  assign sel_779051 = array_index_778974 == array_index_772750 ? add_779050 : sel_779047;
  assign add_779054 = sel_779051 + 8'h01;
  assign sel_779055 = array_index_778974 == array_index_772756 ? add_779054 : sel_779051;
  assign add_779058 = sel_779055 + 8'h01;
  assign sel_779059 = array_index_778974 == array_index_772762 ? add_779058 : sel_779055;
  assign add_779062 = sel_779059 + 8'h01;
  assign sel_779063 = array_index_778974 == array_index_772768 ? add_779062 : sel_779059;
  assign add_779066 = sel_779063 + 8'h01;
  assign sel_779067 = array_index_778974 == array_index_772774 ? add_779066 : sel_779063;
  assign add_779070 = sel_779067 + 8'h01;
  assign sel_779071 = array_index_778974 == array_index_772780 ? add_779070 : sel_779067;
  assign add_779074 = sel_779071 + 8'h01;
  assign sel_779075 = array_index_778974 == array_index_772786 ? add_779074 : sel_779071;
  assign add_779078 = sel_779075 + 8'h01;
  assign sel_779079 = array_index_778974 == array_index_772792 ? add_779078 : sel_779075;
  assign add_779082 = sel_779079 + 8'h01;
  assign sel_779083 = array_index_778974 == array_index_772798 ? add_779082 : sel_779079;
  assign add_779086 = sel_779083 + 8'h01;
  assign sel_779087 = array_index_778974 == array_index_772804 ? add_779086 : sel_779083;
  assign add_779090 = sel_779087 + 8'h01;
  assign sel_779091 = array_index_778974 == array_index_772810 ? add_779090 : sel_779087;
  assign add_779094 = sel_779091 + 8'h01;
  assign sel_779095 = array_index_778974 == array_index_772816 ? add_779094 : sel_779091;
  assign add_779098 = sel_779095 + 8'h01;
  assign sel_779099 = array_index_778974 == array_index_772822 ? add_779098 : sel_779095;
  assign add_779102 = sel_779099 + 8'h01;
  assign sel_779103 = array_index_778974 == array_index_772828 ? add_779102 : sel_779099;
  assign add_779106 = sel_779103 + 8'h01;
  assign sel_779107 = array_index_778974 == array_index_772834 ? add_779106 : sel_779103;
  assign add_779110 = sel_779107 + 8'h01;
  assign sel_779111 = array_index_778974 == array_index_772840 ? add_779110 : sel_779107;
  assign add_779114 = sel_779111 + 8'h01;
  assign sel_779115 = array_index_778974 == array_index_772846 ? add_779114 : sel_779111;
  assign add_779118 = sel_779115 + 8'h01;
  assign sel_779119 = array_index_778974 == array_index_772852 ? add_779118 : sel_779115;
  assign add_779122 = sel_779119 + 8'h01;
  assign sel_779123 = array_index_778974 == array_index_772858 ? add_779122 : sel_779119;
  assign add_779126 = sel_779123 + 8'h01;
  assign sel_779127 = array_index_778974 == array_index_772864 ? add_779126 : sel_779123;
  assign add_779130 = sel_779127 + 8'h01;
  assign sel_779131 = array_index_778974 == array_index_772870 ? add_779130 : sel_779127;
  assign add_779134 = sel_779131 + 8'h01;
  assign sel_779135 = array_index_778974 == array_index_772876 ? add_779134 : sel_779131;
  assign add_779138 = sel_779135 + 8'h01;
  assign sel_779139 = array_index_778974 == array_index_772882 ? add_779138 : sel_779135;
  assign add_779142 = sel_779139 + 8'h01;
  assign sel_779143 = array_index_778974 == array_index_772888 ? add_779142 : sel_779139;
  assign add_779146 = sel_779143 + 8'h01;
  assign sel_779147 = array_index_778974 == array_index_772894 ? add_779146 : sel_779143;
  assign add_779150 = sel_779147 + 8'h01;
  assign sel_779151 = array_index_778974 == array_index_772900 ? add_779150 : sel_779147;
  assign add_779154 = sel_779151 + 8'h01;
  assign sel_779155 = array_index_778974 == array_index_772906 ? add_779154 : sel_779151;
  assign add_779158 = sel_779155 + 8'h01;
  assign sel_779159 = array_index_778974 == array_index_772912 ? add_779158 : sel_779155;
  assign add_779162 = sel_779159 + 8'h01;
  assign sel_779163 = array_index_778974 == array_index_772918 ? add_779162 : sel_779159;
  assign add_779166 = sel_779163 + 8'h01;
  assign sel_779167 = array_index_778974 == array_index_772924 ? add_779166 : sel_779163;
  assign add_779170 = sel_779167 + 8'h01;
  assign sel_779171 = array_index_778974 == array_index_772930 ? add_779170 : sel_779167;
  assign add_779174 = sel_779171 + 8'h01;
  assign sel_779175 = array_index_778974 == array_index_772936 ? add_779174 : sel_779171;
  assign add_779178 = sel_779175 + 8'h01;
  assign sel_779179 = array_index_778974 == array_index_772942 ? add_779178 : sel_779175;
  assign add_779182 = sel_779179 + 8'h01;
  assign sel_779183 = array_index_778974 == array_index_772948 ? add_779182 : sel_779179;
  assign add_779186 = sel_779183 + 8'h01;
  assign sel_779187 = array_index_778974 == array_index_772954 ? add_779186 : sel_779183;
  assign add_779190 = sel_779187 + 8'h01;
  assign sel_779191 = array_index_778974 == array_index_772960 ? add_779190 : sel_779187;
  assign add_779194 = sel_779191 + 8'h01;
  assign sel_779195 = array_index_778974 == array_index_772966 ? add_779194 : sel_779191;
  assign add_779198 = sel_779195 + 8'h01;
  assign sel_779199 = array_index_778974 == array_index_772972 ? add_779198 : sel_779195;
  assign add_779202 = sel_779199 + 8'h01;
  assign sel_779203 = array_index_778974 == array_index_772978 ? add_779202 : sel_779199;
  assign add_779206 = sel_779203 + 8'h01;
  assign sel_779207 = array_index_778974 == array_index_772984 ? add_779206 : sel_779203;
  assign add_779210 = sel_779207 + 8'h01;
  assign sel_779211 = array_index_778974 == array_index_772990 ? add_779210 : sel_779207;
  assign add_779214 = sel_779211 + 8'h01;
  assign sel_779215 = array_index_778974 == array_index_772996 ? add_779214 : sel_779211;
  assign add_779218 = sel_779215 + 8'h01;
  assign sel_779219 = array_index_778974 == array_index_773002 ? add_779218 : sel_779215;
  assign add_779222 = sel_779219 + 8'h01;
  assign sel_779223 = array_index_778974 == array_index_773008 ? add_779222 : sel_779219;
  assign add_779226 = sel_779223 + 8'h01;
  assign sel_779227 = array_index_778974 == array_index_773014 ? add_779226 : sel_779223;
  assign add_779230 = sel_779227 + 8'h01;
  assign sel_779231 = array_index_778974 == array_index_773020 ? add_779230 : sel_779227;
  assign add_779234 = sel_779231 + 8'h01;
  assign sel_779235 = array_index_778974 == array_index_773026 ? add_779234 : sel_779231;
  assign add_779238 = sel_779235 + 8'h01;
  assign sel_779239 = array_index_778974 == array_index_773032 ? add_779238 : sel_779235;
  assign add_779242 = sel_779239 + 8'h01;
  assign sel_779243 = array_index_778974 == array_index_773038 ? add_779242 : sel_779239;
  assign add_779246 = sel_779243 + 8'h01;
  assign sel_779247 = array_index_778974 == array_index_773044 ? add_779246 : sel_779243;
  assign add_779250 = sel_779247 + 8'h01;
  assign sel_779251 = array_index_778974 == array_index_773050 ? add_779250 : sel_779247;
  assign add_779254 = sel_779251 + 8'h01;
  assign sel_779255 = array_index_778974 == array_index_773056 ? add_779254 : sel_779251;
  assign add_779258 = sel_779255 + 8'h01;
  assign sel_779259 = array_index_778974 == array_index_773062 ? add_779258 : sel_779255;
  assign add_779262 = sel_779259 + 8'h01;
  assign sel_779263 = array_index_778974 == array_index_773068 ? add_779262 : sel_779259;
  assign add_779266 = sel_779263 + 8'h01;
  assign sel_779267 = array_index_778974 == array_index_773074 ? add_779266 : sel_779263;
  assign add_779270 = sel_779267 + 8'h01;
  assign sel_779271 = array_index_778974 == array_index_773080 ? add_779270 : sel_779267;
  assign add_779274 = sel_779271 + 8'h01;
  assign sel_779275 = array_index_778974 == array_index_773086 ? add_779274 : sel_779271;
  assign add_779278 = sel_779275 + 8'h01;
  assign sel_779279 = array_index_778974 == array_index_773092 ? add_779278 : sel_779275;
  assign add_779282 = sel_779279 + 8'h01;
  assign sel_779283 = array_index_778974 == array_index_773098 ? add_779282 : sel_779279;
  assign add_779286 = sel_779283 + 8'h01;
  assign sel_779287 = array_index_778974 == array_index_773104 ? add_779286 : sel_779283;
  assign add_779290 = sel_779287 + 8'h01;
  assign sel_779291 = array_index_778974 == array_index_773110 ? add_779290 : sel_779287;
  assign add_779294 = sel_779291 + 8'h01;
  assign sel_779295 = array_index_778974 == array_index_773116 ? add_779294 : sel_779291;
  assign add_779298 = sel_779295 + 8'h01;
  assign sel_779299 = array_index_778974 == array_index_773122 ? add_779298 : sel_779295;
  assign add_779302 = sel_779299 + 8'h01;
  assign sel_779303 = array_index_778974 == array_index_773128 ? add_779302 : sel_779299;
  assign add_779306 = sel_779303 + 8'h01;
  assign sel_779307 = array_index_778974 == array_index_773134 ? add_779306 : sel_779303;
  assign add_779310 = sel_779307 + 8'h01;
  assign sel_779311 = array_index_778974 == array_index_773140 ? add_779310 : sel_779307;
  assign add_779314 = sel_779311 + 8'h01;
  assign sel_779315 = array_index_778974 == array_index_773146 ? add_779314 : sel_779311;
  assign add_779318 = sel_779315 + 8'h01;
  assign sel_779319 = array_index_778974 == array_index_773152 ? add_779318 : sel_779315;
  assign add_779322 = sel_779319 + 8'h01;
  assign sel_779323 = array_index_778974 == array_index_773158 ? add_779322 : sel_779319;
  assign add_779326 = sel_779323 + 8'h01;
  assign sel_779327 = array_index_778974 == array_index_773164 ? add_779326 : sel_779323;
  assign add_779330 = sel_779327 + 8'h01;
  assign sel_779331 = array_index_778974 == array_index_773170 ? add_779330 : sel_779327;
  assign add_779335 = sel_779331 + 8'h01;
  assign array_index_779336 = set1_unflattened[7'h12];
  assign sel_779337 = array_index_778974 == array_index_773176 ? add_779335 : sel_779331;
  assign add_779340 = sel_779337 + 8'h01;
  assign sel_779341 = array_index_779336 == array_index_772632 ? add_779340 : sel_779337;
  assign add_779344 = sel_779341 + 8'h01;
  assign sel_779345 = array_index_779336 == array_index_772636 ? add_779344 : sel_779341;
  assign add_779348 = sel_779345 + 8'h01;
  assign sel_779349 = array_index_779336 == array_index_772644 ? add_779348 : sel_779345;
  assign add_779352 = sel_779349 + 8'h01;
  assign sel_779353 = array_index_779336 == array_index_772652 ? add_779352 : sel_779349;
  assign add_779356 = sel_779353 + 8'h01;
  assign sel_779357 = array_index_779336 == array_index_772660 ? add_779356 : sel_779353;
  assign add_779360 = sel_779357 + 8'h01;
  assign sel_779361 = array_index_779336 == array_index_772668 ? add_779360 : sel_779357;
  assign add_779364 = sel_779361 + 8'h01;
  assign sel_779365 = array_index_779336 == array_index_772676 ? add_779364 : sel_779361;
  assign add_779368 = sel_779365 + 8'h01;
  assign sel_779369 = array_index_779336 == array_index_772684 ? add_779368 : sel_779365;
  assign add_779372 = sel_779369 + 8'h01;
  assign sel_779373 = array_index_779336 == array_index_772690 ? add_779372 : sel_779369;
  assign add_779376 = sel_779373 + 8'h01;
  assign sel_779377 = array_index_779336 == array_index_772696 ? add_779376 : sel_779373;
  assign add_779380 = sel_779377 + 8'h01;
  assign sel_779381 = array_index_779336 == array_index_772702 ? add_779380 : sel_779377;
  assign add_779384 = sel_779381 + 8'h01;
  assign sel_779385 = array_index_779336 == array_index_772708 ? add_779384 : sel_779381;
  assign add_779388 = sel_779385 + 8'h01;
  assign sel_779389 = array_index_779336 == array_index_772714 ? add_779388 : sel_779385;
  assign add_779392 = sel_779389 + 8'h01;
  assign sel_779393 = array_index_779336 == array_index_772720 ? add_779392 : sel_779389;
  assign add_779396 = sel_779393 + 8'h01;
  assign sel_779397 = array_index_779336 == array_index_772726 ? add_779396 : sel_779393;
  assign add_779400 = sel_779397 + 8'h01;
  assign sel_779401 = array_index_779336 == array_index_772732 ? add_779400 : sel_779397;
  assign add_779404 = sel_779401 + 8'h01;
  assign sel_779405 = array_index_779336 == array_index_772738 ? add_779404 : sel_779401;
  assign add_779408 = sel_779405 + 8'h01;
  assign sel_779409 = array_index_779336 == array_index_772744 ? add_779408 : sel_779405;
  assign add_779412 = sel_779409 + 8'h01;
  assign sel_779413 = array_index_779336 == array_index_772750 ? add_779412 : sel_779409;
  assign add_779416 = sel_779413 + 8'h01;
  assign sel_779417 = array_index_779336 == array_index_772756 ? add_779416 : sel_779413;
  assign add_779420 = sel_779417 + 8'h01;
  assign sel_779421 = array_index_779336 == array_index_772762 ? add_779420 : sel_779417;
  assign add_779424 = sel_779421 + 8'h01;
  assign sel_779425 = array_index_779336 == array_index_772768 ? add_779424 : sel_779421;
  assign add_779428 = sel_779425 + 8'h01;
  assign sel_779429 = array_index_779336 == array_index_772774 ? add_779428 : sel_779425;
  assign add_779432 = sel_779429 + 8'h01;
  assign sel_779433 = array_index_779336 == array_index_772780 ? add_779432 : sel_779429;
  assign add_779436 = sel_779433 + 8'h01;
  assign sel_779437 = array_index_779336 == array_index_772786 ? add_779436 : sel_779433;
  assign add_779440 = sel_779437 + 8'h01;
  assign sel_779441 = array_index_779336 == array_index_772792 ? add_779440 : sel_779437;
  assign add_779444 = sel_779441 + 8'h01;
  assign sel_779445 = array_index_779336 == array_index_772798 ? add_779444 : sel_779441;
  assign add_779448 = sel_779445 + 8'h01;
  assign sel_779449 = array_index_779336 == array_index_772804 ? add_779448 : sel_779445;
  assign add_779452 = sel_779449 + 8'h01;
  assign sel_779453 = array_index_779336 == array_index_772810 ? add_779452 : sel_779449;
  assign add_779456 = sel_779453 + 8'h01;
  assign sel_779457 = array_index_779336 == array_index_772816 ? add_779456 : sel_779453;
  assign add_779460 = sel_779457 + 8'h01;
  assign sel_779461 = array_index_779336 == array_index_772822 ? add_779460 : sel_779457;
  assign add_779464 = sel_779461 + 8'h01;
  assign sel_779465 = array_index_779336 == array_index_772828 ? add_779464 : sel_779461;
  assign add_779468 = sel_779465 + 8'h01;
  assign sel_779469 = array_index_779336 == array_index_772834 ? add_779468 : sel_779465;
  assign add_779472 = sel_779469 + 8'h01;
  assign sel_779473 = array_index_779336 == array_index_772840 ? add_779472 : sel_779469;
  assign add_779476 = sel_779473 + 8'h01;
  assign sel_779477 = array_index_779336 == array_index_772846 ? add_779476 : sel_779473;
  assign add_779480 = sel_779477 + 8'h01;
  assign sel_779481 = array_index_779336 == array_index_772852 ? add_779480 : sel_779477;
  assign add_779484 = sel_779481 + 8'h01;
  assign sel_779485 = array_index_779336 == array_index_772858 ? add_779484 : sel_779481;
  assign add_779488 = sel_779485 + 8'h01;
  assign sel_779489 = array_index_779336 == array_index_772864 ? add_779488 : sel_779485;
  assign add_779492 = sel_779489 + 8'h01;
  assign sel_779493 = array_index_779336 == array_index_772870 ? add_779492 : sel_779489;
  assign add_779496 = sel_779493 + 8'h01;
  assign sel_779497 = array_index_779336 == array_index_772876 ? add_779496 : sel_779493;
  assign add_779500 = sel_779497 + 8'h01;
  assign sel_779501 = array_index_779336 == array_index_772882 ? add_779500 : sel_779497;
  assign add_779504 = sel_779501 + 8'h01;
  assign sel_779505 = array_index_779336 == array_index_772888 ? add_779504 : sel_779501;
  assign add_779508 = sel_779505 + 8'h01;
  assign sel_779509 = array_index_779336 == array_index_772894 ? add_779508 : sel_779505;
  assign add_779512 = sel_779509 + 8'h01;
  assign sel_779513 = array_index_779336 == array_index_772900 ? add_779512 : sel_779509;
  assign add_779516 = sel_779513 + 8'h01;
  assign sel_779517 = array_index_779336 == array_index_772906 ? add_779516 : sel_779513;
  assign add_779520 = sel_779517 + 8'h01;
  assign sel_779521 = array_index_779336 == array_index_772912 ? add_779520 : sel_779517;
  assign add_779524 = sel_779521 + 8'h01;
  assign sel_779525 = array_index_779336 == array_index_772918 ? add_779524 : sel_779521;
  assign add_779528 = sel_779525 + 8'h01;
  assign sel_779529 = array_index_779336 == array_index_772924 ? add_779528 : sel_779525;
  assign add_779532 = sel_779529 + 8'h01;
  assign sel_779533 = array_index_779336 == array_index_772930 ? add_779532 : sel_779529;
  assign add_779536 = sel_779533 + 8'h01;
  assign sel_779537 = array_index_779336 == array_index_772936 ? add_779536 : sel_779533;
  assign add_779540 = sel_779537 + 8'h01;
  assign sel_779541 = array_index_779336 == array_index_772942 ? add_779540 : sel_779537;
  assign add_779544 = sel_779541 + 8'h01;
  assign sel_779545 = array_index_779336 == array_index_772948 ? add_779544 : sel_779541;
  assign add_779548 = sel_779545 + 8'h01;
  assign sel_779549 = array_index_779336 == array_index_772954 ? add_779548 : sel_779545;
  assign add_779552 = sel_779549 + 8'h01;
  assign sel_779553 = array_index_779336 == array_index_772960 ? add_779552 : sel_779549;
  assign add_779556 = sel_779553 + 8'h01;
  assign sel_779557 = array_index_779336 == array_index_772966 ? add_779556 : sel_779553;
  assign add_779560 = sel_779557 + 8'h01;
  assign sel_779561 = array_index_779336 == array_index_772972 ? add_779560 : sel_779557;
  assign add_779564 = sel_779561 + 8'h01;
  assign sel_779565 = array_index_779336 == array_index_772978 ? add_779564 : sel_779561;
  assign add_779568 = sel_779565 + 8'h01;
  assign sel_779569 = array_index_779336 == array_index_772984 ? add_779568 : sel_779565;
  assign add_779572 = sel_779569 + 8'h01;
  assign sel_779573 = array_index_779336 == array_index_772990 ? add_779572 : sel_779569;
  assign add_779576 = sel_779573 + 8'h01;
  assign sel_779577 = array_index_779336 == array_index_772996 ? add_779576 : sel_779573;
  assign add_779580 = sel_779577 + 8'h01;
  assign sel_779581 = array_index_779336 == array_index_773002 ? add_779580 : sel_779577;
  assign add_779584 = sel_779581 + 8'h01;
  assign sel_779585 = array_index_779336 == array_index_773008 ? add_779584 : sel_779581;
  assign add_779588 = sel_779585 + 8'h01;
  assign sel_779589 = array_index_779336 == array_index_773014 ? add_779588 : sel_779585;
  assign add_779592 = sel_779589 + 8'h01;
  assign sel_779593 = array_index_779336 == array_index_773020 ? add_779592 : sel_779589;
  assign add_779596 = sel_779593 + 8'h01;
  assign sel_779597 = array_index_779336 == array_index_773026 ? add_779596 : sel_779593;
  assign add_779600 = sel_779597 + 8'h01;
  assign sel_779601 = array_index_779336 == array_index_773032 ? add_779600 : sel_779597;
  assign add_779604 = sel_779601 + 8'h01;
  assign sel_779605 = array_index_779336 == array_index_773038 ? add_779604 : sel_779601;
  assign add_779608 = sel_779605 + 8'h01;
  assign sel_779609 = array_index_779336 == array_index_773044 ? add_779608 : sel_779605;
  assign add_779612 = sel_779609 + 8'h01;
  assign sel_779613 = array_index_779336 == array_index_773050 ? add_779612 : sel_779609;
  assign add_779616 = sel_779613 + 8'h01;
  assign sel_779617 = array_index_779336 == array_index_773056 ? add_779616 : sel_779613;
  assign add_779620 = sel_779617 + 8'h01;
  assign sel_779621 = array_index_779336 == array_index_773062 ? add_779620 : sel_779617;
  assign add_779624 = sel_779621 + 8'h01;
  assign sel_779625 = array_index_779336 == array_index_773068 ? add_779624 : sel_779621;
  assign add_779628 = sel_779625 + 8'h01;
  assign sel_779629 = array_index_779336 == array_index_773074 ? add_779628 : sel_779625;
  assign add_779632 = sel_779629 + 8'h01;
  assign sel_779633 = array_index_779336 == array_index_773080 ? add_779632 : sel_779629;
  assign add_779636 = sel_779633 + 8'h01;
  assign sel_779637 = array_index_779336 == array_index_773086 ? add_779636 : sel_779633;
  assign add_779640 = sel_779637 + 8'h01;
  assign sel_779641 = array_index_779336 == array_index_773092 ? add_779640 : sel_779637;
  assign add_779644 = sel_779641 + 8'h01;
  assign sel_779645 = array_index_779336 == array_index_773098 ? add_779644 : sel_779641;
  assign add_779648 = sel_779645 + 8'h01;
  assign sel_779649 = array_index_779336 == array_index_773104 ? add_779648 : sel_779645;
  assign add_779652 = sel_779649 + 8'h01;
  assign sel_779653 = array_index_779336 == array_index_773110 ? add_779652 : sel_779649;
  assign add_779656 = sel_779653 + 8'h01;
  assign sel_779657 = array_index_779336 == array_index_773116 ? add_779656 : sel_779653;
  assign add_779660 = sel_779657 + 8'h01;
  assign sel_779661 = array_index_779336 == array_index_773122 ? add_779660 : sel_779657;
  assign add_779664 = sel_779661 + 8'h01;
  assign sel_779665 = array_index_779336 == array_index_773128 ? add_779664 : sel_779661;
  assign add_779668 = sel_779665 + 8'h01;
  assign sel_779669 = array_index_779336 == array_index_773134 ? add_779668 : sel_779665;
  assign add_779672 = sel_779669 + 8'h01;
  assign sel_779673 = array_index_779336 == array_index_773140 ? add_779672 : sel_779669;
  assign add_779676 = sel_779673 + 8'h01;
  assign sel_779677 = array_index_779336 == array_index_773146 ? add_779676 : sel_779673;
  assign add_779680 = sel_779677 + 8'h01;
  assign sel_779681 = array_index_779336 == array_index_773152 ? add_779680 : sel_779677;
  assign add_779684 = sel_779681 + 8'h01;
  assign sel_779685 = array_index_779336 == array_index_773158 ? add_779684 : sel_779681;
  assign add_779688 = sel_779685 + 8'h01;
  assign sel_779689 = array_index_779336 == array_index_773164 ? add_779688 : sel_779685;
  assign add_779692 = sel_779689 + 8'h01;
  assign sel_779693 = array_index_779336 == array_index_773170 ? add_779692 : sel_779689;
  assign add_779697 = sel_779693 + 8'h01;
  assign array_index_779698 = set1_unflattened[7'h13];
  assign sel_779699 = array_index_779336 == array_index_773176 ? add_779697 : sel_779693;
  assign add_779702 = sel_779699 + 8'h01;
  assign sel_779703 = array_index_779698 == array_index_772632 ? add_779702 : sel_779699;
  assign add_779706 = sel_779703 + 8'h01;
  assign sel_779707 = array_index_779698 == array_index_772636 ? add_779706 : sel_779703;
  assign add_779710 = sel_779707 + 8'h01;
  assign sel_779711 = array_index_779698 == array_index_772644 ? add_779710 : sel_779707;
  assign add_779714 = sel_779711 + 8'h01;
  assign sel_779715 = array_index_779698 == array_index_772652 ? add_779714 : sel_779711;
  assign add_779718 = sel_779715 + 8'h01;
  assign sel_779719 = array_index_779698 == array_index_772660 ? add_779718 : sel_779715;
  assign add_779722 = sel_779719 + 8'h01;
  assign sel_779723 = array_index_779698 == array_index_772668 ? add_779722 : sel_779719;
  assign add_779726 = sel_779723 + 8'h01;
  assign sel_779727 = array_index_779698 == array_index_772676 ? add_779726 : sel_779723;
  assign add_779730 = sel_779727 + 8'h01;
  assign sel_779731 = array_index_779698 == array_index_772684 ? add_779730 : sel_779727;
  assign add_779734 = sel_779731 + 8'h01;
  assign sel_779735 = array_index_779698 == array_index_772690 ? add_779734 : sel_779731;
  assign add_779738 = sel_779735 + 8'h01;
  assign sel_779739 = array_index_779698 == array_index_772696 ? add_779738 : sel_779735;
  assign add_779742 = sel_779739 + 8'h01;
  assign sel_779743 = array_index_779698 == array_index_772702 ? add_779742 : sel_779739;
  assign add_779746 = sel_779743 + 8'h01;
  assign sel_779747 = array_index_779698 == array_index_772708 ? add_779746 : sel_779743;
  assign add_779750 = sel_779747 + 8'h01;
  assign sel_779751 = array_index_779698 == array_index_772714 ? add_779750 : sel_779747;
  assign add_779754 = sel_779751 + 8'h01;
  assign sel_779755 = array_index_779698 == array_index_772720 ? add_779754 : sel_779751;
  assign add_779758 = sel_779755 + 8'h01;
  assign sel_779759 = array_index_779698 == array_index_772726 ? add_779758 : sel_779755;
  assign add_779762 = sel_779759 + 8'h01;
  assign sel_779763 = array_index_779698 == array_index_772732 ? add_779762 : sel_779759;
  assign add_779766 = sel_779763 + 8'h01;
  assign sel_779767 = array_index_779698 == array_index_772738 ? add_779766 : sel_779763;
  assign add_779770 = sel_779767 + 8'h01;
  assign sel_779771 = array_index_779698 == array_index_772744 ? add_779770 : sel_779767;
  assign add_779774 = sel_779771 + 8'h01;
  assign sel_779775 = array_index_779698 == array_index_772750 ? add_779774 : sel_779771;
  assign add_779778 = sel_779775 + 8'h01;
  assign sel_779779 = array_index_779698 == array_index_772756 ? add_779778 : sel_779775;
  assign add_779782 = sel_779779 + 8'h01;
  assign sel_779783 = array_index_779698 == array_index_772762 ? add_779782 : sel_779779;
  assign add_779786 = sel_779783 + 8'h01;
  assign sel_779787 = array_index_779698 == array_index_772768 ? add_779786 : sel_779783;
  assign add_779790 = sel_779787 + 8'h01;
  assign sel_779791 = array_index_779698 == array_index_772774 ? add_779790 : sel_779787;
  assign add_779794 = sel_779791 + 8'h01;
  assign sel_779795 = array_index_779698 == array_index_772780 ? add_779794 : sel_779791;
  assign add_779798 = sel_779795 + 8'h01;
  assign sel_779799 = array_index_779698 == array_index_772786 ? add_779798 : sel_779795;
  assign add_779802 = sel_779799 + 8'h01;
  assign sel_779803 = array_index_779698 == array_index_772792 ? add_779802 : sel_779799;
  assign add_779806 = sel_779803 + 8'h01;
  assign sel_779807 = array_index_779698 == array_index_772798 ? add_779806 : sel_779803;
  assign add_779810 = sel_779807 + 8'h01;
  assign sel_779811 = array_index_779698 == array_index_772804 ? add_779810 : sel_779807;
  assign add_779814 = sel_779811 + 8'h01;
  assign sel_779815 = array_index_779698 == array_index_772810 ? add_779814 : sel_779811;
  assign add_779818 = sel_779815 + 8'h01;
  assign sel_779819 = array_index_779698 == array_index_772816 ? add_779818 : sel_779815;
  assign add_779822 = sel_779819 + 8'h01;
  assign sel_779823 = array_index_779698 == array_index_772822 ? add_779822 : sel_779819;
  assign add_779826 = sel_779823 + 8'h01;
  assign sel_779827 = array_index_779698 == array_index_772828 ? add_779826 : sel_779823;
  assign add_779830 = sel_779827 + 8'h01;
  assign sel_779831 = array_index_779698 == array_index_772834 ? add_779830 : sel_779827;
  assign add_779834 = sel_779831 + 8'h01;
  assign sel_779835 = array_index_779698 == array_index_772840 ? add_779834 : sel_779831;
  assign add_779838 = sel_779835 + 8'h01;
  assign sel_779839 = array_index_779698 == array_index_772846 ? add_779838 : sel_779835;
  assign add_779842 = sel_779839 + 8'h01;
  assign sel_779843 = array_index_779698 == array_index_772852 ? add_779842 : sel_779839;
  assign add_779846 = sel_779843 + 8'h01;
  assign sel_779847 = array_index_779698 == array_index_772858 ? add_779846 : sel_779843;
  assign add_779850 = sel_779847 + 8'h01;
  assign sel_779851 = array_index_779698 == array_index_772864 ? add_779850 : sel_779847;
  assign add_779854 = sel_779851 + 8'h01;
  assign sel_779855 = array_index_779698 == array_index_772870 ? add_779854 : sel_779851;
  assign add_779858 = sel_779855 + 8'h01;
  assign sel_779859 = array_index_779698 == array_index_772876 ? add_779858 : sel_779855;
  assign add_779862 = sel_779859 + 8'h01;
  assign sel_779863 = array_index_779698 == array_index_772882 ? add_779862 : sel_779859;
  assign add_779866 = sel_779863 + 8'h01;
  assign sel_779867 = array_index_779698 == array_index_772888 ? add_779866 : sel_779863;
  assign add_779870 = sel_779867 + 8'h01;
  assign sel_779871 = array_index_779698 == array_index_772894 ? add_779870 : sel_779867;
  assign add_779874 = sel_779871 + 8'h01;
  assign sel_779875 = array_index_779698 == array_index_772900 ? add_779874 : sel_779871;
  assign add_779878 = sel_779875 + 8'h01;
  assign sel_779879 = array_index_779698 == array_index_772906 ? add_779878 : sel_779875;
  assign add_779882 = sel_779879 + 8'h01;
  assign sel_779883 = array_index_779698 == array_index_772912 ? add_779882 : sel_779879;
  assign add_779886 = sel_779883 + 8'h01;
  assign sel_779887 = array_index_779698 == array_index_772918 ? add_779886 : sel_779883;
  assign add_779890 = sel_779887 + 8'h01;
  assign sel_779891 = array_index_779698 == array_index_772924 ? add_779890 : sel_779887;
  assign add_779894 = sel_779891 + 8'h01;
  assign sel_779895 = array_index_779698 == array_index_772930 ? add_779894 : sel_779891;
  assign add_779898 = sel_779895 + 8'h01;
  assign sel_779899 = array_index_779698 == array_index_772936 ? add_779898 : sel_779895;
  assign add_779902 = sel_779899 + 8'h01;
  assign sel_779903 = array_index_779698 == array_index_772942 ? add_779902 : sel_779899;
  assign add_779906 = sel_779903 + 8'h01;
  assign sel_779907 = array_index_779698 == array_index_772948 ? add_779906 : sel_779903;
  assign add_779910 = sel_779907 + 8'h01;
  assign sel_779911 = array_index_779698 == array_index_772954 ? add_779910 : sel_779907;
  assign add_779914 = sel_779911 + 8'h01;
  assign sel_779915 = array_index_779698 == array_index_772960 ? add_779914 : sel_779911;
  assign add_779918 = sel_779915 + 8'h01;
  assign sel_779919 = array_index_779698 == array_index_772966 ? add_779918 : sel_779915;
  assign add_779922 = sel_779919 + 8'h01;
  assign sel_779923 = array_index_779698 == array_index_772972 ? add_779922 : sel_779919;
  assign add_779926 = sel_779923 + 8'h01;
  assign sel_779927 = array_index_779698 == array_index_772978 ? add_779926 : sel_779923;
  assign add_779930 = sel_779927 + 8'h01;
  assign sel_779931 = array_index_779698 == array_index_772984 ? add_779930 : sel_779927;
  assign add_779934 = sel_779931 + 8'h01;
  assign sel_779935 = array_index_779698 == array_index_772990 ? add_779934 : sel_779931;
  assign add_779938 = sel_779935 + 8'h01;
  assign sel_779939 = array_index_779698 == array_index_772996 ? add_779938 : sel_779935;
  assign add_779942 = sel_779939 + 8'h01;
  assign sel_779943 = array_index_779698 == array_index_773002 ? add_779942 : sel_779939;
  assign add_779946 = sel_779943 + 8'h01;
  assign sel_779947 = array_index_779698 == array_index_773008 ? add_779946 : sel_779943;
  assign add_779950 = sel_779947 + 8'h01;
  assign sel_779951 = array_index_779698 == array_index_773014 ? add_779950 : sel_779947;
  assign add_779954 = sel_779951 + 8'h01;
  assign sel_779955 = array_index_779698 == array_index_773020 ? add_779954 : sel_779951;
  assign add_779958 = sel_779955 + 8'h01;
  assign sel_779959 = array_index_779698 == array_index_773026 ? add_779958 : sel_779955;
  assign add_779962 = sel_779959 + 8'h01;
  assign sel_779963 = array_index_779698 == array_index_773032 ? add_779962 : sel_779959;
  assign add_779966 = sel_779963 + 8'h01;
  assign sel_779967 = array_index_779698 == array_index_773038 ? add_779966 : sel_779963;
  assign add_779970 = sel_779967 + 8'h01;
  assign sel_779971 = array_index_779698 == array_index_773044 ? add_779970 : sel_779967;
  assign add_779974 = sel_779971 + 8'h01;
  assign sel_779975 = array_index_779698 == array_index_773050 ? add_779974 : sel_779971;
  assign add_779978 = sel_779975 + 8'h01;
  assign sel_779979 = array_index_779698 == array_index_773056 ? add_779978 : sel_779975;
  assign add_779982 = sel_779979 + 8'h01;
  assign sel_779983 = array_index_779698 == array_index_773062 ? add_779982 : sel_779979;
  assign add_779986 = sel_779983 + 8'h01;
  assign sel_779987 = array_index_779698 == array_index_773068 ? add_779986 : sel_779983;
  assign add_779990 = sel_779987 + 8'h01;
  assign sel_779991 = array_index_779698 == array_index_773074 ? add_779990 : sel_779987;
  assign add_779994 = sel_779991 + 8'h01;
  assign sel_779995 = array_index_779698 == array_index_773080 ? add_779994 : sel_779991;
  assign add_779998 = sel_779995 + 8'h01;
  assign sel_779999 = array_index_779698 == array_index_773086 ? add_779998 : sel_779995;
  assign add_780002 = sel_779999 + 8'h01;
  assign sel_780003 = array_index_779698 == array_index_773092 ? add_780002 : sel_779999;
  assign add_780006 = sel_780003 + 8'h01;
  assign sel_780007 = array_index_779698 == array_index_773098 ? add_780006 : sel_780003;
  assign add_780010 = sel_780007 + 8'h01;
  assign sel_780011 = array_index_779698 == array_index_773104 ? add_780010 : sel_780007;
  assign add_780014 = sel_780011 + 8'h01;
  assign sel_780015 = array_index_779698 == array_index_773110 ? add_780014 : sel_780011;
  assign add_780018 = sel_780015 + 8'h01;
  assign sel_780019 = array_index_779698 == array_index_773116 ? add_780018 : sel_780015;
  assign add_780022 = sel_780019 + 8'h01;
  assign sel_780023 = array_index_779698 == array_index_773122 ? add_780022 : sel_780019;
  assign add_780026 = sel_780023 + 8'h01;
  assign sel_780027 = array_index_779698 == array_index_773128 ? add_780026 : sel_780023;
  assign add_780030 = sel_780027 + 8'h01;
  assign sel_780031 = array_index_779698 == array_index_773134 ? add_780030 : sel_780027;
  assign add_780034 = sel_780031 + 8'h01;
  assign sel_780035 = array_index_779698 == array_index_773140 ? add_780034 : sel_780031;
  assign add_780038 = sel_780035 + 8'h01;
  assign sel_780039 = array_index_779698 == array_index_773146 ? add_780038 : sel_780035;
  assign add_780042 = sel_780039 + 8'h01;
  assign sel_780043 = array_index_779698 == array_index_773152 ? add_780042 : sel_780039;
  assign add_780046 = sel_780043 + 8'h01;
  assign sel_780047 = array_index_779698 == array_index_773158 ? add_780046 : sel_780043;
  assign add_780050 = sel_780047 + 8'h01;
  assign sel_780051 = array_index_779698 == array_index_773164 ? add_780050 : sel_780047;
  assign add_780054 = sel_780051 + 8'h01;
  assign sel_780055 = array_index_779698 == array_index_773170 ? add_780054 : sel_780051;
  assign add_780059 = sel_780055 + 8'h01;
  assign array_index_780060 = set1_unflattened[7'h14];
  assign sel_780061 = array_index_779698 == array_index_773176 ? add_780059 : sel_780055;
  assign add_780064 = sel_780061 + 8'h01;
  assign sel_780065 = array_index_780060 == array_index_772632 ? add_780064 : sel_780061;
  assign add_780068 = sel_780065 + 8'h01;
  assign sel_780069 = array_index_780060 == array_index_772636 ? add_780068 : sel_780065;
  assign add_780072 = sel_780069 + 8'h01;
  assign sel_780073 = array_index_780060 == array_index_772644 ? add_780072 : sel_780069;
  assign add_780076 = sel_780073 + 8'h01;
  assign sel_780077 = array_index_780060 == array_index_772652 ? add_780076 : sel_780073;
  assign add_780080 = sel_780077 + 8'h01;
  assign sel_780081 = array_index_780060 == array_index_772660 ? add_780080 : sel_780077;
  assign add_780084 = sel_780081 + 8'h01;
  assign sel_780085 = array_index_780060 == array_index_772668 ? add_780084 : sel_780081;
  assign add_780088 = sel_780085 + 8'h01;
  assign sel_780089 = array_index_780060 == array_index_772676 ? add_780088 : sel_780085;
  assign add_780092 = sel_780089 + 8'h01;
  assign sel_780093 = array_index_780060 == array_index_772684 ? add_780092 : sel_780089;
  assign add_780096 = sel_780093 + 8'h01;
  assign sel_780097 = array_index_780060 == array_index_772690 ? add_780096 : sel_780093;
  assign add_780100 = sel_780097 + 8'h01;
  assign sel_780101 = array_index_780060 == array_index_772696 ? add_780100 : sel_780097;
  assign add_780104 = sel_780101 + 8'h01;
  assign sel_780105 = array_index_780060 == array_index_772702 ? add_780104 : sel_780101;
  assign add_780108 = sel_780105 + 8'h01;
  assign sel_780109 = array_index_780060 == array_index_772708 ? add_780108 : sel_780105;
  assign add_780112 = sel_780109 + 8'h01;
  assign sel_780113 = array_index_780060 == array_index_772714 ? add_780112 : sel_780109;
  assign add_780116 = sel_780113 + 8'h01;
  assign sel_780117 = array_index_780060 == array_index_772720 ? add_780116 : sel_780113;
  assign add_780120 = sel_780117 + 8'h01;
  assign sel_780121 = array_index_780060 == array_index_772726 ? add_780120 : sel_780117;
  assign add_780124 = sel_780121 + 8'h01;
  assign sel_780125 = array_index_780060 == array_index_772732 ? add_780124 : sel_780121;
  assign add_780128 = sel_780125 + 8'h01;
  assign sel_780129 = array_index_780060 == array_index_772738 ? add_780128 : sel_780125;
  assign add_780132 = sel_780129 + 8'h01;
  assign sel_780133 = array_index_780060 == array_index_772744 ? add_780132 : sel_780129;
  assign add_780136 = sel_780133 + 8'h01;
  assign sel_780137 = array_index_780060 == array_index_772750 ? add_780136 : sel_780133;
  assign add_780140 = sel_780137 + 8'h01;
  assign sel_780141 = array_index_780060 == array_index_772756 ? add_780140 : sel_780137;
  assign add_780144 = sel_780141 + 8'h01;
  assign sel_780145 = array_index_780060 == array_index_772762 ? add_780144 : sel_780141;
  assign add_780148 = sel_780145 + 8'h01;
  assign sel_780149 = array_index_780060 == array_index_772768 ? add_780148 : sel_780145;
  assign add_780152 = sel_780149 + 8'h01;
  assign sel_780153 = array_index_780060 == array_index_772774 ? add_780152 : sel_780149;
  assign add_780156 = sel_780153 + 8'h01;
  assign sel_780157 = array_index_780060 == array_index_772780 ? add_780156 : sel_780153;
  assign add_780160 = sel_780157 + 8'h01;
  assign sel_780161 = array_index_780060 == array_index_772786 ? add_780160 : sel_780157;
  assign add_780164 = sel_780161 + 8'h01;
  assign sel_780165 = array_index_780060 == array_index_772792 ? add_780164 : sel_780161;
  assign add_780168 = sel_780165 + 8'h01;
  assign sel_780169 = array_index_780060 == array_index_772798 ? add_780168 : sel_780165;
  assign add_780172 = sel_780169 + 8'h01;
  assign sel_780173 = array_index_780060 == array_index_772804 ? add_780172 : sel_780169;
  assign add_780176 = sel_780173 + 8'h01;
  assign sel_780177 = array_index_780060 == array_index_772810 ? add_780176 : sel_780173;
  assign add_780180 = sel_780177 + 8'h01;
  assign sel_780181 = array_index_780060 == array_index_772816 ? add_780180 : sel_780177;
  assign add_780184 = sel_780181 + 8'h01;
  assign sel_780185 = array_index_780060 == array_index_772822 ? add_780184 : sel_780181;
  assign add_780188 = sel_780185 + 8'h01;
  assign sel_780189 = array_index_780060 == array_index_772828 ? add_780188 : sel_780185;
  assign add_780192 = sel_780189 + 8'h01;
  assign sel_780193 = array_index_780060 == array_index_772834 ? add_780192 : sel_780189;
  assign add_780196 = sel_780193 + 8'h01;
  assign sel_780197 = array_index_780060 == array_index_772840 ? add_780196 : sel_780193;
  assign add_780200 = sel_780197 + 8'h01;
  assign sel_780201 = array_index_780060 == array_index_772846 ? add_780200 : sel_780197;
  assign add_780204 = sel_780201 + 8'h01;
  assign sel_780205 = array_index_780060 == array_index_772852 ? add_780204 : sel_780201;
  assign add_780208 = sel_780205 + 8'h01;
  assign sel_780209 = array_index_780060 == array_index_772858 ? add_780208 : sel_780205;
  assign add_780212 = sel_780209 + 8'h01;
  assign sel_780213 = array_index_780060 == array_index_772864 ? add_780212 : sel_780209;
  assign add_780216 = sel_780213 + 8'h01;
  assign sel_780217 = array_index_780060 == array_index_772870 ? add_780216 : sel_780213;
  assign add_780220 = sel_780217 + 8'h01;
  assign sel_780221 = array_index_780060 == array_index_772876 ? add_780220 : sel_780217;
  assign add_780224 = sel_780221 + 8'h01;
  assign sel_780225 = array_index_780060 == array_index_772882 ? add_780224 : sel_780221;
  assign add_780228 = sel_780225 + 8'h01;
  assign sel_780229 = array_index_780060 == array_index_772888 ? add_780228 : sel_780225;
  assign add_780232 = sel_780229 + 8'h01;
  assign sel_780233 = array_index_780060 == array_index_772894 ? add_780232 : sel_780229;
  assign add_780236 = sel_780233 + 8'h01;
  assign sel_780237 = array_index_780060 == array_index_772900 ? add_780236 : sel_780233;
  assign add_780240 = sel_780237 + 8'h01;
  assign sel_780241 = array_index_780060 == array_index_772906 ? add_780240 : sel_780237;
  assign add_780244 = sel_780241 + 8'h01;
  assign sel_780245 = array_index_780060 == array_index_772912 ? add_780244 : sel_780241;
  assign add_780248 = sel_780245 + 8'h01;
  assign sel_780249 = array_index_780060 == array_index_772918 ? add_780248 : sel_780245;
  assign add_780252 = sel_780249 + 8'h01;
  assign sel_780253 = array_index_780060 == array_index_772924 ? add_780252 : sel_780249;
  assign add_780256 = sel_780253 + 8'h01;
  assign sel_780257 = array_index_780060 == array_index_772930 ? add_780256 : sel_780253;
  assign add_780260 = sel_780257 + 8'h01;
  assign sel_780261 = array_index_780060 == array_index_772936 ? add_780260 : sel_780257;
  assign add_780264 = sel_780261 + 8'h01;
  assign sel_780265 = array_index_780060 == array_index_772942 ? add_780264 : sel_780261;
  assign add_780268 = sel_780265 + 8'h01;
  assign sel_780269 = array_index_780060 == array_index_772948 ? add_780268 : sel_780265;
  assign add_780272 = sel_780269 + 8'h01;
  assign sel_780273 = array_index_780060 == array_index_772954 ? add_780272 : sel_780269;
  assign add_780276 = sel_780273 + 8'h01;
  assign sel_780277 = array_index_780060 == array_index_772960 ? add_780276 : sel_780273;
  assign add_780280 = sel_780277 + 8'h01;
  assign sel_780281 = array_index_780060 == array_index_772966 ? add_780280 : sel_780277;
  assign add_780284 = sel_780281 + 8'h01;
  assign sel_780285 = array_index_780060 == array_index_772972 ? add_780284 : sel_780281;
  assign add_780288 = sel_780285 + 8'h01;
  assign sel_780289 = array_index_780060 == array_index_772978 ? add_780288 : sel_780285;
  assign add_780292 = sel_780289 + 8'h01;
  assign sel_780293 = array_index_780060 == array_index_772984 ? add_780292 : sel_780289;
  assign add_780296 = sel_780293 + 8'h01;
  assign sel_780297 = array_index_780060 == array_index_772990 ? add_780296 : sel_780293;
  assign add_780300 = sel_780297 + 8'h01;
  assign sel_780301 = array_index_780060 == array_index_772996 ? add_780300 : sel_780297;
  assign add_780304 = sel_780301 + 8'h01;
  assign sel_780305 = array_index_780060 == array_index_773002 ? add_780304 : sel_780301;
  assign add_780308 = sel_780305 + 8'h01;
  assign sel_780309 = array_index_780060 == array_index_773008 ? add_780308 : sel_780305;
  assign add_780312 = sel_780309 + 8'h01;
  assign sel_780313 = array_index_780060 == array_index_773014 ? add_780312 : sel_780309;
  assign add_780316 = sel_780313 + 8'h01;
  assign sel_780317 = array_index_780060 == array_index_773020 ? add_780316 : sel_780313;
  assign add_780320 = sel_780317 + 8'h01;
  assign sel_780321 = array_index_780060 == array_index_773026 ? add_780320 : sel_780317;
  assign add_780324 = sel_780321 + 8'h01;
  assign sel_780325 = array_index_780060 == array_index_773032 ? add_780324 : sel_780321;
  assign add_780328 = sel_780325 + 8'h01;
  assign sel_780329 = array_index_780060 == array_index_773038 ? add_780328 : sel_780325;
  assign add_780332 = sel_780329 + 8'h01;
  assign sel_780333 = array_index_780060 == array_index_773044 ? add_780332 : sel_780329;
  assign add_780336 = sel_780333 + 8'h01;
  assign sel_780337 = array_index_780060 == array_index_773050 ? add_780336 : sel_780333;
  assign add_780340 = sel_780337 + 8'h01;
  assign sel_780341 = array_index_780060 == array_index_773056 ? add_780340 : sel_780337;
  assign add_780344 = sel_780341 + 8'h01;
  assign sel_780345 = array_index_780060 == array_index_773062 ? add_780344 : sel_780341;
  assign add_780348 = sel_780345 + 8'h01;
  assign sel_780349 = array_index_780060 == array_index_773068 ? add_780348 : sel_780345;
  assign add_780352 = sel_780349 + 8'h01;
  assign sel_780353 = array_index_780060 == array_index_773074 ? add_780352 : sel_780349;
  assign add_780356 = sel_780353 + 8'h01;
  assign sel_780357 = array_index_780060 == array_index_773080 ? add_780356 : sel_780353;
  assign add_780360 = sel_780357 + 8'h01;
  assign sel_780361 = array_index_780060 == array_index_773086 ? add_780360 : sel_780357;
  assign add_780364 = sel_780361 + 8'h01;
  assign sel_780365 = array_index_780060 == array_index_773092 ? add_780364 : sel_780361;
  assign add_780368 = sel_780365 + 8'h01;
  assign sel_780369 = array_index_780060 == array_index_773098 ? add_780368 : sel_780365;
  assign add_780372 = sel_780369 + 8'h01;
  assign sel_780373 = array_index_780060 == array_index_773104 ? add_780372 : sel_780369;
  assign add_780376 = sel_780373 + 8'h01;
  assign sel_780377 = array_index_780060 == array_index_773110 ? add_780376 : sel_780373;
  assign add_780380 = sel_780377 + 8'h01;
  assign sel_780381 = array_index_780060 == array_index_773116 ? add_780380 : sel_780377;
  assign add_780384 = sel_780381 + 8'h01;
  assign sel_780385 = array_index_780060 == array_index_773122 ? add_780384 : sel_780381;
  assign add_780388 = sel_780385 + 8'h01;
  assign sel_780389 = array_index_780060 == array_index_773128 ? add_780388 : sel_780385;
  assign add_780392 = sel_780389 + 8'h01;
  assign sel_780393 = array_index_780060 == array_index_773134 ? add_780392 : sel_780389;
  assign add_780396 = sel_780393 + 8'h01;
  assign sel_780397 = array_index_780060 == array_index_773140 ? add_780396 : sel_780393;
  assign add_780400 = sel_780397 + 8'h01;
  assign sel_780401 = array_index_780060 == array_index_773146 ? add_780400 : sel_780397;
  assign add_780404 = sel_780401 + 8'h01;
  assign sel_780405 = array_index_780060 == array_index_773152 ? add_780404 : sel_780401;
  assign add_780408 = sel_780405 + 8'h01;
  assign sel_780409 = array_index_780060 == array_index_773158 ? add_780408 : sel_780405;
  assign add_780412 = sel_780409 + 8'h01;
  assign sel_780413 = array_index_780060 == array_index_773164 ? add_780412 : sel_780409;
  assign add_780416 = sel_780413 + 8'h01;
  assign sel_780417 = array_index_780060 == array_index_773170 ? add_780416 : sel_780413;
  assign add_780421 = sel_780417 + 8'h01;
  assign array_index_780422 = set1_unflattened[7'h15];
  assign sel_780423 = array_index_780060 == array_index_773176 ? add_780421 : sel_780417;
  assign add_780426 = sel_780423 + 8'h01;
  assign sel_780427 = array_index_780422 == array_index_772632 ? add_780426 : sel_780423;
  assign add_780430 = sel_780427 + 8'h01;
  assign sel_780431 = array_index_780422 == array_index_772636 ? add_780430 : sel_780427;
  assign add_780434 = sel_780431 + 8'h01;
  assign sel_780435 = array_index_780422 == array_index_772644 ? add_780434 : sel_780431;
  assign add_780438 = sel_780435 + 8'h01;
  assign sel_780439 = array_index_780422 == array_index_772652 ? add_780438 : sel_780435;
  assign add_780442 = sel_780439 + 8'h01;
  assign sel_780443 = array_index_780422 == array_index_772660 ? add_780442 : sel_780439;
  assign add_780446 = sel_780443 + 8'h01;
  assign sel_780447 = array_index_780422 == array_index_772668 ? add_780446 : sel_780443;
  assign add_780450 = sel_780447 + 8'h01;
  assign sel_780451 = array_index_780422 == array_index_772676 ? add_780450 : sel_780447;
  assign add_780454 = sel_780451 + 8'h01;
  assign sel_780455 = array_index_780422 == array_index_772684 ? add_780454 : sel_780451;
  assign add_780458 = sel_780455 + 8'h01;
  assign sel_780459 = array_index_780422 == array_index_772690 ? add_780458 : sel_780455;
  assign add_780462 = sel_780459 + 8'h01;
  assign sel_780463 = array_index_780422 == array_index_772696 ? add_780462 : sel_780459;
  assign add_780466 = sel_780463 + 8'h01;
  assign sel_780467 = array_index_780422 == array_index_772702 ? add_780466 : sel_780463;
  assign add_780470 = sel_780467 + 8'h01;
  assign sel_780471 = array_index_780422 == array_index_772708 ? add_780470 : sel_780467;
  assign add_780474 = sel_780471 + 8'h01;
  assign sel_780475 = array_index_780422 == array_index_772714 ? add_780474 : sel_780471;
  assign add_780478 = sel_780475 + 8'h01;
  assign sel_780479 = array_index_780422 == array_index_772720 ? add_780478 : sel_780475;
  assign add_780482 = sel_780479 + 8'h01;
  assign sel_780483 = array_index_780422 == array_index_772726 ? add_780482 : sel_780479;
  assign add_780486 = sel_780483 + 8'h01;
  assign sel_780487 = array_index_780422 == array_index_772732 ? add_780486 : sel_780483;
  assign add_780490 = sel_780487 + 8'h01;
  assign sel_780491 = array_index_780422 == array_index_772738 ? add_780490 : sel_780487;
  assign add_780494 = sel_780491 + 8'h01;
  assign sel_780495 = array_index_780422 == array_index_772744 ? add_780494 : sel_780491;
  assign add_780498 = sel_780495 + 8'h01;
  assign sel_780499 = array_index_780422 == array_index_772750 ? add_780498 : sel_780495;
  assign add_780502 = sel_780499 + 8'h01;
  assign sel_780503 = array_index_780422 == array_index_772756 ? add_780502 : sel_780499;
  assign add_780506 = sel_780503 + 8'h01;
  assign sel_780507 = array_index_780422 == array_index_772762 ? add_780506 : sel_780503;
  assign add_780510 = sel_780507 + 8'h01;
  assign sel_780511 = array_index_780422 == array_index_772768 ? add_780510 : sel_780507;
  assign add_780514 = sel_780511 + 8'h01;
  assign sel_780515 = array_index_780422 == array_index_772774 ? add_780514 : sel_780511;
  assign add_780518 = sel_780515 + 8'h01;
  assign sel_780519 = array_index_780422 == array_index_772780 ? add_780518 : sel_780515;
  assign add_780522 = sel_780519 + 8'h01;
  assign sel_780523 = array_index_780422 == array_index_772786 ? add_780522 : sel_780519;
  assign add_780526 = sel_780523 + 8'h01;
  assign sel_780527 = array_index_780422 == array_index_772792 ? add_780526 : sel_780523;
  assign add_780530 = sel_780527 + 8'h01;
  assign sel_780531 = array_index_780422 == array_index_772798 ? add_780530 : sel_780527;
  assign add_780534 = sel_780531 + 8'h01;
  assign sel_780535 = array_index_780422 == array_index_772804 ? add_780534 : sel_780531;
  assign add_780538 = sel_780535 + 8'h01;
  assign sel_780539 = array_index_780422 == array_index_772810 ? add_780538 : sel_780535;
  assign add_780542 = sel_780539 + 8'h01;
  assign sel_780543 = array_index_780422 == array_index_772816 ? add_780542 : sel_780539;
  assign add_780546 = sel_780543 + 8'h01;
  assign sel_780547 = array_index_780422 == array_index_772822 ? add_780546 : sel_780543;
  assign add_780550 = sel_780547 + 8'h01;
  assign sel_780551 = array_index_780422 == array_index_772828 ? add_780550 : sel_780547;
  assign add_780554 = sel_780551 + 8'h01;
  assign sel_780555 = array_index_780422 == array_index_772834 ? add_780554 : sel_780551;
  assign add_780558 = sel_780555 + 8'h01;
  assign sel_780559 = array_index_780422 == array_index_772840 ? add_780558 : sel_780555;
  assign add_780562 = sel_780559 + 8'h01;
  assign sel_780563 = array_index_780422 == array_index_772846 ? add_780562 : sel_780559;
  assign add_780566 = sel_780563 + 8'h01;
  assign sel_780567 = array_index_780422 == array_index_772852 ? add_780566 : sel_780563;
  assign add_780570 = sel_780567 + 8'h01;
  assign sel_780571 = array_index_780422 == array_index_772858 ? add_780570 : sel_780567;
  assign add_780574 = sel_780571 + 8'h01;
  assign sel_780575 = array_index_780422 == array_index_772864 ? add_780574 : sel_780571;
  assign add_780578 = sel_780575 + 8'h01;
  assign sel_780579 = array_index_780422 == array_index_772870 ? add_780578 : sel_780575;
  assign add_780582 = sel_780579 + 8'h01;
  assign sel_780583 = array_index_780422 == array_index_772876 ? add_780582 : sel_780579;
  assign add_780586 = sel_780583 + 8'h01;
  assign sel_780587 = array_index_780422 == array_index_772882 ? add_780586 : sel_780583;
  assign add_780590 = sel_780587 + 8'h01;
  assign sel_780591 = array_index_780422 == array_index_772888 ? add_780590 : sel_780587;
  assign add_780594 = sel_780591 + 8'h01;
  assign sel_780595 = array_index_780422 == array_index_772894 ? add_780594 : sel_780591;
  assign add_780598 = sel_780595 + 8'h01;
  assign sel_780599 = array_index_780422 == array_index_772900 ? add_780598 : sel_780595;
  assign add_780602 = sel_780599 + 8'h01;
  assign sel_780603 = array_index_780422 == array_index_772906 ? add_780602 : sel_780599;
  assign add_780606 = sel_780603 + 8'h01;
  assign sel_780607 = array_index_780422 == array_index_772912 ? add_780606 : sel_780603;
  assign add_780610 = sel_780607 + 8'h01;
  assign sel_780611 = array_index_780422 == array_index_772918 ? add_780610 : sel_780607;
  assign add_780614 = sel_780611 + 8'h01;
  assign sel_780615 = array_index_780422 == array_index_772924 ? add_780614 : sel_780611;
  assign add_780618 = sel_780615 + 8'h01;
  assign sel_780619 = array_index_780422 == array_index_772930 ? add_780618 : sel_780615;
  assign add_780622 = sel_780619 + 8'h01;
  assign sel_780623 = array_index_780422 == array_index_772936 ? add_780622 : sel_780619;
  assign add_780626 = sel_780623 + 8'h01;
  assign sel_780627 = array_index_780422 == array_index_772942 ? add_780626 : sel_780623;
  assign add_780630 = sel_780627 + 8'h01;
  assign sel_780631 = array_index_780422 == array_index_772948 ? add_780630 : sel_780627;
  assign add_780634 = sel_780631 + 8'h01;
  assign sel_780635 = array_index_780422 == array_index_772954 ? add_780634 : sel_780631;
  assign add_780638 = sel_780635 + 8'h01;
  assign sel_780639 = array_index_780422 == array_index_772960 ? add_780638 : sel_780635;
  assign add_780642 = sel_780639 + 8'h01;
  assign sel_780643 = array_index_780422 == array_index_772966 ? add_780642 : sel_780639;
  assign add_780646 = sel_780643 + 8'h01;
  assign sel_780647 = array_index_780422 == array_index_772972 ? add_780646 : sel_780643;
  assign add_780650 = sel_780647 + 8'h01;
  assign sel_780651 = array_index_780422 == array_index_772978 ? add_780650 : sel_780647;
  assign add_780654 = sel_780651 + 8'h01;
  assign sel_780655 = array_index_780422 == array_index_772984 ? add_780654 : sel_780651;
  assign add_780658 = sel_780655 + 8'h01;
  assign sel_780659 = array_index_780422 == array_index_772990 ? add_780658 : sel_780655;
  assign add_780662 = sel_780659 + 8'h01;
  assign sel_780663 = array_index_780422 == array_index_772996 ? add_780662 : sel_780659;
  assign add_780666 = sel_780663 + 8'h01;
  assign sel_780667 = array_index_780422 == array_index_773002 ? add_780666 : sel_780663;
  assign add_780670 = sel_780667 + 8'h01;
  assign sel_780671 = array_index_780422 == array_index_773008 ? add_780670 : sel_780667;
  assign add_780674 = sel_780671 + 8'h01;
  assign sel_780675 = array_index_780422 == array_index_773014 ? add_780674 : sel_780671;
  assign add_780678 = sel_780675 + 8'h01;
  assign sel_780679 = array_index_780422 == array_index_773020 ? add_780678 : sel_780675;
  assign add_780682 = sel_780679 + 8'h01;
  assign sel_780683 = array_index_780422 == array_index_773026 ? add_780682 : sel_780679;
  assign add_780686 = sel_780683 + 8'h01;
  assign sel_780687 = array_index_780422 == array_index_773032 ? add_780686 : sel_780683;
  assign add_780690 = sel_780687 + 8'h01;
  assign sel_780691 = array_index_780422 == array_index_773038 ? add_780690 : sel_780687;
  assign add_780694 = sel_780691 + 8'h01;
  assign sel_780695 = array_index_780422 == array_index_773044 ? add_780694 : sel_780691;
  assign add_780698 = sel_780695 + 8'h01;
  assign sel_780699 = array_index_780422 == array_index_773050 ? add_780698 : sel_780695;
  assign add_780702 = sel_780699 + 8'h01;
  assign sel_780703 = array_index_780422 == array_index_773056 ? add_780702 : sel_780699;
  assign add_780706 = sel_780703 + 8'h01;
  assign sel_780707 = array_index_780422 == array_index_773062 ? add_780706 : sel_780703;
  assign add_780710 = sel_780707 + 8'h01;
  assign sel_780711 = array_index_780422 == array_index_773068 ? add_780710 : sel_780707;
  assign add_780714 = sel_780711 + 8'h01;
  assign sel_780715 = array_index_780422 == array_index_773074 ? add_780714 : sel_780711;
  assign add_780718 = sel_780715 + 8'h01;
  assign sel_780719 = array_index_780422 == array_index_773080 ? add_780718 : sel_780715;
  assign add_780722 = sel_780719 + 8'h01;
  assign sel_780723 = array_index_780422 == array_index_773086 ? add_780722 : sel_780719;
  assign add_780726 = sel_780723 + 8'h01;
  assign sel_780727 = array_index_780422 == array_index_773092 ? add_780726 : sel_780723;
  assign add_780730 = sel_780727 + 8'h01;
  assign sel_780731 = array_index_780422 == array_index_773098 ? add_780730 : sel_780727;
  assign add_780734 = sel_780731 + 8'h01;
  assign sel_780735 = array_index_780422 == array_index_773104 ? add_780734 : sel_780731;
  assign add_780738 = sel_780735 + 8'h01;
  assign sel_780739 = array_index_780422 == array_index_773110 ? add_780738 : sel_780735;
  assign add_780742 = sel_780739 + 8'h01;
  assign sel_780743 = array_index_780422 == array_index_773116 ? add_780742 : sel_780739;
  assign add_780746 = sel_780743 + 8'h01;
  assign sel_780747 = array_index_780422 == array_index_773122 ? add_780746 : sel_780743;
  assign add_780750 = sel_780747 + 8'h01;
  assign sel_780751 = array_index_780422 == array_index_773128 ? add_780750 : sel_780747;
  assign add_780754 = sel_780751 + 8'h01;
  assign sel_780755 = array_index_780422 == array_index_773134 ? add_780754 : sel_780751;
  assign add_780758 = sel_780755 + 8'h01;
  assign sel_780759 = array_index_780422 == array_index_773140 ? add_780758 : sel_780755;
  assign add_780762 = sel_780759 + 8'h01;
  assign sel_780763 = array_index_780422 == array_index_773146 ? add_780762 : sel_780759;
  assign add_780766 = sel_780763 + 8'h01;
  assign sel_780767 = array_index_780422 == array_index_773152 ? add_780766 : sel_780763;
  assign add_780770 = sel_780767 + 8'h01;
  assign sel_780771 = array_index_780422 == array_index_773158 ? add_780770 : sel_780767;
  assign add_780774 = sel_780771 + 8'h01;
  assign sel_780775 = array_index_780422 == array_index_773164 ? add_780774 : sel_780771;
  assign add_780778 = sel_780775 + 8'h01;
  assign sel_780779 = array_index_780422 == array_index_773170 ? add_780778 : sel_780775;
  assign add_780783 = sel_780779 + 8'h01;
  assign array_index_780784 = set1_unflattened[7'h16];
  assign sel_780785 = array_index_780422 == array_index_773176 ? add_780783 : sel_780779;
  assign add_780788 = sel_780785 + 8'h01;
  assign sel_780789 = array_index_780784 == array_index_772632 ? add_780788 : sel_780785;
  assign add_780792 = sel_780789 + 8'h01;
  assign sel_780793 = array_index_780784 == array_index_772636 ? add_780792 : sel_780789;
  assign add_780796 = sel_780793 + 8'h01;
  assign sel_780797 = array_index_780784 == array_index_772644 ? add_780796 : sel_780793;
  assign add_780800 = sel_780797 + 8'h01;
  assign sel_780801 = array_index_780784 == array_index_772652 ? add_780800 : sel_780797;
  assign add_780804 = sel_780801 + 8'h01;
  assign sel_780805 = array_index_780784 == array_index_772660 ? add_780804 : sel_780801;
  assign add_780808 = sel_780805 + 8'h01;
  assign sel_780809 = array_index_780784 == array_index_772668 ? add_780808 : sel_780805;
  assign add_780812 = sel_780809 + 8'h01;
  assign sel_780813 = array_index_780784 == array_index_772676 ? add_780812 : sel_780809;
  assign add_780816 = sel_780813 + 8'h01;
  assign sel_780817 = array_index_780784 == array_index_772684 ? add_780816 : sel_780813;
  assign add_780820 = sel_780817 + 8'h01;
  assign sel_780821 = array_index_780784 == array_index_772690 ? add_780820 : sel_780817;
  assign add_780824 = sel_780821 + 8'h01;
  assign sel_780825 = array_index_780784 == array_index_772696 ? add_780824 : sel_780821;
  assign add_780828 = sel_780825 + 8'h01;
  assign sel_780829 = array_index_780784 == array_index_772702 ? add_780828 : sel_780825;
  assign add_780832 = sel_780829 + 8'h01;
  assign sel_780833 = array_index_780784 == array_index_772708 ? add_780832 : sel_780829;
  assign add_780836 = sel_780833 + 8'h01;
  assign sel_780837 = array_index_780784 == array_index_772714 ? add_780836 : sel_780833;
  assign add_780840 = sel_780837 + 8'h01;
  assign sel_780841 = array_index_780784 == array_index_772720 ? add_780840 : sel_780837;
  assign add_780844 = sel_780841 + 8'h01;
  assign sel_780845 = array_index_780784 == array_index_772726 ? add_780844 : sel_780841;
  assign add_780848 = sel_780845 + 8'h01;
  assign sel_780849 = array_index_780784 == array_index_772732 ? add_780848 : sel_780845;
  assign add_780852 = sel_780849 + 8'h01;
  assign sel_780853 = array_index_780784 == array_index_772738 ? add_780852 : sel_780849;
  assign add_780856 = sel_780853 + 8'h01;
  assign sel_780857 = array_index_780784 == array_index_772744 ? add_780856 : sel_780853;
  assign add_780860 = sel_780857 + 8'h01;
  assign sel_780861 = array_index_780784 == array_index_772750 ? add_780860 : sel_780857;
  assign add_780864 = sel_780861 + 8'h01;
  assign sel_780865 = array_index_780784 == array_index_772756 ? add_780864 : sel_780861;
  assign add_780868 = sel_780865 + 8'h01;
  assign sel_780869 = array_index_780784 == array_index_772762 ? add_780868 : sel_780865;
  assign add_780872 = sel_780869 + 8'h01;
  assign sel_780873 = array_index_780784 == array_index_772768 ? add_780872 : sel_780869;
  assign add_780876 = sel_780873 + 8'h01;
  assign sel_780877 = array_index_780784 == array_index_772774 ? add_780876 : sel_780873;
  assign add_780880 = sel_780877 + 8'h01;
  assign sel_780881 = array_index_780784 == array_index_772780 ? add_780880 : sel_780877;
  assign add_780884 = sel_780881 + 8'h01;
  assign sel_780885 = array_index_780784 == array_index_772786 ? add_780884 : sel_780881;
  assign add_780888 = sel_780885 + 8'h01;
  assign sel_780889 = array_index_780784 == array_index_772792 ? add_780888 : sel_780885;
  assign add_780892 = sel_780889 + 8'h01;
  assign sel_780893 = array_index_780784 == array_index_772798 ? add_780892 : sel_780889;
  assign add_780896 = sel_780893 + 8'h01;
  assign sel_780897 = array_index_780784 == array_index_772804 ? add_780896 : sel_780893;
  assign add_780900 = sel_780897 + 8'h01;
  assign sel_780901 = array_index_780784 == array_index_772810 ? add_780900 : sel_780897;
  assign add_780904 = sel_780901 + 8'h01;
  assign sel_780905 = array_index_780784 == array_index_772816 ? add_780904 : sel_780901;
  assign add_780908 = sel_780905 + 8'h01;
  assign sel_780909 = array_index_780784 == array_index_772822 ? add_780908 : sel_780905;
  assign add_780912 = sel_780909 + 8'h01;
  assign sel_780913 = array_index_780784 == array_index_772828 ? add_780912 : sel_780909;
  assign add_780916 = sel_780913 + 8'h01;
  assign sel_780917 = array_index_780784 == array_index_772834 ? add_780916 : sel_780913;
  assign add_780920 = sel_780917 + 8'h01;
  assign sel_780921 = array_index_780784 == array_index_772840 ? add_780920 : sel_780917;
  assign add_780924 = sel_780921 + 8'h01;
  assign sel_780925 = array_index_780784 == array_index_772846 ? add_780924 : sel_780921;
  assign add_780928 = sel_780925 + 8'h01;
  assign sel_780929 = array_index_780784 == array_index_772852 ? add_780928 : sel_780925;
  assign add_780932 = sel_780929 + 8'h01;
  assign sel_780933 = array_index_780784 == array_index_772858 ? add_780932 : sel_780929;
  assign add_780936 = sel_780933 + 8'h01;
  assign sel_780937 = array_index_780784 == array_index_772864 ? add_780936 : sel_780933;
  assign add_780940 = sel_780937 + 8'h01;
  assign sel_780941 = array_index_780784 == array_index_772870 ? add_780940 : sel_780937;
  assign add_780944 = sel_780941 + 8'h01;
  assign sel_780945 = array_index_780784 == array_index_772876 ? add_780944 : sel_780941;
  assign add_780948 = sel_780945 + 8'h01;
  assign sel_780949 = array_index_780784 == array_index_772882 ? add_780948 : sel_780945;
  assign add_780952 = sel_780949 + 8'h01;
  assign sel_780953 = array_index_780784 == array_index_772888 ? add_780952 : sel_780949;
  assign add_780956 = sel_780953 + 8'h01;
  assign sel_780957 = array_index_780784 == array_index_772894 ? add_780956 : sel_780953;
  assign add_780960 = sel_780957 + 8'h01;
  assign sel_780961 = array_index_780784 == array_index_772900 ? add_780960 : sel_780957;
  assign add_780964 = sel_780961 + 8'h01;
  assign sel_780965 = array_index_780784 == array_index_772906 ? add_780964 : sel_780961;
  assign add_780968 = sel_780965 + 8'h01;
  assign sel_780969 = array_index_780784 == array_index_772912 ? add_780968 : sel_780965;
  assign add_780972 = sel_780969 + 8'h01;
  assign sel_780973 = array_index_780784 == array_index_772918 ? add_780972 : sel_780969;
  assign add_780976 = sel_780973 + 8'h01;
  assign sel_780977 = array_index_780784 == array_index_772924 ? add_780976 : sel_780973;
  assign add_780980 = sel_780977 + 8'h01;
  assign sel_780981 = array_index_780784 == array_index_772930 ? add_780980 : sel_780977;
  assign add_780984 = sel_780981 + 8'h01;
  assign sel_780985 = array_index_780784 == array_index_772936 ? add_780984 : sel_780981;
  assign add_780988 = sel_780985 + 8'h01;
  assign sel_780989 = array_index_780784 == array_index_772942 ? add_780988 : sel_780985;
  assign add_780992 = sel_780989 + 8'h01;
  assign sel_780993 = array_index_780784 == array_index_772948 ? add_780992 : sel_780989;
  assign add_780996 = sel_780993 + 8'h01;
  assign sel_780997 = array_index_780784 == array_index_772954 ? add_780996 : sel_780993;
  assign add_781000 = sel_780997 + 8'h01;
  assign sel_781001 = array_index_780784 == array_index_772960 ? add_781000 : sel_780997;
  assign add_781004 = sel_781001 + 8'h01;
  assign sel_781005 = array_index_780784 == array_index_772966 ? add_781004 : sel_781001;
  assign add_781008 = sel_781005 + 8'h01;
  assign sel_781009 = array_index_780784 == array_index_772972 ? add_781008 : sel_781005;
  assign add_781012 = sel_781009 + 8'h01;
  assign sel_781013 = array_index_780784 == array_index_772978 ? add_781012 : sel_781009;
  assign add_781016 = sel_781013 + 8'h01;
  assign sel_781017 = array_index_780784 == array_index_772984 ? add_781016 : sel_781013;
  assign add_781020 = sel_781017 + 8'h01;
  assign sel_781021 = array_index_780784 == array_index_772990 ? add_781020 : sel_781017;
  assign add_781024 = sel_781021 + 8'h01;
  assign sel_781025 = array_index_780784 == array_index_772996 ? add_781024 : sel_781021;
  assign add_781028 = sel_781025 + 8'h01;
  assign sel_781029 = array_index_780784 == array_index_773002 ? add_781028 : sel_781025;
  assign add_781032 = sel_781029 + 8'h01;
  assign sel_781033 = array_index_780784 == array_index_773008 ? add_781032 : sel_781029;
  assign add_781036 = sel_781033 + 8'h01;
  assign sel_781037 = array_index_780784 == array_index_773014 ? add_781036 : sel_781033;
  assign add_781040 = sel_781037 + 8'h01;
  assign sel_781041 = array_index_780784 == array_index_773020 ? add_781040 : sel_781037;
  assign add_781044 = sel_781041 + 8'h01;
  assign sel_781045 = array_index_780784 == array_index_773026 ? add_781044 : sel_781041;
  assign add_781048 = sel_781045 + 8'h01;
  assign sel_781049 = array_index_780784 == array_index_773032 ? add_781048 : sel_781045;
  assign add_781052 = sel_781049 + 8'h01;
  assign sel_781053 = array_index_780784 == array_index_773038 ? add_781052 : sel_781049;
  assign add_781056 = sel_781053 + 8'h01;
  assign sel_781057 = array_index_780784 == array_index_773044 ? add_781056 : sel_781053;
  assign add_781060 = sel_781057 + 8'h01;
  assign sel_781061 = array_index_780784 == array_index_773050 ? add_781060 : sel_781057;
  assign add_781064 = sel_781061 + 8'h01;
  assign sel_781065 = array_index_780784 == array_index_773056 ? add_781064 : sel_781061;
  assign add_781068 = sel_781065 + 8'h01;
  assign sel_781069 = array_index_780784 == array_index_773062 ? add_781068 : sel_781065;
  assign add_781072 = sel_781069 + 8'h01;
  assign sel_781073 = array_index_780784 == array_index_773068 ? add_781072 : sel_781069;
  assign add_781076 = sel_781073 + 8'h01;
  assign sel_781077 = array_index_780784 == array_index_773074 ? add_781076 : sel_781073;
  assign add_781080 = sel_781077 + 8'h01;
  assign sel_781081 = array_index_780784 == array_index_773080 ? add_781080 : sel_781077;
  assign add_781084 = sel_781081 + 8'h01;
  assign sel_781085 = array_index_780784 == array_index_773086 ? add_781084 : sel_781081;
  assign add_781088 = sel_781085 + 8'h01;
  assign sel_781089 = array_index_780784 == array_index_773092 ? add_781088 : sel_781085;
  assign add_781092 = sel_781089 + 8'h01;
  assign sel_781093 = array_index_780784 == array_index_773098 ? add_781092 : sel_781089;
  assign add_781096 = sel_781093 + 8'h01;
  assign sel_781097 = array_index_780784 == array_index_773104 ? add_781096 : sel_781093;
  assign add_781100 = sel_781097 + 8'h01;
  assign sel_781101 = array_index_780784 == array_index_773110 ? add_781100 : sel_781097;
  assign add_781104 = sel_781101 + 8'h01;
  assign sel_781105 = array_index_780784 == array_index_773116 ? add_781104 : sel_781101;
  assign add_781108 = sel_781105 + 8'h01;
  assign sel_781109 = array_index_780784 == array_index_773122 ? add_781108 : sel_781105;
  assign add_781112 = sel_781109 + 8'h01;
  assign sel_781113 = array_index_780784 == array_index_773128 ? add_781112 : sel_781109;
  assign add_781116 = sel_781113 + 8'h01;
  assign sel_781117 = array_index_780784 == array_index_773134 ? add_781116 : sel_781113;
  assign add_781120 = sel_781117 + 8'h01;
  assign sel_781121 = array_index_780784 == array_index_773140 ? add_781120 : sel_781117;
  assign add_781124 = sel_781121 + 8'h01;
  assign sel_781125 = array_index_780784 == array_index_773146 ? add_781124 : sel_781121;
  assign add_781128 = sel_781125 + 8'h01;
  assign sel_781129 = array_index_780784 == array_index_773152 ? add_781128 : sel_781125;
  assign add_781132 = sel_781129 + 8'h01;
  assign sel_781133 = array_index_780784 == array_index_773158 ? add_781132 : sel_781129;
  assign add_781136 = sel_781133 + 8'h01;
  assign sel_781137 = array_index_780784 == array_index_773164 ? add_781136 : sel_781133;
  assign add_781140 = sel_781137 + 8'h01;
  assign sel_781141 = array_index_780784 == array_index_773170 ? add_781140 : sel_781137;
  assign add_781145 = sel_781141 + 8'h01;
  assign array_index_781146 = set1_unflattened[7'h17];
  assign sel_781147 = array_index_780784 == array_index_773176 ? add_781145 : sel_781141;
  assign add_781150 = sel_781147 + 8'h01;
  assign sel_781151 = array_index_781146 == array_index_772632 ? add_781150 : sel_781147;
  assign add_781154 = sel_781151 + 8'h01;
  assign sel_781155 = array_index_781146 == array_index_772636 ? add_781154 : sel_781151;
  assign add_781158 = sel_781155 + 8'h01;
  assign sel_781159 = array_index_781146 == array_index_772644 ? add_781158 : sel_781155;
  assign add_781162 = sel_781159 + 8'h01;
  assign sel_781163 = array_index_781146 == array_index_772652 ? add_781162 : sel_781159;
  assign add_781166 = sel_781163 + 8'h01;
  assign sel_781167 = array_index_781146 == array_index_772660 ? add_781166 : sel_781163;
  assign add_781170 = sel_781167 + 8'h01;
  assign sel_781171 = array_index_781146 == array_index_772668 ? add_781170 : sel_781167;
  assign add_781174 = sel_781171 + 8'h01;
  assign sel_781175 = array_index_781146 == array_index_772676 ? add_781174 : sel_781171;
  assign add_781178 = sel_781175 + 8'h01;
  assign sel_781179 = array_index_781146 == array_index_772684 ? add_781178 : sel_781175;
  assign add_781182 = sel_781179 + 8'h01;
  assign sel_781183 = array_index_781146 == array_index_772690 ? add_781182 : sel_781179;
  assign add_781186 = sel_781183 + 8'h01;
  assign sel_781187 = array_index_781146 == array_index_772696 ? add_781186 : sel_781183;
  assign add_781190 = sel_781187 + 8'h01;
  assign sel_781191 = array_index_781146 == array_index_772702 ? add_781190 : sel_781187;
  assign add_781194 = sel_781191 + 8'h01;
  assign sel_781195 = array_index_781146 == array_index_772708 ? add_781194 : sel_781191;
  assign add_781198 = sel_781195 + 8'h01;
  assign sel_781199 = array_index_781146 == array_index_772714 ? add_781198 : sel_781195;
  assign add_781202 = sel_781199 + 8'h01;
  assign sel_781203 = array_index_781146 == array_index_772720 ? add_781202 : sel_781199;
  assign add_781206 = sel_781203 + 8'h01;
  assign sel_781207 = array_index_781146 == array_index_772726 ? add_781206 : sel_781203;
  assign add_781210 = sel_781207 + 8'h01;
  assign sel_781211 = array_index_781146 == array_index_772732 ? add_781210 : sel_781207;
  assign add_781214 = sel_781211 + 8'h01;
  assign sel_781215 = array_index_781146 == array_index_772738 ? add_781214 : sel_781211;
  assign add_781218 = sel_781215 + 8'h01;
  assign sel_781219 = array_index_781146 == array_index_772744 ? add_781218 : sel_781215;
  assign add_781222 = sel_781219 + 8'h01;
  assign sel_781223 = array_index_781146 == array_index_772750 ? add_781222 : sel_781219;
  assign add_781226 = sel_781223 + 8'h01;
  assign sel_781227 = array_index_781146 == array_index_772756 ? add_781226 : sel_781223;
  assign add_781230 = sel_781227 + 8'h01;
  assign sel_781231 = array_index_781146 == array_index_772762 ? add_781230 : sel_781227;
  assign add_781234 = sel_781231 + 8'h01;
  assign sel_781235 = array_index_781146 == array_index_772768 ? add_781234 : sel_781231;
  assign add_781238 = sel_781235 + 8'h01;
  assign sel_781239 = array_index_781146 == array_index_772774 ? add_781238 : sel_781235;
  assign add_781242 = sel_781239 + 8'h01;
  assign sel_781243 = array_index_781146 == array_index_772780 ? add_781242 : sel_781239;
  assign add_781246 = sel_781243 + 8'h01;
  assign sel_781247 = array_index_781146 == array_index_772786 ? add_781246 : sel_781243;
  assign add_781250 = sel_781247 + 8'h01;
  assign sel_781251 = array_index_781146 == array_index_772792 ? add_781250 : sel_781247;
  assign add_781254 = sel_781251 + 8'h01;
  assign sel_781255 = array_index_781146 == array_index_772798 ? add_781254 : sel_781251;
  assign add_781258 = sel_781255 + 8'h01;
  assign sel_781259 = array_index_781146 == array_index_772804 ? add_781258 : sel_781255;
  assign add_781262 = sel_781259 + 8'h01;
  assign sel_781263 = array_index_781146 == array_index_772810 ? add_781262 : sel_781259;
  assign add_781266 = sel_781263 + 8'h01;
  assign sel_781267 = array_index_781146 == array_index_772816 ? add_781266 : sel_781263;
  assign add_781270 = sel_781267 + 8'h01;
  assign sel_781271 = array_index_781146 == array_index_772822 ? add_781270 : sel_781267;
  assign add_781274 = sel_781271 + 8'h01;
  assign sel_781275 = array_index_781146 == array_index_772828 ? add_781274 : sel_781271;
  assign add_781278 = sel_781275 + 8'h01;
  assign sel_781279 = array_index_781146 == array_index_772834 ? add_781278 : sel_781275;
  assign add_781282 = sel_781279 + 8'h01;
  assign sel_781283 = array_index_781146 == array_index_772840 ? add_781282 : sel_781279;
  assign add_781286 = sel_781283 + 8'h01;
  assign sel_781287 = array_index_781146 == array_index_772846 ? add_781286 : sel_781283;
  assign add_781290 = sel_781287 + 8'h01;
  assign sel_781291 = array_index_781146 == array_index_772852 ? add_781290 : sel_781287;
  assign add_781294 = sel_781291 + 8'h01;
  assign sel_781295 = array_index_781146 == array_index_772858 ? add_781294 : sel_781291;
  assign add_781298 = sel_781295 + 8'h01;
  assign sel_781299 = array_index_781146 == array_index_772864 ? add_781298 : sel_781295;
  assign add_781302 = sel_781299 + 8'h01;
  assign sel_781303 = array_index_781146 == array_index_772870 ? add_781302 : sel_781299;
  assign add_781306 = sel_781303 + 8'h01;
  assign sel_781307 = array_index_781146 == array_index_772876 ? add_781306 : sel_781303;
  assign add_781310 = sel_781307 + 8'h01;
  assign sel_781311 = array_index_781146 == array_index_772882 ? add_781310 : sel_781307;
  assign add_781314 = sel_781311 + 8'h01;
  assign sel_781315 = array_index_781146 == array_index_772888 ? add_781314 : sel_781311;
  assign add_781318 = sel_781315 + 8'h01;
  assign sel_781319 = array_index_781146 == array_index_772894 ? add_781318 : sel_781315;
  assign add_781322 = sel_781319 + 8'h01;
  assign sel_781323 = array_index_781146 == array_index_772900 ? add_781322 : sel_781319;
  assign add_781326 = sel_781323 + 8'h01;
  assign sel_781327 = array_index_781146 == array_index_772906 ? add_781326 : sel_781323;
  assign add_781330 = sel_781327 + 8'h01;
  assign sel_781331 = array_index_781146 == array_index_772912 ? add_781330 : sel_781327;
  assign add_781334 = sel_781331 + 8'h01;
  assign sel_781335 = array_index_781146 == array_index_772918 ? add_781334 : sel_781331;
  assign add_781338 = sel_781335 + 8'h01;
  assign sel_781339 = array_index_781146 == array_index_772924 ? add_781338 : sel_781335;
  assign add_781342 = sel_781339 + 8'h01;
  assign sel_781343 = array_index_781146 == array_index_772930 ? add_781342 : sel_781339;
  assign add_781346 = sel_781343 + 8'h01;
  assign sel_781347 = array_index_781146 == array_index_772936 ? add_781346 : sel_781343;
  assign add_781350 = sel_781347 + 8'h01;
  assign sel_781351 = array_index_781146 == array_index_772942 ? add_781350 : sel_781347;
  assign add_781354 = sel_781351 + 8'h01;
  assign sel_781355 = array_index_781146 == array_index_772948 ? add_781354 : sel_781351;
  assign add_781358 = sel_781355 + 8'h01;
  assign sel_781359 = array_index_781146 == array_index_772954 ? add_781358 : sel_781355;
  assign add_781362 = sel_781359 + 8'h01;
  assign sel_781363 = array_index_781146 == array_index_772960 ? add_781362 : sel_781359;
  assign add_781366 = sel_781363 + 8'h01;
  assign sel_781367 = array_index_781146 == array_index_772966 ? add_781366 : sel_781363;
  assign add_781370 = sel_781367 + 8'h01;
  assign sel_781371 = array_index_781146 == array_index_772972 ? add_781370 : sel_781367;
  assign add_781374 = sel_781371 + 8'h01;
  assign sel_781375 = array_index_781146 == array_index_772978 ? add_781374 : sel_781371;
  assign add_781378 = sel_781375 + 8'h01;
  assign sel_781379 = array_index_781146 == array_index_772984 ? add_781378 : sel_781375;
  assign add_781382 = sel_781379 + 8'h01;
  assign sel_781383 = array_index_781146 == array_index_772990 ? add_781382 : sel_781379;
  assign add_781386 = sel_781383 + 8'h01;
  assign sel_781387 = array_index_781146 == array_index_772996 ? add_781386 : sel_781383;
  assign add_781390 = sel_781387 + 8'h01;
  assign sel_781391 = array_index_781146 == array_index_773002 ? add_781390 : sel_781387;
  assign add_781394 = sel_781391 + 8'h01;
  assign sel_781395 = array_index_781146 == array_index_773008 ? add_781394 : sel_781391;
  assign add_781398 = sel_781395 + 8'h01;
  assign sel_781399 = array_index_781146 == array_index_773014 ? add_781398 : sel_781395;
  assign add_781402 = sel_781399 + 8'h01;
  assign sel_781403 = array_index_781146 == array_index_773020 ? add_781402 : sel_781399;
  assign add_781406 = sel_781403 + 8'h01;
  assign sel_781407 = array_index_781146 == array_index_773026 ? add_781406 : sel_781403;
  assign add_781410 = sel_781407 + 8'h01;
  assign sel_781411 = array_index_781146 == array_index_773032 ? add_781410 : sel_781407;
  assign add_781414 = sel_781411 + 8'h01;
  assign sel_781415 = array_index_781146 == array_index_773038 ? add_781414 : sel_781411;
  assign add_781418 = sel_781415 + 8'h01;
  assign sel_781419 = array_index_781146 == array_index_773044 ? add_781418 : sel_781415;
  assign add_781422 = sel_781419 + 8'h01;
  assign sel_781423 = array_index_781146 == array_index_773050 ? add_781422 : sel_781419;
  assign add_781426 = sel_781423 + 8'h01;
  assign sel_781427 = array_index_781146 == array_index_773056 ? add_781426 : sel_781423;
  assign add_781430 = sel_781427 + 8'h01;
  assign sel_781431 = array_index_781146 == array_index_773062 ? add_781430 : sel_781427;
  assign add_781434 = sel_781431 + 8'h01;
  assign sel_781435 = array_index_781146 == array_index_773068 ? add_781434 : sel_781431;
  assign add_781438 = sel_781435 + 8'h01;
  assign sel_781439 = array_index_781146 == array_index_773074 ? add_781438 : sel_781435;
  assign add_781442 = sel_781439 + 8'h01;
  assign sel_781443 = array_index_781146 == array_index_773080 ? add_781442 : sel_781439;
  assign add_781446 = sel_781443 + 8'h01;
  assign sel_781447 = array_index_781146 == array_index_773086 ? add_781446 : sel_781443;
  assign add_781450 = sel_781447 + 8'h01;
  assign sel_781451 = array_index_781146 == array_index_773092 ? add_781450 : sel_781447;
  assign add_781454 = sel_781451 + 8'h01;
  assign sel_781455 = array_index_781146 == array_index_773098 ? add_781454 : sel_781451;
  assign add_781458 = sel_781455 + 8'h01;
  assign sel_781459 = array_index_781146 == array_index_773104 ? add_781458 : sel_781455;
  assign add_781462 = sel_781459 + 8'h01;
  assign sel_781463 = array_index_781146 == array_index_773110 ? add_781462 : sel_781459;
  assign add_781466 = sel_781463 + 8'h01;
  assign sel_781467 = array_index_781146 == array_index_773116 ? add_781466 : sel_781463;
  assign add_781470 = sel_781467 + 8'h01;
  assign sel_781471 = array_index_781146 == array_index_773122 ? add_781470 : sel_781467;
  assign add_781474 = sel_781471 + 8'h01;
  assign sel_781475 = array_index_781146 == array_index_773128 ? add_781474 : sel_781471;
  assign add_781478 = sel_781475 + 8'h01;
  assign sel_781479 = array_index_781146 == array_index_773134 ? add_781478 : sel_781475;
  assign add_781482 = sel_781479 + 8'h01;
  assign sel_781483 = array_index_781146 == array_index_773140 ? add_781482 : sel_781479;
  assign add_781486 = sel_781483 + 8'h01;
  assign sel_781487 = array_index_781146 == array_index_773146 ? add_781486 : sel_781483;
  assign add_781490 = sel_781487 + 8'h01;
  assign sel_781491 = array_index_781146 == array_index_773152 ? add_781490 : sel_781487;
  assign add_781494 = sel_781491 + 8'h01;
  assign sel_781495 = array_index_781146 == array_index_773158 ? add_781494 : sel_781491;
  assign add_781498 = sel_781495 + 8'h01;
  assign sel_781499 = array_index_781146 == array_index_773164 ? add_781498 : sel_781495;
  assign add_781502 = sel_781499 + 8'h01;
  assign sel_781503 = array_index_781146 == array_index_773170 ? add_781502 : sel_781499;
  assign add_781507 = sel_781503 + 8'h01;
  assign array_index_781508 = set1_unflattened[7'h18];
  assign sel_781509 = array_index_781146 == array_index_773176 ? add_781507 : sel_781503;
  assign add_781512 = sel_781509 + 8'h01;
  assign sel_781513 = array_index_781508 == array_index_772632 ? add_781512 : sel_781509;
  assign add_781516 = sel_781513 + 8'h01;
  assign sel_781517 = array_index_781508 == array_index_772636 ? add_781516 : sel_781513;
  assign add_781520 = sel_781517 + 8'h01;
  assign sel_781521 = array_index_781508 == array_index_772644 ? add_781520 : sel_781517;
  assign add_781524 = sel_781521 + 8'h01;
  assign sel_781525 = array_index_781508 == array_index_772652 ? add_781524 : sel_781521;
  assign add_781528 = sel_781525 + 8'h01;
  assign sel_781529 = array_index_781508 == array_index_772660 ? add_781528 : sel_781525;
  assign add_781532 = sel_781529 + 8'h01;
  assign sel_781533 = array_index_781508 == array_index_772668 ? add_781532 : sel_781529;
  assign add_781536 = sel_781533 + 8'h01;
  assign sel_781537 = array_index_781508 == array_index_772676 ? add_781536 : sel_781533;
  assign add_781540 = sel_781537 + 8'h01;
  assign sel_781541 = array_index_781508 == array_index_772684 ? add_781540 : sel_781537;
  assign add_781544 = sel_781541 + 8'h01;
  assign sel_781545 = array_index_781508 == array_index_772690 ? add_781544 : sel_781541;
  assign add_781548 = sel_781545 + 8'h01;
  assign sel_781549 = array_index_781508 == array_index_772696 ? add_781548 : sel_781545;
  assign add_781552 = sel_781549 + 8'h01;
  assign sel_781553 = array_index_781508 == array_index_772702 ? add_781552 : sel_781549;
  assign add_781556 = sel_781553 + 8'h01;
  assign sel_781557 = array_index_781508 == array_index_772708 ? add_781556 : sel_781553;
  assign add_781560 = sel_781557 + 8'h01;
  assign sel_781561 = array_index_781508 == array_index_772714 ? add_781560 : sel_781557;
  assign add_781564 = sel_781561 + 8'h01;
  assign sel_781565 = array_index_781508 == array_index_772720 ? add_781564 : sel_781561;
  assign add_781568 = sel_781565 + 8'h01;
  assign sel_781569 = array_index_781508 == array_index_772726 ? add_781568 : sel_781565;
  assign add_781572 = sel_781569 + 8'h01;
  assign sel_781573 = array_index_781508 == array_index_772732 ? add_781572 : sel_781569;
  assign add_781576 = sel_781573 + 8'h01;
  assign sel_781577 = array_index_781508 == array_index_772738 ? add_781576 : sel_781573;
  assign add_781580 = sel_781577 + 8'h01;
  assign sel_781581 = array_index_781508 == array_index_772744 ? add_781580 : sel_781577;
  assign add_781584 = sel_781581 + 8'h01;
  assign sel_781585 = array_index_781508 == array_index_772750 ? add_781584 : sel_781581;
  assign add_781588 = sel_781585 + 8'h01;
  assign sel_781589 = array_index_781508 == array_index_772756 ? add_781588 : sel_781585;
  assign add_781592 = sel_781589 + 8'h01;
  assign sel_781593 = array_index_781508 == array_index_772762 ? add_781592 : sel_781589;
  assign add_781596 = sel_781593 + 8'h01;
  assign sel_781597 = array_index_781508 == array_index_772768 ? add_781596 : sel_781593;
  assign add_781600 = sel_781597 + 8'h01;
  assign sel_781601 = array_index_781508 == array_index_772774 ? add_781600 : sel_781597;
  assign add_781604 = sel_781601 + 8'h01;
  assign sel_781605 = array_index_781508 == array_index_772780 ? add_781604 : sel_781601;
  assign add_781608 = sel_781605 + 8'h01;
  assign sel_781609 = array_index_781508 == array_index_772786 ? add_781608 : sel_781605;
  assign add_781612 = sel_781609 + 8'h01;
  assign sel_781613 = array_index_781508 == array_index_772792 ? add_781612 : sel_781609;
  assign add_781616 = sel_781613 + 8'h01;
  assign sel_781617 = array_index_781508 == array_index_772798 ? add_781616 : sel_781613;
  assign add_781620 = sel_781617 + 8'h01;
  assign sel_781621 = array_index_781508 == array_index_772804 ? add_781620 : sel_781617;
  assign add_781624 = sel_781621 + 8'h01;
  assign sel_781625 = array_index_781508 == array_index_772810 ? add_781624 : sel_781621;
  assign add_781628 = sel_781625 + 8'h01;
  assign sel_781629 = array_index_781508 == array_index_772816 ? add_781628 : sel_781625;
  assign add_781632 = sel_781629 + 8'h01;
  assign sel_781633 = array_index_781508 == array_index_772822 ? add_781632 : sel_781629;
  assign add_781636 = sel_781633 + 8'h01;
  assign sel_781637 = array_index_781508 == array_index_772828 ? add_781636 : sel_781633;
  assign add_781640 = sel_781637 + 8'h01;
  assign sel_781641 = array_index_781508 == array_index_772834 ? add_781640 : sel_781637;
  assign add_781644 = sel_781641 + 8'h01;
  assign sel_781645 = array_index_781508 == array_index_772840 ? add_781644 : sel_781641;
  assign add_781648 = sel_781645 + 8'h01;
  assign sel_781649 = array_index_781508 == array_index_772846 ? add_781648 : sel_781645;
  assign add_781652 = sel_781649 + 8'h01;
  assign sel_781653 = array_index_781508 == array_index_772852 ? add_781652 : sel_781649;
  assign add_781656 = sel_781653 + 8'h01;
  assign sel_781657 = array_index_781508 == array_index_772858 ? add_781656 : sel_781653;
  assign add_781660 = sel_781657 + 8'h01;
  assign sel_781661 = array_index_781508 == array_index_772864 ? add_781660 : sel_781657;
  assign add_781664 = sel_781661 + 8'h01;
  assign sel_781665 = array_index_781508 == array_index_772870 ? add_781664 : sel_781661;
  assign add_781668 = sel_781665 + 8'h01;
  assign sel_781669 = array_index_781508 == array_index_772876 ? add_781668 : sel_781665;
  assign add_781672 = sel_781669 + 8'h01;
  assign sel_781673 = array_index_781508 == array_index_772882 ? add_781672 : sel_781669;
  assign add_781676 = sel_781673 + 8'h01;
  assign sel_781677 = array_index_781508 == array_index_772888 ? add_781676 : sel_781673;
  assign add_781680 = sel_781677 + 8'h01;
  assign sel_781681 = array_index_781508 == array_index_772894 ? add_781680 : sel_781677;
  assign add_781684 = sel_781681 + 8'h01;
  assign sel_781685 = array_index_781508 == array_index_772900 ? add_781684 : sel_781681;
  assign add_781688 = sel_781685 + 8'h01;
  assign sel_781689 = array_index_781508 == array_index_772906 ? add_781688 : sel_781685;
  assign add_781692 = sel_781689 + 8'h01;
  assign sel_781693 = array_index_781508 == array_index_772912 ? add_781692 : sel_781689;
  assign add_781696 = sel_781693 + 8'h01;
  assign sel_781697 = array_index_781508 == array_index_772918 ? add_781696 : sel_781693;
  assign add_781700 = sel_781697 + 8'h01;
  assign sel_781701 = array_index_781508 == array_index_772924 ? add_781700 : sel_781697;
  assign add_781704 = sel_781701 + 8'h01;
  assign sel_781705 = array_index_781508 == array_index_772930 ? add_781704 : sel_781701;
  assign add_781708 = sel_781705 + 8'h01;
  assign sel_781709 = array_index_781508 == array_index_772936 ? add_781708 : sel_781705;
  assign add_781712 = sel_781709 + 8'h01;
  assign sel_781713 = array_index_781508 == array_index_772942 ? add_781712 : sel_781709;
  assign add_781716 = sel_781713 + 8'h01;
  assign sel_781717 = array_index_781508 == array_index_772948 ? add_781716 : sel_781713;
  assign add_781720 = sel_781717 + 8'h01;
  assign sel_781721 = array_index_781508 == array_index_772954 ? add_781720 : sel_781717;
  assign add_781724 = sel_781721 + 8'h01;
  assign sel_781725 = array_index_781508 == array_index_772960 ? add_781724 : sel_781721;
  assign add_781728 = sel_781725 + 8'h01;
  assign sel_781729 = array_index_781508 == array_index_772966 ? add_781728 : sel_781725;
  assign add_781732 = sel_781729 + 8'h01;
  assign sel_781733 = array_index_781508 == array_index_772972 ? add_781732 : sel_781729;
  assign add_781736 = sel_781733 + 8'h01;
  assign sel_781737 = array_index_781508 == array_index_772978 ? add_781736 : sel_781733;
  assign add_781740 = sel_781737 + 8'h01;
  assign sel_781741 = array_index_781508 == array_index_772984 ? add_781740 : sel_781737;
  assign add_781744 = sel_781741 + 8'h01;
  assign sel_781745 = array_index_781508 == array_index_772990 ? add_781744 : sel_781741;
  assign add_781748 = sel_781745 + 8'h01;
  assign sel_781749 = array_index_781508 == array_index_772996 ? add_781748 : sel_781745;
  assign add_781752 = sel_781749 + 8'h01;
  assign sel_781753 = array_index_781508 == array_index_773002 ? add_781752 : sel_781749;
  assign add_781756 = sel_781753 + 8'h01;
  assign sel_781757 = array_index_781508 == array_index_773008 ? add_781756 : sel_781753;
  assign add_781760 = sel_781757 + 8'h01;
  assign sel_781761 = array_index_781508 == array_index_773014 ? add_781760 : sel_781757;
  assign add_781764 = sel_781761 + 8'h01;
  assign sel_781765 = array_index_781508 == array_index_773020 ? add_781764 : sel_781761;
  assign add_781768 = sel_781765 + 8'h01;
  assign sel_781769 = array_index_781508 == array_index_773026 ? add_781768 : sel_781765;
  assign add_781772 = sel_781769 + 8'h01;
  assign sel_781773 = array_index_781508 == array_index_773032 ? add_781772 : sel_781769;
  assign add_781776 = sel_781773 + 8'h01;
  assign sel_781777 = array_index_781508 == array_index_773038 ? add_781776 : sel_781773;
  assign add_781780 = sel_781777 + 8'h01;
  assign sel_781781 = array_index_781508 == array_index_773044 ? add_781780 : sel_781777;
  assign add_781784 = sel_781781 + 8'h01;
  assign sel_781785 = array_index_781508 == array_index_773050 ? add_781784 : sel_781781;
  assign add_781788 = sel_781785 + 8'h01;
  assign sel_781789 = array_index_781508 == array_index_773056 ? add_781788 : sel_781785;
  assign add_781792 = sel_781789 + 8'h01;
  assign sel_781793 = array_index_781508 == array_index_773062 ? add_781792 : sel_781789;
  assign add_781796 = sel_781793 + 8'h01;
  assign sel_781797 = array_index_781508 == array_index_773068 ? add_781796 : sel_781793;
  assign add_781800 = sel_781797 + 8'h01;
  assign sel_781801 = array_index_781508 == array_index_773074 ? add_781800 : sel_781797;
  assign add_781804 = sel_781801 + 8'h01;
  assign sel_781805 = array_index_781508 == array_index_773080 ? add_781804 : sel_781801;
  assign add_781808 = sel_781805 + 8'h01;
  assign sel_781809 = array_index_781508 == array_index_773086 ? add_781808 : sel_781805;
  assign add_781812 = sel_781809 + 8'h01;
  assign sel_781813 = array_index_781508 == array_index_773092 ? add_781812 : sel_781809;
  assign add_781816 = sel_781813 + 8'h01;
  assign sel_781817 = array_index_781508 == array_index_773098 ? add_781816 : sel_781813;
  assign add_781820 = sel_781817 + 8'h01;
  assign sel_781821 = array_index_781508 == array_index_773104 ? add_781820 : sel_781817;
  assign add_781824 = sel_781821 + 8'h01;
  assign sel_781825 = array_index_781508 == array_index_773110 ? add_781824 : sel_781821;
  assign add_781828 = sel_781825 + 8'h01;
  assign sel_781829 = array_index_781508 == array_index_773116 ? add_781828 : sel_781825;
  assign add_781832 = sel_781829 + 8'h01;
  assign sel_781833 = array_index_781508 == array_index_773122 ? add_781832 : sel_781829;
  assign add_781836 = sel_781833 + 8'h01;
  assign sel_781837 = array_index_781508 == array_index_773128 ? add_781836 : sel_781833;
  assign add_781840 = sel_781837 + 8'h01;
  assign sel_781841 = array_index_781508 == array_index_773134 ? add_781840 : sel_781837;
  assign add_781844 = sel_781841 + 8'h01;
  assign sel_781845 = array_index_781508 == array_index_773140 ? add_781844 : sel_781841;
  assign add_781848 = sel_781845 + 8'h01;
  assign sel_781849 = array_index_781508 == array_index_773146 ? add_781848 : sel_781845;
  assign add_781852 = sel_781849 + 8'h01;
  assign sel_781853 = array_index_781508 == array_index_773152 ? add_781852 : sel_781849;
  assign add_781856 = sel_781853 + 8'h01;
  assign sel_781857 = array_index_781508 == array_index_773158 ? add_781856 : sel_781853;
  assign add_781860 = sel_781857 + 8'h01;
  assign sel_781861 = array_index_781508 == array_index_773164 ? add_781860 : sel_781857;
  assign add_781864 = sel_781861 + 8'h01;
  assign sel_781865 = array_index_781508 == array_index_773170 ? add_781864 : sel_781861;
  assign add_781869 = sel_781865 + 8'h01;
  assign array_index_781870 = set1_unflattened[7'h19];
  assign sel_781871 = array_index_781508 == array_index_773176 ? add_781869 : sel_781865;
  assign add_781874 = sel_781871 + 8'h01;
  assign sel_781875 = array_index_781870 == array_index_772632 ? add_781874 : sel_781871;
  assign add_781878 = sel_781875 + 8'h01;
  assign sel_781879 = array_index_781870 == array_index_772636 ? add_781878 : sel_781875;
  assign add_781882 = sel_781879 + 8'h01;
  assign sel_781883 = array_index_781870 == array_index_772644 ? add_781882 : sel_781879;
  assign add_781886 = sel_781883 + 8'h01;
  assign sel_781887 = array_index_781870 == array_index_772652 ? add_781886 : sel_781883;
  assign add_781890 = sel_781887 + 8'h01;
  assign sel_781891 = array_index_781870 == array_index_772660 ? add_781890 : sel_781887;
  assign add_781894 = sel_781891 + 8'h01;
  assign sel_781895 = array_index_781870 == array_index_772668 ? add_781894 : sel_781891;
  assign add_781898 = sel_781895 + 8'h01;
  assign sel_781899 = array_index_781870 == array_index_772676 ? add_781898 : sel_781895;
  assign add_781902 = sel_781899 + 8'h01;
  assign sel_781903 = array_index_781870 == array_index_772684 ? add_781902 : sel_781899;
  assign add_781906 = sel_781903 + 8'h01;
  assign sel_781907 = array_index_781870 == array_index_772690 ? add_781906 : sel_781903;
  assign add_781910 = sel_781907 + 8'h01;
  assign sel_781911 = array_index_781870 == array_index_772696 ? add_781910 : sel_781907;
  assign add_781914 = sel_781911 + 8'h01;
  assign sel_781915 = array_index_781870 == array_index_772702 ? add_781914 : sel_781911;
  assign add_781918 = sel_781915 + 8'h01;
  assign sel_781919 = array_index_781870 == array_index_772708 ? add_781918 : sel_781915;
  assign add_781922 = sel_781919 + 8'h01;
  assign sel_781923 = array_index_781870 == array_index_772714 ? add_781922 : sel_781919;
  assign add_781926 = sel_781923 + 8'h01;
  assign sel_781927 = array_index_781870 == array_index_772720 ? add_781926 : sel_781923;
  assign add_781930 = sel_781927 + 8'h01;
  assign sel_781931 = array_index_781870 == array_index_772726 ? add_781930 : sel_781927;
  assign add_781934 = sel_781931 + 8'h01;
  assign sel_781935 = array_index_781870 == array_index_772732 ? add_781934 : sel_781931;
  assign add_781938 = sel_781935 + 8'h01;
  assign sel_781939 = array_index_781870 == array_index_772738 ? add_781938 : sel_781935;
  assign add_781942 = sel_781939 + 8'h01;
  assign sel_781943 = array_index_781870 == array_index_772744 ? add_781942 : sel_781939;
  assign add_781946 = sel_781943 + 8'h01;
  assign sel_781947 = array_index_781870 == array_index_772750 ? add_781946 : sel_781943;
  assign add_781950 = sel_781947 + 8'h01;
  assign sel_781951 = array_index_781870 == array_index_772756 ? add_781950 : sel_781947;
  assign add_781954 = sel_781951 + 8'h01;
  assign sel_781955 = array_index_781870 == array_index_772762 ? add_781954 : sel_781951;
  assign add_781958 = sel_781955 + 8'h01;
  assign sel_781959 = array_index_781870 == array_index_772768 ? add_781958 : sel_781955;
  assign add_781962 = sel_781959 + 8'h01;
  assign sel_781963 = array_index_781870 == array_index_772774 ? add_781962 : sel_781959;
  assign add_781966 = sel_781963 + 8'h01;
  assign sel_781967 = array_index_781870 == array_index_772780 ? add_781966 : sel_781963;
  assign add_781970 = sel_781967 + 8'h01;
  assign sel_781971 = array_index_781870 == array_index_772786 ? add_781970 : sel_781967;
  assign add_781974 = sel_781971 + 8'h01;
  assign sel_781975 = array_index_781870 == array_index_772792 ? add_781974 : sel_781971;
  assign add_781978 = sel_781975 + 8'h01;
  assign sel_781979 = array_index_781870 == array_index_772798 ? add_781978 : sel_781975;
  assign add_781982 = sel_781979 + 8'h01;
  assign sel_781983 = array_index_781870 == array_index_772804 ? add_781982 : sel_781979;
  assign add_781986 = sel_781983 + 8'h01;
  assign sel_781987 = array_index_781870 == array_index_772810 ? add_781986 : sel_781983;
  assign add_781990 = sel_781987 + 8'h01;
  assign sel_781991 = array_index_781870 == array_index_772816 ? add_781990 : sel_781987;
  assign add_781994 = sel_781991 + 8'h01;
  assign sel_781995 = array_index_781870 == array_index_772822 ? add_781994 : sel_781991;
  assign add_781998 = sel_781995 + 8'h01;
  assign sel_781999 = array_index_781870 == array_index_772828 ? add_781998 : sel_781995;
  assign add_782002 = sel_781999 + 8'h01;
  assign sel_782003 = array_index_781870 == array_index_772834 ? add_782002 : sel_781999;
  assign add_782006 = sel_782003 + 8'h01;
  assign sel_782007 = array_index_781870 == array_index_772840 ? add_782006 : sel_782003;
  assign add_782010 = sel_782007 + 8'h01;
  assign sel_782011 = array_index_781870 == array_index_772846 ? add_782010 : sel_782007;
  assign add_782014 = sel_782011 + 8'h01;
  assign sel_782015 = array_index_781870 == array_index_772852 ? add_782014 : sel_782011;
  assign add_782018 = sel_782015 + 8'h01;
  assign sel_782019 = array_index_781870 == array_index_772858 ? add_782018 : sel_782015;
  assign add_782022 = sel_782019 + 8'h01;
  assign sel_782023 = array_index_781870 == array_index_772864 ? add_782022 : sel_782019;
  assign add_782026 = sel_782023 + 8'h01;
  assign sel_782027 = array_index_781870 == array_index_772870 ? add_782026 : sel_782023;
  assign add_782030 = sel_782027 + 8'h01;
  assign sel_782031 = array_index_781870 == array_index_772876 ? add_782030 : sel_782027;
  assign add_782034 = sel_782031 + 8'h01;
  assign sel_782035 = array_index_781870 == array_index_772882 ? add_782034 : sel_782031;
  assign add_782038 = sel_782035 + 8'h01;
  assign sel_782039 = array_index_781870 == array_index_772888 ? add_782038 : sel_782035;
  assign add_782042 = sel_782039 + 8'h01;
  assign sel_782043 = array_index_781870 == array_index_772894 ? add_782042 : sel_782039;
  assign add_782046 = sel_782043 + 8'h01;
  assign sel_782047 = array_index_781870 == array_index_772900 ? add_782046 : sel_782043;
  assign add_782050 = sel_782047 + 8'h01;
  assign sel_782051 = array_index_781870 == array_index_772906 ? add_782050 : sel_782047;
  assign add_782054 = sel_782051 + 8'h01;
  assign sel_782055 = array_index_781870 == array_index_772912 ? add_782054 : sel_782051;
  assign add_782058 = sel_782055 + 8'h01;
  assign sel_782059 = array_index_781870 == array_index_772918 ? add_782058 : sel_782055;
  assign add_782062 = sel_782059 + 8'h01;
  assign sel_782063 = array_index_781870 == array_index_772924 ? add_782062 : sel_782059;
  assign add_782066 = sel_782063 + 8'h01;
  assign sel_782067 = array_index_781870 == array_index_772930 ? add_782066 : sel_782063;
  assign add_782070 = sel_782067 + 8'h01;
  assign sel_782071 = array_index_781870 == array_index_772936 ? add_782070 : sel_782067;
  assign add_782074 = sel_782071 + 8'h01;
  assign sel_782075 = array_index_781870 == array_index_772942 ? add_782074 : sel_782071;
  assign add_782078 = sel_782075 + 8'h01;
  assign sel_782079 = array_index_781870 == array_index_772948 ? add_782078 : sel_782075;
  assign add_782082 = sel_782079 + 8'h01;
  assign sel_782083 = array_index_781870 == array_index_772954 ? add_782082 : sel_782079;
  assign add_782086 = sel_782083 + 8'h01;
  assign sel_782087 = array_index_781870 == array_index_772960 ? add_782086 : sel_782083;
  assign add_782090 = sel_782087 + 8'h01;
  assign sel_782091 = array_index_781870 == array_index_772966 ? add_782090 : sel_782087;
  assign add_782094 = sel_782091 + 8'h01;
  assign sel_782095 = array_index_781870 == array_index_772972 ? add_782094 : sel_782091;
  assign add_782098 = sel_782095 + 8'h01;
  assign sel_782099 = array_index_781870 == array_index_772978 ? add_782098 : sel_782095;
  assign add_782102 = sel_782099 + 8'h01;
  assign sel_782103 = array_index_781870 == array_index_772984 ? add_782102 : sel_782099;
  assign add_782106 = sel_782103 + 8'h01;
  assign sel_782107 = array_index_781870 == array_index_772990 ? add_782106 : sel_782103;
  assign add_782110 = sel_782107 + 8'h01;
  assign sel_782111 = array_index_781870 == array_index_772996 ? add_782110 : sel_782107;
  assign add_782114 = sel_782111 + 8'h01;
  assign sel_782115 = array_index_781870 == array_index_773002 ? add_782114 : sel_782111;
  assign add_782118 = sel_782115 + 8'h01;
  assign sel_782119 = array_index_781870 == array_index_773008 ? add_782118 : sel_782115;
  assign add_782122 = sel_782119 + 8'h01;
  assign sel_782123 = array_index_781870 == array_index_773014 ? add_782122 : sel_782119;
  assign add_782126 = sel_782123 + 8'h01;
  assign sel_782127 = array_index_781870 == array_index_773020 ? add_782126 : sel_782123;
  assign add_782130 = sel_782127 + 8'h01;
  assign sel_782131 = array_index_781870 == array_index_773026 ? add_782130 : sel_782127;
  assign add_782134 = sel_782131 + 8'h01;
  assign sel_782135 = array_index_781870 == array_index_773032 ? add_782134 : sel_782131;
  assign add_782138 = sel_782135 + 8'h01;
  assign sel_782139 = array_index_781870 == array_index_773038 ? add_782138 : sel_782135;
  assign add_782142 = sel_782139 + 8'h01;
  assign sel_782143 = array_index_781870 == array_index_773044 ? add_782142 : sel_782139;
  assign add_782146 = sel_782143 + 8'h01;
  assign sel_782147 = array_index_781870 == array_index_773050 ? add_782146 : sel_782143;
  assign add_782150 = sel_782147 + 8'h01;
  assign sel_782151 = array_index_781870 == array_index_773056 ? add_782150 : sel_782147;
  assign add_782154 = sel_782151 + 8'h01;
  assign sel_782155 = array_index_781870 == array_index_773062 ? add_782154 : sel_782151;
  assign add_782158 = sel_782155 + 8'h01;
  assign sel_782159 = array_index_781870 == array_index_773068 ? add_782158 : sel_782155;
  assign add_782162 = sel_782159 + 8'h01;
  assign sel_782163 = array_index_781870 == array_index_773074 ? add_782162 : sel_782159;
  assign add_782166 = sel_782163 + 8'h01;
  assign sel_782167 = array_index_781870 == array_index_773080 ? add_782166 : sel_782163;
  assign add_782170 = sel_782167 + 8'h01;
  assign sel_782171 = array_index_781870 == array_index_773086 ? add_782170 : sel_782167;
  assign add_782174 = sel_782171 + 8'h01;
  assign sel_782175 = array_index_781870 == array_index_773092 ? add_782174 : sel_782171;
  assign add_782178 = sel_782175 + 8'h01;
  assign sel_782179 = array_index_781870 == array_index_773098 ? add_782178 : sel_782175;
  assign add_782182 = sel_782179 + 8'h01;
  assign sel_782183 = array_index_781870 == array_index_773104 ? add_782182 : sel_782179;
  assign add_782186 = sel_782183 + 8'h01;
  assign sel_782187 = array_index_781870 == array_index_773110 ? add_782186 : sel_782183;
  assign add_782190 = sel_782187 + 8'h01;
  assign sel_782191 = array_index_781870 == array_index_773116 ? add_782190 : sel_782187;
  assign add_782194 = sel_782191 + 8'h01;
  assign sel_782195 = array_index_781870 == array_index_773122 ? add_782194 : sel_782191;
  assign add_782198 = sel_782195 + 8'h01;
  assign sel_782199 = array_index_781870 == array_index_773128 ? add_782198 : sel_782195;
  assign add_782202 = sel_782199 + 8'h01;
  assign sel_782203 = array_index_781870 == array_index_773134 ? add_782202 : sel_782199;
  assign add_782206 = sel_782203 + 8'h01;
  assign sel_782207 = array_index_781870 == array_index_773140 ? add_782206 : sel_782203;
  assign add_782210 = sel_782207 + 8'h01;
  assign sel_782211 = array_index_781870 == array_index_773146 ? add_782210 : sel_782207;
  assign add_782214 = sel_782211 + 8'h01;
  assign sel_782215 = array_index_781870 == array_index_773152 ? add_782214 : sel_782211;
  assign add_782218 = sel_782215 + 8'h01;
  assign sel_782219 = array_index_781870 == array_index_773158 ? add_782218 : sel_782215;
  assign add_782222 = sel_782219 + 8'h01;
  assign sel_782223 = array_index_781870 == array_index_773164 ? add_782222 : sel_782219;
  assign add_782226 = sel_782223 + 8'h01;
  assign sel_782227 = array_index_781870 == array_index_773170 ? add_782226 : sel_782223;
  assign add_782231 = sel_782227 + 8'h01;
  assign array_index_782232 = set1_unflattened[7'h1a];
  assign sel_782233 = array_index_781870 == array_index_773176 ? add_782231 : sel_782227;
  assign add_782236 = sel_782233 + 8'h01;
  assign sel_782237 = array_index_782232 == array_index_772632 ? add_782236 : sel_782233;
  assign add_782240 = sel_782237 + 8'h01;
  assign sel_782241 = array_index_782232 == array_index_772636 ? add_782240 : sel_782237;
  assign add_782244 = sel_782241 + 8'h01;
  assign sel_782245 = array_index_782232 == array_index_772644 ? add_782244 : sel_782241;
  assign add_782248 = sel_782245 + 8'h01;
  assign sel_782249 = array_index_782232 == array_index_772652 ? add_782248 : sel_782245;
  assign add_782252 = sel_782249 + 8'h01;
  assign sel_782253 = array_index_782232 == array_index_772660 ? add_782252 : sel_782249;
  assign add_782256 = sel_782253 + 8'h01;
  assign sel_782257 = array_index_782232 == array_index_772668 ? add_782256 : sel_782253;
  assign add_782260 = sel_782257 + 8'h01;
  assign sel_782261 = array_index_782232 == array_index_772676 ? add_782260 : sel_782257;
  assign add_782264 = sel_782261 + 8'h01;
  assign sel_782265 = array_index_782232 == array_index_772684 ? add_782264 : sel_782261;
  assign add_782268 = sel_782265 + 8'h01;
  assign sel_782269 = array_index_782232 == array_index_772690 ? add_782268 : sel_782265;
  assign add_782272 = sel_782269 + 8'h01;
  assign sel_782273 = array_index_782232 == array_index_772696 ? add_782272 : sel_782269;
  assign add_782276 = sel_782273 + 8'h01;
  assign sel_782277 = array_index_782232 == array_index_772702 ? add_782276 : sel_782273;
  assign add_782280 = sel_782277 + 8'h01;
  assign sel_782281 = array_index_782232 == array_index_772708 ? add_782280 : sel_782277;
  assign add_782284 = sel_782281 + 8'h01;
  assign sel_782285 = array_index_782232 == array_index_772714 ? add_782284 : sel_782281;
  assign add_782288 = sel_782285 + 8'h01;
  assign sel_782289 = array_index_782232 == array_index_772720 ? add_782288 : sel_782285;
  assign add_782292 = sel_782289 + 8'h01;
  assign sel_782293 = array_index_782232 == array_index_772726 ? add_782292 : sel_782289;
  assign add_782296 = sel_782293 + 8'h01;
  assign sel_782297 = array_index_782232 == array_index_772732 ? add_782296 : sel_782293;
  assign add_782300 = sel_782297 + 8'h01;
  assign sel_782301 = array_index_782232 == array_index_772738 ? add_782300 : sel_782297;
  assign add_782304 = sel_782301 + 8'h01;
  assign sel_782305 = array_index_782232 == array_index_772744 ? add_782304 : sel_782301;
  assign add_782308 = sel_782305 + 8'h01;
  assign sel_782309 = array_index_782232 == array_index_772750 ? add_782308 : sel_782305;
  assign add_782312 = sel_782309 + 8'h01;
  assign sel_782313 = array_index_782232 == array_index_772756 ? add_782312 : sel_782309;
  assign add_782316 = sel_782313 + 8'h01;
  assign sel_782317 = array_index_782232 == array_index_772762 ? add_782316 : sel_782313;
  assign add_782320 = sel_782317 + 8'h01;
  assign sel_782321 = array_index_782232 == array_index_772768 ? add_782320 : sel_782317;
  assign add_782324 = sel_782321 + 8'h01;
  assign sel_782325 = array_index_782232 == array_index_772774 ? add_782324 : sel_782321;
  assign add_782328 = sel_782325 + 8'h01;
  assign sel_782329 = array_index_782232 == array_index_772780 ? add_782328 : sel_782325;
  assign add_782332 = sel_782329 + 8'h01;
  assign sel_782333 = array_index_782232 == array_index_772786 ? add_782332 : sel_782329;
  assign add_782336 = sel_782333 + 8'h01;
  assign sel_782337 = array_index_782232 == array_index_772792 ? add_782336 : sel_782333;
  assign add_782340 = sel_782337 + 8'h01;
  assign sel_782341 = array_index_782232 == array_index_772798 ? add_782340 : sel_782337;
  assign add_782344 = sel_782341 + 8'h01;
  assign sel_782345 = array_index_782232 == array_index_772804 ? add_782344 : sel_782341;
  assign add_782348 = sel_782345 + 8'h01;
  assign sel_782349 = array_index_782232 == array_index_772810 ? add_782348 : sel_782345;
  assign add_782352 = sel_782349 + 8'h01;
  assign sel_782353 = array_index_782232 == array_index_772816 ? add_782352 : sel_782349;
  assign add_782356 = sel_782353 + 8'h01;
  assign sel_782357 = array_index_782232 == array_index_772822 ? add_782356 : sel_782353;
  assign add_782360 = sel_782357 + 8'h01;
  assign sel_782361 = array_index_782232 == array_index_772828 ? add_782360 : sel_782357;
  assign add_782364 = sel_782361 + 8'h01;
  assign sel_782365 = array_index_782232 == array_index_772834 ? add_782364 : sel_782361;
  assign add_782368 = sel_782365 + 8'h01;
  assign sel_782369 = array_index_782232 == array_index_772840 ? add_782368 : sel_782365;
  assign add_782372 = sel_782369 + 8'h01;
  assign sel_782373 = array_index_782232 == array_index_772846 ? add_782372 : sel_782369;
  assign add_782376 = sel_782373 + 8'h01;
  assign sel_782377 = array_index_782232 == array_index_772852 ? add_782376 : sel_782373;
  assign add_782380 = sel_782377 + 8'h01;
  assign sel_782381 = array_index_782232 == array_index_772858 ? add_782380 : sel_782377;
  assign add_782384 = sel_782381 + 8'h01;
  assign sel_782385 = array_index_782232 == array_index_772864 ? add_782384 : sel_782381;
  assign add_782388 = sel_782385 + 8'h01;
  assign sel_782389 = array_index_782232 == array_index_772870 ? add_782388 : sel_782385;
  assign add_782392 = sel_782389 + 8'h01;
  assign sel_782393 = array_index_782232 == array_index_772876 ? add_782392 : sel_782389;
  assign add_782396 = sel_782393 + 8'h01;
  assign sel_782397 = array_index_782232 == array_index_772882 ? add_782396 : sel_782393;
  assign add_782400 = sel_782397 + 8'h01;
  assign sel_782401 = array_index_782232 == array_index_772888 ? add_782400 : sel_782397;
  assign add_782404 = sel_782401 + 8'h01;
  assign sel_782405 = array_index_782232 == array_index_772894 ? add_782404 : sel_782401;
  assign add_782408 = sel_782405 + 8'h01;
  assign sel_782409 = array_index_782232 == array_index_772900 ? add_782408 : sel_782405;
  assign add_782412 = sel_782409 + 8'h01;
  assign sel_782413 = array_index_782232 == array_index_772906 ? add_782412 : sel_782409;
  assign add_782416 = sel_782413 + 8'h01;
  assign sel_782417 = array_index_782232 == array_index_772912 ? add_782416 : sel_782413;
  assign add_782420 = sel_782417 + 8'h01;
  assign sel_782421 = array_index_782232 == array_index_772918 ? add_782420 : sel_782417;
  assign add_782424 = sel_782421 + 8'h01;
  assign sel_782425 = array_index_782232 == array_index_772924 ? add_782424 : sel_782421;
  assign add_782428 = sel_782425 + 8'h01;
  assign sel_782429 = array_index_782232 == array_index_772930 ? add_782428 : sel_782425;
  assign add_782432 = sel_782429 + 8'h01;
  assign sel_782433 = array_index_782232 == array_index_772936 ? add_782432 : sel_782429;
  assign add_782436 = sel_782433 + 8'h01;
  assign sel_782437 = array_index_782232 == array_index_772942 ? add_782436 : sel_782433;
  assign add_782440 = sel_782437 + 8'h01;
  assign sel_782441 = array_index_782232 == array_index_772948 ? add_782440 : sel_782437;
  assign add_782444 = sel_782441 + 8'h01;
  assign sel_782445 = array_index_782232 == array_index_772954 ? add_782444 : sel_782441;
  assign add_782448 = sel_782445 + 8'h01;
  assign sel_782449 = array_index_782232 == array_index_772960 ? add_782448 : sel_782445;
  assign add_782452 = sel_782449 + 8'h01;
  assign sel_782453 = array_index_782232 == array_index_772966 ? add_782452 : sel_782449;
  assign add_782456 = sel_782453 + 8'h01;
  assign sel_782457 = array_index_782232 == array_index_772972 ? add_782456 : sel_782453;
  assign add_782460 = sel_782457 + 8'h01;
  assign sel_782461 = array_index_782232 == array_index_772978 ? add_782460 : sel_782457;
  assign add_782464 = sel_782461 + 8'h01;
  assign sel_782465 = array_index_782232 == array_index_772984 ? add_782464 : sel_782461;
  assign add_782468 = sel_782465 + 8'h01;
  assign sel_782469 = array_index_782232 == array_index_772990 ? add_782468 : sel_782465;
  assign add_782472 = sel_782469 + 8'h01;
  assign sel_782473 = array_index_782232 == array_index_772996 ? add_782472 : sel_782469;
  assign add_782476 = sel_782473 + 8'h01;
  assign sel_782477 = array_index_782232 == array_index_773002 ? add_782476 : sel_782473;
  assign add_782480 = sel_782477 + 8'h01;
  assign sel_782481 = array_index_782232 == array_index_773008 ? add_782480 : sel_782477;
  assign add_782484 = sel_782481 + 8'h01;
  assign sel_782485 = array_index_782232 == array_index_773014 ? add_782484 : sel_782481;
  assign add_782488 = sel_782485 + 8'h01;
  assign sel_782489 = array_index_782232 == array_index_773020 ? add_782488 : sel_782485;
  assign add_782492 = sel_782489 + 8'h01;
  assign sel_782493 = array_index_782232 == array_index_773026 ? add_782492 : sel_782489;
  assign add_782496 = sel_782493 + 8'h01;
  assign sel_782497 = array_index_782232 == array_index_773032 ? add_782496 : sel_782493;
  assign add_782500 = sel_782497 + 8'h01;
  assign sel_782501 = array_index_782232 == array_index_773038 ? add_782500 : sel_782497;
  assign add_782504 = sel_782501 + 8'h01;
  assign sel_782505 = array_index_782232 == array_index_773044 ? add_782504 : sel_782501;
  assign add_782508 = sel_782505 + 8'h01;
  assign sel_782509 = array_index_782232 == array_index_773050 ? add_782508 : sel_782505;
  assign add_782512 = sel_782509 + 8'h01;
  assign sel_782513 = array_index_782232 == array_index_773056 ? add_782512 : sel_782509;
  assign add_782516 = sel_782513 + 8'h01;
  assign sel_782517 = array_index_782232 == array_index_773062 ? add_782516 : sel_782513;
  assign add_782520 = sel_782517 + 8'h01;
  assign sel_782521 = array_index_782232 == array_index_773068 ? add_782520 : sel_782517;
  assign add_782524 = sel_782521 + 8'h01;
  assign sel_782525 = array_index_782232 == array_index_773074 ? add_782524 : sel_782521;
  assign add_782528 = sel_782525 + 8'h01;
  assign sel_782529 = array_index_782232 == array_index_773080 ? add_782528 : sel_782525;
  assign add_782532 = sel_782529 + 8'h01;
  assign sel_782533 = array_index_782232 == array_index_773086 ? add_782532 : sel_782529;
  assign add_782536 = sel_782533 + 8'h01;
  assign sel_782537 = array_index_782232 == array_index_773092 ? add_782536 : sel_782533;
  assign add_782540 = sel_782537 + 8'h01;
  assign sel_782541 = array_index_782232 == array_index_773098 ? add_782540 : sel_782537;
  assign add_782544 = sel_782541 + 8'h01;
  assign sel_782545 = array_index_782232 == array_index_773104 ? add_782544 : sel_782541;
  assign add_782548 = sel_782545 + 8'h01;
  assign sel_782549 = array_index_782232 == array_index_773110 ? add_782548 : sel_782545;
  assign add_782552 = sel_782549 + 8'h01;
  assign sel_782553 = array_index_782232 == array_index_773116 ? add_782552 : sel_782549;
  assign add_782556 = sel_782553 + 8'h01;
  assign sel_782557 = array_index_782232 == array_index_773122 ? add_782556 : sel_782553;
  assign add_782560 = sel_782557 + 8'h01;
  assign sel_782561 = array_index_782232 == array_index_773128 ? add_782560 : sel_782557;
  assign add_782564 = sel_782561 + 8'h01;
  assign sel_782565 = array_index_782232 == array_index_773134 ? add_782564 : sel_782561;
  assign add_782568 = sel_782565 + 8'h01;
  assign sel_782569 = array_index_782232 == array_index_773140 ? add_782568 : sel_782565;
  assign add_782572 = sel_782569 + 8'h01;
  assign sel_782573 = array_index_782232 == array_index_773146 ? add_782572 : sel_782569;
  assign add_782576 = sel_782573 + 8'h01;
  assign sel_782577 = array_index_782232 == array_index_773152 ? add_782576 : sel_782573;
  assign add_782580 = sel_782577 + 8'h01;
  assign sel_782581 = array_index_782232 == array_index_773158 ? add_782580 : sel_782577;
  assign add_782584 = sel_782581 + 8'h01;
  assign sel_782585 = array_index_782232 == array_index_773164 ? add_782584 : sel_782581;
  assign add_782588 = sel_782585 + 8'h01;
  assign sel_782589 = array_index_782232 == array_index_773170 ? add_782588 : sel_782585;
  assign add_782593 = sel_782589 + 8'h01;
  assign array_index_782594 = set1_unflattened[7'h1b];
  assign sel_782595 = array_index_782232 == array_index_773176 ? add_782593 : sel_782589;
  assign add_782598 = sel_782595 + 8'h01;
  assign sel_782599 = array_index_782594 == array_index_772632 ? add_782598 : sel_782595;
  assign add_782602 = sel_782599 + 8'h01;
  assign sel_782603 = array_index_782594 == array_index_772636 ? add_782602 : sel_782599;
  assign add_782606 = sel_782603 + 8'h01;
  assign sel_782607 = array_index_782594 == array_index_772644 ? add_782606 : sel_782603;
  assign add_782610 = sel_782607 + 8'h01;
  assign sel_782611 = array_index_782594 == array_index_772652 ? add_782610 : sel_782607;
  assign add_782614 = sel_782611 + 8'h01;
  assign sel_782615 = array_index_782594 == array_index_772660 ? add_782614 : sel_782611;
  assign add_782618 = sel_782615 + 8'h01;
  assign sel_782619 = array_index_782594 == array_index_772668 ? add_782618 : sel_782615;
  assign add_782622 = sel_782619 + 8'h01;
  assign sel_782623 = array_index_782594 == array_index_772676 ? add_782622 : sel_782619;
  assign add_782626 = sel_782623 + 8'h01;
  assign sel_782627 = array_index_782594 == array_index_772684 ? add_782626 : sel_782623;
  assign add_782630 = sel_782627 + 8'h01;
  assign sel_782631 = array_index_782594 == array_index_772690 ? add_782630 : sel_782627;
  assign add_782634 = sel_782631 + 8'h01;
  assign sel_782635 = array_index_782594 == array_index_772696 ? add_782634 : sel_782631;
  assign add_782638 = sel_782635 + 8'h01;
  assign sel_782639 = array_index_782594 == array_index_772702 ? add_782638 : sel_782635;
  assign add_782642 = sel_782639 + 8'h01;
  assign sel_782643 = array_index_782594 == array_index_772708 ? add_782642 : sel_782639;
  assign add_782646 = sel_782643 + 8'h01;
  assign sel_782647 = array_index_782594 == array_index_772714 ? add_782646 : sel_782643;
  assign add_782650 = sel_782647 + 8'h01;
  assign sel_782651 = array_index_782594 == array_index_772720 ? add_782650 : sel_782647;
  assign add_782654 = sel_782651 + 8'h01;
  assign sel_782655 = array_index_782594 == array_index_772726 ? add_782654 : sel_782651;
  assign add_782658 = sel_782655 + 8'h01;
  assign sel_782659 = array_index_782594 == array_index_772732 ? add_782658 : sel_782655;
  assign add_782662 = sel_782659 + 8'h01;
  assign sel_782663 = array_index_782594 == array_index_772738 ? add_782662 : sel_782659;
  assign add_782666 = sel_782663 + 8'h01;
  assign sel_782667 = array_index_782594 == array_index_772744 ? add_782666 : sel_782663;
  assign add_782670 = sel_782667 + 8'h01;
  assign sel_782671 = array_index_782594 == array_index_772750 ? add_782670 : sel_782667;
  assign add_782674 = sel_782671 + 8'h01;
  assign sel_782675 = array_index_782594 == array_index_772756 ? add_782674 : sel_782671;
  assign add_782678 = sel_782675 + 8'h01;
  assign sel_782679 = array_index_782594 == array_index_772762 ? add_782678 : sel_782675;
  assign add_782682 = sel_782679 + 8'h01;
  assign sel_782683 = array_index_782594 == array_index_772768 ? add_782682 : sel_782679;
  assign add_782686 = sel_782683 + 8'h01;
  assign sel_782687 = array_index_782594 == array_index_772774 ? add_782686 : sel_782683;
  assign add_782690 = sel_782687 + 8'h01;
  assign sel_782691 = array_index_782594 == array_index_772780 ? add_782690 : sel_782687;
  assign add_782694 = sel_782691 + 8'h01;
  assign sel_782695 = array_index_782594 == array_index_772786 ? add_782694 : sel_782691;
  assign add_782698 = sel_782695 + 8'h01;
  assign sel_782699 = array_index_782594 == array_index_772792 ? add_782698 : sel_782695;
  assign add_782702 = sel_782699 + 8'h01;
  assign sel_782703 = array_index_782594 == array_index_772798 ? add_782702 : sel_782699;
  assign add_782706 = sel_782703 + 8'h01;
  assign sel_782707 = array_index_782594 == array_index_772804 ? add_782706 : sel_782703;
  assign add_782710 = sel_782707 + 8'h01;
  assign sel_782711 = array_index_782594 == array_index_772810 ? add_782710 : sel_782707;
  assign add_782714 = sel_782711 + 8'h01;
  assign sel_782715 = array_index_782594 == array_index_772816 ? add_782714 : sel_782711;
  assign add_782718 = sel_782715 + 8'h01;
  assign sel_782719 = array_index_782594 == array_index_772822 ? add_782718 : sel_782715;
  assign add_782722 = sel_782719 + 8'h01;
  assign sel_782723 = array_index_782594 == array_index_772828 ? add_782722 : sel_782719;
  assign add_782726 = sel_782723 + 8'h01;
  assign sel_782727 = array_index_782594 == array_index_772834 ? add_782726 : sel_782723;
  assign add_782730 = sel_782727 + 8'h01;
  assign sel_782731 = array_index_782594 == array_index_772840 ? add_782730 : sel_782727;
  assign add_782734 = sel_782731 + 8'h01;
  assign sel_782735 = array_index_782594 == array_index_772846 ? add_782734 : sel_782731;
  assign add_782738 = sel_782735 + 8'h01;
  assign sel_782739 = array_index_782594 == array_index_772852 ? add_782738 : sel_782735;
  assign add_782742 = sel_782739 + 8'h01;
  assign sel_782743 = array_index_782594 == array_index_772858 ? add_782742 : sel_782739;
  assign add_782746 = sel_782743 + 8'h01;
  assign sel_782747 = array_index_782594 == array_index_772864 ? add_782746 : sel_782743;
  assign add_782750 = sel_782747 + 8'h01;
  assign sel_782751 = array_index_782594 == array_index_772870 ? add_782750 : sel_782747;
  assign add_782754 = sel_782751 + 8'h01;
  assign sel_782755 = array_index_782594 == array_index_772876 ? add_782754 : sel_782751;
  assign add_782758 = sel_782755 + 8'h01;
  assign sel_782759 = array_index_782594 == array_index_772882 ? add_782758 : sel_782755;
  assign add_782762 = sel_782759 + 8'h01;
  assign sel_782763 = array_index_782594 == array_index_772888 ? add_782762 : sel_782759;
  assign add_782766 = sel_782763 + 8'h01;
  assign sel_782767 = array_index_782594 == array_index_772894 ? add_782766 : sel_782763;
  assign add_782770 = sel_782767 + 8'h01;
  assign sel_782771 = array_index_782594 == array_index_772900 ? add_782770 : sel_782767;
  assign add_782774 = sel_782771 + 8'h01;
  assign sel_782775 = array_index_782594 == array_index_772906 ? add_782774 : sel_782771;
  assign add_782778 = sel_782775 + 8'h01;
  assign sel_782779 = array_index_782594 == array_index_772912 ? add_782778 : sel_782775;
  assign add_782782 = sel_782779 + 8'h01;
  assign sel_782783 = array_index_782594 == array_index_772918 ? add_782782 : sel_782779;
  assign add_782786 = sel_782783 + 8'h01;
  assign sel_782787 = array_index_782594 == array_index_772924 ? add_782786 : sel_782783;
  assign add_782790 = sel_782787 + 8'h01;
  assign sel_782791 = array_index_782594 == array_index_772930 ? add_782790 : sel_782787;
  assign add_782794 = sel_782791 + 8'h01;
  assign sel_782795 = array_index_782594 == array_index_772936 ? add_782794 : sel_782791;
  assign add_782798 = sel_782795 + 8'h01;
  assign sel_782799 = array_index_782594 == array_index_772942 ? add_782798 : sel_782795;
  assign add_782802 = sel_782799 + 8'h01;
  assign sel_782803 = array_index_782594 == array_index_772948 ? add_782802 : sel_782799;
  assign add_782806 = sel_782803 + 8'h01;
  assign sel_782807 = array_index_782594 == array_index_772954 ? add_782806 : sel_782803;
  assign add_782810 = sel_782807 + 8'h01;
  assign sel_782811 = array_index_782594 == array_index_772960 ? add_782810 : sel_782807;
  assign add_782814 = sel_782811 + 8'h01;
  assign sel_782815 = array_index_782594 == array_index_772966 ? add_782814 : sel_782811;
  assign add_782818 = sel_782815 + 8'h01;
  assign sel_782819 = array_index_782594 == array_index_772972 ? add_782818 : sel_782815;
  assign add_782822 = sel_782819 + 8'h01;
  assign sel_782823 = array_index_782594 == array_index_772978 ? add_782822 : sel_782819;
  assign add_782826 = sel_782823 + 8'h01;
  assign sel_782827 = array_index_782594 == array_index_772984 ? add_782826 : sel_782823;
  assign add_782830 = sel_782827 + 8'h01;
  assign sel_782831 = array_index_782594 == array_index_772990 ? add_782830 : sel_782827;
  assign add_782834 = sel_782831 + 8'h01;
  assign sel_782835 = array_index_782594 == array_index_772996 ? add_782834 : sel_782831;
  assign add_782838 = sel_782835 + 8'h01;
  assign sel_782839 = array_index_782594 == array_index_773002 ? add_782838 : sel_782835;
  assign add_782842 = sel_782839 + 8'h01;
  assign sel_782843 = array_index_782594 == array_index_773008 ? add_782842 : sel_782839;
  assign add_782846 = sel_782843 + 8'h01;
  assign sel_782847 = array_index_782594 == array_index_773014 ? add_782846 : sel_782843;
  assign add_782850 = sel_782847 + 8'h01;
  assign sel_782851 = array_index_782594 == array_index_773020 ? add_782850 : sel_782847;
  assign add_782854 = sel_782851 + 8'h01;
  assign sel_782855 = array_index_782594 == array_index_773026 ? add_782854 : sel_782851;
  assign add_782858 = sel_782855 + 8'h01;
  assign sel_782859 = array_index_782594 == array_index_773032 ? add_782858 : sel_782855;
  assign add_782862 = sel_782859 + 8'h01;
  assign sel_782863 = array_index_782594 == array_index_773038 ? add_782862 : sel_782859;
  assign add_782866 = sel_782863 + 8'h01;
  assign sel_782867 = array_index_782594 == array_index_773044 ? add_782866 : sel_782863;
  assign add_782870 = sel_782867 + 8'h01;
  assign sel_782871 = array_index_782594 == array_index_773050 ? add_782870 : sel_782867;
  assign add_782874 = sel_782871 + 8'h01;
  assign sel_782875 = array_index_782594 == array_index_773056 ? add_782874 : sel_782871;
  assign add_782878 = sel_782875 + 8'h01;
  assign sel_782879 = array_index_782594 == array_index_773062 ? add_782878 : sel_782875;
  assign add_782882 = sel_782879 + 8'h01;
  assign sel_782883 = array_index_782594 == array_index_773068 ? add_782882 : sel_782879;
  assign add_782886 = sel_782883 + 8'h01;
  assign sel_782887 = array_index_782594 == array_index_773074 ? add_782886 : sel_782883;
  assign add_782890 = sel_782887 + 8'h01;
  assign sel_782891 = array_index_782594 == array_index_773080 ? add_782890 : sel_782887;
  assign add_782894 = sel_782891 + 8'h01;
  assign sel_782895 = array_index_782594 == array_index_773086 ? add_782894 : sel_782891;
  assign add_782898 = sel_782895 + 8'h01;
  assign sel_782899 = array_index_782594 == array_index_773092 ? add_782898 : sel_782895;
  assign add_782902 = sel_782899 + 8'h01;
  assign sel_782903 = array_index_782594 == array_index_773098 ? add_782902 : sel_782899;
  assign add_782906 = sel_782903 + 8'h01;
  assign sel_782907 = array_index_782594 == array_index_773104 ? add_782906 : sel_782903;
  assign add_782910 = sel_782907 + 8'h01;
  assign sel_782911 = array_index_782594 == array_index_773110 ? add_782910 : sel_782907;
  assign add_782914 = sel_782911 + 8'h01;
  assign sel_782915 = array_index_782594 == array_index_773116 ? add_782914 : sel_782911;
  assign add_782918 = sel_782915 + 8'h01;
  assign sel_782919 = array_index_782594 == array_index_773122 ? add_782918 : sel_782915;
  assign add_782922 = sel_782919 + 8'h01;
  assign sel_782923 = array_index_782594 == array_index_773128 ? add_782922 : sel_782919;
  assign add_782926 = sel_782923 + 8'h01;
  assign sel_782927 = array_index_782594 == array_index_773134 ? add_782926 : sel_782923;
  assign add_782930 = sel_782927 + 8'h01;
  assign sel_782931 = array_index_782594 == array_index_773140 ? add_782930 : sel_782927;
  assign add_782934 = sel_782931 + 8'h01;
  assign sel_782935 = array_index_782594 == array_index_773146 ? add_782934 : sel_782931;
  assign add_782938 = sel_782935 + 8'h01;
  assign sel_782939 = array_index_782594 == array_index_773152 ? add_782938 : sel_782935;
  assign add_782942 = sel_782939 + 8'h01;
  assign sel_782943 = array_index_782594 == array_index_773158 ? add_782942 : sel_782939;
  assign add_782946 = sel_782943 + 8'h01;
  assign sel_782947 = array_index_782594 == array_index_773164 ? add_782946 : sel_782943;
  assign add_782950 = sel_782947 + 8'h01;
  assign sel_782951 = array_index_782594 == array_index_773170 ? add_782950 : sel_782947;
  assign add_782955 = sel_782951 + 8'h01;
  assign array_index_782956 = set1_unflattened[7'h1c];
  assign sel_782957 = array_index_782594 == array_index_773176 ? add_782955 : sel_782951;
  assign add_782960 = sel_782957 + 8'h01;
  assign sel_782961 = array_index_782956 == array_index_772632 ? add_782960 : sel_782957;
  assign add_782964 = sel_782961 + 8'h01;
  assign sel_782965 = array_index_782956 == array_index_772636 ? add_782964 : sel_782961;
  assign add_782968 = sel_782965 + 8'h01;
  assign sel_782969 = array_index_782956 == array_index_772644 ? add_782968 : sel_782965;
  assign add_782972 = sel_782969 + 8'h01;
  assign sel_782973 = array_index_782956 == array_index_772652 ? add_782972 : sel_782969;
  assign add_782976 = sel_782973 + 8'h01;
  assign sel_782977 = array_index_782956 == array_index_772660 ? add_782976 : sel_782973;
  assign add_782980 = sel_782977 + 8'h01;
  assign sel_782981 = array_index_782956 == array_index_772668 ? add_782980 : sel_782977;
  assign add_782984 = sel_782981 + 8'h01;
  assign sel_782985 = array_index_782956 == array_index_772676 ? add_782984 : sel_782981;
  assign add_782988 = sel_782985 + 8'h01;
  assign sel_782989 = array_index_782956 == array_index_772684 ? add_782988 : sel_782985;
  assign add_782992 = sel_782989 + 8'h01;
  assign sel_782993 = array_index_782956 == array_index_772690 ? add_782992 : sel_782989;
  assign add_782996 = sel_782993 + 8'h01;
  assign sel_782997 = array_index_782956 == array_index_772696 ? add_782996 : sel_782993;
  assign add_783000 = sel_782997 + 8'h01;
  assign sel_783001 = array_index_782956 == array_index_772702 ? add_783000 : sel_782997;
  assign add_783004 = sel_783001 + 8'h01;
  assign sel_783005 = array_index_782956 == array_index_772708 ? add_783004 : sel_783001;
  assign add_783008 = sel_783005 + 8'h01;
  assign sel_783009 = array_index_782956 == array_index_772714 ? add_783008 : sel_783005;
  assign add_783012 = sel_783009 + 8'h01;
  assign sel_783013 = array_index_782956 == array_index_772720 ? add_783012 : sel_783009;
  assign add_783016 = sel_783013 + 8'h01;
  assign sel_783017 = array_index_782956 == array_index_772726 ? add_783016 : sel_783013;
  assign add_783020 = sel_783017 + 8'h01;
  assign sel_783021 = array_index_782956 == array_index_772732 ? add_783020 : sel_783017;
  assign add_783024 = sel_783021 + 8'h01;
  assign sel_783025 = array_index_782956 == array_index_772738 ? add_783024 : sel_783021;
  assign add_783028 = sel_783025 + 8'h01;
  assign sel_783029 = array_index_782956 == array_index_772744 ? add_783028 : sel_783025;
  assign add_783032 = sel_783029 + 8'h01;
  assign sel_783033 = array_index_782956 == array_index_772750 ? add_783032 : sel_783029;
  assign add_783036 = sel_783033 + 8'h01;
  assign sel_783037 = array_index_782956 == array_index_772756 ? add_783036 : sel_783033;
  assign add_783040 = sel_783037 + 8'h01;
  assign sel_783041 = array_index_782956 == array_index_772762 ? add_783040 : sel_783037;
  assign add_783044 = sel_783041 + 8'h01;
  assign sel_783045 = array_index_782956 == array_index_772768 ? add_783044 : sel_783041;
  assign add_783048 = sel_783045 + 8'h01;
  assign sel_783049 = array_index_782956 == array_index_772774 ? add_783048 : sel_783045;
  assign add_783052 = sel_783049 + 8'h01;
  assign sel_783053 = array_index_782956 == array_index_772780 ? add_783052 : sel_783049;
  assign add_783056 = sel_783053 + 8'h01;
  assign sel_783057 = array_index_782956 == array_index_772786 ? add_783056 : sel_783053;
  assign add_783060 = sel_783057 + 8'h01;
  assign sel_783061 = array_index_782956 == array_index_772792 ? add_783060 : sel_783057;
  assign add_783064 = sel_783061 + 8'h01;
  assign sel_783065 = array_index_782956 == array_index_772798 ? add_783064 : sel_783061;
  assign add_783068 = sel_783065 + 8'h01;
  assign sel_783069 = array_index_782956 == array_index_772804 ? add_783068 : sel_783065;
  assign add_783072 = sel_783069 + 8'h01;
  assign sel_783073 = array_index_782956 == array_index_772810 ? add_783072 : sel_783069;
  assign add_783076 = sel_783073 + 8'h01;
  assign sel_783077 = array_index_782956 == array_index_772816 ? add_783076 : sel_783073;
  assign add_783080 = sel_783077 + 8'h01;
  assign sel_783081 = array_index_782956 == array_index_772822 ? add_783080 : sel_783077;
  assign add_783084 = sel_783081 + 8'h01;
  assign sel_783085 = array_index_782956 == array_index_772828 ? add_783084 : sel_783081;
  assign add_783088 = sel_783085 + 8'h01;
  assign sel_783089 = array_index_782956 == array_index_772834 ? add_783088 : sel_783085;
  assign add_783092 = sel_783089 + 8'h01;
  assign sel_783093 = array_index_782956 == array_index_772840 ? add_783092 : sel_783089;
  assign add_783096 = sel_783093 + 8'h01;
  assign sel_783097 = array_index_782956 == array_index_772846 ? add_783096 : sel_783093;
  assign add_783100 = sel_783097 + 8'h01;
  assign sel_783101 = array_index_782956 == array_index_772852 ? add_783100 : sel_783097;
  assign add_783104 = sel_783101 + 8'h01;
  assign sel_783105 = array_index_782956 == array_index_772858 ? add_783104 : sel_783101;
  assign add_783108 = sel_783105 + 8'h01;
  assign sel_783109 = array_index_782956 == array_index_772864 ? add_783108 : sel_783105;
  assign add_783112 = sel_783109 + 8'h01;
  assign sel_783113 = array_index_782956 == array_index_772870 ? add_783112 : sel_783109;
  assign add_783116 = sel_783113 + 8'h01;
  assign sel_783117 = array_index_782956 == array_index_772876 ? add_783116 : sel_783113;
  assign add_783120 = sel_783117 + 8'h01;
  assign sel_783121 = array_index_782956 == array_index_772882 ? add_783120 : sel_783117;
  assign add_783124 = sel_783121 + 8'h01;
  assign sel_783125 = array_index_782956 == array_index_772888 ? add_783124 : sel_783121;
  assign add_783128 = sel_783125 + 8'h01;
  assign sel_783129 = array_index_782956 == array_index_772894 ? add_783128 : sel_783125;
  assign add_783132 = sel_783129 + 8'h01;
  assign sel_783133 = array_index_782956 == array_index_772900 ? add_783132 : sel_783129;
  assign add_783136 = sel_783133 + 8'h01;
  assign sel_783137 = array_index_782956 == array_index_772906 ? add_783136 : sel_783133;
  assign add_783140 = sel_783137 + 8'h01;
  assign sel_783141 = array_index_782956 == array_index_772912 ? add_783140 : sel_783137;
  assign add_783144 = sel_783141 + 8'h01;
  assign sel_783145 = array_index_782956 == array_index_772918 ? add_783144 : sel_783141;
  assign add_783148 = sel_783145 + 8'h01;
  assign sel_783149 = array_index_782956 == array_index_772924 ? add_783148 : sel_783145;
  assign add_783152 = sel_783149 + 8'h01;
  assign sel_783153 = array_index_782956 == array_index_772930 ? add_783152 : sel_783149;
  assign add_783156 = sel_783153 + 8'h01;
  assign sel_783157 = array_index_782956 == array_index_772936 ? add_783156 : sel_783153;
  assign add_783160 = sel_783157 + 8'h01;
  assign sel_783161 = array_index_782956 == array_index_772942 ? add_783160 : sel_783157;
  assign add_783164 = sel_783161 + 8'h01;
  assign sel_783165 = array_index_782956 == array_index_772948 ? add_783164 : sel_783161;
  assign add_783168 = sel_783165 + 8'h01;
  assign sel_783169 = array_index_782956 == array_index_772954 ? add_783168 : sel_783165;
  assign add_783172 = sel_783169 + 8'h01;
  assign sel_783173 = array_index_782956 == array_index_772960 ? add_783172 : sel_783169;
  assign add_783176 = sel_783173 + 8'h01;
  assign sel_783177 = array_index_782956 == array_index_772966 ? add_783176 : sel_783173;
  assign add_783180 = sel_783177 + 8'h01;
  assign sel_783181 = array_index_782956 == array_index_772972 ? add_783180 : sel_783177;
  assign add_783184 = sel_783181 + 8'h01;
  assign sel_783185 = array_index_782956 == array_index_772978 ? add_783184 : sel_783181;
  assign add_783188 = sel_783185 + 8'h01;
  assign sel_783189 = array_index_782956 == array_index_772984 ? add_783188 : sel_783185;
  assign add_783192 = sel_783189 + 8'h01;
  assign sel_783193 = array_index_782956 == array_index_772990 ? add_783192 : sel_783189;
  assign add_783196 = sel_783193 + 8'h01;
  assign sel_783197 = array_index_782956 == array_index_772996 ? add_783196 : sel_783193;
  assign add_783200 = sel_783197 + 8'h01;
  assign sel_783201 = array_index_782956 == array_index_773002 ? add_783200 : sel_783197;
  assign add_783204 = sel_783201 + 8'h01;
  assign sel_783205 = array_index_782956 == array_index_773008 ? add_783204 : sel_783201;
  assign add_783208 = sel_783205 + 8'h01;
  assign sel_783209 = array_index_782956 == array_index_773014 ? add_783208 : sel_783205;
  assign add_783212 = sel_783209 + 8'h01;
  assign sel_783213 = array_index_782956 == array_index_773020 ? add_783212 : sel_783209;
  assign add_783216 = sel_783213 + 8'h01;
  assign sel_783217 = array_index_782956 == array_index_773026 ? add_783216 : sel_783213;
  assign add_783220 = sel_783217 + 8'h01;
  assign sel_783221 = array_index_782956 == array_index_773032 ? add_783220 : sel_783217;
  assign add_783224 = sel_783221 + 8'h01;
  assign sel_783225 = array_index_782956 == array_index_773038 ? add_783224 : sel_783221;
  assign add_783228 = sel_783225 + 8'h01;
  assign sel_783229 = array_index_782956 == array_index_773044 ? add_783228 : sel_783225;
  assign add_783232 = sel_783229 + 8'h01;
  assign sel_783233 = array_index_782956 == array_index_773050 ? add_783232 : sel_783229;
  assign add_783236 = sel_783233 + 8'h01;
  assign sel_783237 = array_index_782956 == array_index_773056 ? add_783236 : sel_783233;
  assign add_783240 = sel_783237 + 8'h01;
  assign sel_783241 = array_index_782956 == array_index_773062 ? add_783240 : sel_783237;
  assign add_783244 = sel_783241 + 8'h01;
  assign sel_783245 = array_index_782956 == array_index_773068 ? add_783244 : sel_783241;
  assign add_783248 = sel_783245 + 8'h01;
  assign sel_783249 = array_index_782956 == array_index_773074 ? add_783248 : sel_783245;
  assign add_783252 = sel_783249 + 8'h01;
  assign sel_783253 = array_index_782956 == array_index_773080 ? add_783252 : sel_783249;
  assign add_783256 = sel_783253 + 8'h01;
  assign sel_783257 = array_index_782956 == array_index_773086 ? add_783256 : sel_783253;
  assign add_783260 = sel_783257 + 8'h01;
  assign sel_783261 = array_index_782956 == array_index_773092 ? add_783260 : sel_783257;
  assign add_783264 = sel_783261 + 8'h01;
  assign sel_783265 = array_index_782956 == array_index_773098 ? add_783264 : sel_783261;
  assign add_783268 = sel_783265 + 8'h01;
  assign sel_783269 = array_index_782956 == array_index_773104 ? add_783268 : sel_783265;
  assign add_783272 = sel_783269 + 8'h01;
  assign sel_783273 = array_index_782956 == array_index_773110 ? add_783272 : sel_783269;
  assign add_783276 = sel_783273 + 8'h01;
  assign sel_783277 = array_index_782956 == array_index_773116 ? add_783276 : sel_783273;
  assign add_783280 = sel_783277 + 8'h01;
  assign sel_783281 = array_index_782956 == array_index_773122 ? add_783280 : sel_783277;
  assign add_783284 = sel_783281 + 8'h01;
  assign sel_783285 = array_index_782956 == array_index_773128 ? add_783284 : sel_783281;
  assign add_783288 = sel_783285 + 8'h01;
  assign sel_783289 = array_index_782956 == array_index_773134 ? add_783288 : sel_783285;
  assign add_783292 = sel_783289 + 8'h01;
  assign sel_783293 = array_index_782956 == array_index_773140 ? add_783292 : sel_783289;
  assign add_783296 = sel_783293 + 8'h01;
  assign sel_783297 = array_index_782956 == array_index_773146 ? add_783296 : sel_783293;
  assign add_783300 = sel_783297 + 8'h01;
  assign sel_783301 = array_index_782956 == array_index_773152 ? add_783300 : sel_783297;
  assign add_783304 = sel_783301 + 8'h01;
  assign sel_783305 = array_index_782956 == array_index_773158 ? add_783304 : sel_783301;
  assign add_783308 = sel_783305 + 8'h01;
  assign sel_783309 = array_index_782956 == array_index_773164 ? add_783308 : sel_783305;
  assign add_783312 = sel_783309 + 8'h01;
  assign sel_783313 = array_index_782956 == array_index_773170 ? add_783312 : sel_783309;
  assign add_783317 = sel_783313 + 8'h01;
  assign array_index_783318 = set1_unflattened[7'h1d];
  assign sel_783319 = array_index_782956 == array_index_773176 ? add_783317 : sel_783313;
  assign add_783322 = sel_783319 + 8'h01;
  assign sel_783323 = array_index_783318 == array_index_772632 ? add_783322 : sel_783319;
  assign add_783326 = sel_783323 + 8'h01;
  assign sel_783327 = array_index_783318 == array_index_772636 ? add_783326 : sel_783323;
  assign add_783330 = sel_783327 + 8'h01;
  assign sel_783331 = array_index_783318 == array_index_772644 ? add_783330 : sel_783327;
  assign add_783334 = sel_783331 + 8'h01;
  assign sel_783335 = array_index_783318 == array_index_772652 ? add_783334 : sel_783331;
  assign add_783338 = sel_783335 + 8'h01;
  assign sel_783339 = array_index_783318 == array_index_772660 ? add_783338 : sel_783335;
  assign add_783342 = sel_783339 + 8'h01;
  assign sel_783343 = array_index_783318 == array_index_772668 ? add_783342 : sel_783339;
  assign add_783346 = sel_783343 + 8'h01;
  assign sel_783347 = array_index_783318 == array_index_772676 ? add_783346 : sel_783343;
  assign add_783350 = sel_783347 + 8'h01;
  assign sel_783351 = array_index_783318 == array_index_772684 ? add_783350 : sel_783347;
  assign add_783354 = sel_783351 + 8'h01;
  assign sel_783355 = array_index_783318 == array_index_772690 ? add_783354 : sel_783351;
  assign add_783358 = sel_783355 + 8'h01;
  assign sel_783359 = array_index_783318 == array_index_772696 ? add_783358 : sel_783355;
  assign add_783362 = sel_783359 + 8'h01;
  assign sel_783363 = array_index_783318 == array_index_772702 ? add_783362 : sel_783359;
  assign add_783366 = sel_783363 + 8'h01;
  assign sel_783367 = array_index_783318 == array_index_772708 ? add_783366 : sel_783363;
  assign add_783370 = sel_783367 + 8'h01;
  assign sel_783371 = array_index_783318 == array_index_772714 ? add_783370 : sel_783367;
  assign add_783374 = sel_783371 + 8'h01;
  assign sel_783375 = array_index_783318 == array_index_772720 ? add_783374 : sel_783371;
  assign add_783378 = sel_783375 + 8'h01;
  assign sel_783379 = array_index_783318 == array_index_772726 ? add_783378 : sel_783375;
  assign add_783382 = sel_783379 + 8'h01;
  assign sel_783383 = array_index_783318 == array_index_772732 ? add_783382 : sel_783379;
  assign add_783386 = sel_783383 + 8'h01;
  assign sel_783387 = array_index_783318 == array_index_772738 ? add_783386 : sel_783383;
  assign add_783390 = sel_783387 + 8'h01;
  assign sel_783391 = array_index_783318 == array_index_772744 ? add_783390 : sel_783387;
  assign add_783394 = sel_783391 + 8'h01;
  assign sel_783395 = array_index_783318 == array_index_772750 ? add_783394 : sel_783391;
  assign add_783398 = sel_783395 + 8'h01;
  assign sel_783399 = array_index_783318 == array_index_772756 ? add_783398 : sel_783395;
  assign add_783402 = sel_783399 + 8'h01;
  assign sel_783403 = array_index_783318 == array_index_772762 ? add_783402 : sel_783399;
  assign add_783406 = sel_783403 + 8'h01;
  assign sel_783407 = array_index_783318 == array_index_772768 ? add_783406 : sel_783403;
  assign add_783410 = sel_783407 + 8'h01;
  assign sel_783411 = array_index_783318 == array_index_772774 ? add_783410 : sel_783407;
  assign add_783414 = sel_783411 + 8'h01;
  assign sel_783415 = array_index_783318 == array_index_772780 ? add_783414 : sel_783411;
  assign add_783418 = sel_783415 + 8'h01;
  assign sel_783419 = array_index_783318 == array_index_772786 ? add_783418 : sel_783415;
  assign add_783422 = sel_783419 + 8'h01;
  assign sel_783423 = array_index_783318 == array_index_772792 ? add_783422 : sel_783419;
  assign add_783426 = sel_783423 + 8'h01;
  assign sel_783427 = array_index_783318 == array_index_772798 ? add_783426 : sel_783423;
  assign add_783430 = sel_783427 + 8'h01;
  assign sel_783431 = array_index_783318 == array_index_772804 ? add_783430 : sel_783427;
  assign add_783434 = sel_783431 + 8'h01;
  assign sel_783435 = array_index_783318 == array_index_772810 ? add_783434 : sel_783431;
  assign add_783438 = sel_783435 + 8'h01;
  assign sel_783439 = array_index_783318 == array_index_772816 ? add_783438 : sel_783435;
  assign add_783442 = sel_783439 + 8'h01;
  assign sel_783443 = array_index_783318 == array_index_772822 ? add_783442 : sel_783439;
  assign add_783446 = sel_783443 + 8'h01;
  assign sel_783447 = array_index_783318 == array_index_772828 ? add_783446 : sel_783443;
  assign add_783450 = sel_783447 + 8'h01;
  assign sel_783451 = array_index_783318 == array_index_772834 ? add_783450 : sel_783447;
  assign add_783454 = sel_783451 + 8'h01;
  assign sel_783455 = array_index_783318 == array_index_772840 ? add_783454 : sel_783451;
  assign add_783458 = sel_783455 + 8'h01;
  assign sel_783459 = array_index_783318 == array_index_772846 ? add_783458 : sel_783455;
  assign add_783462 = sel_783459 + 8'h01;
  assign sel_783463 = array_index_783318 == array_index_772852 ? add_783462 : sel_783459;
  assign add_783466 = sel_783463 + 8'h01;
  assign sel_783467 = array_index_783318 == array_index_772858 ? add_783466 : sel_783463;
  assign add_783470 = sel_783467 + 8'h01;
  assign sel_783471 = array_index_783318 == array_index_772864 ? add_783470 : sel_783467;
  assign add_783474 = sel_783471 + 8'h01;
  assign sel_783475 = array_index_783318 == array_index_772870 ? add_783474 : sel_783471;
  assign add_783478 = sel_783475 + 8'h01;
  assign sel_783479 = array_index_783318 == array_index_772876 ? add_783478 : sel_783475;
  assign add_783482 = sel_783479 + 8'h01;
  assign sel_783483 = array_index_783318 == array_index_772882 ? add_783482 : sel_783479;
  assign add_783486 = sel_783483 + 8'h01;
  assign sel_783487 = array_index_783318 == array_index_772888 ? add_783486 : sel_783483;
  assign add_783490 = sel_783487 + 8'h01;
  assign sel_783491 = array_index_783318 == array_index_772894 ? add_783490 : sel_783487;
  assign add_783494 = sel_783491 + 8'h01;
  assign sel_783495 = array_index_783318 == array_index_772900 ? add_783494 : sel_783491;
  assign add_783498 = sel_783495 + 8'h01;
  assign sel_783499 = array_index_783318 == array_index_772906 ? add_783498 : sel_783495;
  assign add_783502 = sel_783499 + 8'h01;
  assign sel_783503 = array_index_783318 == array_index_772912 ? add_783502 : sel_783499;
  assign add_783506 = sel_783503 + 8'h01;
  assign sel_783507 = array_index_783318 == array_index_772918 ? add_783506 : sel_783503;
  assign add_783510 = sel_783507 + 8'h01;
  assign sel_783511 = array_index_783318 == array_index_772924 ? add_783510 : sel_783507;
  assign add_783514 = sel_783511 + 8'h01;
  assign sel_783515 = array_index_783318 == array_index_772930 ? add_783514 : sel_783511;
  assign add_783518 = sel_783515 + 8'h01;
  assign sel_783519 = array_index_783318 == array_index_772936 ? add_783518 : sel_783515;
  assign add_783522 = sel_783519 + 8'h01;
  assign sel_783523 = array_index_783318 == array_index_772942 ? add_783522 : sel_783519;
  assign add_783526 = sel_783523 + 8'h01;
  assign sel_783527 = array_index_783318 == array_index_772948 ? add_783526 : sel_783523;
  assign add_783530 = sel_783527 + 8'h01;
  assign sel_783531 = array_index_783318 == array_index_772954 ? add_783530 : sel_783527;
  assign add_783534 = sel_783531 + 8'h01;
  assign sel_783535 = array_index_783318 == array_index_772960 ? add_783534 : sel_783531;
  assign add_783538 = sel_783535 + 8'h01;
  assign sel_783539 = array_index_783318 == array_index_772966 ? add_783538 : sel_783535;
  assign add_783542 = sel_783539 + 8'h01;
  assign sel_783543 = array_index_783318 == array_index_772972 ? add_783542 : sel_783539;
  assign add_783546 = sel_783543 + 8'h01;
  assign sel_783547 = array_index_783318 == array_index_772978 ? add_783546 : sel_783543;
  assign add_783550 = sel_783547 + 8'h01;
  assign sel_783551 = array_index_783318 == array_index_772984 ? add_783550 : sel_783547;
  assign add_783554 = sel_783551 + 8'h01;
  assign sel_783555 = array_index_783318 == array_index_772990 ? add_783554 : sel_783551;
  assign add_783558 = sel_783555 + 8'h01;
  assign sel_783559 = array_index_783318 == array_index_772996 ? add_783558 : sel_783555;
  assign add_783562 = sel_783559 + 8'h01;
  assign sel_783563 = array_index_783318 == array_index_773002 ? add_783562 : sel_783559;
  assign add_783566 = sel_783563 + 8'h01;
  assign sel_783567 = array_index_783318 == array_index_773008 ? add_783566 : sel_783563;
  assign add_783570 = sel_783567 + 8'h01;
  assign sel_783571 = array_index_783318 == array_index_773014 ? add_783570 : sel_783567;
  assign add_783574 = sel_783571 + 8'h01;
  assign sel_783575 = array_index_783318 == array_index_773020 ? add_783574 : sel_783571;
  assign add_783578 = sel_783575 + 8'h01;
  assign sel_783579 = array_index_783318 == array_index_773026 ? add_783578 : sel_783575;
  assign add_783582 = sel_783579 + 8'h01;
  assign sel_783583 = array_index_783318 == array_index_773032 ? add_783582 : sel_783579;
  assign add_783586 = sel_783583 + 8'h01;
  assign sel_783587 = array_index_783318 == array_index_773038 ? add_783586 : sel_783583;
  assign add_783590 = sel_783587 + 8'h01;
  assign sel_783591 = array_index_783318 == array_index_773044 ? add_783590 : sel_783587;
  assign add_783594 = sel_783591 + 8'h01;
  assign sel_783595 = array_index_783318 == array_index_773050 ? add_783594 : sel_783591;
  assign add_783598 = sel_783595 + 8'h01;
  assign sel_783599 = array_index_783318 == array_index_773056 ? add_783598 : sel_783595;
  assign add_783602 = sel_783599 + 8'h01;
  assign sel_783603 = array_index_783318 == array_index_773062 ? add_783602 : sel_783599;
  assign add_783606 = sel_783603 + 8'h01;
  assign sel_783607 = array_index_783318 == array_index_773068 ? add_783606 : sel_783603;
  assign add_783610 = sel_783607 + 8'h01;
  assign sel_783611 = array_index_783318 == array_index_773074 ? add_783610 : sel_783607;
  assign add_783614 = sel_783611 + 8'h01;
  assign sel_783615 = array_index_783318 == array_index_773080 ? add_783614 : sel_783611;
  assign add_783618 = sel_783615 + 8'h01;
  assign sel_783619 = array_index_783318 == array_index_773086 ? add_783618 : sel_783615;
  assign add_783622 = sel_783619 + 8'h01;
  assign sel_783623 = array_index_783318 == array_index_773092 ? add_783622 : sel_783619;
  assign add_783626 = sel_783623 + 8'h01;
  assign sel_783627 = array_index_783318 == array_index_773098 ? add_783626 : sel_783623;
  assign add_783630 = sel_783627 + 8'h01;
  assign sel_783631 = array_index_783318 == array_index_773104 ? add_783630 : sel_783627;
  assign add_783634 = sel_783631 + 8'h01;
  assign sel_783635 = array_index_783318 == array_index_773110 ? add_783634 : sel_783631;
  assign add_783638 = sel_783635 + 8'h01;
  assign sel_783639 = array_index_783318 == array_index_773116 ? add_783638 : sel_783635;
  assign add_783642 = sel_783639 + 8'h01;
  assign sel_783643 = array_index_783318 == array_index_773122 ? add_783642 : sel_783639;
  assign add_783646 = sel_783643 + 8'h01;
  assign sel_783647 = array_index_783318 == array_index_773128 ? add_783646 : sel_783643;
  assign add_783650 = sel_783647 + 8'h01;
  assign sel_783651 = array_index_783318 == array_index_773134 ? add_783650 : sel_783647;
  assign add_783654 = sel_783651 + 8'h01;
  assign sel_783655 = array_index_783318 == array_index_773140 ? add_783654 : sel_783651;
  assign add_783658 = sel_783655 + 8'h01;
  assign sel_783659 = array_index_783318 == array_index_773146 ? add_783658 : sel_783655;
  assign add_783662 = sel_783659 + 8'h01;
  assign sel_783663 = array_index_783318 == array_index_773152 ? add_783662 : sel_783659;
  assign add_783666 = sel_783663 + 8'h01;
  assign sel_783667 = array_index_783318 == array_index_773158 ? add_783666 : sel_783663;
  assign add_783670 = sel_783667 + 8'h01;
  assign sel_783671 = array_index_783318 == array_index_773164 ? add_783670 : sel_783667;
  assign add_783674 = sel_783671 + 8'h01;
  assign sel_783675 = array_index_783318 == array_index_773170 ? add_783674 : sel_783671;
  assign add_783679 = sel_783675 + 8'h01;
  assign array_index_783680 = set1_unflattened[7'h1e];
  assign sel_783681 = array_index_783318 == array_index_773176 ? add_783679 : sel_783675;
  assign add_783684 = sel_783681 + 8'h01;
  assign sel_783685 = array_index_783680 == array_index_772632 ? add_783684 : sel_783681;
  assign add_783688 = sel_783685 + 8'h01;
  assign sel_783689 = array_index_783680 == array_index_772636 ? add_783688 : sel_783685;
  assign add_783692 = sel_783689 + 8'h01;
  assign sel_783693 = array_index_783680 == array_index_772644 ? add_783692 : sel_783689;
  assign add_783696 = sel_783693 + 8'h01;
  assign sel_783697 = array_index_783680 == array_index_772652 ? add_783696 : sel_783693;
  assign add_783700 = sel_783697 + 8'h01;
  assign sel_783701 = array_index_783680 == array_index_772660 ? add_783700 : sel_783697;
  assign add_783704 = sel_783701 + 8'h01;
  assign sel_783705 = array_index_783680 == array_index_772668 ? add_783704 : sel_783701;
  assign add_783708 = sel_783705 + 8'h01;
  assign sel_783709 = array_index_783680 == array_index_772676 ? add_783708 : sel_783705;
  assign add_783712 = sel_783709 + 8'h01;
  assign sel_783713 = array_index_783680 == array_index_772684 ? add_783712 : sel_783709;
  assign add_783716 = sel_783713 + 8'h01;
  assign sel_783717 = array_index_783680 == array_index_772690 ? add_783716 : sel_783713;
  assign add_783720 = sel_783717 + 8'h01;
  assign sel_783721 = array_index_783680 == array_index_772696 ? add_783720 : sel_783717;
  assign add_783724 = sel_783721 + 8'h01;
  assign sel_783725 = array_index_783680 == array_index_772702 ? add_783724 : sel_783721;
  assign add_783728 = sel_783725 + 8'h01;
  assign sel_783729 = array_index_783680 == array_index_772708 ? add_783728 : sel_783725;
  assign add_783732 = sel_783729 + 8'h01;
  assign sel_783733 = array_index_783680 == array_index_772714 ? add_783732 : sel_783729;
  assign add_783736 = sel_783733 + 8'h01;
  assign sel_783737 = array_index_783680 == array_index_772720 ? add_783736 : sel_783733;
  assign add_783740 = sel_783737 + 8'h01;
  assign sel_783741 = array_index_783680 == array_index_772726 ? add_783740 : sel_783737;
  assign add_783744 = sel_783741 + 8'h01;
  assign sel_783745 = array_index_783680 == array_index_772732 ? add_783744 : sel_783741;
  assign add_783748 = sel_783745 + 8'h01;
  assign sel_783749 = array_index_783680 == array_index_772738 ? add_783748 : sel_783745;
  assign add_783752 = sel_783749 + 8'h01;
  assign sel_783753 = array_index_783680 == array_index_772744 ? add_783752 : sel_783749;
  assign add_783756 = sel_783753 + 8'h01;
  assign sel_783757 = array_index_783680 == array_index_772750 ? add_783756 : sel_783753;
  assign add_783760 = sel_783757 + 8'h01;
  assign sel_783761 = array_index_783680 == array_index_772756 ? add_783760 : sel_783757;
  assign add_783764 = sel_783761 + 8'h01;
  assign sel_783765 = array_index_783680 == array_index_772762 ? add_783764 : sel_783761;
  assign add_783768 = sel_783765 + 8'h01;
  assign sel_783769 = array_index_783680 == array_index_772768 ? add_783768 : sel_783765;
  assign add_783772 = sel_783769 + 8'h01;
  assign sel_783773 = array_index_783680 == array_index_772774 ? add_783772 : sel_783769;
  assign add_783776 = sel_783773 + 8'h01;
  assign sel_783777 = array_index_783680 == array_index_772780 ? add_783776 : sel_783773;
  assign add_783780 = sel_783777 + 8'h01;
  assign sel_783781 = array_index_783680 == array_index_772786 ? add_783780 : sel_783777;
  assign add_783784 = sel_783781 + 8'h01;
  assign sel_783785 = array_index_783680 == array_index_772792 ? add_783784 : sel_783781;
  assign add_783788 = sel_783785 + 8'h01;
  assign sel_783789 = array_index_783680 == array_index_772798 ? add_783788 : sel_783785;
  assign add_783792 = sel_783789 + 8'h01;
  assign sel_783793 = array_index_783680 == array_index_772804 ? add_783792 : sel_783789;
  assign add_783796 = sel_783793 + 8'h01;
  assign sel_783797 = array_index_783680 == array_index_772810 ? add_783796 : sel_783793;
  assign add_783800 = sel_783797 + 8'h01;
  assign sel_783801 = array_index_783680 == array_index_772816 ? add_783800 : sel_783797;
  assign add_783804 = sel_783801 + 8'h01;
  assign sel_783805 = array_index_783680 == array_index_772822 ? add_783804 : sel_783801;
  assign add_783808 = sel_783805 + 8'h01;
  assign sel_783809 = array_index_783680 == array_index_772828 ? add_783808 : sel_783805;
  assign add_783812 = sel_783809 + 8'h01;
  assign sel_783813 = array_index_783680 == array_index_772834 ? add_783812 : sel_783809;
  assign add_783816 = sel_783813 + 8'h01;
  assign sel_783817 = array_index_783680 == array_index_772840 ? add_783816 : sel_783813;
  assign add_783820 = sel_783817 + 8'h01;
  assign sel_783821 = array_index_783680 == array_index_772846 ? add_783820 : sel_783817;
  assign add_783824 = sel_783821 + 8'h01;
  assign sel_783825 = array_index_783680 == array_index_772852 ? add_783824 : sel_783821;
  assign add_783828 = sel_783825 + 8'h01;
  assign sel_783829 = array_index_783680 == array_index_772858 ? add_783828 : sel_783825;
  assign add_783832 = sel_783829 + 8'h01;
  assign sel_783833 = array_index_783680 == array_index_772864 ? add_783832 : sel_783829;
  assign add_783836 = sel_783833 + 8'h01;
  assign sel_783837 = array_index_783680 == array_index_772870 ? add_783836 : sel_783833;
  assign add_783840 = sel_783837 + 8'h01;
  assign sel_783841 = array_index_783680 == array_index_772876 ? add_783840 : sel_783837;
  assign add_783844 = sel_783841 + 8'h01;
  assign sel_783845 = array_index_783680 == array_index_772882 ? add_783844 : sel_783841;
  assign add_783848 = sel_783845 + 8'h01;
  assign sel_783849 = array_index_783680 == array_index_772888 ? add_783848 : sel_783845;
  assign add_783852 = sel_783849 + 8'h01;
  assign sel_783853 = array_index_783680 == array_index_772894 ? add_783852 : sel_783849;
  assign add_783856 = sel_783853 + 8'h01;
  assign sel_783857 = array_index_783680 == array_index_772900 ? add_783856 : sel_783853;
  assign add_783860 = sel_783857 + 8'h01;
  assign sel_783861 = array_index_783680 == array_index_772906 ? add_783860 : sel_783857;
  assign add_783864 = sel_783861 + 8'h01;
  assign sel_783865 = array_index_783680 == array_index_772912 ? add_783864 : sel_783861;
  assign add_783868 = sel_783865 + 8'h01;
  assign sel_783869 = array_index_783680 == array_index_772918 ? add_783868 : sel_783865;
  assign add_783872 = sel_783869 + 8'h01;
  assign sel_783873 = array_index_783680 == array_index_772924 ? add_783872 : sel_783869;
  assign add_783876 = sel_783873 + 8'h01;
  assign sel_783877 = array_index_783680 == array_index_772930 ? add_783876 : sel_783873;
  assign add_783880 = sel_783877 + 8'h01;
  assign sel_783881 = array_index_783680 == array_index_772936 ? add_783880 : sel_783877;
  assign add_783884 = sel_783881 + 8'h01;
  assign sel_783885 = array_index_783680 == array_index_772942 ? add_783884 : sel_783881;
  assign add_783888 = sel_783885 + 8'h01;
  assign sel_783889 = array_index_783680 == array_index_772948 ? add_783888 : sel_783885;
  assign add_783892 = sel_783889 + 8'h01;
  assign sel_783893 = array_index_783680 == array_index_772954 ? add_783892 : sel_783889;
  assign add_783896 = sel_783893 + 8'h01;
  assign sel_783897 = array_index_783680 == array_index_772960 ? add_783896 : sel_783893;
  assign add_783900 = sel_783897 + 8'h01;
  assign sel_783901 = array_index_783680 == array_index_772966 ? add_783900 : sel_783897;
  assign add_783904 = sel_783901 + 8'h01;
  assign sel_783905 = array_index_783680 == array_index_772972 ? add_783904 : sel_783901;
  assign add_783908 = sel_783905 + 8'h01;
  assign sel_783909 = array_index_783680 == array_index_772978 ? add_783908 : sel_783905;
  assign add_783912 = sel_783909 + 8'h01;
  assign sel_783913 = array_index_783680 == array_index_772984 ? add_783912 : sel_783909;
  assign add_783916 = sel_783913 + 8'h01;
  assign sel_783917 = array_index_783680 == array_index_772990 ? add_783916 : sel_783913;
  assign add_783920 = sel_783917 + 8'h01;
  assign sel_783921 = array_index_783680 == array_index_772996 ? add_783920 : sel_783917;
  assign add_783924 = sel_783921 + 8'h01;
  assign sel_783925 = array_index_783680 == array_index_773002 ? add_783924 : sel_783921;
  assign add_783928 = sel_783925 + 8'h01;
  assign sel_783929 = array_index_783680 == array_index_773008 ? add_783928 : sel_783925;
  assign add_783932 = sel_783929 + 8'h01;
  assign sel_783933 = array_index_783680 == array_index_773014 ? add_783932 : sel_783929;
  assign add_783936 = sel_783933 + 8'h01;
  assign sel_783937 = array_index_783680 == array_index_773020 ? add_783936 : sel_783933;
  assign add_783940 = sel_783937 + 8'h01;
  assign sel_783941 = array_index_783680 == array_index_773026 ? add_783940 : sel_783937;
  assign add_783944 = sel_783941 + 8'h01;
  assign sel_783945 = array_index_783680 == array_index_773032 ? add_783944 : sel_783941;
  assign add_783948 = sel_783945 + 8'h01;
  assign sel_783949 = array_index_783680 == array_index_773038 ? add_783948 : sel_783945;
  assign add_783952 = sel_783949 + 8'h01;
  assign sel_783953 = array_index_783680 == array_index_773044 ? add_783952 : sel_783949;
  assign add_783956 = sel_783953 + 8'h01;
  assign sel_783957 = array_index_783680 == array_index_773050 ? add_783956 : sel_783953;
  assign add_783960 = sel_783957 + 8'h01;
  assign sel_783961 = array_index_783680 == array_index_773056 ? add_783960 : sel_783957;
  assign add_783964 = sel_783961 + 8'h01;
  assign sel_783965 = array_index_783680 == array_index_773062 ? add_783964 : sel_783961;
  assign add_783968 = sel_783965 + 8'h01;
  assign sel_783969 = array_index_783680 == array_index_773068 ? add_783968 : sel_783965;
  assign add_783972 = sel_783969 + 8'h01;
  assign sel_783973 = array_index_783680 == array_index_773074 ? add_783972 : sel_783969;
  assign add_783976 = sel_783973 + 8'h01;
  assign sel_783977 = array_index_783680 == array_index_773080 ? add_783976 : sel_783973;
  assign add_783980 = sel_783977 + 8'h01;
  assign sel_783981 = array_index_783680 == array_index_773086 ? add_783980 : sel_783977;
  assign add_783984 = sel_783981 + 8'h01;
  assign sel_783985 = array_index_783680 == array_index_773092 ? add_783984 : sel_783981;
  assign add_783988 = sel_783985 + 8'h01;
  assign sel_783989 = array_index_783680 == array_index_773098 ? add_783988 : sel_783985;
  assign add_783992 = sel_783989 + 8'h01;
  assign sel_783993 = array_index_783680 == array_index_773104 ? add_783992 : sel_783989;
  assign add_783996 = sel_783993 + 8'h01;
  assign sel_783997 = array_index_783680 == array_index_773110 ? add_783996 : sel_783993;
  assign add_784000 = sel_783997 + 8'h01;
  assign sel_784001 = array_index_783680 == array_index_773116 ? add_784000 : sel_783997;
  assign add_784004 = sel_784001 + 8'h01;
  assign sel_784005 = array_index_783680 == array_index_773122 ? add_784004 : sel_784001;
  assign add_784008 = sel_784005 + 8'h01;
  assign sel_784009 = array_index_783680 == array_index_773128 ? add_784008 : sel_784005;
  assign add_784012 = sel_784009 + 8'h01;
  assign sel_784013 = array_index_783680 == array_index_773134 ? add_784012 : sel_784009;
  assign add_784016 = sel_784013 + 8'h01;
  assign sel_784017 = array_index_783680 == array_index_773140 ? add_784016 : sel_784013;
  assign add_784020 = sel_784017 + 8'h01;
  assign sel_784021 = array_index_783680 == array_index_773146 ? add_784020 : sel_784017;
  assign add_784024 = sel_784021 + 8'h01;
  assign sel_784025 = array_index_783680 == array_index_773152 ? add_784024 : sel_784021;
  assign add_784028 = sel_784025 + 8'h01;
  assign sel_784029 = array_index_783680 == array_index_773158 ? add_784028 : sel_784025;
  assign add_784032 = sel_784029 + 8'h01;
  assign sel_784033 = array_index_783680 == array_index_773164 ? add_784032 : sel_784029;
  assign add_784036 = sel_784033 + 8'h01;
  assign sel_784037 = array_index_783680 == array_index_773170 ? add_784036 : sel_784033;
  assign add_784041 = sel_784037 + 8'h01;
  assign array_index_784042 = set1_unflattened[7'h1f];
  assign sel_784043 = array_index_783680 == array_index_773176 ? add_784041 : sel_784037;
  assign add_784046 = sel_784043 + 8'h01;
  assign sel_784047 = array_index_784042 == array_index_772632 ? add_784046 : sel_784043;
  assign add_784050 = sel_784047 + 8'h01;
  assign sel_784051 = array_index_784042 == array_index_772636 ? add_784050 : sel_784047;
  assign add_784054 = sel_784051 + 8'h01;
  assign sel_784055 = array_index_784042 == array_index_772644 ? add_784054 : sel_784051;
  assign add_784058 = sel_784055 + 8'h01;
  assign sel_784059 = array_index_784042 == array_index_772652 ? add_784058 : sel_784055;
  assign add_784062 = sel_784059 + 8'h01;
  assign sel_784063 = array_index_784042 == array_index_772660 ? add_784062 : sel_784059;
  assign add_784066 = sel_784063 + 8'h01;
  assign sel_784067 = array_index_784042 == array_index_772668 ? add_784066 : sel_784063;
  assign add_784070 = sel_784067 + 8'h01;
  assign sel_784071 = array_index_784042 == array_index_772676 ? add_784070 : sel_784067;
  assign add_784074 = sel_784071 + 8'h01;
  assign sel_784075 = array_index_784042 == array_index_772684 ? add_784074 : sel_784071;
  assign add_784078 = sel_784075 + 8'h01;
  assign sel_784079 = array_index_784042 == array_index_772690 ? add_784078 : sel_784075;
  assign add_784082 = sel_784079 + 8'h01;
  assign sel_784083 = array_index_784042 == array_index_772696 ? add_784082 : sel_784079;
  assign add_784086 = sel_784083 + 8'h01;
  assign sel_784087 = array_index_784042 == array_index_772702 ? add_784086 : sel_784083;
  assign add_784090 = sel_784087 + 8'h01;
  assign sel_784091 = array_index_784042 == array_index_772708 ? add_784090 : sel_784087;
  assign add_784094 = sel_784091 + 8'h01;
  assign sel_784095 = array_index_784042 == array_index_772714 ? add_784094 : sel_784091;
  assign add_784098 = sel_784095 + 8'h01;
  assign sel_784099 = array_index_784042 == array_index_772720 ? add_784098 : sel_784095;
  assign add_784102 = sel_784099 + 8'h01;
  assign sel_784103 = array_index_784042 == array_index_772726 ? add_784102 : sel_784099;
  assign add_784106 = sel_784103 + 8'h01;
  assign sel_784107 = array_index_784042 == array_index_772732 ? add_784106 : sel_784103;
  assign add_784110 = sel_784107 + 8'h01;
  assign sel_784111 = array_index_784042 == array_index_772738 ? add_784110 : sel_784107;
  assign add_784114 = sel_784111 + 8'h01;
  assign sel_784115 = array_index_784042 == array_index_772744 ? add_784114 : sel_784111;
  assign add_784118 = sel_784115 + 8'h01;
  assign sel_784119 = array_index_784042 == array_index_772750 ? add_784118 : sel_784115;
  assign add_784122 = sel_784119 + 8'h01;
  assign sel_784123 = array_index_784042 == array_index_772756 ? add_784122 : sel_784119;
  assign add_784126 = sel_784123 + 8'h01;
  assign sel_784127 = array_index_784042 == array_index_772762 ? add_784126 : sel_784123;
  assign add_784130 = sel_784127 + 8'h01;
  assign sel_784131 = array_index_784042 == array_index_772768 ? add_784130 : sel_784127;
  assign add_784134 = sel_784131 + 8'h01;
  assign sel_784135 = array_index_784042 == array_index_772774 ? add_784134 : sel_784131;
  assign add_784138 = sel_784135 + 8'h01;
  assign sel_784139 = array_index_784042 == array_index_772780 ? add_784138 : sel_784135;
  assign add_784142 = sel_784139 + 8'h01;
  assign sel_784143 = array_index_784042 == array_index_772786 ? add_784142 : sel_784139;
  assign add_784146 = sel_784143 + 8'h01;
  assign sel_784147 = array_index_784042 == array_index_772792 ? add_784146 : sel_784143;
  assign add_784150 = sel_784147 + 8'h01;
  assign sel_784151 = array_index_784042 == array_index_772798 ? add_784150 : sel_784147;
  assign add_784154 = sel_784151 + 8'h01;
  assign sel_784155 = array_index_784042 == array_index_772804 ? add_784154 : sel_784151;
  assign add_784158 = sel_784155 + 8'h01;
  assign sel_784159 = array_index_784042 == array_index_772810 ? add_784158 : sel_784155;
  assign add_784162 = sel_784159 + 8'h01;
  assign sel_784163 = array_index_784042 == array_index_772816 ? add_784162 : sel_784159;
  assign add_784166 = sel_784163 + 8'h01;
  assign sel_784167 = array_index_784042 == array_index_772822 ? add_784166 : sel_784163;
  assign add_784170 = sel_784167 + 8'h01;
  assign sel_784171 = array_index_784042 == array_index_772828 ? add_784170 : sel_784167;
  assign add_784174 = sel_784171 + 8'h01;
  assign sel_784175 = array_index_784042 == array_index_772834 ? add_784174 : sel_784171;
  assign add_784178 = sel_784175 + 8'h01;
  assign sel_784179 = array_index_784042 == array_index_772840 ? add_784178 : sel_784175;
  assign add_784182 = sel_784179 + 8'h01;
  assign sel_784183 = array_index_784042 == array_index_772846 ? add_784182 : sel_784179;
  assign add_784186 = sel_784183 + 8'h01;
  assign sel_784187 = array_index_784042 == array_index_772852 ? add_784186 : sel_784183;
  assign add_784190 = sel_784187 + 8'h01;
  assign sel_784191 = array_index_784042 == array_index_772858 ? add_784190 : sel_784187;
  assign add_784194 = sel_784191 + 8'h01;
  assign sel_784195 = array_index_784042 == array_index_772864 ? add_784194 : sel_784191;
  assign add_784198 = sel_784195 + 8'h01;
  assign sel_784199 = array_index_784042 == array_index_772870 ? add_784198 : sel_784195;
  assign add_784202 = sel_784199 + 8'h01;
  assign sel_784203 = array_index_784042 == array_index_772876 ? add_784202 : sel_784199;
  assign add_784206 = sel_784203 + 8'h01;
  assign sel_784207 = array_index_784042 == array_index_772882 ? add_784206 : sel_784203;
  assign add_784210 = sel_784207 + 8'h01;
  assign sel_784211 = array_index_784042 == array_index_772888 ? add_784210 : sel_784207;
  assign add_784214 = sel_784211 + 8'h01;
  assign sel_784215 = array_index_784042 == array_index_772894 ? add_784214 : sel_784211;
  assign add_784218 = sel_784215 + 8'h01;
  assign sel_784219 = array_index_784042 == array_index_772900 ? add_784218 : sel_784215;
  assign add_784222 = sel_784219 + 8'h01;
  assign sel_784223 = array_index_784042 == array_index_772906 ? add_784222 : sel_784219;
  assign add_784226 = sel_784223 + 8'h01;
  assign sel_784227 = array_index_784042 == array_index_772912 ? add_784226 : sel_784223;
  assign add_784230 = sel_784227 + 8'h01;
  assign sel_784231 = array_index_784042 == array_index_772918 ? add_784230 : sel_784227;
  assign add_784234 = sel_784231 + 8'h01;
  assign sel_784235 = array_index_784042 == array_index_772924 ? add_784234 : sel_784231;
  assign add_784238 = sel_784235 + 8'h01;
  assign sel_784239 = array_index_784042 == array_index_772930 ? add_784238 : sel_784235;
  assign add_784242 = sel_784239 + 8'h01;
  assign sel_784243 = array_index_784042 == array_index_772936 ? add_784242 : sel_784239;
  assign add_784246 = sel_784243 + 8'h01;
  assign sel_784247 = array_index_784042 == array_index_772942 ? add_784246 : sel_784243;
  assign add_784250 = sel_784247 + 8'h01;
  assign sel_784251 = array_index_784042 == array_index_772948 ? add_784250 : sel_784247;
  assign add_784254 = sel_784251 + 8'h01;
  assign sel_784255 = array_index_784042 == array_index_772954 ? add_784254 : sel_784251;
  assign add_784258 = sel_784255 + 8'h01;
  assign sel_784259 = array_index_784042 == array_index_772960 ? add_784258 : sel_784255;
  assign add_784262 = sel_784259 + 8'h01;
  assign sel_784263 = array_index_784042 == array_index_772966 ? add_784262 : sel_784259;
  assign add_784266 = sel_784263 + 8'h01;
  assign sel_784267 = array_index_784042 == array_index_772972 ? add_784266 : sel_784263;
  assign add_784270 = sel_784267 + 8'h01;
  assign sel_784271 = array_index_784042 == array_index_772978 ? add_784270 : sel_784267;
  assign add_784274 = sel_784271 + 8'h01;
  assign sel_784275 = array_index_784042 == array_index_772984 ? add_784274 : sel_784271;
  assign add_784278 = sel_784275 + 8'h01;
  assign sel_784279 = array_index_784042 == array_index_772990 ? add_784278 : sel_784275;
  assign add_784282 = sel_784279 + 8'h01;
  assign sel_784283 = array_index_784042 == array_index_772996 ? add_784282 : sel_784279;
  assign add_784286 = sel_784283 + 8'h01;
  assign sel_784287 = array_index_784042 == array_index_773002 ? add_784286 : sel_784283;
  assign add_784290 = sel_784287 + 8'h01;
  assign sel_784291 = array_index_784042 == array_index_773008 ? add_784290 : sel_784287;
  assign add_784294 = sel_784291 + 8'h01;
  assign sel_784295 = array_index_784042 == array_index_773014 ? add_784294 : sel_784291;
  assign add_784298 = sel_784295 + 8'h01;
  assign sel_784299 = array_index_784042 == array_index_773020 ? add_784298 : sel_784295;
  assign add_784302 = sel_784299 + 8'h01;
  assign sel_784303 = array_index_784042 == array_index_773026 ? add_784302 : sel_784299;
  assign add_784306 = sel_784303 + 8'h01;
  assign sel_784307 = array_index_784042 == array_index_773032 ? add_784306 : sel_784303;
  assign add_784310 = sel_784307 + 8'h01;
  assign sel_784311 = array_index_784042 == array_index_773038 ? add_784310 : sel_784307;
  assign add_784314 = sel_784311 + 8'h01;
  assign sel_784315 = array_index_784042 == array_index_773044 ? add_784314 : sel_784311;
  assign add_784318 = sel_784315 + 8'h01;
  assign sel_784319 = array_index_784042 == array_index_773050 ? add_784318 : sel_784315;
  assign add_784322 = sel_784319 + 8'h01;
  assign sel_784323 = array_index_784042 == array_index_773056 ? add_784322 : sel_784319;
  assign add_784326 = sel_784323 + 8'h01;
  assign sel_784327 = array_index_784042 == array_index_773062 ? add_784326 : sel_784323;
  assign add_784330 = sel_784327 + 8'h01;
  assign sel_784331 = array_index_784042 == array_index_773068 ? add_784330 : sel_784327;
  assign add_784334 = sel_784331 + 8'h01;
  assign sel_784335 = array_index_784042 == array_index_773074 ? add_784334 : sel_784331;
  assign add_784338 = sel_784335 + 8'h01;
  assign sel_784339 = array_index_784042 == array_index_773080 ? add_784338 : sel_784335;
  assign add_784342 = sel_784339 + 8'h01;
  assign sel_784343 = array_index_784042 == array_index_773086 ? add_784342 : sel_784339;
  assign add_784346 = sel_784343 + 8'h01;
  assign sel_784347 = array_index_784042 == array_index_773092 ? add_784346 : sel_784343;
  assign add_784350 = sel_784347 + 8'h01;
  assign sel_784351 = array_index_784042 == array_index_773098 ? add_784350 : sel_784347;
  assign add_784354 = sel_784351 + 8'h01;
  assign sel_784355 = array_index_784042 == array_index_773104 ? add_784354 : sel_784351;
  assign add_784358 = sel_784355 + 8'h01;
  assign sel_784359 = array_index_784042 == array_index_773110 ? add_784358 : sel_784355;
  assign add_784362 = sel_784359 + 8'h01;
  assign sel_784363 = array_index_784042 == array_index_773116 ? add_784362 : sel_784359;
  assign add_784366 = sel_784363 + 8'h01;
  assign sel_784367 = array_index_784042 == array_index_773122 ? add_784366 : sel_784363;
  assign add_784370 = sel_784367 + 8'h01;
  assign sel_784371 = array_index_784042 == array_index_773128 ? add_784370 : sel_784367;
  assign add_784374 = sel_784371 + 8'h01;
  assign sel_784375 = array_index_784042 == array_index_773134 ? add_784374 : sel_784371;
  assign add_784378 = sel_784375 + 8'h01;
  assign sel_784379 = array_index_784042 == array_index_773140 ? add_784378 : sel_784375;
  assign add_784382 = sel_784379 + 8'h01;
  assign sel_784383 = array_index_784042 == array_index_773146 ? add_784382 : sel_784379;
  assign add_784386 = sel_784383 + 8'h01;
  assign sel_784387 = array_index_784042 == array_index_773152 ? add_784386 : sel_784383;
  assign add_784390 = sel_784387 + 8'h01;
  assign sel_784391 = array_index_784042 == array_index_773158 ? add_784390 : sel_784387;
  assign add_784394 = sel_784391 + 8'h01;
  assign sel_784395 = array_index_784042 == array_index_773164 ? add_784394 : sel_784391;
  assign add_784398 = sel_784395 + 8'h01;
  assign sel_784399 = array_index_784042 == array_index_773170 ? add_784398 : sel_784395;
  assign add_784403 = sel_784399 + 8'h01;
  assign array_index_784404 = set1_unflattened[7'h20];
  assign sel_784405 = array_index_784042 == array_index_773176 ? add_784403 : sel_784399;
  assign add_784408 = sel_784405 + 8'h01;
  assign sel_784409 = array_index_784404 == array_index_772632 ? add_784408 : sel_784405;
  assign add_784412 = sel_784409 + 8'h01;
  assign sel_784413 = array_index_784404 == array_index_772636 ? add_784412 : sel_784409;
  assign add_784416 = sel_784413 + 8'h01;
  assign sel_784417 = array_index_784404 == array_index_772644 ? add_784416 : sel_784413;
  assign add_784420 = sel_784417 + 8'h01;
  assign sel_784421 = array_index_784404 == array_index_772652 ? add_784420 : sel_784417;
  assign add_784424 = sel_784421 + 8'h01;
  assign sel_784425 = array_index_784404 == array_index_772660 ? add_784424 : sel_784421;
  assign add_784428 = sel_784425 + 8'h01;
  assign sel_784429 = array_index_784404 == array_index_772668 ? add_784428 : sel_784425;
  assign add_784432 = sel_784429 + 8'h01;
  assign sel_784433 = array_index_784404 == array_index_772676 ? add_784432 : sel_784429;
  assign add_784436 = sel_784433 + 8'h01;
  assign sel_784437 = array_index_784404 == array_index_772684 ? add_784436 : sel_784433;
  assign add_784440 = sel_784437 + 8'h01;
  assign sel_784441 = array_index_784404 == array_index_772690 ? add_784440 : sel_784437;
  assign add_784444 = sel_784441 + 8'h01;
  assign sel_784445 = array_index_784404 == array_index_772696 ? add_784444 : sel_784441;
  assign add_784448 = sel_784445 + 8'h01;
  assign sel_784449 = array_index_784404 == array_index_772702 ? add_784448 : sel_784445;
  assign add_784452 = sel_784449 + 8'h01;
  assign sel_784453 = array_index_784404 == array_index_772708 ? add_784452 : sel_784449;
  assign add_784456 = sel_784453 + 8'h01;
  assign sel_784457 = array_index_784404 == array_index_772714 ? add_784456 : sel_784453;
  assign add_784460 = sel_784457 + 8'h01;
  assign sel_784461 = array_index_784404 == array_index_772720 ? add_784460 : sel_784457;
  assign add_784464 = sel_784461 + 8'h01;
  assign sel_784465 = array_index_784404 == array_index_772726 ? add_784464 : sel_784461;
  assign add_784468 = sel_784465 + 8'h01;
  assign sel_784469 = array_index_784404 == array_index_772732 ? add_784468 : sel_784465;
  assign add_784472 = sel_784469 + 8'h01;
  assign sel_784473 = array_index_784404 == array_index_772738 ? add_784472 : sel_784469;
  assign add_784476 = sel_784473 + 8'h01;
  assign sel_784477 = array_index_784404 == array_index_772744 ? add_784476 : sel_784473;
  assign add_784480 = sel_784477 + 8'h01;
  assign sel_784481 = array_index_784404 == array_index_772750 ? add_784480 : sel_784477;
  assign add_784484 = sel_784481 + 8'h01;
  assign sel_784485 = array_index_784404 == array_index_772756 ? add_784484 : sel_784481;
  assign add_784488 = sel_784485 + 8'h01;
  assign sel_784489 = array_index_784404 == array_index_772762 ? add_784488 : sel_784485;
  assign add_784492 = sel_784489 + 8'h01;
  assign sel_784493 = array_index_784404 == array_index_772768 ? add_784492 : sel_784489;
  assign add_784496 = sel_784493 + 8'h01;
  assign sel_784497 = array_index_784404 == array_index_772774 ? add_784496 : sel_784493;
  assign add_784500 = sel_784497 + 8'h01;
  assign sel_784501 = array_index_784404 == array_index_772780 ? add_784500 : sel_784497;
  assign add_784504 = sel_784501 + 8'h01;
  assign sel_784505 = array_index_784404 == array_index_772786 ? add_784504 : sel_784501;
  assign add_784508 = sel_784505 + 8'h01;
  assign sel_784509 = array_index_784404 == array_index_772792 ? add_784508 : sel_784505;
  assign add_784512 = sel_784509 + 8'h01;
  assign sel_784513 = array_index_784404 == array_index_772798 ? add_784512 : sel_784509;
  assign add_784516 = sel_784513 + 8'h01;
  assign sel_784517 = array_index_784404 == array_index_772804 ? add_784516 : sel_784513;
  assign add_784520 = sel_784517 + 8'h01;
  assign sel_784521 = array_index_784404 == array_index_772810 ? add_784520 : sel_784517;
  assign add_784524 = sel_784521 + 8'h01;
  assign sel_784525 = array_index_784404 == array_index_772816 ? add_784524 : sel_784521;
  assign add_784528 = sel_784525 + 8'h01;
  assign sel_784529 = array_index_784404 == array_index_772822 ? add_784528 : sel_784525;
  assign add_784532 = sel_784529 + 8'h01;
  assign sel_784533 = array_index_784404 == array_index_772828 ? add_784532 : sel_784529;
  assign add_784536 = sel_784533 + 8'h01;
  assign sel_784537 = array_index_784404 == array_index_772834 ? add_784536 : sel_784533;
  assign add_784540 = sel_784537 + 8'h01;
  assign sel_784541 = array_index_784404 == array_index_772840 ? add_784540 : sel_784537;
  assign add_784544 = sel_784541 + 8'h01;
  assign sel_784545 = array_index_784404 == array_index_772846 ? add_784544 : sel_784541;
  assign add_784548 = sel_784545 + 8'h01;
  assign sel_784549 = array_index_784404 == array_index_772852 ? add_784548 : sel_784545;
  assign add_784552 = sel_784549 + 8'h01;
  assign sel_784553 = array_index_784404 == array_index_772858 ? add_784552 : sel_784549;
  assign add_784556 = sel_784553 + 8'h01;
  assign sel_784557 = array_index_784404 == array_index_772864 ? add_784556 : sel_784553;
  assign add_784560 = sel_784557 + 8'h01;
  assign sel_784561 = array_index_784404 == array_index_772870 ? add_784560 : sel_784557;
  assign add_784564 = sel_784561 + 8'h01;
  assign sel_784565 = array_index_784404 == array_index_772876 ? add_784564 : sel_784561;
  assign add_784568 = sel_784565 + 8'h01;
  assign sel_784569 = array_index_784404 == array_index_772882 ? add_784568 : sel_784565;
  assign add_784572 = sel_784569 + 8'h01;
  assign sel_784573 = array_index_784404 == array_index_772888 ? add_784572 : sel_784569;
  assign add_784576 = sel_784573 + 8'h01;
  assign sel_784577 = array_index_784404 == array_index_772894 ? add_784576 : sel_784573;
  assign add_784580 = sel_784577 + 8'h01;
  assign sel_784581 = array_index_784404 == array_index_772900 ? add_784580 : sel_784577;
  assign add_784584 = sel_784581 + 8'h01;
  assign sel_784585 = array_index_784404 == array_index_772906 ? add_784584 : sel_784581;
  assign add_784588 = sel_784585 + 8'h01;
  assign sel_784589 = array_index_784404 == array_index_772912 ? add_784588 : sel_784585;
  assign add_784592 = sel_784589 + 8'h01;
  assign sel_784593 = array_index_784404 == array_index_772918 ? add_784592 : sel_784589;
  assign add_784596 = sel_784593 + 8'h01;
  assign sel_784597 = array_index_784404 == array_index_772924 ? add_784596 : sel_784593;
  assign add_784600 = sel_784597 + 8'h01;
  assign sel_784601 = array_index_784404 == array_index_772930 ? add_784600 : sel_784597;
  assign add_784604 = sel_784601 + 8'h01;
  assign sel_784605 = array_index_784404 == array_index_772936 ? add_784604 : sel_784601;
  assign add_784608 = sel_784605 + 8'h01;
  assign sel_784609 = array_index_784404 == array_index_772942 ? add_784608 : sel_784605;
  assign add_784612 = sel_784609 + 8'h01;
  assign sel_784613 = array_index_784404 == array_index_772948 ? add_784612 : sel_784609;
  assign add_784616 = sel_784613 + 8'h01;
  assign sel_784617 = array_index_784404 == array_index_772954 ? add_784616 : sel_784613;
  assign add_784620 = sel_784617 + 8'h01;
  assign sel_784621 = array_index_784404 == array_index_772960 ? add_784620 : sel_784617;
  assign add_784624 = sel_784621 + 8'h01;
  assign sel_784625 = array_index_784404 == array_index_772966 ? add_784624 : sel_784621;
  assign add_784628 = sel_784625 + 8'h01;
  assign sel_784629 = array_index_784404 == array_index_772972 ? add_784628 : sel_784625;
  assign add_784632 = sel_784629 + 8'h01;
  assign sel_784633 = array_index_784404 == array_index_772978 ? add_784632 : sel_784629;
  assign add_784636 = sel_784633 + 8'h01;
  assign sel_784637 = array_index_784404 == array_index_772984 ? add_784636 : sel_784633;
  assign add_784640 = sel_784637 + 8'h01;
  assign sel_784641 = array_index_784404 == array_index_772990 ? add_784640 : sel_784637;
  assign add_784644 = sel_784641 + 8'h01;
  assign sel_784645 = array_index_784404 == array_index_772996 ? add_784644 : sel_784641;
  assign add_784648 = sel_784645 + 8'h01;
  assign sel_784649 = array_index_784404 == array_index_773002 ? add_784648 : sel_784645;
  assign add_784652 = sel_784649 + 8'h01;
  assign sel_784653 = array_index_784404 == array_index_773008 ? add_784652 : sel_784649;
  assign add_784656 = sel_784653 + 8'h01;
  assign sel_784657 = array_index_784404 == array_index_773014 ? add_784656 : sel_784653;
  assign add_784660 = sel_784657 + 8'h01;
  assign sel_784661 = array_index_784404 == array_index_773020 ? add_784660 : sel_784657;
  assign add_784664 = sel_784661 + 8'h01;
  assign sel_784665 = array_index_784404 == array_index_773026 ? add_784664 : sel_784661;
  assign add_784668 = sel_784665 + 8'h01;
  assign sel_784669 = array_index_784404 == array_index_773032 ? add_784668 : sel_784665;
  assign add_784672 = sel_784669 + 8'h01;
  assign sel_784673 = array_index_784404 == array_index_773038 ? add_784672 : sel_784669;
  assign add_784676 = sel_784673 + 8'h01;
  assign sel_784677 = array_index_784404 == array_index_773044 ? add_784676 : sel_784673;
  assign add_784680 = sel_784677 + 8'h01;
  assign sel_784681 = array_index_784404 == array_index_773050 ? add_784680 : sel_784677;
  assign add_784684 = sel_784681 + 8'h01;
  assign sel_784685 = array_index_784404 == array_index_773056 ? add_784684 : sel_784681;
  assign add_784688 = sel_784685 + 8'h01;
  assign sel_784689 = array_index_784404 == array_index_773062 ? add_784688 : sel_784685;
  assign add_784692 = sel_784689 + 8'h01;
  assign sel_784693 = array_index_784404 == array_index_773068 ? add_784692 : sel_784689;
  assign add_784696 = sel_784693 + 8'h01;
  assign sel_784697 = array_index_784404 == array_index_773074 ? add_784696 : sel_784693;
  assign add_784700 = sel_784697 + 8'h01;
  assign sel_784701 = array_index_784404 == array_index_773080 ? add_784700 : sel_784697;
  assign add_784704 = sel_784701 + 8'h01;
  assign sel_784705 = array_index_784404 == array_index_773086 ? add_784704 : sel_784701;
  assign add_784708 = sel_784705 + 8'h01;
  assign sel_784709 = array_index_784404 == array_index_773092 ? add_784708 : sel_784705;
  assign add_784712 = sel_784709 + 8'h01;
  assign sel_784713 = array_index_784404 == array_index_773098 ? add_784712 : sel_784709;
  assign add_784716 = sel_784713 + 8'h01;
  assign sel_784717 = array_index_784404 == array_index_773104 ? add_784716 : sel_784713;
  assign add_784720 = sel_784717 + 8'h01;
  assign sel_784721 = array_index_784404 == array_index_773110 ? add_784720 : sel_784717;
  assign add_784724 = sel_784721 + 8'h01;
  assign sel_784725 = array_index_784404 == array_index_773116 ? add_784724 : sel_784721;
  assign add_784728 = sel_784725 + 8'h01;
  assign sel_784729 = array_index_784404 == array_index_773122 ? add_784728 : sel_784725;
  assign add_784732 = sel_784729 + 8'h01;
  assign sel_784733 = array_index_784404 == array_index_773128 ? add_784732 : sel_784729;
  assign add_784736 = sel_784733 + 8'h01;
  assign sel_784737 = array_index_784404 == array_index_773134 ? add_784736 : sel_784733;
  assign add_784740 = sel_784737 + 8'h01;
  assign sel_784741 = array_index_784404 == array_index_773140 ? add_784740 : sel_784737;
  assign add_784744 = sel_784741 + 8'h01;
  assign sel_784745 = array_index_784404 == array_index_773146 ? add_784744 : sel_784741;
  assign add_784748 = sel_784745 + 8'h01;
  assign sel_784749 = array_index_784404 == array_index_773152 ? add_784748 : sel_784745;
  assign add_784752 = sel_784749 + 8'h01;
  assign sel_784753 = array_index_784404 == array_index_773158 ? add_784752 : sel_784749;
  assign add_784756 = sel_784753 + 8'h01;
  assign sel_784757 = array_index_784404 == array_index_773164 ? add_784756 : sel_784753;
  assign add_784760 = sel_784757 + 8'h01;
  assign sel_784761 = array_index_784404 == array_index_773170 ? add_784760 : sel_784757;
  assign add_784765 = sel_784761 + 8'h01;
  assign array_index_784766 = set1_unflattened[7'h21];
  assign sel_784767 = array_index_784404 == array_index_773176 ? add_784765 : sel_784761;
  assign add_784770 = sel_784767 + 8'h01;
  assign sel_784771 = array_index_784766 == array_index_772632 ? add_784770 : sel_784767;
  assign add_784774 = sel_784771 + 8'h01;
  assign sel_784775 = array_index_784766 == array_index_772636 ? add_784774 : sel_784771;
  assign add_784778 = sel_784775 + 8'h01;
  assign sel_784779 = array_index_784766 == array_index_772644 ? add_784778 : sel_784775;
  assign add_784782 = sel_784779 + 8'h01;
  assign sel_784783 = array_index_784766 == array_index_772652 ? add_784782 : sel_784779;
  assign add_784786 = sel_784783 + 8'h01;
  assign sel_784787 = array_index_784766 == array_index_772660 ? add_784786 : sel_784783;
  assign add_784790 = sel_784787 + 8'h01;
  assign sel_784791 = array_index_784766 == array_index_772668 ? add_784790 : sel_784787;
  assign add_784794 = sel_784791 + 8'h01;
  assign sel_784795 = array_index_784766 == array_index_772676 ? add_784794 : sel_784791;
  assign add_784798 = sel_784795 + 8'h01;
  assign sel_784799 = array_index_784766 == array_index_772684 ? add_784798 : sel_784795;
  assign add_784802 = sel_784799 + 8'h01;
  assign sel_784803 = array_index_784766 == array_index_772690 ? add_784802 : sel_784799;
  assign add_784806 = sel_784803 + 8'h01;
  assign sel_784807 = array_index_784766 == array_index_772696 ? add_784806 : sel_784803;
  assign add_784810 = sel_784807 + 8'h01;
  assign sel_784811 = array_index_784766 == array_index_772702 ? add_784810 : sel_784807;
  assign add_784814 = sel_784811 + 8'h01;
  assign sel_784815 = array_index_784766 == array_index_772708 ? add_784814 : sel_784811;
  assign add_784818 = sel_784815 + 8'h01;
  assign sel_784819 = array_index_784766 == array_index_772714 ? add_784818 : sel_784815;
  assign add_784822 = sel_784819 + 8'h01;
  assign sel_784823 = array_index_784766 == array_index_772720 ? add_784822 : sel_784819;
  assign add_784826 = sel_784823 + 8'h01;
  assign sel_784827 = array_index_784766 == array_index_772726 ? add_784826 : sel_784823;
  assign add_784830 = sel_784827 + 8'h01;
  assign sel_784831 = array_index_784766 == array_index_772732 ? add_784830 : sel_784827;
  assign add_784834 = sel_784831 + 8'h01;
  assign sel_784835 = array_index_784766 == array_index_772738 ? add_784834 : sel_784831;
  assign add_784838 = sel_784835 + 8'h01;
  assign sel_784839 = array_index_784766 == array_index_772744 ? add_784838 : sel_784835;
  assign add_784842 = sel_784839 + 8'h01;
  assign sel_784843 = array_index_784766 == array_index_772750 ? add_784842 : sel_784839;
  assign add_784846 = sel_784843 + 8'h01;
  assign sel_784847 = array_index_784766 == array_index_772756 ? add_784846 : sel_784843;
  assign add_784850 = sel_784847 + 8'h01;
  assign sel_784851 = array_index_784766 == array_index_772762 ? add_784850 : sel_784847;
  assign add_784854 = sel_784851 + 8'h01;
  assign sel_784855 = array_index_784766 == array_index_772768 ? add_784854 : sel_784851;
  assign add_784858 = sel_784855 + 8'h01;
  assign sel_784859 = array_index_784766 == array_index_772774 ? add_784858 : sel_784855;
  assign add_784862 = sel_784859 + 8'h01;
  assign sel_784863 = array_index_784766 == array_index_772780 ? add_784862 : sel_784859;
  assign add_784866 = sel_784863 + 8'h01;
  assign sel_784867 = array_index_784766 == array_index_772786 ? add_784866 : sel_784863;
  assign add_784870 = sel_784867 + 8'h01;
  assign sel_784871 = array_index_784766 == array_index_772792 ? add_784870 : sel_784867;
  assign add_784874 = sel_784871 + 8'h01;
  assign sel_784875 = array_index_784766 == array_index_772798 ? add_784874 : sel_784871;
  assign add_784878 = sel_784875 + 8'h01;
  assign sel_784879 = array_index_784766 == array_index_772804 ? add_784878 : sel_784875;
  assign add_784882 = sel_784879 + 8'h01;
  assign sel_784883 = array_index_784766 == array_index_772810 ? add_784882 : sel_784879;
  assign add_784886 = sel_784883 + 8'h01;
  assign sel_784887 = array_index_784766 == array_index_772816 ? add_784886 : sel_784883;
  assign add_784890 = sel_784887 + 8'h01;
  assign sel_784891 = array_index_784766 == array_index_772822 ? add_784890 : sel_784887;
  assign add_784894 = sel_784891 + 8'h01;
  assign sel_784895 = array_index_784766 == array_index_772828 ? add_784894 : sel_784891;
  assign add_784898 = sel_784895 + 8'h01;
  assign sel_784899 = array_index_784766 == array_index_772834 ? add_784898 : sel_784895;
  assign add_784902 = sel_784899 + 8'h01;
  assign sel_784903 = array_index_784766 == array_index_772840 ? add_784902 : sel_784899;
  assign add_784906 = sel_784903 + 8'h01;
  assign sel_784907 = array_index_784766 == array_index_772846 ? add_784906 : sel_784903;
  assign add_784910 = sel_784907 + 8'h01;
  assign sel_784911 = array_index_784766 == array_index_772852 ? add_784910 : sel_784907;
  assign add_784914 = sel_784911 + 8'h01;
  assign sel_784915 = array_index_784766 == array_index_772858 ? add_784914 : sel_784911;
  assign add_784918 = sel_784915 + 8'h01;
  assign sel_784919 = array_index_784766 == array_index_772864 ? add_784918 : sel_784915;
  assign add_784922 = sel_784919 + 8'h01;
  assign sel_784923 = array_index_784766 == array_index_772870 ? add_784922 : sel_784919;
  assign add_784926 = sel_784923 + 8'h01;
  assign sel_784927 = array_index_784766 == array_index_772876 ? add_784926 : sel_784923;
  assign add_784930 = sel_784927 + 8'h01;
  assign sel_784931 = array_index_784766 == array_index_772882 ? add_784930 : sel_784927;
  assign add_784934 = sel_784931 + 8'h01;
  assign sel_784935 = array_index_784766 == array_index_772888 ? add_784934 : sel_784931;
  assign add_784938 = sel_784935 + 8'h01;
  assign sel_784939 = array_index_784766 == array_index_772894 ? add_784938 : sel_784935;
  assign add_784942 = sel_784939 + 8'h01;
  assign sel_784943 = array_index_784766 == array_index_772900 ? add_784942 : sel_784939;
  assign add_784946 = sel_784943 + 8'h01;
  assign sel_784947 = array_index_784766 == array_index_772906 ? add_784946 : sel_784943;
  assign add_784950 = sel_784947 + 8'h01;
  assign sel_784951 = array_index_784766 == array_index_772912 ? add_784950 : sel_784947;
  assign add_784954 = sel_784951 + 8'h01;
  assign sel_784955 = array_index_784766 == array_index_772918 ? add_784954 : sel_784951;
  assign add_784958 = sel_784955 + 8'h01;
  assign sel_784959 = array_index_784766 == array_index_772924 ? add_784958 : sel_784955;
  assign add_784962 = sel_784959 + 8'h01;
  assign sel_784963 = array_index_784766 == array_index_772930 ? add_784962 : sel_784959;
  assign add_784966 = sel_784963 + 8'h01;
  assign sel_784967 = array_index_784766 == array_index_772936 ? add_784966 : sel_784963;
  assign add_784970 = sel_784967 + 8'h01;
  assign sel_784971 = array_index_784766 == array_index_772942 ? add_784970 : sel_784967;
  assign add_784974 = sel_784971 + 8'h01;
  assign sel_784975 = array_index_784766 == array_index_772948 ? add_784974 : sel_784971;
  assign add_784978 = sel_784975 + 8'h01;
  assign sel_784979 = array_index_784766 == array_index_772954 ? add_784978 : sel_784975;
  assign add_784982 = sel_784979 + 8'h01;
  assign sel_784983 = array_index_784766 == array_index_772960 ? add_784982 : sel_784979;
  assign add_784986 = sel_784983 + 8'h01;
  assign sel_784987 = array_index_784766 == array_index_772966 ? add_784986 : sel_784983;
  assign add_784990 = sel_784987 + 8'h01;
  assign sel_784991 = array_index_784766 == array_index_772972 ? add_784990 : sel_784987;
  assign add_784994 = sel_784991 + 8'h01;
  assign sel_784995 = array_index_784766 == array_index_772978 ? add_784994 : sel_784991;
  assign add_784998 = sel_784995 + 8'h01;
  assign sel_784999 = array_index_784766 == array_index_772984 ? add_784998 : sel_784995;
  assign add_785002 = sel_784999 + 8'h01;
  assign sel_785003 = array_index_784766 == array_index_772990 ? add_785002 : sel_784999;
  assign add_785006 = sel_785003 + 8'h01;
  assign sel_785007 = array_index_784766 == array_index_772996 ? add_785006 : sel_785003;
  assign add_785010 = sel_785007 + 8'h01;
  assign sel_785011 = array_index_784766 == array_index_773002 ? add_785010 : sel_785007;
  assign add_785014 = sel_785011 + 8'h01;
  assign sel_785015 = array_index_784766 == array_index_773008 ? add_785014 : sel_785011;
  assign add_785018 = sel_785015 + 8'h01;
  assign sel_785019 = array_index_784766 == array_index_773014 ? add_785018 : sel_785015;
  assign add_785022 = sel_785019 + 8'h01;
  assign sel_785023 = array_index_784766 == array_index_773020 ? add_785022 : sel_785019;
  assign add_785026 = sel_785023 + 8'h01;
  assign sel_785027 = array_index_784766 == array_index_773026 ? add_785026 : sel_785023;
  assign add_785030 = sel_785027 + 8'h01;
  assign sel_785031 = array_index_784766 == array_index_773032 ? add_785030 : sel_785027;
  assign add_785034 = sel_785031 + 8'h01;
  assign sel_785035 = array_index_784766 == array_index_773038 ? add_785034 : sel_785031;
  assign add_785038 = sel_785035 + 8'h01;
  assign sel_785039 = array_index_784766 == array_index_773044 ? add_785038 : sel_785035;
  assign add_785042 = sel_785039 + 8'h01;
  assign sel_785043 = array_index_784766 == array_index_773050 ? add_785042 : sel_785039;
  assign add_785046 = sel_785043 + 8'h01;
  assign sel_785047 = array_index_784766 == array_index_773056 ? add_785046 : sel_785043;
  assign add_785050 = sel_785047 + 8'h01;
  assign sel_785051 = array_index_784766 == array_index_773062 ? add_785050 : sel_785047;
  assign add_785054 = sel_785051 + 8'h01;
  assign sel_785055 = array_index_784766 == array_index_773068 ? add_785054 : sel_785051;
  assign add_785058 = sel_785055 + 8'h01;
  assign sel_785059 = array_index_784766 == array_index_773074 ? add_785058 : sel_785055;
  assign add_785062 = sel_785059 + 8'h01;
  assign sel_785063 = array_index_784766 == array_index_773080 ? add_785062 : sel_785059;
  assign add_785066 = sel_785063 + 8'h01;
  assign sel_785067 = array_index_784766 == array_index_773086 ? add_785066 : sel_785063;
  assign add_785070 = sel_785067 + 8'h01;
  assign sel_785071 = array_index_784766 == array_index_773092 ? add_785070 : sel_785067;
  assign add_785074 = sel_785071 + 8'h01;
  assign sel_785075 = array_index_784766 == array_index_773098 ? add_785074 : sel_785071;
  assign add_785078 = sel_785075 + 8'h01;
  assign sel_785079 = array_index_784766 == array_index_773104 ? add_785078 : sel_785075;
  assign add_785082 = sel_785079 + 8'h01;
  assign sel_785083 = array_index_784766 == array_index_773110 ? add_785082 : sel_785079;
  assign add_785086 = sel_785083 + 8'h01;
  assign sel_785087 = array_index_784766 == array_index_773116 ? add_785086 : sel_785083;
  assign add_785090 = sel_785087 + 8'h01;
  assign sel_785091 = array_index_784766 == array_index_773122 ? add_785090 : sel_785087;
  assign add_785094 = sel_785091 + 8'h01;
  assign sel_785095 = array_index_784766 == array_index_773128 ? add_785094 : sel_785091;
  assign add_785098 = sel_785095 + 8'h01;
  assign sel_785099 = array_index_784766 == array_index_773134 ? add_785098 : sel_785095;
  assign add_785102 = sel_785099 + 8'h01;
  assign sel_785103 = array_index_784766 == array_index_773140 ? add_785102 : sel_785099;
  assign add_785106 = sel_785103 + 8'h01;
  assign sel_785107 = array_index_784766 == array_index_773146 ? add_785106 : sel_785103;
  assign add_785110 = sel_785107 + 8'h01;
  assign sel_785111 = array_index_784766 == array_index_773152 ? add_785110 : sel_785107;
  assign add_785114 = sel_785111 + 8'h01;
  assign sel_785115 = array_index_784766 == array_index_773158 ? add_785114 : sel_785111;
  assign add_785118 = sel_785115 + 8'h01;
  assign sel_785119 = array_index_784766 == array_index_773164 ? add_785118 : sel_785115;
  assign add_785122 = sel_785119 + 8'h01;
  assign sel_785123 = array_index_784766 == array_index_773170 ? add_785122 : sel_785119;
  assign add_785127 = sel_785123 + 8'h01;
  assign array_index_785128 = set1_unflattened[7'h22];
  assign sel_785129 = array_index_784766 == array_index_773176 ? add_785127 : sel_785123;
  assign add_785132 = sel_785129 + 8'h01;
  assign sel_785133 = array_index_785128 == array_index_772632 ? add_785132 : sel_785129;
  assign add_785136 = sel_785133 + 8'h01;
  assign sel_785137 = array_index_785128 == array_index_772636 ? add_785136 : sel_785133;
  assign add_785140 = sel_785137 + 8'h01;
  assign sel_785141 = array_index_785128 == array_index_772644 ? add_785140 : sel_785137;
  assign add_785144 = sel_785141 + 8'h01;
  assign sel_785145 = array_index_785128 == array_index_772652 ? add_785144 : sel_785141;
  assign add_785148 = sel_785145 + 8'h01;
  assign sel_785149 = array_index_785128 == array_index_772660 ? add_785148 : sel_785145;
  assign add_785152 = sel_785149 + 8'h01;
  assign sel_785153 = array_index_785128 == array_index_772668 ? add_785152 : sel_785149;
  assign add_785156 = sel_785153 + 8'h01;
  assign sel_785157 = array_index_785128 == array_index_772676 ? add_785156 : sel_785153;
  assign add_785160 = sel_785157 + 8'h01;
  assign sel_785161 = array_index_785128 == array_index_772684 ? add_785160 : sel_785157;
  assign add_785164 = sel_785161 + 8'h01;
  assign sel_785165 = array_index_785128 == array_index_772690 ? add_785164 : sel_785161;
  assign add_785168 = sel_785165 + 8'h01;
  assign sel_785169 = array_index_785128 == array_index_772696 ? add_785168 : sel_785165;
  assign add_785172 = sel_785169 + 8'h01;
  assign sel_785173 = array_index_785128 == array_index_772702 ? add_785172 : sel_785169;
  assign add_785176 = sel_785173 + 8'h01;
  assign sel_785177 = array_index_785128 == array_index_772708 ? add_785176 : sel_785173;
  assign add_785180 = sel_785177 + 8'h01;
  assign sel_785181 = array_index_785128 == array_index_772714 ? add_785180 : sel_785177;
  assign add_785184 = sel_785181 + 8'h01;
  assign sel_785185 = array_index_785128 == array_index_772720 ? add_785184 : sel_785181;
  assign add_785188 = sel_785185 + 8'h01;
  assign sel_785189 = array_index_785128 == array_index_772726 ? add_785188 : sel_785185;
  assign add_785192 = sel_785189 + 8'h01;
  assign sel_785193 = array_index_785128 == array_index_772732 ? add_785192 : sel_785189;
  assign add_785196 = sel_785193 + 8'h01;
  assign sel_785197 = array_index_785128 == array_index_772738 ? add_785196 : sel_785193;
  assign add_785200 = sel_785197 + 8'h01;
  assign sel_785201 = array_index_785128 == array_index_772744 ? add_785200 : sel_785197;
  assign add_785204 = sel_785201 + 8'h01;
  assign sel_785205 = array_index_785128 == array_index_772750 ? add_785204 : sel_785201;
  assign add_785208 = sel_785205 + 8'h01;
  assign sel_785209 = array_index_785128 == array_index_772756 ? add_785208 : sel_785205;
  assign add_785212 = sel_785209 + 8'h01;
  assign sel_785213 = array_index_785128 == array_index_772762 ? add_785212 : sel_785209;
  assign add_785216 = sel_785213 + 8'h01;
  assign sel_785217 = array_index_785128 == array_index_772768 ? add_785216 : sel_785213;
  assign add_785220 = sel_785217 + 8'h01;
  assign sel_785221 = array_index_785128 == array_index_772774 ? add_785220 : sel_785217;
  assign add_785224 = sel_785221 + 8'h01;
  assign sel_785225 = array_index_785128 == array_index_772780 ? add_785224 : sel_785221;
  assign add_785228 = sel_785225 + 8'h01;
  assign sel_785229 = array_index_785128 == array_index_772786 ? add_785228 : sel_785225;
  assign add_785232 = sel_785229 + 8'h01;
  assign sel_785233 = array_index_785128 == array_index_772792 ? add_785232 : sel_785229;
  assign add_785236 = sel_785233 + 8'h01;
  assign sel_785237 = array_index_785128 == array_index_772798 ? add_785236 : sel_785233;
  assign add_785240 = sel_785237 + 8'h01;
  assign sel_785241 = array_index_785128 == array_index_772804 ? add_785240 : sel_785237;
  assign add_785244 = sel_785241 + 8'h01;
  assign sel_785245 = array_index_785128 == array_index_772810 ? add_785244 : sel_785241;
  assign add_785248 = sel_785245 + 8'h01;
  assign sel_785249 = array_index_785128 == array_index_772816 ? add_785248 : sel_785245;
  assign add_785252 = sel_785249 + 8'h01;
  assign sel_785253 = array_index_785128 == array_index_772822 ? add_785252 : sel_785249;
  assign add_785256 = sel_785253 + 8'h01;
  assign sel_785257 = array_index_785128 == array_index_772828 ? add_785256 : sel_785253;
  assign add_785260 = sel_785257 + 8'h01;
  assign sel_785261 = array_index_785128 == array_index_772834 ? add_785260 : sel_785257;
  assign add_785264 = sel_785261 + 8'h01;
  assign sel_785265 = array_index_785128 == array_index_772840 ? add_785264 : sel_785261;
  assign add_785268 = sel_785265 + 8'h01;
  assign sel_785269 = array_index_785128 == array_index_772846 ? add_785268 : sel_785265;
  assign add_785272 = sel_785269 + 8'h01;
  assign sel_785273 = array_index_785128 == array_index_772852 ? add_785272 : sel_785269;
  assign add_785276 = sel_785273 + 8'h01;
  assign sel_785277 = array_index_785128 == array_index_772858 ? add_785276 : sel_785273;
  assign add_785280 = sel_785277 + 8'h01;
  assign sel_785281 = array_index_785128 == array_index_772864 ? add_785280 : sel_785277;
  assign add_785284 = sel_785281 + 8'h01;
  assign sel_785285 = array_index_785128 == array_index_772870 ? add_785284 : sel_785281;
  assign add_785288 = sel_785285 + 8'h01;
  assign sel_785289 = array_index_785128 == array_index_772876 ? add_785288 : sel_785285;
  assign add_785292 = sel_785289 + 8'h01;
  assign sel_785293 = array_index_785128 == array_index_772882 ? add_785292 : sel_785289;
  assign add_785296 = sel_785293 + 8'h01;
  assign sel_785297 = array_index_785128 == array_index_772888 ? add_785296 : sel_785293;
  assign add_785300 = sel_785297 + 8'h01;
  assign sel_785301 = array_index_785128 == array_index_772894 ? add_785300 : sel_785297;
  assign add_785304 = sel_785301 + 8'h01;
  assign sel_785305 = array_index_785128 == array_index_772900 ? add_785304 : sel_785301;
  assign add_785308 = sel_785305 + 8'h01;
  assign sel_785309 = array_index_785128 == array_index_772906 ? add_785308 : sel_785305;
  assign add_785312 = sel_785309 + 8'h01;
  assign sel_785313 = array_index_785128 == array_index_772912 ? add_785312 : sel_785309;
  assign add_785316 = sel_785313 + 8'h01;
  assign sel_785317 = array_index_785128 == array_index_772918 ? add_785316 : sel_785313;
  assign add_785320 = sel_785317 + 8'h01;
  assign sel_785321 = array_index_785128 == array_index_772924 ? add_785320 : sel_785317;
  assign add_785324 = sel_785321 + 8'h01;
  assign sel_785325 = array_index_785128 == array_index_772930 ? add_785324 : sel_785321;
  assign add_785328 = sel_785325 + 8'h01;
  assign sel_785329 = array_index_785128 == array_index_772936 ? add_785328 : sel_785325;
  assign add_785332 = sel_785329 + 8'h01;
  assign sel_785333 = array_index_785128 == array_index_772942 ? add_785332 : sel_785329;
  assign add_785336 = sel_785333 + 8'h01;
  assign sel_785337 = array_index_785128 == array_index_772948 ? add_785336 : sel_785333;
  assign add_785340 = sel_785337 + 8'h01;
  assign sel_785341 = array_index_785128 == array_index_772954 ? add_785340 : sel_785337;
  assign add_785344 = sel_785341 + 8'h01;
  assign sel_785345 = array_index_785128 == array_index_772960 ? add_785344 : sel_785341;
  assign add_785348 = sel_785345 + 8'h01;
  assign sel_785349 = array_index_785128 == array_index_772966 ? add_785348 : sel_785345;
  assign add_785352 = sel_785349 + 8'h01;
  assign sel_785353 = array_index_785128 == array_index_772972 ? add_785352 : sel_785349;
  assign add_785356 = sel_785353 + 8'h01;
  assign sel_785357 = array_index_785128 == array_index_772978 ? add_785356 : sel_785353;
  assign add_785360 = sel_785357 + 8'h01;
  assign sel_785361 = array_index_785128 == array_index_772984 ? add_785360 : sel_785357;
  assign add_785364 = sel_785361 + 8'h01;
  assign sel_785365 = array_index_785128 == array_index_772990 ? add_785364 : sel_785361;
  assign add_785368 = sel_785365 + 8'h01;
  assign sel_785369 = array_index_785128 == array_index_772996 ? add_785368 : sel_785365;
  assign add_785372 = sel_785369 + 8'h01;
  assign sel_785373 = array_index_785128 == array_index_773002 ? add_785372 : sel_785369;
  assign add_785376 = sel_785373 + 8'h01;
  assign sel_785377 = array_index_785128 == array_index_773008 ? add_785376 : sel_785373;
  assign add_785380 = sel_785377 + 8'h01;
  assign sel_785381 = array_index_785128 == array_index_773014 ? add_785380 : sel_785377;
  assign add_785384 = sel_785381 + 8'h01;
  assign sel_785385 = array_index_785128 == array_index_773020 ? add_785384 : sel_785381;
  assign add_785388 = sel_785385 + 8'h01;
  assign sel_785389 = array_index_785128 == array_index_773026 ? add_785388 : sel_785385;
  assign add_785392 = sel_785389 + 8'h01;
  assign sel_785393 = array_index_785128 == array_index_773032 ? add_785392 : sel_785389;
  assign add_785396 = sel_785393 + 8'h01;
  assign sel_785397 = array_index_785128 == array_index_773038 ? add_785396 : sel_785393;
  assign add_785400 = sel_785397 + 8'h01;
  assign sel_785401 = array_index_785128 == array_index_773044 ? add_785400 : sel_785397;
  assign add_785404 = sel_785401 + 8'h01;
  assign sel_785405 = array_index_785128 == array_index_773050 ? add_785404 : sel_785401;
  assign add_785408 = sel_785405 + 8'h01;
  assign sel_785409 = array_index_785128 == array_index_773056 ? add_785408 : sel_785405;
  assign add_785412 = sel_785409 + 8'h01;
  assign sel_785413 = array_index_785128 == array_index_773062 ? add_785412 : sel_785409;
  assign add_785416 = sel_785413 + 8'h01;
  assign sel_785417 = array_index_785128 == array_index_773068 ? add_785416 : sel_785413;
  assign add_785420 = sel_785417 + 8'h01;
  assign sel_785421 = array_index_785128 == array_index_773074 ? add_785420 : sel_785417;
  assign add_785424 = sel_785421 + 8'h01;
  assign sel_785425 = array_index_785128 == array_index_773080 ? add_785424 : sel_785421;
  assign add_785428 = sel_785425 + 8'h01;
  assign sel_785429 = array_index_785128 == array_index_773086 ? add_785428 : sel_785425;
  assign add_785432 = sel_785429 + 8'h01;
  assign sel_785433 = array_index_785128 == array_index_773092 ? add_785432 : sel_785429;
  assign add_785436 = sel_785433 + 8'h01;
  assign sel_785437 = array_index_785128 == array_index_773098 ? add_785436 : sel_785433;
  assign add_785440 = sel_785437 + 8'h01;
  assign sel_785441 = array_index_785128 == array_index_773104 ? add_785440 : sel_785437;
  assign add_785444 = sel_785441 + 8'h01;
  assign sel_785445 = array_index_785128 == array_index_773110 ? add_785444 : sel_785441;
  assign add_785448 = sel_785445 + 8'h01;
  assign sel_785449 = array_index_785128 == array_index_773116 ? add_785448 : sel_785445;
  assign add_785452 = sel_785449 + 8'h01;
  assign sel_785453 = array_index_785128 == array_index_773122 ? add_785452 : sel_785449;
  assign add_785456 = sel_785453 + 8'h01;
  assign sel_785457 = array_index_785128 == array_index_773128 ? add_785456 : sel_785453;
  assign add_785460 = sel_785457 + 8'h01;
  assign sel_785461 = array_index_785128 == array_index_773134 ? add_785460 : sel_785457;
  assign add_785464 = sel_785461 + 8'h01;
  assign sel_785465 = array_index_785128 == array_index_773140 ? add_785464 : sel_785461;
  assign add_785468 = sel_785465 + 8'h01;
  assign sel_785469 = array_index_785128 == array_index_773146 ? add_785468 : sel_785465;
  assign add_785472 = sel_785469 + 8'h01;
  assign sel_785473 = array_index_785128 == array_index_773152 ? add_785472 : sel_785469;
  assign add_785476 = sel_785473 + 8'h01;
  assign sel_785477 = array_index_785128 == array_index_773158 ? add_785476 : sel_785473;
  assign add_785480 = sel_785477 + 8'h01;
  assign sel_785481 = array_index_785128 == array_index_773164 ? add_785480 : sel_785477;
  assign add_785484 = sel_785481 + 8'h01;
  assign sel_785485 = array_index_785128 == array_index_773170 ? add_785484 : sel_785481;
  assign add_785489 = sel_785485 + 8'h01;
  assign array_index_785490 = set1_unflattened[7'h23];
  assign sel_785491 = array_index_785128 == array_index_773176 ? add_785489 : sel_785485;
  assign add_785494 = sel_785491 + 8'h01;
  assign sel_785495 = array_index_785490 == array_index_772632 ? add_785494 : sel_785491;
  assign add_785498 = sel_785495 + 8'h01;
  assign sel_785499 = array_index_785490 == array_index_772636 ? add_785498 : sel_785495;
  assign add_785502 = sel_785499 + 8'h01;
  assign sel_785503 = array_index_785490 == array_index_772644 ? add_785502 : sel_785499;
  assign add_785506 = sel_785503 + 8'h01;
  assign sel_785507 = array_index_785490 == array_index_772652 ? add_785506 : sel_785503;
  assign add_785510 = sel_785507 + 8'h01;
  assign sel_785511 = array_index_785490 == array_index_772660 ? add_785510 : sel_785507;
  assign add_785514 = sel_785511 + 8'h01;
  assign sel_785515 = array_index_785490 == array_index_772668 ? add_785514 : sel_785511;
  assign add_785518 = sel_785515 + 8'h01;
  assign sel_785519 = array_index_785490 == array_index_772676 ? add_785518 : sel_785515;
  assign add_785522 = sel_785519 + 8'h01;
  assign sel_785523 = array_index_785490 == array_index_772684 ? add_785522 : sel_785519;
  assign add_785526 = sel_785523 + 8'h01;
  assign sel_785527 = array_index_785490 == array_index_772690 ? add_785526 : sel_785523;
  assign add_785530 = sel_785527 + 8'h01;
  assign sel_785531 = array_index_785490 == array_index_772696 ? add_785530 : sel_785527;
  assign add_785534 = sel_785531 + 8'h01;
  assign sel_785535 = array_index_785490 == array_index_772702 ? add_785534 : sel_785531;
  assign add_785538 = sel_785535 + 8'h01;
  assign sel_785539 = array_index_785490 == array_index_772708 ? add_785538 : sel_785535;
  assign add_785542 = sel_785539 + 8'h01;
  assign sel_785543 = array_index_785490 == array_index_772714 ? add_785542 : sel_785539;
  assign add_785546 = sel_785543 + 8'h01;
  assign sel_785547 = array_index_785490 == array_index_772720 ? add_785546 : sel_785543;
  assign add_785550 = sel_785547 + 8'h01;
  assign sel_785551 = array_index_785490 == array_index_772726 ? add_785550 : sel_785547;
  assign add_785554 = sel_785551 + 8'h01;
  assign sel_785555 = array_index_785490 == array_index_772732 ? add_785554 : sel_785551;
  assign add_785558 = sel_785555 + 8'h01;
  assign sel_785559 = array_index_785490 == array_index_772738 ? add_785558 : sel_785555;
  assign add_785562 = sel_785559 + 8'h01;
  assign sel_785563 = array_index_785490 == array_index_772744 ? add_785562 : sel_785559;
  assign add_785566 = sel_785563 + 8'h01;
  assign sel_785567 = array_index_785490 == array_index_772750 ? add_785566 : sel_785563;
  assign add_785570 = sel_785567 + 8'h01;
  assign sel_785571 = array_index_785490 == array_index_772756 ? add_785570 : sel_785567;
  assign add_785574 = sel_785571 + 8'h01;
  assign sel_785575 = array_index_785490 == array_index_772762 ? add_785574 : sel_785571;
  assign add_785578 = sel_785575 + 8'h01;
  assign sel_785579 = array_index_785490 == array_index_772768 ? add_785578 : sel_785575;
  assign add_785582 = sel_785579 + 8'h01;
  assign sel_785583 = array_index_785490 == array_index_772774 ? add_785582 : sel_785579;
  assign add_785586 = sel_785583 + 8'h01;
  assign sel_785587 = array_index_785490 == array_index_772780 ? add_785586 : sel_785583;
  assign add_785590 = sel_785587 + 8'h01;
  assign sel_785591 = array_index_785490 == array_index_772786 ? add_785590 : sel_785587;
  assign add_785594 = sel_785591 + 8'h01;
  assign sel_785595 = array_index_785490 == array_index_772792 ? add_785594 : sel_785591;
  assign add_785598 = sel_785595 + 8'h01;
  assign sel_785599 = array_index_785490 == array_index_772798 ? add_785598 : sel_785595;
  assign add_785602 = sel_785599 + 8'h01;
  assign sel_785603 = array_index_785490 == array_index_772804 ? add_785602 : sel_785599;
  assign add_785606 = sel_785603 + 8'h01;
  assign sel_785607 = array_index_785490 == array_index_772810 ? add_785606 : sel_785603;
  assign add_785610 = sel_785607 + 8'h01;
  assign sel_785611 = array_index_785490 == array_index_772816 ? add_785610 : sel_785607;
  assign add_785614 = sel_785611 + 8'h01;
  assign sel_785615 = array_index_785490 == array_index_772822 ? add_785614 : sel_785611;
  assign add_785618 = sel_785615 + 8'h01;
  assign sel_785619 = array_index_785490 == array_index_772828 ? add_785618 : sel_785615;
  assign add_785622 = sel_785619 + 8'h01;
  assign sel_785623 = array_index_785490 == array_index_772834 ? add_785622 : sel_785619;
  assign add_785626 = sel_785623 + 8'h01;
  assign sel_785627 = array_index_785490 == array_index_772840 ? add_785626 : sel_785623;
  assign add_785630 = sel_785627 + 8'h01;
  assign sel_785631 = array_index_785490 == array_index_772846 ? add_785630 : sel_785627;
  assign add_785634 = sel_785631 + 8'h01;
  assign sel_785635 = array_index_785490 == array_index_772852 ? add_785634 : sel_785631;
  assign add_785638 = sel_785635 + 8'h01;
  assign sel_785639 = array_index_785490 == array_index_772858 ? add_785638 : sel_785635;
  assign add_785642 = sel_785639 + 8'h01;
  assign sel_785643 = array_index_785490 == array_index_772864 ? add_785642 : sel_785639;
  assign add_785646 = sel_785643 + 8'h01;
  assign sel_785647 = array_index_785490 == array_index_772870 ? add_785646 : sel_785643;
  assign add_785650 = sel_785647 + 8'h01;
  assign sel_785651 = array_index_785490 == array_index_772876 ? add_785650 : sel_785647;
  assign add_785654 = sel_785651 + 8'h01;
  assign sel_785655 = array_index_785490 == array_index_772882 ? add_785654 : sel_785651;
  assign add_785658 = sel_785655 + 8'h01;
  assign sel_785659 = array_index_785490 == array_index_772888 ? add_785658 : sel_785655;
  assign add_785662 = sel_785659 + 8'h01;
  assign sel_785663 = array_index_785490 == array_index_772894 ? add_785662 : sel_785659;
  assign add_785666 = sel_785663 + 8'h01;
  assign sel_785667 = array_index_785490 == array_index_772900 ? add_785666 : sel_785663;
  assign add_785670 = sel_785667 + 8'h01;
  assign sel_785671 = array_index_785490 == array_index_772906 ? add_785670 : sel_785667;
  assign add_785674 = sel_785671 + 8'h01;
  assign sel_785675 = array_index_785490 == array_index_772912 ? add_785674 : sel_785671;
  assign add_785678 = sel_785675 + 8'h01;
  assign sel_785679 = array_index_785490 == array_index_772918 ? add_785678 : sel_785675;
  assign add_785682 = sel_785679 + 8'h01;
  assign sel_785683 = array_index_785490 == array_index_772924 ? add_785682 : sel_785679;
  assign add_785686 = sel_785683 + 8'h01;
  assign sel_785687 = array_index_785490 == array_index_772930 ? add_785686 : sel_785683;
  assign add_785690 = sel_785687 + 8'h01;
  assign sel_785691 = array_index_785490 == array_index_772936 ? add_785690 : sel_785687;
  assign add_785694 = sel_785691 + 8'h01;
  assign sel_785695 = array_index_785490 == array_index_772942 ? add_785694 : sel_785691;
  assign add_785698 = sel_785695 + 8'h01;
  assign sel_785699 = array_index_785490 == array_index_772948 ? add_785698 : sel_785695;
  assign add_785702 = sel_785699 + 8'h01;
  assign sel_785703 = array_index_785490 == array_index_772954 ? add_785702 : sel_785699;
  assign add_785706 = sel_785703 + 8'h01;
  assign sel_785707 = array_index_785490 == array_index_772960 ? add_785706 : sel_785703;
  assign add_785710 = sel_785707 + 8'h01;
  assign sel_785711 = array_index_785490 == array_index_772966 ? add_785710 : sel_785707;
  assign add_785714 = sel_785711 + 8'h01;
  assign sel_785715 = array_index_785490 == array_index_772972 ? add_785714 : sel_785711;
  assign add_785718 = sel_785715 + 8'h01;
  assign sel_785719 = array_index_785490 == array_index_772978 ? add_785718 : sel_785715;
  assign add_785722 = sel_785719 + 8'h01;
  assign sel_785723 = array_index_785490 == array_index_772984 ? add_785722 : sel_785719;
  assign add_785726 = sel_785723 + 8'h01;
  assign sel_785727 = array_index_785490 == array_index_772990 ? add_785726 : sel_785723;
  assign add_785730 = sel_785727 + 8'h01;
  assign sel_785731 = array_index_785490 == array_index_772996 ? add_785730 : sel_785727;
  assign add_785734 = sel_785731 + 8'h01;
  assign sel_785735 = array_index_785490 == array_index_773002 ? add_785734 : sel_785731;
  assign add_785738 = sel_785735 + 8'h01;
  assign sel_785739 = array_index_785490 == array_index_773008 ? add_785738 : sel_785735;
  assign add_785742 = sel_785739 + 8'h01;
  assign sel_785743 = array_index_785490 == array_index_773014 ? add_785742 : sel_785739;
  assign add_785746 = sel_785743 + 8'h01;
  assign sel_785747 = array_index_785490 == array_index_773020 ? add_785746 : sel_785743;
  assign add_785750 = sel_785747 + 8'h01;
  assign sel_785751 = array_index_785490 == array_index_773026 ? add_785750 : sel_785747;
  assign add_785754 = sel_785751 + 8'h01;
  assign sel_785755 = array_index_785490 == array_index_773032 ? add_785754 : sel_785751;
  assign add_785758 = sel_785755 + 8'h01;
  assign sel_785759 = array_index_785490 == array_index_773038 ? add_785758 : sel_785755;
  assign add_785762 = sel_785759 + 8'h01;
  assign sel_785763 = array_index_785490 == array_index_773044 ? add_785762 : sel_785759;
  assign add_785766 = sel_785763 + 8'h01;
  assign sel_785767 = array_index_785490 == array_index_773050 ? add_785766 : sel_785763;
  assign add_785770 = sel_785767 + 8'h01;
  assign sel_785771 = array_index_785490 == array_index_773056 ? add_785770 : sel_785767;
  assign add_785774 = sel_785771 + 8'h01;
  assign sel_785775 = array_index_785490 == array_index_773062 ? add_785774 : sel_785771;
  assign add_785778 = sel_785775 + 8'h01;
  assign sel_785779 = array_index_785490 == array_index_773068 ? add_785778 : sel_785775;
  assign add_785782 = sel_785779 + 8'h01;
  assign sel_785783 = array_index_785490 == array_index_773074 ? add_785782 : sel_785779;
  assign add_785786 = sel_785783 + 8'h01;
  assign sel_785787 = array_index_785490 == array_index_773080 ? add_785786 : sel_785783;
  assign add_785790 = sel_785787 + 8'h01;
  assign sel_785791 = array_index_785490 == array_index_773086 ? add_785790 : sel_785787;
  assign add_785794 = sel_785791 + 8'h01;
  assign sel_785795 = array_index_785490 == array_index_773092 ? add_785794 : sel_785791;
  assign add_785798 = sel_785795 + 8'h01;
  assign sel_785799 = array_index_785490 == array_index_773098 ? add_785798 : sel_785795;
  assign add_785802 = sel_785799 + 8'h01;
  assign sel_785803 = array_index_785490 == array_index_773104 ? add_785802 : sel_785799;
  assign add_785806 = sel_785803 + 8'h01;
  assign sel_785807 = array_index_785490 == array_index_773110 ? add_785806 : sel_785803;
  assign add_785810 = sel_785807 + 8'h01;
  assign sel_785811 = array_index_785490 == array_index_773116 ? add_785810 : sel_785807;
  assign add_785814 = sel_785811 + 8'h01;
  assign sel_785815 = array_index_785490 == array_index_773122 ? add_785814 : sel_785811;
  assign add_785818 = sel_785815 + 8'h01;
  assign sel_785819 = array_index_785490 == array_index_773128 ? add_785818 : sel_785815;
  assign add_785822 = sel_785819 + 8'h01;
  assign sel_785823 = array_index_785490 == array_index_773134 ? add_785822 : sel_785819;
  assign add_785826 = sel_785823 + 8'h01;
  assign sel_785827 = array_index_785490 == array_index_773140 ? add_785826 : sel_785823;
  assign add_785830 = sel_785827 + 8'h01;
  assign sel_785831 = array_index_785490 == array_index_773146 ? add_785830 : sel_785827;
  assign add_785834 = sel_785831 + 8'h01;
  assign sel_785835 = array_index_785490 == array_index_773152 ? add_785834 : sel_785831;
  assign add_785838 = sel_785835 + 8'h01;
  assign sel_785839 = array_index_785490 == array_index_773158 ? add_785838 : sel_785835;
  assign add_785842 = sel_785839 + 8'h01;
  assign sel_785843 = array_index_785490 == array_index_773164 ? add_785842 : sel_785839;
  assign add_785846 = sel_785843 + 8'h01;
  assign sel_785847 = array_index_785490 == array_index_773170 ? add_785846 : sel_785843;
  assign add_785851 = sel_785847 + 8'h01;
  assign array_index_785852 = set1_unflattened[7'h24];
  assign sel_785853 = array_index_785490 == array_index_773176 ? add_785851 : sel_785847;
  assign add_785856 = sel_785853 + 8'h01;
  assign sel_785857 = array_index_785852 == array_index_772632 ? add_785856 : sel_785853;
  assign add_785860 = sel_785857 + 8'h01;
  assign sel_785861 = array_index_785852 == array_index_772636 ? add_785860 : sel_785857;
  assign add_785864 = sel_785861 + 8'h01;
  assign sel_785865 = array_index_785852 == array_index_772644 ? add_785864 : sel_785861;
  assign add_785868 = sel_785865 + 8'h01;
  assign sel_785869 = array_index_785852 == array_index_772652 ? add_785868 : sel_785865;
  assign add_785872 = sel_785869 + 8'h01;
  assign sel_785873 = array_index_785852 == array_index_772660 ? add_785872 : sel_785869;
  assign add_785876 = sel_785873 + 8'h01;
  assign sel_785877 = array_index_785852 == array_index_772668 ? add_785876 : sel_785873;
  assign add_785880 = sel_785877 + 8'h01;
  assign sel_785881 = array_index_785852 == array_index_772676 ? add_785880 : sel_785877;
  assign add_785884 = sel_785881 + 8'h01;
  assign sel_785885 = array_index_785852 == array_index_772684 ? add_785884 : sel_785881;
  assign add_785888 = sel_785885 + 8'h01;
  assign sel_785889 = array_index_785852 == array_index_772690 ? add_785888 : sel_785885;
  assign add_785892 = sel_785889 + 8'h01;
  assign sel_785893 = array_index_785852 == array_index_772696 ? add_785892 : sel_785889;
  assign add_785896 = sel_785893 + 8'h01;
  assign sel_785897 = array_index_785852 == array_index_772702 ? add_785896 : sel_785893;
  assign add_785900 = sel_785897 + 8'h01;
  assign sel_785901 = array_index_785852 == array_index_772708 ? add_785900 : sel_785897;
  assign add_785904 = sel_785901 + 8'h01;
  assign sel_785905 = array_index_785852 == array_index_772714 ? add_785904 : sel_785901;
  assign add_785908 = sel_785905 + 8'h01;
  assign sel_785909 = array_index_785852 == array_index_772720 ? add_785908 : sel_785905;
  assign add_785912 = sel_785909 + 8'h01;
  assign sel_785913 = array_index_785852 == array_index_772726 ? add_785912 : sel_785909;
  assign add_785916 = sel_785913 + 8'h01;
  assign sel_785917 = array_index_785852 == array_index_772732 ? add_785916 : sel_785913;
  assign add_785920 = sel_785917 + 8'h01;
  assign sel_785921 = array_index_785852 == array_index_772738 ? add_785920 : sel_785917;
  assign add_785924 = sel_785921 + 8'h01;
  assign sel_785925 = array_index_785852 == array_index_772744 ? add_785924 : sel_785921;
  assign add_785928 = sel_785925 + 8'h01;
  assign sel_785929 = array_index_785852 == array_index_772750 ? add_785928 : sel_785925;
  assign add_785932 = sel_785929 + 8'h01;
  assign sel_785933 = array_index_785852 == array_index_772756 ? add_785932 : sel_785929;
  assign add_785936 = sel_785933 + 8'h01;
  assign sel_785937 = array_index_785852 == array_index_772762 ? add_785936 : sel_785933;
  assign add_785940 = sel_785937 + 8'h01;
  assign sel_785941 = array_index_785852 == array_index_772768 ? add_785940 : sel_785937;
  assign add_785944 = sel_785941 + 8'h01;
  assign sel_785945 = array_index_785852 == array_index_772774 ? add_785944 : sel_785941;
  assign add_785948 = sel_785945 + 8'h01;
  assign sel_785949 = array_index_785852 == array_index_772780 ? add_785948 : sel_785945;
  assign add_785952 = sel_785949 + 8'h01;
  assign sel_785953 = array_index_785852 == array_index_772786 ? add_785952 : sel_785949;
  assign add_785956 = sel_785953 + 8'h01;
  assign sel_785957 = array_index_785852 == array_index_772792 ? add_785956 : sel_785953;
  assign add_785960 = sel_785957 + 8'h01;
  assign sel_785961 = array_index_785852 == array_index_772798 ? add_785960 : sel_785957;
  assign add_785964 = sel_785961 + 8'h01;
  assign sel_785965 = array_index_785852 == array_index_772804 ? add_785964 : sel_785961;
  assign add_785968 = sel_785965 + 8'h01;
  assign sel_785969 = array_index_785852 == array_index_772810 ? add_785968 : sel_785965;
  assign add_785972 = sel_785969 + 8'h01;
  assign sel_785973 = array_index_785852 == array_index_772816 ? add_785972 : sel_785969;
  assign add_785976 = sel_785973 + 8'h01;
  assign sel_785977 = array_index_785852 == array_index_772822 ? add_785976 : sel_785973;
  assign add_785980 = sel_785977 + 8'h01;
  assign sel_785981 = array_index_785852 == array_index_772828 ? add_785980 : sel_785977;
  assign add_785984 = sel_785981 + 8'h01;
  assign sel_785985 = array_index_785852 == array_index_772834 ? add_785984 : sel_785981;
  assign add_785988 = sel_785985 + 8'h01;
  assign sel_785989 = array_index_785852 == array_index_772840 ? add_785988 : sel_785985;
  assign add_785992 = sel_785989 + 8'h01;
  assign sel_785993 = array_index_785852 == array_index_772846 ? add_785992 : sel_785989;
  assign add_785996 = sel_785993 + 8'h01;
  assign sel_785997 = array_index_785852 == array_index_772852 ? add_785996 : sel_785993;
  assign add_786000 = sel_785997 + 8'h01;
  assign sel_786001 = array_index_785852 == array_index_772858 ? add_786000 : sel_785997;
  assign add_786004 = sel_786001 + 8'h01;
  assign sel_786005 = array_index_785852 == array_index_772864 ? add_786004 : sel_786001;
  assign add_786008 = sel_786005 + 8'h01;
  assign sel_786009 = array_index_785852 == array_index_772870 ? add_786008 : sel_786005;
  assign add_786012 = sel_786009 + 8'h01;
  assign sel_786013 = array_index_785852 == array_index_772876 ? add_786012 : sel_786009;
  assign add_786016 = sel_786013 + 8'h01;
  assign sel_786017 = array_index_785852 == array_index_772882 ? add_786016 : sel_786013;
  assign add_786020 = sel_786017 + 8'h01;
  assign sel_786021 = array_index_785852 == array_index_772888 ? add_786020 : sel_786017;
  assign add_786024 = sel_786021 + 8'h01;
  assign sel_786025 = array_index_785852 == array_index_772894 ? add_786024 : sel_786021;
  assign add_786028 = sel_786025 + 8'h01;
  assign sel_786029 = array_index_785852 == array_index_772900 ? add_786028 : sel_786025;
  assign add_786032 = sel_786029 + 8'h01;
  assign sel_786033 = array_index_785852 == array_index_772906 ? add_786032 : sel_786029;
  assign add_786036 = sel_786033 + 8'h01;
  assign sel_786037 = array_index_785852 == array_index_772912 ? add_786036 : sel_786033;
  assign add_786040 = sel_786037 + 8'h01;
  assign sel_786041 = array_index_785852 == array_index_772918 ? add_786040 : sel_786037;
  assign add_786044 = sel_786041 + 8'h01;
  assign sel_786045 = array_index_785852 == array_index_772924 ? add_786044 : sel_786041;
  assign add_786048 = sel_786045 + 8'h01;
  assign sel_786049 = array_index_785852 == array_index_772930 ? add_786048 : sel_786045;
  assign add_786052 = sel_786049 + 8'h01;
  assign sel_786053 = array_index_785852 == array_index_772936 ? add_786052 : sel_786049;
  assign add_786056 = sel_786053 + 8'h01;
  assign sel_786057 = array_index_785852 == array_index_772942 ? add_786056 : sel_786053;
  assign add_786060 = sel_786057 + 8'h01;
  assign sel_786061 = array_index_785852 == array_index_772948 ? add_786060 : sel_786057;
  assign add_786064 = sel_786061 + 8'h01;
  assign sel_786065 = array_index_785852 == array_index_772954 ? add_786064 : sel_786061;
  assign add_786068 = sel_786065 + 8'h01;
  assign sel_786069 = array_index_785852 == array_index_772960 ? add_786068 : sel_786065;
  assign add_786072 = sel_786069 + 8'h01;
  assign sel_786073 = array_index_785852 == array_index_772966 ? add_786072 : sel_786069;
  assign add_786076 = sel_786073 + 8'h01;
  assign sel_786077 = array_index_785852 == array_index_772972 ? add_786076 : sel_786073;
  assign add_786080 = sel_786077 + 8'h01;
  assign sel_786081 = array_index_785852 == array_index_772978 ? add_786080 : sel_786077;
  assign add_786084 = sel_786081 + 8'h01;
  assign sel_786085 = array_index_785852 == array_index_772984 ? add_786084 : sel_786081;
  assign add_786088 = sel_786085 + 8'h01;
  assign sel_786089 = array_index_785852 == array_index_772990 ? add_786088 : sel_786085;
  assign add_786092 = sel_786089 + 8'h01;
  assign sel_786093 = array_index_785852 == array_index_772996 ? add_786092 : sel_786089;
  assign add_786096 = sel_786093 + 8'h01;
  assign sel_786097 = array_index_785852 == array_index_773002 ? add_786096 : sel_786093;
  assign add_786100 = sel_786097 + 8'h01;
  assign sel_786101 = array_index_785852 == array_index_773008 ? add_786100 : sel_786097;
  assign add_786104 = sel_786101 + 8'h01;
  assign sel_786105 = array_index_785852 == array_index_773014 ? add_786104 : sel_786101;
  assign add_786108 = sel_786105 + 8'h01;
  assign sel_786109 = array_index_785852 == array_index_773020 ? add_786108 : sel_786105;
  assign add_786112 = sel_786109 + 8'h01;
  assign sel_786113 = array_index_785852 == array_index_773026 ? add_786112 : sel_786109;
  assign add_786116 = sel_786113 + 8'h01;
  assign sel_786117 = array_index_785852 == array_index_773032 ? add_786116 : sel_786113;
  assign add_786120 = sel_786117 + 8'h01;
  assign sel_786121 = array_index_785852 == array_index_773038 ? add_786120 : sel_786117;
  assign add_786124 = sel_786121 + 8'h01;
  assign sel_786125 = array_index_785852 == array_index_773044 ? add_786124 : sel_786121;
  assign add_786128 = sel_786125 + 8'h01;
  assign sel_786129 = array_index_785852 == array_index_773050 ? add_786128 : sel_786125;
  assign add_786132 = sel_786129 + 8'h01;
  assign sel_786133 = array_index_785852 == array_index_773056 ? add_786132 : sel_786129;
  assign add_786136 = sel_786133 + 8'h01;
  assign sel_786137 = array_index_785852 == array_index_773062 ? add_786136 : sel_786133;
  assign add_786140 = sel_786137 + 8'h01;
  assign sel_786141 = array_index_785852 == array_index_773068 ? add_786140 : sel_786137;
  assign add_786144 = sel_786141 + 8'h01;
  assign sel_786145 = array_index_785852 == array_index_773074 ? add_786144 : sel_786141;
  assign add_786148 = sel_786145 + 8'h01;
  assign sel_786149 = array_index_785852 == array_index_773080 ? add_786148 : sel_786145;
  assign add_786152 = sel_786149 + 8'h01;
  assign sel_786153 = array_index_785852 == array_index_773086 ? add_786152 : sel_786149;
  assign add_786156 = sel_786153 + 8'h01;
  assign sel_786157 = array_index_785852 == array_index_773092 ? add_786156 : sel_786153;
  assign add_786160 = sel_786157 + 8'h01;
  assign sel_786161 = array_index_785852 == array_index_773098 ? add_786160 : sel_786157;
  assign add_786164 = sel_786161 + 8'h01;
  assign sel_786165 = array_index_785852 == array_index_773104 ? add_786164 : sel_786161;
  assign add_786168 = sel_786165 + 8'h01;
  assign sel_786169 = array_index_785852 == array_index_773110 ? add_786168 : sel_786165;
  assign add_786172 = sel_786169 + 8'h01;
  assign sel_786173 = array_index_785852 == array_index_773116 ? add_786172 : sel_786169;
  assign add_786176 = sel_786173 + 8'h01;
  assign sel_786177 = array_index_785852 == array_index_773122 ? add_786176 : sel_786173;
  assign add_786180 = sel_786177 + 8'h01;
  assign sel_786181 = array_index_785852 == array_index_773128 ? add_786180 : sel_786177;
  assign add_786184 = sel_786181 + 8'h01;
  assign sel_786185 = array_index_785852 == array_index_773134 ? add_786184 : sel_786181;
  assign add_786188 = sel_786185 + 8'h01;
  assign sel_786189 = array_index_785852 == array_index_773140 ? add_786188 : sel_786185;
  assign add_786192 = sel_786189 + 8'h01;
  assign sel_786193 = array_index_785852 == array_index_773146 ? add_786192 : sel_786189;
  assign add_786196 = sel_786193 + 8'h01;
  assign sel_786197 = array_index_785852 == array_index_773152 ? add_786196 : sel_786193;
  assign add_786200 = sel_786197 + 8'h01;
  assign sel_786201 = array_index_785852 == array_index_773158 ? add_786200 : sel_786197;
  assign add_786204 = sel_786201 + 8'h01;
  assign sel_786205 = array_index_785852 == array_index_773164 ? add_786204 : sel_786201;
  assign add_786208 = sel_786205 + 8'h01;
  assign sel_786209 = array_index_785852 == array_index_773170 ? add_786208 : sel_786205;
  assign add_786213 = sel_786209 + 8'h01;
  assign array_index_786214 = set1_unflattened[7'h25];
  assign sel_786215 = array_index_785852 == array_index_773176 ? add_786213 : sel_786209;
  assign add_786218 = sel_786215 + 8'h01;
  assign sel_786219 = array_index_786214 == array_index_772632 ? add_786218 : sel_786215;
  assign add_786222 = sel_786219 + 8'h01;
  assign sel_786223 = array_index_786214 == array_index_772636 ? add_786222 : sel_786219;
  assign add_786226 = sel_786223 + 8'h01;
  assign sel_786227 = array_index_786214 == array_index_772644 ? add_786226 : sel_786223;
  assign add_786230 = sel_786227 + 8'h01;
  assign sel_786231 = array_index_786214 == array_index_772652 ? add_786230 : sel_786227;
  assign add_786234 = sel_786231 + 8'h01;
  assign sel_786235 = array_index_786214 == array_index_772660 ? add_786234 : sel_786231;
  assign add_786238 = sel_786235 + 8'h01;
  assign sel_786239 = array_index_786214 == array_index_772668 ? add_786238 : sel_786235;
  assign add_786242 = sel_786239 + 8'h01;
  assign sel_786243 = array_index_786214 == array_index_772676 ? add_786242 : sel_786239;
  assign add_786246 = sel_786243 + 8'h01;
  assign sel_786247 = array_index_786214 == array_index_772684 ? add_786246 : sel_786243;
  assign add_786250 = sel_786247 + 8'h01;
  assign sel_786251 = array_index_786214 == array_index_772690 ? add_786250 : sel_786247;
  assign add_786254 = sel_786251 + 8'h01;
  assign sel_786255 = array_index_786214 == array_index_772696 ? add_786254 : sel_786251;
  assign add_786258 = sel_786255 + 8'h01;
  assign sel_786259 = array_index_786214 == array_index_772702 ? add_786258 : sel_786255;
  assign add_786262 = sel_786259 + 8'h01;
  assign sel_786263 = array_index_786214 == array_index_772708 ? add_786262 : sel_786259;
  assign add_786266 = sel_786263 + 8'h01;
  assign sel_786267 = array_index_786214 == array_index_772714 ? add_786266 : sel_786263;
  assign add_786270 = sel_786267 + 8'h01;
  assign sel_786271 = array_index_786214 == array_index_772720 ? add_786270 : sel_786267;
  assign add_786274 = sel_786271 + 8'h01;
  assign sel_786275 = array_index_786214 == array_index_772726 ? add_786274 : sel_786271;
  assign add_786278 = sel_786275 + 8'h01;
  assign sel_786279 = array_index_786214 == array_index_772732 ? add_786278 : sel_786275;
  assign add_786282 = sel_786279 + 8'h01;
  assign sel_786283 = array_index_786214 == array_index_772738 ? add_786282 : sel_786279;
  assign add_786286 = sel_786283 + 8'h01;
  assign sel_786287 = array_index_786214 == array_index_772744 ? add_786286 : sel_786283;
  assign add_786290 = sel_786287 + 8'h01;
  assign sel_786291 = array_index_786214 == array_index_772750 ? add_786290 : sel_786287;
  assign add_786294 = sel_786291 + 8'h01;
  assign sel_786295 = array_index_786214 == array_index_772756 ? add_786294 : sel_786291;
  assign add_786298 = sel_786295 + 8'h01;
  assign sel_786299 = array_index_786214 == array_index_772762 ? add_786298 : sel_786295;
  assign add_786302 = sel_786299 + 8'h01;
  assign sel_786303 = array_index_786214 == array_index_772768 ? add_786302 : sel_786299;
  assign add_786306 = sel_786303 + 8'h01;
  assign sel_786307 = array_index_786214 == array_index_772774 ? add_786306 : sel_786303;
  assign add_786310 = sel_786307 + 8'h01;
  assign sel_786311 = array_index_786214 == array_index_772780 ? add_786310 : sel_786307;
  assign add_786314 = sel_786311 + 8'h01;
  assign sel_786315 = array_index_786214 == array_index_772786 ? add_786314 : sel_786311;
  assign add_786318 = sel_786315 + 8'h01;
  assign sel_786319 = array_index_786214 == array_index_772792 ? add_786318 : sel_786315;
  assign add_786322 = sel_786319 + 8'h01;
  assign sel_786323 = array_index_786214 == array_index_772798 ? add_786322 : sel_786319;
  assign add_786326 = sel_786323 + 8'h01;
  assign sel_786327 = array_index_786214 == array_index_772804 ? add_786326 : sel_786323;
  assign add_786330 = sel_786327 + 8'h01;
  assign sel_786331 = array_index_786214 == array_index_772810 ? add_786330 : sel_786327;
  assign add_786334 = sel_786331 + 8'h01;
  assign sel_786335 = array_index_786214 == array_index_772816 ? add_786334 : sel_786331;
  assign add_786338 = sel_786335 + 8'h01;
  assign sel_786339 = array_index_786214 == array_index_772822 ? add_786338 : sel_786335;
  assign add_786342 = sel_786339 + 8'h01;
  assign sel_786343 = array_index_786214 == array_index_772828 ? add_786342 : sel_786339;
  assign add_786346 = sel_786343 + 8'h01;
  assign sel_786347 = array_index_786214 == array_index_772834 ? add_786346 : sel_786343;
  assign add_786350 = sel_786347 + 8'h01;
  assign sel_786351 = array_index_786214 == array_index_772840 ? add_786350 : sel_786347;
  assign add_786354 = sel_786351 + 8'h01;
  assign sel_786355 = array_index_786214 == array_index_772846 ? add_786354 : sel_786351;
  assign add_786358 = sel_786355 + 8'h01;
  assign sel_786359 = array_index_786214 == array_index_772852 ? add_786358 : sel_786355;
  assign add_786362 = sel_786359 + 8'h01;
  assign sel_786363 = array_index_786214 == array_index_772858 ? add_786362 : sel_786359;
  assign add_786366 = sel_786363 + 8'h01;
  assign sel_786367 = array_index_786214 == array_index_772864 ? add_786366 : sel_786363;
  assign add_786370 = sel_786367 + 8'h01;
  assign sel_786371 = array_index_786214 == array_index_772870 ? add_786370 : sel_786367;
  assign add_786374 = sel_786371 + 8'h01;
  assign sel_786375 = array_index_786214 == array_index_772876 ? add_786374 : sel_786371;
  assign add_786378 = sel_786375 + 8'h01;
  assign sel_786379 = array_index_786214 == array_index_772882 ? add_786378 : sel_786375;
  assign add_786382 = sel_786379 + 8'h01;
  assign sel_786383 = array_index_786214 == array_index_772888 ? add_786382 : sel_786379;
  assign add_786386 = sel_786383 + 8'h01;
  assign sel_786387 = array_index_786214 == array_index_772894 ? add_786386 : sel_786383;
  assign add_786390 = sel_786387 + 8'h01;
  assign sel_786391 = array_index_786214 == array_index_772900 ? add_786390 : sel_786387;
  assign add_786394 = sel_786391 + 8'h01;
  assign sel_786395 = array_index_786214 == array_index_772906 ? add_786394 : sel_786391;
  assign add_786398 = sel_786395 + 8'h01;
  assign sel_786399 = array_index_786214 == array_index_772912 ? add_786398 : sel_786395;
  assign add_786402 = sel_786399 + 8'h01;
  assign sel_786403 = array_index_786214 == array_index_772918 ? add_786402 : sel_786399;
  assign add_786406 = sel_786403 + 8'h01;
  assign sel_786407 = array_index_786214 == array_index_772924 ? add_786406 : sel_786403;
  assign add_786410 = sel_786407 + 8'h01;
  assign sel_786411 = array_index_786214 == array_index_772930 ? add_786410 : sel_786407;
  assign add_786414 = sel_786411 + 8'h01;
  assign sel_786415 = array_index_786214 == array_index_772936 ? add_786414 : sel_786411;
  assign add_786418 = sel_786415 + 8'h01;
  assign sel_786419 = array_index_786214 == array_index_772942 ? add_786418 : sel_786415;
  assign add_786422 = sel_786419 + 8'h01;
  assign sel_786423 = array_index_786214 == array_index_772948 ? add_786422 : sel_786419;
  assign add_786426 = sel_786423 + 8'h01;
  assign sel_786427 = array_index_786214 == array_index_772954 ? add_786426 : sel_786423;
  assign add_786430 = sel_786427 + 8'h01;
  assign sel_786431 = array_index_786214 == array_index_772960 ? add_786430 : sel_786427;
  assign add_786434 = sel_786431 + 8'h01;
  assign sel_786435 = array_index_786214 == array_index_772966 ? add_786434 : sel_786431;
  assign add_786438 = sel_786435 + 8'h01;
  assign sel_786439 = array_index_786214 == array_index_772972 ? add_786438 : sel_786435;
  assign add_786442 = sel_786439 + 8'h01;
  assign sel_786443 = array_index_786214 == array_index_772978 ? add_786442 : sel_786439;
  assign add_786446 = sel_786443 + 8'h01;
  assign sel_786447 = array_index_786214 == array_index_772984 ? add_786446 : sel_786443;
  assign add_786450 = sel_786447 + 8'h01;
  assign sel_786451 = array_index_786214 == array_index_772990 ? add_786450 : sel_786447;
  assign add_786454 = sel_786451 + 8'h01;
  assign sel_786455 = array_index_786214 == array_index_772996 ? add_786454 : sel_786451;
  assign add_786458 = sel_786455 + 8'h01;
  assign sel_786459 = array_index_786214 == array_index_773002 ? add_786458 : sel_786455;
  assign add_786462 = sel_786459 + 8'h01;
  assign sel_786463 = array_index_786214 == array_index_773008 ? add_786462 : sel_786459;
  assign add_786466 = sel_786463 + 8'h01;
  assign sel_786467 = array_index_786214 == array_index_773014 ? add_786466 : sel_786463;
  assign add_786470 = sel_786467 + 8'h01;
  assign sel_786471 = array_index_786214 == array_index_773020 ? add_786470 : sel_786467;
  assign add_786474 = sel_786471 + 8'h01;
  assign sel_786475 = array_index_786214 == array_index_773026 ? add_786474 : sel_786471;
  assign add_786478 = sel_786475 + 8'h01;
  assign sel_786479 = array_index_786214 == array_index_773032 ? add_786478 : sel_786475;
  assign add_786482 = sel_786479 + 8'h01;
  assign sel_786483 = array_index_786214 == array_index_773038 ? add_786482 : sel_786479;
  assign add_786486 = sel_786483 + 8'h01;
  assign sel_786487 = array_index_786214 == array_index_773044 ? add_786486 : sel_786483;
  assign add_786490 = sel_786487 + 8'h01;
  assign sel_786491 = array_index_786214 == array_index_773050 ? add_786490 : sel_786487;
  assign add_786494 = sel_786491 + 8'h01;
  assign sel_786495 = array_index_786214 == array_index_773056 ? add_786494 : sel_786491;
  assign add_786498 = sel_786495 + 8'h01;
  assign sel_786499 = array_index_786214 == array_index_773062 ? add_786498 : sel_786495;
  assign add_786502 = sel_786499 + 8'h01;
  assign sel_786503 = array_index_786214 == array_index_773068 ? add_786502 : sel_786499;
  assign add_786506 = sel_786503 + 8'h01;
  assign sel_786507 = array_index_786214 == array_index_773074 ? add_786506 : sel_786503;
  assign add_786510 = sel_786507 + 8'h01;
  assign sel_786511 = array_index_786214 == array_index_773080 ? add_786510 : sel_786507;
  assign add_786514 = sel_786511 + 8'h01;
  assign sel_786515 = array_index_786214 == array_index_773086 ? add_786514 : sel_786511;
  assign add_786518 = sel_786515 + 8'h01;
  assign sel_786519 = array_index_786214 == array_index_773092 ? add_786518 : sel_786515;
  assign add_786522 = sel_786519 + 8'h01;
  assign sel_786523 = array_index_786214 == array_index_773098 ? add_786522 : sel_786519;
  assign add_786526 = sel_786523 + 8'h01;
  assign sel_786527 = array_index_786214 == array_index_773104 ? add_786526 : sel_786523;
  assign add_786530 = sel_786527 + 8'h01;
  assign sel_786531 = array_index_786214 == array_index_773110 ? add_786530 : sel_786527;
  assign add_786534 = sel_786531 + 8'h01;
  assign sel_786535 = array_index_786214 == array_index_773116 ? add_786534 : sel_786531;
  assign add_786538 = sel_786535 + 8'h01;
  assign sel_786539 = array_index_786214 == array_index_773122 ? add_786538 : sel_786535;
  assign add_786542 = sel_786539 + 8'h01;
  assign sel_786543 = array_index_786214 == array_index_773128 ? add_786542 : sel_786539;
  assign add_786546 = sel_786543 + 8'h01;
  assign sel_786547 = array_index_786214 == array_index_773134 ? add_786546 : sel_786543;
  assign add_786550 = sel_786547 + 8'h01;
  assign sel_786551 = array_index_786214 == array_index_773140 ? add_786550 : sel_786547;
  assign add_786554 = sel_786551 + 8'h01;
  assign sel_786555 = array_index_786214 == array_index_773146 ? add_786554 : sel_786551;
  assign add_786558 = sel_786555 + 8'h01;
  assign sel_786559 = array_index_786214 == array_index_773152 ? add_786558 : sel_786555;
  assign add_786562 = sel_786559 + 8'h01;
  assign sel_786563 = array_index_786214 == array_index_773158 ? add_786562 : sel_786559;
  assign add_786566 = sel_786563 + 8'h01;
  assign sel_786567 = array_index_786214 == array_index_773164 ? add_786566 : sel_786563;
  assign add_786570 = sel_786567 + 8'h01;
  assign sel_786571 = array_index_786214 == array_index_773170 ? add_786570 : sel_786567;
  assign add_786575 = sel_786571 + 8'h01;
  assign array_index_786576 = set1_unflattened[7'h26];
  assign sel_786577 = array_index_786214 == array_index_773176 ? add_786575 : sel_786571;
  assign add_786580 = sel_786577 + 8'h01;
  assign sel_786581 = array_index_786576 == array_index_772632 ? add_786580 : sel_786577;
  assign add_786584 = sel_786581 + 8'h01;
  assign sel_786585 = array_index_786576 == array_index_772636 ? add_786584 : sel_786581;
  assign add_786588 = sel_786585 + 8'h01;
  assign sel_786589 = array_index_786576 == array_index_772644 ? add_786588 : sel_786585;
  assign add_786592 = sel_786589 + 8'h01;
  assign sel_786593 = array_index_786576 == array_index_772652 ? add_786592 : sel_786589;
  assign add_786596 = sel_786593 + 8'h01;
  assign sel_786597 = array_index_786576 == array_index_772660 ? add_786596 : sel_786593;
  assign add_786600 = sel_786597 + 8'h01;
  assign sel_786601 = array_index_786576 == array_index_772668 ? add_786600 : sel_786597;
  assign add_786604 = sel_786601 + 8'h01;
  assign sel_786605 = array_index_786576 == array_index_772676 ? add_786604 : sel_786601;
  assign add_786608 = sel_786605 + 8'h01;
  assign sel_786609 = array_index_786576 == array_index_772684 ? add_786608 : sel_786605;
  assign add_786612 = sel_786609 + 8'h01;
  assign sel_786613 = array_index_786576 == array_index_772690 ? add_786612 : sel_786609;
  assign add_786616 = sel_786613 + 8'h01;
  assign sel_786617 = array_index_786576 == array_index_772696 ? add_786616 : sel_786613;
  assign add_786620 = sel_786617 + 8'h01;
  assign sel_786621 = array_index_786576 == array_index_772702 ? add_786620 : sel_786617;
  assign add_786624 = sel_786621 + 8'h01;
  assign sel_786625 = array_index_786576 == array_index_772708 ? add_786624 : sel_786621;
  assign add_786628 = sel_786625 + 8'h01;
  assign sel_786629 = array_index_786576 == array_index_772714 ? add_786628 : sel_786625;
  assign add_786632 = sel_786629 + 8'h01;
  assign sel_786633 = array_index_786576 == array_index_772720 ? add_786632 : sel_786629;
  assign add_786636 = sel_786633 + 8'h01;
  assign sel_786637 = array_index_786576 == array_index_772726 ? add_786636 : sel_786633;
  assign add_786640 = sel_786637 + 8'h01;
  assign sel_786641 = array_index_786576 == array_index_772732 ? add_786640 : sel_786637;
  assign add_786644 = sel_786641 + 8'h01;
  assign sel_786645 = array_index_786576 == array_index_772738 ? add_786644 : sel_786641;
  assign add_786648 = sel_786645 + 8'h01;
  assign sel_786649 = array_index_786576 == array_index_772744 ? add_786648 : sel_786645;
  assign add_786652 = sel_786649 + 8'h01;
  assign sel_786653 = array_index_786576 == array_index_772750 ? add_786652 : sel_786649;
  assign add_786656 = sel_786653 + 8'h01;
  assign sel_786657 = array_index_786576 == array_index_772756 ? add_786656 : sel_786653;
  assign add_786660 = sel_786657 + 8'h01;
  assign sel_786661 = array_index_786576 == array_index_772762 ? add_786660 : sel_786657;
  assign add_786664 = sel_786661 + 8'h01;
  assign sel_786665 = array_index_786576 == array_index_772768 ? add_786664 : sel_786661;
  assign add_786668 = sel_786665 + 8'h01;
  assign sel_786669 = array_index_786576 == array_index_772774 ? add_786668 : sel_786665;
  assign add_786672 = sel_786669 + 8'h01;
  assign sel_786673 = array_index_786576 == array_index_772780 ? add_786672 : sel_786669;
  assign add_786676 = sel_786673 + 8'h01;
  assign sel_786677 = array_index_786576 == array_index_772786 ? add_786676 : sel_786673;
  assign add_786680 = sel_786677 + 8'h01;
  assign sel_786681 = array_index_786576 == array_index_772792 ? add_786680 : sel_786677;
  assign add_786684 = sel_786681 + 8'h01;
  assign sel_786685 = array_index_786576 == array_index_772798 ? add_786684 : sel_786681;
  assign add_786688 = sel_786685 + 8'h01;
  assign sel_786689 = array_index_786576 == array_index_772804 ? add_786688 : sel_786685;
  assign add_786692 = sel_786689 + 8'h01;
  assign sel_786693 = array_index_786576 == array_index_772810 ? add_786692 : sel_786689;
  assign add_786696 = sel_786693 + 8'h01;
  assign sel_786697 = array_index_786576 == array_index_772816 ? add_786696 : sel_786693;
  assign add_786700 = sel_786697 + 8'h01;
  assign sel_786701 = array_index_786576 == array_index_772822 ? add_786700 : sel_786697;
  assign add_786704 = sel_786701 + 8'h01;
  assign sel_786705 = array_index_786576 == array_index_772828 ? add_786704 : sel_786701;
  assign add_786708 = sel_786705 + 8'h01;
  assign sel_786709 = array_index_786576 == array_index_772834 ? add_786708 : sel_786705;
  assign add_786712 = sel_786709 + 8'h01;
  assign sel_786713 = array_index_786576 == array_index_772840 ? add_786712 : sel_786709;
  assign add_786716 = sel_786713 + 8'h01;
  assign sel_786717 = array_index_786576 == array_index_772846 ? add_786716 : sel_786713;
  assign add_786720 = sel_786717 + 8'h01;
  assign sel_786721 = array_index_786576 == array_index_772852 ? add_786720 : sel_786717;
  assign add_786724 = sel_786721 + 8'h01;
  assign sel_786725 = array_index_786576 == array_index_772858 ? add_786724 : sel_786721;
  assign add_786728 = sel_786725 + 8'h01;
  assign sel_786729 = array_index_786576 == array_index_772864 ? add_786728 : sel_786725;
  assign add_786732 = sel_786729 + 8'h01;
  assign sel_786733 = array_index_786576 == array_index_772870 ? add_786732 : sel_786729;
  assign add_786736 = sel_786733 + 8'h01;
  assign sel_786737 = array_index_786576 == array_index_772876 ? add_786736 : sel_786733;
  assign add_786740 = sel_786737 + 8'h01;
  assign sel_786741 = array_index_786576 == array_index_772882 ? add_786740 : sel_786737;
  assign add_786744 = sel_786741 + 8'h01;
  assign sel_786745 = array_index_786576 == array_index_772888 ? add_786744 : sel_786741;
  assign add_786748 = sel_786745 + 8'h01;
  assign sel_786749 = array_index_786576 == array_index_772894 ? add_786748 : sel_786745;
  assign add_786752 = sel_786749 + 8'h01;
  assign sel_786753 = array_index_786576 == array_index_772900 ? add_786752 : sel_786749;
  assign add_786756 = sel_786753 + 8'h01;
  assign sel_786757 = array_index_786576 == array_index_772906 ? add_786756 : sel_786753;
  assign add_786760 = sel_786757 + 8'h01;
  assign sel_786761 = array_index_786576 == array_index_772912 ? add_786760 : sel_786757;
  assign add_786764 = sel_786761 + 8'h01;
  assign sel_786765 = array_index_786576 == array_index_772918 ? add_786764 : sel_786761;
  assign add_786768 = sel_786765 + 8'h01;
  assign sel_786769 = array_index_786576 == array_index_772924 ? add_786768 : sel_786765;
  assign add_786772 = sel_786769 + 8'h01;
  assign sel_786773 = array_index_786576 == array_index_772930 ? add_786772 : sel_786769;
  assign add_786776 = sel_786773 + 8'h01;
  assign sel_786777 = array_index_786576 == array_index_772936 ? add_786776 : sel_786773;
  assign add_786780 = sel_786777 + 8'h01;
  assign sel_786781 = array_index_786576 == array_index_772942 ? add_786780 : sel_786777;
  assign add_786784 = sel_786781 + 8'h01;
  assign sel_786785 = array_index_786576 == array_index_772948 ? add_786784 : sel_786781;
  assign add_786788 = sel_786785 + 8'h01;
  assign sel_786789 = array_index_786576 == array_index_772954 ? add_786788 : sel_786785;
  assign add_786792 = sel_786789 + 8'h01;
  assign sel_786793 = array_index_786576 == array_index_772960 ? add_786792 : sel_786789;
  assign add_786796 = sel_786793 + 8'h01;
  assign sel_786797 = array_index_786576 == array_index_772966 ? add_786796 : sel_786793;
  assign add_786800 = sel_786797 + 8'h01;
  assign sel_786801 = array_index_786576 == array_index_772972 ? add_786800 : sel_786797;
  assign add_786804 = sel_786801 + 8'h01;
  assign sel_786805 = array_index_786576 == array_index_772978 ? add_786804 : sel_786801;
  assign add_786808 = sel_786805 + 8'h01;
  assign sel_786809 = array_index_786576 == array_index_772984 ? add_786808 : sel_786805;
  assign add_786812 = sel_786809 + 8'h01;
  assign sel_786813 = array_index_786576 == array_index_772990 ? add_786812 : sel_786809;
  assign add_786816 = sel_786813 + 8'h01;
  assign sel_786817 = array_index_786576 == array_index_772996 ? add_786816 : sel_786813;
  assign add_786820 = sel_786817 + 8'h01;
  assign sel_786821 = array_index_786576 == array_index_773002 ? add_786820 : sel_786817;
  assign add_786824 = sel_786821 + 8'h01;
  assign sel_786825 = array_index_786576 == array_index_773008 ? add_786824 : sel_786821;
  assign add_786828 = sel_786825 + 8'h01;
  assign sel_786829 = array_index_786576 == array_index_773014 ? add_786828 : sel_786825;
  assign add_786832 = sel_786829 + 8'h01;
  assign sel_786833 = array_index_786576 == array_index_773020 ? add_786832 : sel_786829;
  assign add_786836 = sel_786833 + 8'h01;
  assign sel_786837 = array_index_786576 == array_index_773026 ? add_786836 : sel_786833;
  assign add_786840 = sel_786837 + 8'h01;
  assign sel_786841 = array_index_786576 == array_index_773032 ? add_786840 : sel_786837;
  assign add_786844 = sel_786841 + 8'h01;
  assign sel_786845 = array_index_786576 == array_index_773038 ? add_786844 : sel_786841;
  assign add_786848 = sel_786845 + 8'h01;
  assign sel_786849 = array_index_786576 == array_index_773044 ? add_786848 : sel_786845;
  assign add_786852 = sel_786849 + 8'h01;
  assign sel_786853 = array_index_786576 == array_index_773050 ? add_786852 : sel_786849;
  assign add_786856 = sel_786853 + 8'h01;
  assign sel_786857 = array_index_786576 == array_index_773056 ? add_786856 : sel_786853;
  assign add_786860 = sel_786857 + 8'h01;
  assign sel_786861 = array_index_786576 == array_index_773062 ? add_786860 : sel_786857;
  assign add_786864 = sel_786861 + 8'h01;
  assign sel_786865 = array_index_786576 == array_index_773068 ? add_786864 : sel_786861;
  assign add_786868 = sel_786865 + 8'h01;
  assign sel_786869 = array_index_786576 == array_index_773074 ? add_786868 : sel_786865;
  assign add_786872 = sel_786869 + 8'h01;
  assign sel_786873 = array_index_786576 == array_index_773080 ? add_786872 : sel_786869;
  assign add_786876 = sel_786873 + 8'h01;
  assign sel_786877 = array_index_786576 == array_index_773086 ? add_786876 : sel_786873;
  assign add_786880 = sel_786877 + 8'h01;
  assign sel_786881 = array_index_786576 == array_index_773092 ? add_786880 : sel_786877;
  assign add_786884 = sel_786881 + 8'h01;
  assign sel_786885 = array_index_786576 == array_index_773098 ? add_786884 : sel_786881;
  assign add_786888 = sel_786885 + 8'h01;
  assign sel_786889 = array_index_786576 == array_index_773104 ? add_786888 : sel_786885;
  assign add_786892 = sel_786889 + 8'h01;
  assign sel_786893 = array_index_786576 == array_index_773110 ? add_786892 : sel_786889;
  assign add_786896 = sel_786893 + 8'h01;
  assign sel_786897 = array_index_786576 == array_index_773116 ? add_786896 : sel_786893;
  assign add_786900 = sel_786897 + 8'h01;
  assign sel_786901 = array_index_786576 == array_index_773122 ? add_786900 : sel_786897;
  assign add_786904 = sel_786901 + 8'h01;
  assign sel_786905 = array_index_786576 == array_index_773128 ? add_786904 : sel_786901;
  assign add_786908 = sel_786905 + 8'h01;
  assign sel_786909 = array_index_786576 == array_index_773134 ? add_786908 : sel_786905;
  assign add_786912 = sel_786909 + 8'h01;
  assign sel_786913 = array_index_786576 == array_index_773140 ? add_786912 : sel_786909;
  assign add_786916 = sel_786913 + 8'h01;
  assign sel_786917 = array_index_786576 == array_index_773146 ? add_786916 : sel_786913;
  assign add_786920 = sel_786917 + 8'h01;
  assign sel_786921 = array_index_786576 == array_index_773152 ? add_786920 : sel_786917;
  assign add_786924 = sel_786921 + 8'h01;
  assign sel_786925 = array_index_786576 == array_index_773158 ? add_786924 : sel_786921;
  assign add_786928 = sel_786925 + 8'h01;
  assign sel_786929 = array_index_786576 == array_index_773164 ? add_786928 : sel_786925;
  assign add_786932 = sel_786929 + 8'h01;
  assign sel_786933 = array_index_786576 == array_index_773170 ? add_786932 : sel_786929;
  assign add_786937 = sel_786933 + 8'h01;
  assign array_index_786938 = set1_unflattened[7'h27];
  assign sel_786939 = array_index_786576 == array_index_773176 ? add_786937 : sel_786933;
  assign add_786942 = sel_786939 + 8'h01;
  assign sel_786943 = array_index_786938 == array_index_772632 ? add_786942 : sel_786939;
  assign add_786946 = sel_786943 + 8'h01;
  assign sel_786947 = array_index_786938 == array_index_772636 ? add_786946 : sel_786943;
  assign add_786950 = sel_786947 + 8'h01;
  assign sel_786951 = array_index_786938 == array_index_772644 ? add_786950 : sel_786947;
  assign add_786954 = sel_786951 + 8'h01;
  assign sel_786955 = array_index_786938 == array_index_772652 ? add_786954 : sel_786951;
  assign add_786958 = sel_786955 + 8'h01;
  assign sel_786959 = array_index_786938 == array_index_772660 ? add_786958 : sel_786955;
  assign add_786962 = sel_786959 + 8'h01;
  assign sel_786963 = array_index_786938 == array_index_772668 ? add_786962 : sel_786959;
  assign add_786966 = sel_786963 + 8'h01;
  assign sel_786967 = array_index_786938 == array_index_772676 ? add_786966 : sel_786963;
  assign add_786970 = sel_786967 + 8'h01;
  assign sel_786971 = array_index_786938 == array_index_772684 ? add_786970 : sel_786967;
  assign add_786974 = sel_786971 + 8'h01;
  assign sel_786975 = array_index_786938 == array_index_772690 ? add_786974 : sel_786971;
  assign add_786978 = sel_786975 + 8'h01;
  assign sel_786979 = array_index_786938 == array_index_772696 ? add_786978 : sel_786975;
  assign add_786982 = sel_786979 + 8'h01;
  assign sel_786983 = array_index_786938 == array_index_772702 ? add_786982 : sel_786979;
  assign add_786986 = sel_786983 + 8'h01;
  assign sel_786987 = array_index_786938 == array_index_772708 ? add_786986 : sel_786983;
  assign add_786990 = sel_786987 + 8'h01;
  assign sel_786991 = array_index_786938 == array_index_772714 ? add_786990 : sel_786987;
  assign add_786994 = sel_786991 + 8'h01;
  assign sel_786995 = array_index_786938 == array_index_772720 ? add_786994 : sel_786991;
  assign add_786998 = sel_786995 + 8'h01;
  assign sel_786999 = array_index_786938 == array_index_772726 ? add_786998 : sel_786995;
  assign add_787002 = sel_786999 + 8'h01;
  assign sel_787003 = array_index_786938 == array_index_772732 ? add_787002 : sel_786999;
  assign add_787006 = sel_787003 + 8'h01;
  assign sel_787007 = array_index_786938 == array_index_772738 ? add_787006 : sel_787003;
  assign add_787010 = sel_787007 + 8'h01;
  assign sel_787011 = array_index_786938 == array_index_772744 ? add_787010 : sel_787007;
  assign add_787014 = sel_787011 + 8'h01;
  assign sel_787015 = array_index_786938 == array_index_772750 ? add_787014 : sel_787011;
  assign add_787018 = sel_787015 + 8'h01;
  assign sel_787019 = array_index_786938 == array_index_772756 ? add_787018 : sel_787015;
  assign add_787022 = sel_787019 + 8'h01;
  assign sel_787023 = array_index_786938 == array_index_772762 ? add_787022 : sel_787019;
  assign add_787026 = sel_787023 + 8'h01;
  assign sel_787027 = array_index_786938 == array_index_772768 ? add_787026 : sel_787023;
  assign add_787030 = sel_787027 + 8'h01;
  assign sel_787031 = array_index_786938 == array_index_772774 ? add_787030 : sel_787027;
  assign add_787034 = sel_787031 + 8'h01;
  assign sel_787035 = array_index_786938 == array_index_772780 ? add_787034 : sel_787031;
  assign add_787038 = sel_787035 + 8'h01;
  assign sel_787039 = array_index_786938 == array_index_772786 ? add_787038 : sel_787035;
  assign add_787042 = sel_787039 + 8'h01;
  assign sel_787043 = array_index_786938 == array_index_772792 ? add_787042 : sel_787039;
  assign add_787046 = sel_787043 + 8'h01;
  assign sel_787047 = array_index_786938 == array_index_772798 ? add_787046 : sel_787043;
  assign add_787050 = sel_787047 + 8'h01;
  assign sel_787051 = array_index_786938 == array_index_772804 ? add_787050 : sel_787047;
  assign add_787054 = sel_787051 + 8'h01;
  assign sel_787055 = array_index_786938 == array_index_772810 ? add_787054 : sel_787051;
  assign add_787058 = sel_787055 + 8'h01;
  assign sel_787059 = array_index_786938 == array_index_772816 ? add_787058 : sel_787055;
  assign add_787062 = sel_787059 + 8'h01;
  assign sel_787063 = array_index_786938 == array_index_772822 ? add_787062 : sel_787059;
  assign add_787066 = sel_787063 + 8'h01;
  assign sel_787067 = array_index_786938 == array_index_772828 ? add_787066 : sel_787063;
  assign add_787070 = sel_787067 + 8'h01;
  assign sel_787071 = array_index_786938 == array_index_772834 ? add_787070 : sel_787067;
  assign add_787074 = sel_787071 + 8'h01;
  assign sel_787075 = array_index_786938 == array_index_772840 ? add_787074 : sel_787071;
  assign add_787078 = sel_787075 + 8'h01;
  assign sel_787079 = array_index_786938 == array_index_772846 ? add_787078 : sel_787075;
  assign add_787082 = sel_787079 + 8'h01;
  assign sel_787083 = array_index_786938 == array_index_772852 ? add_787082 : sel_787079;
  assign add_787086 = sel_787083 + 8'h01;
  assign sel_787087 = array_index_786938 == array_index_772858 ? add_787086 : sel_787083;
  assign add_787090 = sel_787087 + 8'h01;
  assign sel_787091 = array_index_786938 == array_index_772864 ? add_787090 : sel_787087;
  assign add_787094 = sel_787091 + 8'h01;
  assign sel_787095 = array_index_786938 == array_index_772870 ? add_787094 : sel_787091;
  assign add_787098 = sel_787095 + 8'h01;
  assign sel_787099 = array_index_786938 == array_index_772876 ? add_787098 : sel_787095;
  assign add_787102 = sel_787099 + 8'h01;
  assign sel_787103 = array_index_786938 == array_index_772882 ? add_787102 : sel_787099;
  assign add_787106 = sel_787103 + 8'h01;
  assign sel_787107 = array_index_786938 == array_index_772888 ? add_787106 : sel_787103;
  assign add_787110 = sel_787107 + 8'h01;
  assign sel_787111 = array_index_786938 == array_index_772894 ? add_787110 : sel_787107;
  assign add_787114 = sel_787111 + 8'h01;
  assign sel_787115 = array_index_786938 == array_index_772900 ? add_787114 : sel_787111;
  assign add_787118 = sel_787115 + 8'h01;
  assign sel_787119 = array_index_786938 == array_index_772906 ? add_787118 : sel_787115;
  assign add_787122 = sel_787119 + 8'h01;
  assign sel_787123 = array_index_786938 == array_index_772912 ? add_787122 : sel_787119;
  assign add_787126 = sel_787123 + 8'h01;
  assign sel_787127 = array_index_786938 == array_index_772918 ? add_787126 : sel_787123;
  assign add_787130 = sel_787127 + 8'h01;
  assign sel_787131 = array_index_786938 == array_index_772924 ? add_787130 : sel_787127;
  assign add_787134 = sel_787131 + 8'h01;
  assign sel_787135 = array_index_786938 == array_index_772930 ? add_787134 : sel_787131;
  assign add_787138 = sel_787135 + 8'h01;
  assign sel_787139 = array_index_786938 == array_index_772936 ? add_787138 : sel_787135;
  assign add_787142 = sel_787139 + 8'h01;
  assign sel_787143 = array_index_786938 == array_index_772942 ? add_787142 : sel_787139;
  assign add_787146 = sel_787143 + 8'h01;
  assign sel_787147 = array_index_786938 == array_index_772948 ? add_787146 : sel_787143;
  assign add_787150 = sel_787147 + 8'h01;
  assign sel_787151 = array_index_786938 == array_index_772954 ? add_787150 : sel_787147;
  assign add_787154 = sel_787151 + 8'h01;
  assign sel_787155 = array_index_786938 == array_index_772960 ? add_787154 : sel_787151;
  assign add_787158 = sel_787155 + 8'h01;
  assign sel_787159 = array_index_786938 == array_index_772966 ? add_787158 : sel_787155;
  assign add_787162 = sel_787159 + 8'h01;
  assign sel_787163 = array_index_786938 == array_index_772972 ? add_787162 : sel_787159;
  assign add_787166 = sel_787163 + 8'h01;
  assign sel_787167 = array_index_786938 == array_index_772978 ? add_787166 : sel_787163;
  assign add_787170 = sel_787167 + 8'h01;
  assign sel_787171 = array_index_786938 == array_index_772984 ? add_787170 : sel_787167;
  assign add_787174 = sel_787171 + 8'h01;
  assign sel_787175 = array_index_786938 == array_index_772990 ? add_787174 : sel_787171;
  assign add_787178 = sel_787175 + 8'h01;
  assign sel_787179 = array_index_786938 == array_index_772996 ? add_787178 : sel_787175;
  assign add_787182 = sel_787179 + 8'h01;
  assign sel_787183 = array_index_786938 == array_index_773002 ? add_787182 : sel_787179;
  assign add_787186 = sel_787183 + 8'h01;
  assign sel_787187 = array_index_786938 == array_index_773008 ? add_787186 : sel_787183;
  assign add_787190 = sel_787187 + 8'h01;
  assign sel_787191 = array_index_786938 == array_index_773014 ? add_787190 : sel_787187;
  assign add_787194 = sel_787191 + 8'h01;
  assign sel_787195 = array_index_786938 == array_index_773020 ? add_787194 : sel_787191;
  assign add_787198 = sel_787195 + 8'h01;
  assign sel_787199 = array_index_786938 == array_index_773026 ? add_787198 : sel_787195;
  assign add_787202 = sel_787199 + 8'h01;
  assign sel_787203 = array_index_786938 == array_index_773032 ? add_787202 : sel_787199;
  assign add_787206 = sel_787203 + 8'h01;
  assign sel_787207 = array_index_786938 == array_index_773038 ? add_787206 : sel_787203;
  assign add_787210 = sel_787207 + 8'h01;
  assign sel_787211 = array_index_786938 == array_index_773044 ? add_787210 : sel_787207;
  assign add_787214 = sel_787211 + 8'h01;
  assign sel_787215 = array_index_786938 == array_index_773050 ? add_787214 : sel_787211;
  assign add_787218 = sel_787215 + 8'h01;
  assign sel_787219 = array_index_786938 == array_index_773056 ? add_787218 : sel_787215;
  assign add_787222 = sel_787219 + 8'h01;
  assign sel_787223 = array_index_786938 == array_index_773062 ? add_787222 : sel_787219;
  assign add_787226 = sel_787223 + 8'h01;
  assign sel_787227 = array_index_786938 == array_index_773068 ? add_787226 : sel_787223;
  assign add_787230 = sel_787227 + 8'h01;
  assign sel_787231 = array_index_786938 == array_index_773074 ? add_787230 : sel_787227;
  assign add_787234 = sel_787231 + 8'h01;
  assign sel_787235 = array_index_786938 == array_index_773080 ? add_787234 : sel_787231;
  assign add_787238 = sel_787235 + 8'h01;
  assign sel_787239 = array_index_786938 == array_index_773086 ? add_787238 : sel_787235;
  assign add_787242 = sel_787239 + 8'h01;
  assign sel_787243 = array_index_786938 == array_index_773092 ? add_787242 : sel_787239;
  assign add_787246 = sel_787243 + 8'h01;
  assign sel_787247 = array_index_786938 == array_index_773098 ? add_787246 : sel_787243;
  assign add_787250 = sel_787247 + 8'h01;
  assign sel_787251 = array_index_786938 == array_index_773104 ? add_787250 : sel_787247;
  assign add_787254 = sel_787251 + 8'h01;
  assign sel_787255 = array_index_786938 == array_index_773110 ? add_787254 : sel_787251;
  assign add_787258 = sel_787255 + 8'h01;
  assign sel_787259 = array_index_786938 == array_index_773116 ? add_787258 : sel_787255;
  assign add_787262 = sel_787259 + 8'h01;
  assign sel_787263 = array_index_786938 == array_index_773122 ? add_787262 : sel_787259;
  assign add_787266 = sel_787263 + 8'h01;
  assign sel_787267 = array_index_786938 == array_index_773128 ? add_787266 : sel_787263;
  assign add_787270 = sel_787267 + 8'h01;
  assign sel_787271 = array_index_786938 == array_index_773134 ? add_787270 : sel_787267;
  assign add_787274 = sel_787271 + 8'h01;
  assign sel_787275 = array_index_786938 == array_index_773140 ? add_787274 : sel_787271;
  assign add_787278 = sel_787275 + 8'h01;
  assign sel_787279 = array_index_786938 == array_index_773146 ? add_787278 : sel_787275;
  assign add_787282 = sel_787279 + 8'h01;
  assign sel_787283 = array_index_786938 == array_index_773152 ? add_787282 : sel_787279;
  assign add_787286 = sel_787283 + 8'h01;
  assign sel_787287 = array_index_786938 == array_index_773158 ? add_787286 : sel_787283;
  assign add_787290 = sel_787287 + 8'h01;
  assign sel_787291 = array_index_786938 == array_index_773164 ? add_787290 : sel_787287;
  assign add_787294 = sel_787291 + 8'h01;
  assign sel_787295 = array_index_786938 == array_index_773170 ? add_787294 : sel_787291;
  assign add_787299 = sel_787295 + 8'h01;
  assign array_index_787300 = set1_unflattened[7'h28];
  assign sel_787301 = array_index_786938 == array_index_773176 ? add_787299 : sel_787295;
  assign add_787304 = sel_787301 + 8'h01;
  assign sel_787305 = array_index_787300 == array_index_772632 ? add_787304 : sel_787301;
  assign add_787308 = sel_787305 + 8'h01;
  assign sel_787309 = array_index_787300 == array_index_772636 ? add_787308 : sel_787305;
  assign add_787312 = sel_787309 + 8'h01;
  assign sel_787313 = array_index_787300 == array_index_772644 ? add_787312 : sel_787309;
  assign add_787316 = sel_787313 + 8'h01;
  assign sel_787317 = array_index_787300 == array_index_772652 ? add_787316 : sel_787313;
  assign add_787320 = sel_787317 + 8'h01;
  assign sel_787321 = array_index_787300 == array_index_772660 ? add_787320 : sel_787317;
  assign add_787324 = sel_787321 + 8'h01;
  assign sel_787325 = array_index_787300 == array_index_772668 ? add_787324 : sel_787321;
  assign add_787328 = sel_787325 + 8'h01;
  assign sel_787329 = array_index_787300 == array_index_772676 ? add_787328 : sel_787325;
  assign add_787332 = sel_787329 + 8'h01;
  assign sel_787333 = array_index_787300 == array_index_772684 ? add_787332 : sel_787329;
  assign add_787336 = sel_787333 + 8'h01;
  assign sel_787337 = array_index_787300 == array_index_772690 ? add_787336 : sel_787333;
  assign add_787340 = sel_787337 + 8'h01;
  assign sel_787341 = array_index_787300 == array_index_772696 ? add_787340 : sel_787337;
  assign add_787344 = sel_787341 + 8'h01;
  assign sel_787345 = array_index_787300 == array_index_772702 ? add_787344 : sel_787341;
  assign add_787348 = sel_787345 + 8'h01;
  assign sel_787349 = array_index_787300 == array_index_772708 ? add_787348 : sel_787345;
  assign add_787352 = sel_787349 + 8'h01;
  assign sel_787353 = array_index_787300 == array_index_772714 ? add_787352 : sel_787349;
  assign add_787356 = sel_787353 + 8'h01;
  assign sel_787357 = array_index_787300 == array_index_772720 ? add_787356 : sel_787353;
  assign add_787360 = sel_787357 + 8'h01;
  assign sel_787361 = array_index_787300 == array_index_772726 ? add_787360 : sel_787357;
  assign add_787364 = sel_787361 + 8'h01;
  assign sel_787365 = array_index_787300 == array_index_772732 ? add_787364 : sel_787361;
  assign add_787368 = sel_787365 + 8'h01;
  assign sel_787369 = array_index_787300 == array_index_772738 ? add_787368 : sel_787365;
  assign add_787372 = sel_787369 + 8'h01;
  assign sel_787373 = array_index_787300 == array_index_772744 ? add_787372 : sel_787369;
  assign add_787376 = sel_787373 + 8'h01;
  assign sel_787377 = array_index_787300 == array_index_772750 ? add_787376 : sel_787373;
  assign add_787380 = sel_787377 + 8'h01;
  assign sel_787381 = array_index_787300 == array_index_772756 ? add_787380 : sel_787377;
  assign add_787384 = sel_787381 + 8'h01;
  assign sel_787385 = array_index_787300 == array_index_772762 ? add_787384 : sel_787381;
  assign add_787388 = sel_787385 + 8'h01;
  assign sel_787389 = array_index_787300 == array_index_772768 ? add_787388 : sel_787385;
  assign add_787392 = sel_787389 + 8'h01;
  assign sel_787393 = array_index_787300 == array_index_772774 ? add_787392 : sel_787389;
  assign add_787396 = sel_787393 + 8'h01;
  assign sel_787397 = array_index_787300 == array_index_772780 ? add_787396 : sel_787393;
  assign add_787400 = sel_787397 + 8'h01;
  assign sel_787401 = array_index_787300 == array_index_772786 ? add_787400 : sel_787397;
  assign add_787404 = sel_787401 + 8'h01;
  assign sel_787405 = array_index_787300 == array_index_772792 ? add_787404 : sel_787401;
  assign add_787408 = sel_787405 + 8'h01;
  assign sel_787409 = array_index_787300 == array_index_772798 ? add_787408 : sel_787405;
  assign add_787412 = sel_787409 + 8'h01;
  assign sel_787413 = array_index_787300 == array_index_772804 ? add_787412 : sel_787409;
  assign add_787416 = sel_787413 + 8'h01;
  assign sel_787417 = array_index_787300 == array_index_772810 ? add_787416 : sel_787413;
  assign add_787420 = sel_787417 + 8'h01;
  assign sel_787421 = array_index_787300 == array_index_772816 ? add_787420 : sel_787417;
  assign add_787424 = sel_787421 + 8'h01;
  assign sel_787425 = array_index_787300 == array_index_772822 ? add_787424 : sel_787421;
  assign add_787428 = sel_787425 + 8'h01;
  assign sel_787429 = array_index_787300 == array_index_772828 ? add_787428 : sel_787425;
  assign add_787432 = sel_787429 + 8'h01;
  assign sel_787433 = array_index_787300 == array_index_772834 ? add_787432 : sel_787429;
  assign add_787436 = sel_787433 + 8'h01;
  assign sel_787437 = array_index_787300 == array_index_772840 ? add_787436 : sel_787433;
  assign add_787440 = sel_787437 + 8'h01;
  assign sel_787441 = array_index_787300 == array_index_772846 ? add_787440 : sel_787437;
  assign add_787444 = sel_787441 + 8'h01;
  assign sel_787445 = array_index_787300 == array_index_772852 ? add_787444 : sel_787441;
  assign add_787448 = sel_787445 + 8'h01;
  assign sel_787449 = array_index_787300 == array_index_772858 ? add_787448 : sel_787445;
  assign add_787452 = sel_787449 + 8'h01;
  assign sel_787453 = array_index_787300 == array_index_772864 ? add_787452 : sel_787449;
  assign add_787456 = sel_787453 + 8'h01;
  assign sel_787457 = array_index_787300 == array_index_772870 ? add_787456 : sel_787453;
  assign add_787460 = sel_787457 + 8'h01;
  assign sel_787461 = array_index_787300 == array_index_772876 ? add_787460 : sel_787457;
  assign add_787464 = sel_787461 + 8'h01;
  assign sel_787465 = array_index_787300 == array_index_772882 ? add_787464 : sel_787461;
  assign add_787468 = sel_787465 + 8'h01;
  assign sel_787469 = array_index_787300 == array_index_772888 ? add_787468 : sel_787465;
  assign add_787472 = sel_787469 + 8'h01;
  assign sel_787473 = array_index_787300 == array_index_772894 ? add_787472 : sel_787469;
  assign add_787476 = sel_787473 + 8'h01;
  assign sel_787477 = array_index_787300 == array_index_772900 ? add_787476 : sel_787473;
  assign add_787480 = sel_787477 + 8'h01;
  assign sel_787481 = array_index_787300 == array_index_772906 ? add_787480 : sel_787477;
  assign add_787484 = sel_787481 + 8'h01;
  assign sel_787485 = array_index_787300 == array_index_772912 ? add_787484 : sel_787481;
  assign add_787488 = sel_787485 + 8'h01;
  assign sel_787489 = array_index_787300 == array_index_772918 ? add_787488 : sel_787485;
  assign add_787492 = sel_787489 + 8'h01;
  assign sel_787493 = array_index_787300 == array_index_772924 ? add_787492 : sel_787489;
  assign add_787496 = sel_787493 + 8'h01;
  assign sel_787497 = array_index_787300 == array_index_772930 ? add_787496 : sel_787493;
  assign add_787500 = sel_787497 + 8'h01;
  assign sel_787501 = array_index_787300 == array_index_772936 ? add_787500 : sel_787497;
  assign add_787504 = sel_787501 + 8'h01;
  assign sel_787505 = array_index_787300 == array_index_772942 ? add_787504 : sel_787501;
  assign add_787508 = sel_787505 + 8'h01;
  assign sel_787509 = array_index_787300 == array_index_772948 ? add_787508 : sel_787505;
  assign add_787512 = sel_787509 + 8'h01;
  assign sel_787513 = array_index_787300 == array_index_772954 ? add_787512 : sel_787509;
  assign add_787516 = sel_787513 + 8'h01;
  assign sel_787517 = array_index_787300 == array_index_772960 ? add_787516 : sel_787513;
  assign add_787520 = sel_787517 + 8'h01;
  assign sel_787521 = array_index_787300 == array_index_772966 ? add_787520 : sel_787517;
  assign add_787524 = sel_787521 + 8'h01;
  assign sel_787525 = array_index_787300 == array_index_772972 ? add_787524 : sel_787521;
  assign add_787528 = sel_787525 + 8'h01;
  assign sel_787529 = array_index_787300 == array_index_772978 ? add_787528 : sel_787525;
  assign add_787532 = sel_787529 + 8'h01;
  assign sel_787533 = array_index_787300 == array_index_772984 ? add_787532 : sel_787529;
  assign add_787536 = sel_787533 + 8'h01;
  assign sel_787537 = array_index_787300 == array_index_772990 ? add_787536 : sel_787533;
  assign add_787540 = sel_787537 + 8'h01;
  assign sel_787541 = array_index_787300 == array_index_772996 ? add_787540 : sel_787537;
  assign add_787544 = sel_787541 + 8'h01;
  assign sel_787545 = array_index_787300 == array_index_773002 ? add_787544 : sel_787541;
  assign add_787548 = sel_787545 + 8'h01;
  assign sel_787549 = array_index_787300 == array_index_773008 ? add_787548 : sel_787545;
  assign add_787552 = sel_787549 + 8'h01;
  assign sel_787553 = array_index_787300 == array_index_773014 ? add_787552 : sel_787549;
  assign add_787556 = sel_787553 + 8'h01;
  assign sel_787557 = array_index_787300 == array_index_773020 ? add_787556 : sel_787553;
  assign add_787560 = sel_787557 + 8'h01;
  assign sel_787561 = array_index_787300 == array_index_773026 ? add_787560 : sel_787557;
  assign add_787564 = sel_787561 + 8'h01;
  assign sel_787565 = array_index_787300 == array_index_773032 ? add_787564 : sel_787561;
  assign add_787568 = sel_787565 + 8'h01;
  assign sel_787569 = array_index_787300 == array_index_773038 ? add_787568 : sel_787565;
  assign add_787572 = sel_787569 + 8'h01;
  assign sel_787573 = array_index_787300 == array_index_773044 ? add_787572 : sel_787569;
  assign add_787576 = sel_787573 + 8'h01;
  assign sel_787577 = array_index_787300 == array_index_773050 ? add_787576 : sel_787573;
  assign add_787580 = sel_787577 + 8'h01;
  assign sel_787581 = array_index_787300 == array_index_773056 ? add_787580 : sel_787577;
  assign add_787584 = sel_787581 + 8'h01;
  assign sel_787585 = array_index_787300 == array_index_773062 ? add_787584 : sel_787581;
  assign add_787588 = sel_787585 + 8'h01;
  assign sel_787589 = array_index_787300 == array_index_773068 ? add_787588 : sel_787585;
  assign add_787592 = sel_787589 + 8'h01;
  assign sel_787593 = array_index_787300 == array_index_773074 ? add_787592 : sel_787589;
  assign add_787596 = sel_787593 + 8'h01;
  assign sel_787597 = array_index_787300 == array_index_773080 ? add_787596 : sel_787593;
  assign add_787600 = sel_787597 + 8'h01;
  assign sel_787601 = array_index_787300 == array_index_773086 ? add_787600 : sel_787597;
  assign add_787604 = sel_787601 + 8'h01;
  assign sel_787605 = array_index_787300 == array_index_773092 ? add_787604 : sel_787601;
  assign add_787608 = sel_787605 + 8'h01;
  assign sel_787609 = array_index_787300 == array_index_773098 ? add_787608 : sel_787605;
  assign add_787612 = sel_787609 + 8'h01;
  assign sel_787613 = array_index_787300 == array_index_773104 ? add_787612 : sel_787609;
  assign add_787616 = sel_787613 + 8'h01;
  assign sel_787617 = array_index_787300 == array_index_773110 ? add_787616 : sel_787613;
  assign add_787620 = sel_787617 + 8'h01;
  assign sel_787621 = array_index_787300 == array_index_773116 ? add_787620 : sel_787617;
  assign add_787624 = sel_787621 + 8'h01;
  assign sel_787625 = array_index_787300 == array_index_773122 ? add_787624 : sel_787621;
  assign add_787628 = sel_787625 + 8'h01;
  assign sel_787629 = array_index_787300 == array_index_773128 ? add_787628 : sel_787625;
  assign add_787632 = sel_787629 + 8'h01;
  assign sel_787633 = array_index_787300 == array_index_773134 ? add_787632 : sel_787629;
  assign add_787636 = sel_787633 + 8'h01;
  assign sel_787637 = array_index_787300 == array_index_773140 ? add_787636 : sel_787633;
  assign add_787640 = sel_787637 + 8'h01;
  assign sel_787641 = array_index_787300 == array_index_773146 ? add_787640 : sel_787637;
  assign add_787644 = sel_787641 + 8'h01;
  assign sel_787645 = array_index_787300 == array_index_773152 ? add_787644 : sel_787641;
  assign add_787648 = sel_787645 + 8'h01;
  assign sel_787649 = array_index_787300 == array_index_773158 ? add_787648 : sel_787645;
  assign add_787652 = sel_787649 + 8'h01;
  assign sel_787653 = array_index_787300 == array_index_773164 ? add_787652 : sel_787649;
  assign add_787656 = sel_787653 + 8'h01;
  assign sel_787657 = array_index_787300 == array_index_773170 ? add_787656 : sel_787653;
  assign add_787661 = sel_787657 + 8'h01;
  assign array_index_787662 = set1_unflattened[7'h29];
  assign sel_787663 = array_index_787300 == array_index_773176 ? add_787661 : sel_787657;
  assign add_787666 = sel_787663 + 8'h01;
  assign sel_787667 = array_index_787662 == array_index_772632 ? add_787666 : sel_787663;
  assign add_787670 = sel_787667 + 8'h01;
  assign sel_787671 = array_index_787662 == array_index_772636 ? add_787670 : sel_787667;
  assign add_787674 = sel_787671 + 8'h01;
  assign sel_787675 = array_index_787662 == array_index_772644 ? add_787674 : sel_787671;
  assign add_787678 = sel_787675 + 8'h01;
  assign sel_787679 = array_index_787662 == array_index_772652 ? add_787678 : sel_787675;
  assign add_787682 = sel_787679 + 8'h01;
  assign sel_787683 = array_index_787662 == array_index_772660 ? add_787682 : sel_787679;
  assign add_787686 = sel_787683 + 8'h01;
  assign sel_787687 = array_index_787662 == array_index_772668 ? add_787686 : sel_787683;
  assign add_787690 = sel_787687 + 8'h01;
  assign sel_787691 = array_index_787662 == array_index_772676 ? add_787690 : sel_787687;
  assign add_787694 = sel_787691 + 8'h01;
  assign sel_787695 = array_index_787662 == array_index_772684 ? add_787694 : sel_787691;
  assign add_787698 = sel_787695 + 8'h01;
  assign sel_787699 = array_index_787662 == array_index_772690 ? add_787698 : sel_787695;
  assign add_787702 = sel_787699 + 8'h01;
  assign sel_787703 = array_index_787662 == array_index_772696 ? add_787702 : sel_787699;
  assign add_787706 = sel_787703 + 8'h01;
  assign sel_787707 = array_index_787662 == array_index_772702 ? add_787706 : sel_787703;
  assign add_787710 = sel_787707 + 8'h01;
  assign sel_787711 = array_index_787662 == array_index_772708 ? add_787710 : sel_787707;
  assign add_787714 = sel_787711 + 8'h01;
  assign sel_787715 = array_index_787662 == array_index_772714 ? add_787714 : sel_787711;
  assign add_787718 = sel_787715 + 8'h01;
  assign sel_787719 = array_index_787662 == array_index_772720 ? add_787718 : sel_787715;
  assign add_787722 = sel_787719 + 8'h01;
  assign sel_787723 = array_index_787662 == array_index_772726 ? add_787722 : sel_787719;
  assign add_787726 = sel_787723 + 8'h01;
  assign sel_787727 = array_index_787662 == array_index_772732 ? add_787726 : sel_787723;
  assign add_787730 = sel_787727 + 8'h01;
  assign sel_787731 = array_index_787662 == array_index_772738 ? add_787730 : sel_787727;
  assign add_787734 = sel_787731 + 8'h01;
  assign sel_787735 = array_index_787662 == array_index_772744 ? add_787734 : sel_787731;
  assign add_787738 = sel_787735 + 8'h01;
  assign sel_787739 = array_index_787662 == array_index_772750 ? add_787738 : sel_787735;
  assign add_787742 = sel_787739 + 8'h01;
  assign sel_787743 = array_index_787662 == array_index_772756 ? add_787742 : sel_787739;
  assign add_787746 = sel_787743 + 8'h01;
  assign sel_787747 = array_index_787662 == array_index_772762 ? add_787746 : sel_787743;
  assign add_787750 = sel_787747 + 8'h01;
  assign sel_787751 = array_index_787662 == array_index_772768 ? add_787750 : sel_787747;
  assign add_787754 = sel_787751 + 8'h01;
  assign sel_787755 = array_index_787662 == array_index_772774 ? add_787754 : sel_787751;
  assign add_787758 = sel_787755 + 8'h01;
  assign sel_787759 = array_index_787662 == array_index_772780 ? add_787758 : sel_787755;
  assign add_787762 = sel_787759 + 8'h01;
  assign sel_787763 = array_index_787662 == array_index_772786 ? add_787762 : sel_787759;
  assign add_787766 = sel_787763 + 8'h01;
  assign sel_787767 = array_index_787662 == array_index_772792 ? add_787766 : sel_787763;
  assign add_787770 = sel_787767 + 8'h01;
  assign sel_787771 = array_index_787662 == array_index_772798 ? add_787770 : sel_787767;
  assign add_787774 = sel_787771 + 8'h01;
  assign sel_787775 = array_index_787662 == array_index_772804 ? add_787774 : sel_787771;
  assign add_787778 = sel_787775 + 8'h01;
  assign sel_787779 = array_index_787662 == array_index_772810 ? add_787778 : sel_787775;
  assign add_787782 = sel_787779 + 8'h01;
  assign sel_787783 = array_index_787662 == array_index_772816 ? add_787782 : sel_787779;
  assign add_787786 = sel_787783 + 8'h01;
  assign sel_787787 = array_index_787662 == array_index_772822 ? add_787786 : sel_787783;
  assign add_787790 = sel_787787 + 8'h01;
  assign sel_787791 = array_index_787662 == array_index_772828 ? add_787790 : sel_787787;
  assign add_787794 = sel_787791 + 8'h01;
  assign sel_787795 = array_index_787662 == array_index_772834 ? add_787794 : sel_787791;
  assign add_787798 = sel_787795 + 8'h01;
  assign sel_787799 = array_index_787662 == array_index_772840 ? add_787798 : sel_787795;
  assign add_787802 = sel_787799 + 8'h01;
  assign sel_787803 = array_index_787662 == array_index_772846 ? add_787802 : sel_787799;
  assign add_787806 = sel_787803 + 8'h01;
  assign sel_787807 = array_index_787662 == array_index_772852 ? add_787806 : sel_787803;
  assign add_787810 = sel_787807 + 8'h01;
  assign sel_787811 = array_index_787662 == array_index_772858 ? add_787810 : sel_787807;
  assign add_787814 = sel_787811 + 8'h01;
  assign sel_787815 = array_index_787662 == array_index_772864 ? add_787814 : sel_787811;
  assign add_787818 = sel_787815 + 8'h01;
  assign sel_787819 = array_index_787662 == array_index_772870 ? add_787818 : sel_787815;
  assign add_787822 = sel_787819 + 8'h01;
  assign sel_787823 = array_index_787662 == array_index_772876 ? add_787822 : sel_787819;
  assign add_787826 = sel_787823 + 8'h01;
  assign sel_787827 = array_index_787662 == array_index_772882 ? add_787826 : sel_787823;
  assign add_787830 = sel_787827 + 8'h01;
  assign sel_787831 = array_index_787662 == array_index_772888 ? add_787830 : sel_787827;
  assign add_787834 = sel_787831 + 8'h01;
  assign sel_787835 = array_index_787662 == array_index_772894 ? add_787834 : sel_787831;
  assign add_787838 = sel_787835 + 8'h01;
  assign sel_787839 = array_index_787662 == array_index_772900 ? add_787838 : sel_787835;
  assign add_787842 = sel_787839 + 8'h01;
  assign sel_787843 = array_index_787662 == array_index_772906 ? add_787842 : sel_787839;
  assign add_787846 = sel_787843 + 8'h01;
  assign sel_787847 = array_index_787662 == array_index_772912 ? add_787846 : sel_787843;
  assign add_787850 = sel_787847 + 8'h01;
  assign sel_787851 = array_index_787662 == array_index_772918 ? add_787850 : sel_787847;
  assign add_787854 = sel_787851 + 8'h01;
  assign sel_787855 = array_index_787662 == array_index_772924 ? add_787854 : sel_787851;
  assign add_787858 = sel_787855 + 8'h01;
  assign sel_787859 = array_index_787662 == array_index_772930 ? add_787858 : sel_787855;
  assign add_787862 = sel_787859 + 8'h01;
  assign sel_787863 = array_index_787662 == array_index_772936 ? add_787862 : sel_787859;
  assign add_787866 = sel_787863 + 8'h01;
  assign sel_787867 = array_index_787662 == array_index_772942 ? add_787866 : sel_787863;
  assign add_787870 = sel_787867 + 8'h01;
  assign sel_787871 = array_index_787662 == array_index_772948 ? add_787870 : sel_787867;
  assign add_787874 = sel_787871 + 8'h01;
  assign sel_787875 = array_index_787662 == array_index_772954 ? add_787874 : sel_787871;
  assign add_787878 = sel_787875 + 8'h01;
  assign sel_787879 = array_index_787662 == array_index_772960 ? add_787878 : sel_787875;
  assign add_787882 = sel_787879 + 8'h01;
  assign sel_787883 = array_index_787662 == array_index_772966 ? add_787882 : sel_787879;
  assign add_787886 = sel_787883 + 8'h01;
  assign sel_787887 = array_index_787662 == array_index_772972 ? add_787886 : sel_787883;
  assign add_787890 = sel_787887 + 8'h01;
  assign sel_787891 = array_index_787662 == array_index_772978 ? add_787890 : sel_787887;
  assign add_787894 = sel_787891 + 8'h01;
  assign sel_787895 = array_index_787662 == array_index_772984 ? add_787894 : sel_787891;
  assign add_787898 = sel_787895 + 8'h01;
  assign sel_787899 = array_index_787662 == array_index_772990 ? add_787898 : sel_787895;
  assign add_787902 = sel_787899 + 8'h01;
  assign sel_787903 = array_index_787662 == array_index_772996 ? add_787902 : sel_787899;
  assign add_787906 = sel_787903 + 8'h01;
  assign sel_787907 = array_index_787662 == array_index_773002 ? add_787906 : sel_787903;
  assign add_787910 = sel_787907 + 8'h01;
  assign sel_787911 = array_index_787662 == array_index_773008 ? add_787910 : sel_787907;
  assign add_787914 = sel_787911 + 8'h01;
  assign sel_787915 = array_index_787662 == array_index_773014 ? add_787914 : sel_787911;
  assign add_787918 = sel_787915 + 8'h01;
  assign sel_787919 = array_index_787662 == array_index_773020 ? add_787918 : sel_787915;
  assign add_787922 = sel_787919 + 8'h01;
  assign sel_787923 = array_index_787662 == array_index_773026 ? add_787922 : sel_787919;
  assign add_787926 = sel_787923 + 8'h01;
  assign sel_787927 = array_index_787662 == array_index_773032 ? add_787926 : sel_787923;
  assign add_787930 = sel_787927 + 8'h01;
  assign sel_787931 = array_index_787662 == array_index_773038 ? add_787930 : sel_787927;
  assign add_787934 = sel_787931 + 8'h01;
  assign sel_787935 = array_index_787662 == array_index_773044 ? add_787934 : sel_787931;
  assign add_787938 = sel_787935 + 8'h01;
  assign sel_787939 = array_index_787662 == array_index_773050 ? add_787938 : sel_787935;
  assign add_787942 = sel_787939 + 8'h01;
  assign sel_787943 = array_index_787662 == array_index_773056 ? add_787942 : sel_787939;
  assign add_787946 = sel_787943 + 8'h01;
  assign sel_787947 = array_index_787662 == array_index_773062 ? add_787946 : sel_787943;
  assign add_787950 = sel_787947 + 8'h01;
  assign sel_787951 = array_index_787662 == array_index_773068 ? add_787950 : sel_787947;
  assign add_787954 = sel_787951 + 8'h01;
  assign sel_787955 = array_index_787662 == array_index_773074 ? add_787954 : sel_787951;
  assign add_787958 = sel_787955 + 8'h01;
  assign sel_787959 = array_index_787662 == array_index_773080 ? add_787958 : sel_787955;
  assign add_787962 = sel_787959 + 8'h01;
  assign sel_787963 = array_index_787662 == array_index_773086 ? add_787962 : sel_787959;
  assign add_787966 = sel_787963 + 8'h01;
  assign sel_787967 = array_index_787662 == array_index_773092 ? add_787966 : sel_787963;
  assign add_787970 = sel_787967 + 8'h01;
  assign sel_787971 = array_index_787662 == array_index_773098 ? add_787970 : sel_787967;
  assign add_787974 = sel_787971 + 8'h01;
  assign sel_787975 = array_index_787662 == array_index_773104 ? add_787974 : sel_787971;
  assign add_787978 = sel_787975 + 8'h01;
  assign sel_787979 = array_index_787662 == array_index_773110 ? add_787978 : sel_787975;
  assign add_787982 = sel_787979 + 8'h01;
  assign sel_787983 = array_index_787662 == array_index_773116 ? add_787982 : sel_787979;
  assign add_787986 = sel_787983 + 8'h01;
  assign sel_787987 = array_index_787662 == array_index_773122 ? add_787986 : sel_787983;
  assign add_787990 = sel_787987 + 8'h01;
  assign sel_787991 = array_index_787662 == array_index_773128 ? add_787990 : sel_787987;
  assign add_787994 = sel_787991 + 8'h01;
  assign sel_787995 = array_index_787662 == array_index_773134 ? add_787994 : sel_787991;
  assign add_787998 = sel_787995 + 8'h01;
  assign sel_787999 = array_index_787662 == array_index_773140 ? add_787998 : sel_787995;
  assign add_788002 = sel_787999 + 8'h01;
  assign sel_788003 = array_index_787662 == array_index_773146 ? add_788002 : sel_787999;
  assign add_788006 = sel_788003 + 8'h01;
  assign sel_788007 = array_index_787662 == array_index_773152 ? add_788006 : sel_788003;
  assign add_788010 = sel_788007 + 8'h01;
  assign sel_788011 = array_index_787662 == array_index_773158 ? add_788010 : sel_788007;
  assign add_788014 = sel_788011 + 8'h01;
  assign sel_788015 = array_index_787662 == array_index_773164 ? add_788014 : sel_788011;
  assign add_788018 = sel_788015 + 8'h01;
  assign sel_788019 = array_index_787662 == array_index_773170 ? add_788018 : sel_788015;
  assign add_788023 = sel_788019 + 8'h01;
  assign array_index_788024 = set1_unflattened[7'h2a];
  assign sel_788025 = array_index_787662 == array_index_773176 ? add_788023 : sel_788019;
  assign add_788028 = sel_788025 + 8'h01;
  assign sel_788029 = array_index_788024 == array_index_772632 ? add_788028 : sel_788025;
  assign add_788032 = sel_788029 + 8'h01;
  assign sel_788033 = array_index_788024 == array_index_772636 ? add_788032 : sel_788029;
  assign add_788036 = sel_788033 + 8'h01;
  assign sel_788037 = array_index_788024 == array_index_772644 ? add_788036 : sel_788033;
  assign add_788040 = sel_788037 + 8'h01;
  assign sel_788041 = array_index_788024 == array_index_772652 ? add_788040 : sel_788037;
  assign add_788044 = sel_788041 + 8'h01;
  assign sel_788045 = array_index_788024 == array_index_772660 ? add_788044 : sel_788041;
  assign add_788048 = sel_788045 + 8'h01;
  assign sel_788049 = array_index_788024 == array_index_772668 ? add_788048 : sel_788045;
  assign add_788052 = sel_788049 + 8'h01;
  assign sel_788053 = array_index_788024 == array_index_772676 ? add_788052 : sel_788049;
  assign add_788056 = sel_788053 + 8'h01;
  assign sel_788057 = array_index_788024 == array_index_772684 ? add_788056 : sel_788053;
  assign add_788060 = sel_788057 + 8'h01;
  assign sel_788061 = array_index_788024 == array_index_772690 ? add_788060 : sel_788057;
  assign add_788064 = sel_788061 + 8'h01;
  assign sel_788065 = array_index_788024 == array_index_772696 ? add_788064 : sel_788061;
  assign add_788068 = sel_788065 + 8'h01;
  assign sel_788069 = array_index_788024 == array_index_772702 ? add_788068 : sel_788065;
  assign add_788072 = sel_788069 + 8'h01;
  assign sel_788073 = array_index_788024 == array_index_772708 ? add_788072 : sel_788069;
  assign add_788076 = sel_788073 + 8'h01;
  assign sel_788077 = array_index_788024 == array_index_772714 ? add_788076 : sel_788073;
  assign add_788080 = sel_788077 + 8'h01;
  assign sel_788081 = array_index_788024 == array_index_772720 ? add_788080 : sel_788077;
  assign add_788084 = sel_788081 + 8'h01;
  assign sel_788085 = array_index_788024 == array_index_772726 ? add_788084 : sel_788081;
  assign add_788088 = sel_788085 + 8'h01;
  assign sel_788089 = array_index_788024 == array_index_772732 ? add_788088 : sel_788085;
  assign add_788092 = sel_788089 + 8'h01;
  assign sel_788093 = array_index_788024 == array_index_772738 ? add_788092 : sel_788089;
  assign add_788096 = sel_788093 + 8'h01;
  assign sel_788097 = array_index_788024 == array_index_772744 ? add_788096 : sel_788093;
  assign add_788100 = sel_788097 + 8'h01;
  assign sel_788101 = array_index_788024 == array_index_772750 ? add_788100 : sel_788097;
  assign add_788104 = sel_788101 + 8'h01;
  assign sel_788105 = array_index_788024 == array_index_772756 ? add_788104 : sel_788101;
  assign add_788108 = sel_788105 + 8'h01;
  assign sel_788109 = array_index_788024 == array_index_772762 ? add_788108 : sel_788105;
  assign add_788112 = sel_788109 + 8'h01;
  assign sel_788113 = array_index_788024 == array_index_772768 ? add_788112 : sel_788109;
  assign add_788116 = sel_788113 + 8'h01;
  assign sel_788117 = array_index_788024 == array_index_772774 ? add_788116 : sel_788113;
  assign add_788120 = sel_788117 + 8'h01;
  assign sel_788121 = array_index_788024 == array_index_772780 ? add_788120 : sel_788117;
  assign add_788124 = sel_788121 + 8'h01;
  assign sel_788125 = array_index_788024 == array_index_772786 ? add_788124 : sel_788121;
  assign add_788128 = sel_788125 + 8'h01;
  assign sel_788129 = array_index_788024 == array_index_772792 ? add_788128 : sel_788125;
  assign add_788132 = sel_788129 + 8'h01;
  assign sel_788133 = array_index_788024 == array_index_772798 ? add_788132 : sel_788129;
  assign add_788136 = sel_788133 + 8'h01;
  assign sel_788137 = array_index_788024 == array_index_772804 ? add_788136 : sel_788133;
  assign add_788140 = sel_788137 + 8'h01;
  assign sel_788141 = array_index_788024 == array_index_772810 ? add_788140 : sel_788137;
  assign add_788144 = sel_788141 + 8'h01;
  assign sel_788145 = array_index_788024 == array_index_772816 ? add_788144 : sel_788141;
  assign add_788148 = sel_788145 + 8'h01;
  assign sel_788149 = array_index_788024 == array_index_772822 ? add_788148 : sel_788145;
  assign add_788152 = sel_788149 + 8'h01;
  assign sel_788153 = array_index_788024 == array_index_772828 ? add_788152 : sel_788149;
  assign add_788156 = sel_788153 + 8'h01;
  assign sel_788157 = array_index_788024 == array_index_772834 ? add_788156 : sel_788153;
  assign add_788160 = sel_788157 + 8'h01;
  assign sel_788161 = array_index_788024 == array_index_772840 ? add_788160 : sel_788157;
  assign add_788164 = sel_788161 + 8'h01;
  assign sel_788165 = array_index_788024 == array_index_772846 ? add_788164 : sel_788161;
  assign add_788168 = sel_788165 + 8'h01;
  assign sel_788169 = array_index_788024 == array_index_772852 ? add_788168 : sel_788165;
  assign add_788172 = sel_788169 + 8'h01;
  assign sel_788173 = array_index_788024 == array_index_772858 ? add_788172 : sel_788169;
  assign add_788176 = sel_788173 + 8'h01;
  assign sel_788177 = array_index_788024 == array_index_772864 ? add_788176 : sel_788173;
  assign add_788180 = sel_788177 + 8'h01;
  assign sel_788181 = array_index_788024 == array_index_772870 ? add_788180 : sel_788177;
  assign add_788184 = sel_788181 + 8'h01;
  assign sel_788185 = array_index_788024 == array_index_772876 ? add_788184 : sel_788181;
  assign add_788188 = sel_788185 + 8'h01;
  assign sel_788189 = array_index_788024 == array_index_772882 ? add_788188 : sel_788185;
  assign add_788192 = sel_788189 + 8'h01;
  assign sel_788193 = array_index_788024 == array_index_772888 ? add_788192 : sel_788189;
  assign add_788196 = sel_788193 + 8'h01;
  assign sel_788197 = array_index_788024 == array_index_772894 ? add_788196 : sel_788193;
  assign add_788200 = sel_788197 + 8'h01;
  assign sel_788201 = array_index_788024 == array_index_772900 ? add_788200 : sel_788197;
  assign add_788204 = sel_788201 + 8'h01;
  assign sel_788205 = array_index_788024 == array_index_772906 ? add_788204 : sel_788201;
  assign add_788208 = sel_788205 + 8'h01;
  assign sel_788209 = array_index_788024 == array_index_772912 ? add_788208 : sel_788205;
  assign add_788212 = sel_788209 + 8'h01;
  assign sel_788213 = array_index_788024 == array_index_772918 ? add_788212 : sel_788209;
  assign add_788216 = sel_788213 + 8'h01;
  assign sel_788217 = array_index_788024 == array_index_772924 ? add_788216 : sel_788213;
  assign add_788220 = sel_788217 + 8'h01;
  assign sel_788221 = array_index_788024 == array_index_772930 ? add_788220 : sel_788217;
  assign add_788224 = sel_788221 + 8'h01;
  assign sel_788225 = array_index_788024 == array_index_772936 ? add_788224 : sel_788221;
  assign add_788228 = sel_788225 + 8'h01;
  assign sel_788229 = array_index_788024 == array_index_772942 ? add_788228 : sel_788225;
  assign add_788232 = sel_788229 + 8'h01;
  assign sel_788233 = array_index_788024 == array_index_772948 ? add_788232 : sel_788229;
  assign add_788236 = sel_788233 + 8'h01;
  assign sel_788237 = array_index_788024 == array_index_772954 ? add_788236 : sel_788233;
  assign add_788240 = sel_788237 + 8'h01;
  assign sel_788241 = array_index_788024 == array_index_772960 ? add_788240 : sel_788237;
  assign add_788244 = sel_788241 + 8'h01;
  assign sel_788245 = array_index_788024 == array_index_772966 ? add_788244 : sel_788241;
  assign add_788248 = sel_788245 + 8'h01;
  assign sel_788249 = array_index_788024 == array_index_772972 ? add_788248 : sel_788245;
  assign add_788252 = sel_788249 + 8'h01;
  assign sel_788253 = array_index_788024 == array_index_772978 ? add_788252 : sel_788249;
  assign add_788256 = sel_788253 + 8'h01;
  assign sel_788257 = array_index_788024 == array_index_772984 ? add_788256 : sel_788253;
  assign add_788260 = sel_788257 + 8'h01;
  assign sel_788261 = array_index_788024 == array_index_772990 ? add_788260 : sel_788257;
  assign add_788264 = sel_788261 + 8'h01;
  assign sel_788265 = array_index_788024 == array_index_772996 ? add_788264 : sel_788261;
  assign add_788268 = sel_788265 + 8'h01;
  assign sel_788269 = array_index_788024 == array_index_773002 ? add_788268 : sel_788265;
  assign add_788272 = sel_788269 + 8'h01;
  assign sel_788273 = array_index_788024 == array_index_773008 ? add_788272 : sel_788269;
  assign add_788276 = sel_788273 + 8'h01;
  assign sel_788277 = array_index_788024 == array_index_773014 ? add_788276 : sel_788273;
  assign add_788280 = sel_788277 + 8'h01;
  assign sel_788281 = array_index_788024 == array_index_773020 ? add_788280 : sel_788277;
  assign add_788284 = sel_788281 + 8'h01;
  assign sel_788285 = array_index_788024 == array_index_773026 ? add_788284 : sel_788281;
  assign add_788288 = sel_788285 + 8'h01;
  assign sel_788289 = array_index_788024 == array_index_773032 ? add_788288 : sel_788285;
  assign add_788292 = sel_788289 + 8'h01;
  assign sel_788293 = array_index_788024 == array_index_773038 ? add_788292 : sel_788289;
  assign add_788296 = sel_788293 + 8'h01;
  assign sel_788297 = array_index_788024 == array_index_773044 ? add_788296 : sel_788293;
  assign add_788300 = sel_788297 + 8'h01;
  assign sel_788301 = array_index_788024 == array_index_773050 ? add_788300 : sel_788297;
  assign add_788304 = sel_788301 + 8'h01;
  assign sel_788305 = array_index_788024 == array_index_773056 ? add_788304 : sel_788301;
  assign add_788308 = sel_788305 + 8'h01;
  assign sel_788309 = array_index_788024 == array_index_773062 ? add_788308 : sel_788305;
  assign add_788312 = sel_788309 + 8'h01;
  assign sel_788313 = array_index_788024 == array_index_773068 ? add_788312 : sel_788309;
  assign add_788316 = sel_788313 + 8'h01;
  assign sel_788317 = array_index_788024 == array_index_773074 ? add_788316 : sel_788313;
  assign add_788320 = sel_788317 + 8'h01;
  assign sel_788321 = array_index_788024 == array_index_773080 ? add_788320 : sel_788317;
  assign add_788324 = sel_788321 + 8'h01;
  assign sel_788325 = array_index_788024 == array_index_773086 ? add_788324 : sel_788321;
  assign add_788328 = sel_788325 + 8'h01;
  assign sel_788329 = array_index_788024 == array_index_773092 ? add_788328 : sel_788325;
  assign add_788332 = sel_788329 + 8'h01;
  assign sel_788333 = array_index_788024 == array_index_773098 ? add_788332 : sel_788329;
  assign add_788336 = sel_788333 + 8'h01;
  assign sel_788337 = array_index_788024 == array_index_773104 ? add_788336 : sel_788333;
  assign add_788340 = sel_788337 + 8'h01;
  assign sel_788341 = array_index_788024 == array_index_773110 ? add_788340 : sel_788337;
  assign add_788344 = sel_788341 + 8'h01;
  assign sel_788345 = array_index_788024 == array_index_773116 ? add_788344 : sel_788341;
  assign add_788348 = sel_788345 + 8'h01;
  assign sel_788349 = array_index_788024 == array_index_773122 ? add_788348 : sel_788345;
  assign add_788352 = sel_788349 + 8'h01;
  assign sel_788353 = array_index_788024 == array_index_773128 ? add_788352 : sel_788349;
  assign add_788356 = sel_788353 + 8'h01;
  assign sel_788357 = array_index_788024 == array_index_773134 ? add_788356 : sel_788353;
  assign add_788360 = sel_788357 + 8'h01;
  assign sel_788361 = array_index_788024 == array_index_773140 ? add_788360 : sel_788357;
  assign add_788364 = sel_788361 + 8'h01;
  assign sel_788365 = array_index_788024 == array_index_773146 ? add_788364 : sel_788361;
  assign add_788368 = sel_788365 + 8'h01;
  assign sel_788369 = array_index_788024 == array_index_773152 ? add_788368 : sel_788365;
  assign add_788372 = sel_788369 + 8'h01;
  assign sel_788373 = array_index_788024 == array_index_773158 ? add_788372 : sel_788369;
  assign add_788376 = sel_788373 + 8'h01;
  assign sel_788377 = array_index_788024 == array_index_773164 ? add_788376 : sel_788373;
  assign add_788380 = sel_788377 + 8'h01;
  assign sel_788381 = array_index_788024 == array_index_773170 ? add_788380 : sel_788377;
  assign add_788385 = sel_788381 + 8'h01;
  assign array_index_788386 = set1_unflattened[7'h2b];
  assign sel_788387 = array_index_788024 == array_index_773176 ? add_788385 : sel_788381;
  assign add_788390 = sel_788387 + 8'h01;
  assign sel_788391 = array_index_788386 == array_index_772632 ? add_788390 : sel_788387;
  assign add_788394 = sel_788391 + 8'h01;
  assign sel_788395 = array_index_788386 == array_index_772636 ? add_788394 : sel_788391;
  assign add_788398 = sel_788395 + 8'h01;
  assign sel_788399 = array_index_788386 == array_index_772644 ? add_788398 : sel_788395;
  assign add_788402 = sel_788399 + 8'h01;
  assign sel_788403 = array_index_788386 == array_index_772652 ? add_788402 : sel_788399;
  assign add_788406 = sel_788403 + 8'h01;
  assign sel_788407 = array_index_788386 == array_index_772660 ? add_788406 : sel_788403;
  assign add_788410 = sel_788407 + 8'h01;
  assign sel_788411 = array_index_788386 == array_index_772668 ? add_788410 : sel_788407;
  assign add_788414 = sel_788411 + 8'h01;
  assign sel_788415 = array_index_788386 == array_index_772676 ? add_788414 : sel_788411;
  assign add_788418 = sel_788415 + 8'h01;
  assign sel_788419 = array_index_788386 == array_index_772684 ? add_788418 : sel_788415;
  assign add_788422 = sel_788419 + 8'h01;
  assign sel_788423 = array_index_788386 == array_index_772690 ? add_788422 : sel_788419;
  assign add_788426 = sel_788423 + 8'h01;
  assign sel_788427 = array_index_788386 == array_index_772696 ? add_788426 : sel_788423;
  assign add_788430 = sel_788427 + 8'h01;
  assign sel_788431 = array_index_788386 == array_index_772702 ? add_788430 : sel_788427;
  assign add_788434 = sel_788431 + 8'h01;
  assign sel_788435 = array_index_788386 == array_index_772708 ? add_788434 : sel_788431;
  assign add_788438 = sel_788435 + 8'h01;
  assign sel_788439 = array_index_788386 == array_index_772714 ? add_788438 : sel_788435;
  assign add_788442 = sel_788439 + 8'h01;
  assign sel_788443 = array_index_788386 == array_index_772720 ? add_788442 : sel_788439;
  assign add_788446 = sel_788443 + 8'h01;
  assign sel_788447 = array_index_788386 == array_index_772726 ? add_788446 : sel_788443;
  assign add_788450 = sel_788447 + 8'h01;
  assign sel_788451 = array_index_788386 == array_index_772732 ? add_788450 : sel_788447;
  assign add_788454 = sel_788451 + 8'h01;
  assign sel_788455 = array_index_788386 == array_index_772738 ? add_788454 : sel_788451;
  assign add_788458 = sel_788455 + 8'h01;
  assign sel_788459 = array_index_788386 == array_index_772744 ? add_788458 : sel_788455;
  assign add_788462 = sel_788459 + 8'h01;
  assign sel_788463 = array_index_788386 == array_index_772750 ? add_788462 : sel_788459;
  assign add_788466 = sel_788463 + 8'h01;
  assign sel_788467 = array_index_788386 == array_index_772756 ? add_788466 : sel_788463;
  assign add_788470 = sel_788467 + 8'h01;
  assign sel_788471 = array_index_788386 == array_index_772762 ? add_788470 : sel_788467;
  assign add_788474 = sel_788471 + 8'h01;
  assign sel_788475 = array_index_788386 == array_index_772768 ? add_788474 : sel_788471;
  assign add_788478 = sel_788475 + 8'h01;
  assign sel_788479 = array_index_788386 == array_index_772774 ? add_788478 : sel_788475;
  assign add_788482 = sel_788479 + 8'h01;
  assign sel_788483 = array_index_788386 == array_index_772780 ? add_788482 : sel_788479;
  assign add_788486 = sel_788483 + 8'h01;
  assign sel_788487 = array_index_788386 == array_index_772786 ? add_788486 : sel_788483;
  assign add_788490 = sel_788487 + 8'h01;
  assign sel_788491 = array_index_788386 == array_index_772792 ? add_788490 : sel_788487;
  assign add_788494 = sel_788491 + 8'h01;
  assign sel_788495 = array_index_788386 == array_index_772798 ? add_788494 : sel_788491;
  assign add_788498 = sel_788495 + 8'h01;
  assign sel_788499 = array_index_788386 == array_index_772804 ? add_788498 : sel_788495;
  assign add_788502 = sel_788499 + 8'h01;
  assign sel_788503 = array_index_788386 == array_index_772810 ? add_788502 : sel_788499;
  assign add_788506 = sel_788503 + 8'h01;
  assign sel_788507 = array_index_788386 == array_index_772816 ? add_788506 : sel_788503;
  assign add_788510 = sel_788507 + 8'h01;
  assign sel_788511 = array_index_788386 == array_index_772822 ? add_788510 : sel_788507;
  assign add_788514 = sel_788511 + 8'h01;
  assign sel_788515 = array_index_788386 == array_index_772828 ? add_788514 : sel_788511;
  assign add_788518 = sel_788515 + 8'h01;
  assign sel_788519 = array_index_788386 == array_index_772834 ? add_788518 : sel_788515;
  assign add_788522 = sel_788519 + 8'h01;
  assign sel_788523 = array_index_788386 == array_index_772840 ? add_788522 : sel_788519;
  assign add_788526 = sel_788523 + 8'h01;
  assign sel_788527 = array_index_788386 == array_index_772846 ? add_788526 : sel_788523;
  assign add_788530 = sel_788527 + 8'h01;
  assign sel_788531 = array_index_788386 == array_index_772852 ? add_788530 : sel_788527;
  assign add_788534 = sel_788531 + 8'h01;
  assign sel_788535 = array_index_788386 == array_index_772858 ? add_788534 : sel_788531;
  assign add_788538 = sel_788535 + 8'h01;
  assign sel_788539 = array_index_788386 == array_index_772864 ? add_788538 : sel_788535;
  assign add_788542 = sel_788539 + 8'h01;
  assign sel_788543 = array_index_788386 == array_index_772870 ? add_788542 : sel_788539;
  assign add_788546 = sel_788543 + 8'h01;
  assign sel_788547 = array_index_788386 == array_index_772876 ? add_788546 : sel_788543;
  assign add_788550 = sel_788547 + 8'h01;
  assign sel_788551 = array_index_788386 == array_index_772882 ? add_788550 : sel_788547;
  assign add_788554 = sel_788551 + 8'h01;
  assign sel_788555 = array_index_788386 == array_index_772888 ? add_788554 : sel_788551;
  assign add_788558 = sel_788555 + 8'h01;
  assign sel_788559 = array_index_788386 == array_index_772894 ? add_788558 : sel_788555;
  assign add_788562 = sel_788559 + 8'h01;
  assign sel_788563 = array_index_788386 == array_index_772900 ? add_788562 : sel_788559;
  assign add_788566 = sel_788563 + 8'h01;
  assign sel_788567 = array_index_788386 == array_index_772906 ? add_788566 : sel_788563;
  assign add_788570 = sel_788567 + 8'h01;
  assign sel_788571 = array_index_788386 == array_index_772912 ? add_788570 : sel_788567;
  assign add_788574 = sel_788571 + 8'h01;
  assign sel_788575 = array_index_788386 == array_index_772918 ? add_788574 : sel_788571;
  assign add_788578 = sel_788575 + 8'h01;
  assign sel_788579 = array_index_788386 == array_index_772924 ? add_788578 : sel_788575;
  assign add_788582 = sel_788579 + 8'h01;
  assign sel_788583 = array_index_788386 == array_index_772930 ? add_788582 : sel_788579;
  assign add_788586 = sel_788583 + 8'h01;
  assign sel_788587 = array_index_788386 == array_index_772936 ? add_788586 : sel_788583;
  assign add_788590 = sel_788587 + 8'h01;
  assign sel_788591 = array_index_788386 == array_index_772942 ? add_788590 : sel_788587;
  assign add_788594 = sel_788591 + 8'h01;
  assign sel_788595 = array_index_788386 == array_index_772948 ? add_788594 : sel_788591;
  assign add_788598 = sel_788595 + 8'h01;
  assign sel_788599 = array_index_788386 == array_index_772954 ? add_788598 : sel_788595;
  assign add_788602 = sel_788599 + 8'h01;
  assign sel_788603 = array_index_788386 == array_index_772960 ? add_788602 : sel_788599;
  assign add_788606 = sel_788603 + 8'h01;
  assign sel_788607 = array_index_788386 == array_index_772966 ? add_788606 : sel_788603;
  assign add_788610 = sel_788607 + 8'h01;
  assign sel_788611 = array_index_788386 == array_index_772972 ? add_788610 : sel_788607;
  assign add_788614 = sel_788611 + 8'h01;
  assign sel_788615 = array_index_788386 == array_index_772978 ? add_788614 : sel_788611;
  assign add_788618 = sel_788615 + 8'h01;
  assign sel_788619 = array_index_788386 == array_index_772984 ? add_788618 : sel_788615;
  assign add_788622 = sel_788619 + 8'h01;
  assign sel_788623 = array_index_788386 == array_index_772990 ? add_788622 : sel_788619;
  assign add_788626 = sel_788623 + 8'h01;
  assign sel_788627 = array_index_788386 == array_index_772996 ? add_788626 : sel_788623;
  assign add_788630 = sel_788627 + 8'h01;
  assign sel_788631 = array_index_788386 == array_index_773002 ? add_788630 : sel_788627;
  assign add_788634 = sel_788631 + 8'h01;
  assign sel_788635 = array_index_788386 == array_index_773008 ? add_788634 : sel_788631;
  assign add_788638 = sel_788635 + 8'h01;
  assign sel_788639 = array_index_788386 == array_index_773014 ? add_788638 : sel_788635;
  assign add_788642 = sel_788639 + 8'h01;
  assign sel_788643 = array_index_788386 == array_index_773020 ? add_788642 : sel_788639;
  assign add_788646 = sel_788643 + 8'h01;
  assign sel_788647 = array_index_788386 == array_index_773026 ? add_788646 : sel_788643;
  assign add_788650 = sel_788647 + 8'h01;
  assign sel_788651 = array_index_788386 == array_index_773032 ? add_788650 : sel_788647;
  assign add_788654 = sel_788651 + 8'h01;
  assign sel_788655 = array_index_788386 == array_index_773038 ? add_788654 : sel_788651;
  assign add_788658 = sel_788655 + 8'h01;
  assign sel_788659 = array_index_788386 == array_index_773044 ? add_788658 : sel_788655;
  assign add_788662 = sel_788659 + 8'h01;
  assign sel_788663 = array_index_788386 == array_index_773050 ? add_788662 : sel_788659;
  assign add_788666 = sel_788663 + 8'h01;
  assign sel_788667 = array_index_788386 == array_index_773056 ? add_788666 : sel_788663;
  assign add_788670 = sel_788667 + 8'h01;
  assign sel_788671 = array_index_788386 == array_index_773062 ? add_788670 : sel_788667;
  assign add_788674 = sel_788671 + 8'h01;
  assign sel_788675 = array_index_788386 == array_index_773068 ? add_788674 : sel_788671;
  assign add_788678 = sel_788675 + 8'h01;
  assign sel_788679 = array_index_788386 == array_index_773074 ? add_788678 : sel_788675;
  assign add_788682 = sel_788679 + 8'h01;
  assign sel_788683 = array_index_788386 == array_index_773080 ? add_788682 : sel_788679;
  assign add_788686 = sel_788683 + 8'h01;
  assign sel_788687 = array_index_788386 == array_index_773086 ? add_788686 : sel_788683;
  assign add_788690 = sel_788687 + 8'h01;
  assign sel_788691 = array_index_788386 == array_index_773092 ? add_788690 : sel_788687;
  assign add_788694 = sel_788691 + 8'h01;
  assign sel_788695 = array_index_788386 == array_index_773098 ? add_788694 : sel_788691;
  assign add_788698 = sel_788695 + 8'h01;
  assign sel_788699 = array_index_788386 == array_index_773104 ? add_788698 : sel_788695;
  assign add_788702 = sel_788699 + 8'h01;
  assign sel_788703 = array_index_788386 == array_index_773110 ? add_788702 : sel_788699;
  assign add_788706 = sel_788703 + 8'h01;
  assign sel_788707 = array_index_788386 == array_index_773116 ? add_788706 : sel_788703;
  assign add_788710 = sel_788707 + 8'h01;
  assign sel_788711 = array_index_788386 == array_index_773122 ? add_788710 : sel_788707;
  assign add_788714 = sel_788711 + 8'h01;
  assign sel_788715 = array_index_788386 == array_index_773128 ? add_788714 : sel_788711;
  assign add_788718 = sel_788715 + 8'h01;
  assign sel_788719 = array_index_788386 == array_index_773134 ? add_788718 : sel_788715;
  assign add_788722 = sel_788719 + 8'h01;
  assign sel_788723 = array_index_788386 == array_index_773140 ? add_788722 : sel_788719;
  assign add_788726 = sel_788723 + 8'h01;
  assign sel_788727 = array_index_788386 == array_index_773146 ? add_788726 : sel_788723;
  assign add_788730 = sel_788727 + 8'h01;
  assign sel_788731 = array_index_788386 == array_index_773152 ? add_788730 : sel_788727;
  assign add_788734 = sel_788731 + 8'h01;
  assign sel_788735 = array_index_788386 == array_index_773158 ? add_788734 : sel_788731;
  assign add_788738 = sel_788735 + 8'h01;
  assign sel_788739 = array_index_788386 == array_index_773164 ? add_788738 : sel_788735;
  assign add_788742 = sel_788739 + 8'h01;
  assign sel_788743 = array_index_788386 == array_index_773170 ? add_788742 : sel_788739;
  assign add_788747 = sel_788743 + 8'h01;
  assign array_index_788748 = set1_unflattened[7'h2c];
  assign sel_788749 = array_index_788386 == array_index_773176 ? add_788747 : sel_788743;
  assign add_788752 = sel_788749 + 8'h01;
  assign sel_788753 = array_index_788748 == array_index_772632 ? add_788752 : sel_788749;
  assign add_788756 = sel_788753 + 8'h01;
  assign sel_788757 = array_index_788748 == array_index_772636 ? add_788756 : sel_788753;
  assign add_788760 = sel_788757 + 8'h01;
  assign sel_788761 = array_index_788748 == array_index_772644 ? add_788760 : sel_788757;
  assign add_788764 = sel_788761 + 8'h01;
  assign sel_788765 = array_index_788748 == array_index_772652 ? add_788764 : sel_788761;
  assign add_788768 = sel_788765 + 8'h01;
  assign sel_788769 = array_index_788748 == array_index_772660 ? add_788768 : sel_788765;
  assign add_788772 = sel_788769 + 8'h01;
  assign sel_788773 = array_index_788748 == array_index_772668 ? add_788772 : sel_788769;
  assign add_788776 = sel_788773 + 8'h01;
  assign sel_788777 = array_index_788748 == array_index_772676 ? add_788776 : sel_788773;
  assign add_788780 = sel_788777 + 8'h01;
  assign sel_788781 = array_index_788748 == array_index_772684 ? add_788780 : sel_788777;
  assign add_788784 = sel_788781 + 8'h01;
  assign sel_788785 = array_index_788748 == array_index_772690 ? add_788784 : sel_788781;
  assign add_788788 = sel_788785 + 8'h01;
  assign sel_788789 = array_index_788748 == array_index_772696 ? add_788788 : sel_788785;
  assign add_788792 = sel_788789 + 8'h01;
  assign sel_788793 = array_index_788748 == array_index_772702 ? add_788792 : sel_788789;
  assign add_788796 = sel_788793 + 8'h01;
  assign sel_788797 = array_index_788748 == array_index_772708 ? add_788796 : sel_788793;
  assign add_788800 = sel_788797 + 8'h01;
  assign sel_788801 = array_index_788748 == array_index_772714 ? add_788800 : sel_788797;
  assign add_788804 = sel_788801 + 8'h01;
  assign sel_788805 = array_index_788748 == array_index_772720 ? add_788804 : sel_788801;
  assign add_788808 = sel_788805 + 8'h01;
  assign sel_788809 = array_index_788748 == array_index_772726 ? add_788808 : sel_788805;
  assign add_788812 = sel_788809 + 8'h01;
  assign sel_788813 = array_index_788748 == array_index_772732 ? add_788812 : sel_788809;
  assign add_788816 = sel_788813 + 8'h01;
  assign sel_788817 = array_index_788748 == array_index_772738 ? add_788816 : sel_788813;
  assign add_788820 = sel_788817 + 8'h01;
  assign sel_788821 = array_index_788748 == array_index_772744 ? add_788820 : sel_788817;
  assign add_788824 = sel_788821 + 8'h01;
  assign sel_788825 = array_index_788748 == array_index_772750 ? add_788824 : sel_788821;
  assign add_788828 = sel_788825 + 8'h01;
  assign sel_788829 = array_index_788748 == array_index_772756 ? add_788828 : sel_788825;
  assign add_788832 = sel_788829 + 8'h01;
  assign sel_788833 = array_index_788748 == array_index_772762 ? add_788832 : sel_788829;
  assign add_788836 = sel_788833 + 8'h01;
  assign sel_788837 = array_index_788748 == array_index_772768 ? add_788836 : sel_788833;
  assign add_788840 = sel_788837 + 8'h01;
  assign sel_788841 = array_index_788748 == array_index_772774 ? add_788840 : sel_788837;
  assign add_788844 = sel_788841 + 8'h01;
  assign sel_788845 = array_index_788748 == array_index_772780 ? add_788844 : sel_788841;
  assign add_788848 = sel_788845 + 8'h01;
  assign sel_788849 = array_index_788748 == array_index_772786 ? add_788848 : sel_788845;
  assign add_788852 = sel_788849 + 8'h01;
  assign sel_788853 = array_index_788748 == array_index_772792 ? add_788852 : sel_788849;
  assign add_788856 = sel_788853 + 8'h01;
  assign sel_788857 = array_index_788748 == array_index_772798 ? add_788856 : sel_788853;
  assign add_788860 = sel_788857 + 8'h01;
  assign sel_788861 = array_index_788748 == array_index_772804 ? add_788860 : sel_788857;
  assign add_788864 = sel_788861 + 8'h01;
  assign sel_788865 = array_index_788748 == array_index_772810 ? add_788864 : sel_788861;
  assign add_788868 = sel_788865 + 8'h01;
  assign sel_788869 = array_index_788748 == array_index_772816 ? add_788868 : sel_788865;
  assign add_788872 = sel_788869 + 8'h01;
  assign sel_788873 = array_index_788748 == array_index_772822 ? add_788872 : sel_788869;
  assign add_788876 = sel_788873 + 8'h01;
  assign sel_788877 = array_index_788748 == array_index_772828 ? add_788876 : sel_788873;
  assign add_788880 = sel_788877 + 8'h01;
  assign sel_788881 = array_index_788748 == array_index_772834 ? add_788880 : sel_788877;
  assign add_788884 = sel_788881 + 8'h01;
  assign sel_788885 = array_index_788748 == array_index_772840 ? add_788884 : sel_788881;
  assign add_788888 = sel_788885 + 8'h01;
  assign sel_788889 = array_index_788748 == array_index_772846 ? add_788888 : sel_788885;
  assign add_788892 = sel_788889 + 8'h01;
  assign sel_788893 = array_index_788748 == array_index_772852 ? add_788892 : sel_788889;
  assign add_788896 = sel_788893 + 8'h01;
  assign sel_788897 = array_index_788748 == array_index_772858 ? add_788896 : sel_788893;
  assign add_788900 = sel_788897 + 8'h01;
  assign sel_788901 = array_index_788748 == array_index_772864 ? add_788900 : sel_788897;
  assign add_788904 = sel_788901 + 8'h01;
  assign sel_788905 = array_index_788748 == array_index_772870 ? add_788904 : sel_788901;
  assign add_788908 = sel_788905 + 8'h01;
  assign sel_788909 = array_index_788748 == array_index_772876 ? add_788908 : sel_788905;
  assign add_788912 = sel_788909 + 8'h01;
  assign sel_788913 = array_index_788748 == array_index_772882 ? add_788912 : sel_788909;
  assign add_788916 = sel_788913 + 8'h01;
  assign sel_788917 = array_index_788748 == array_index_772888 ? add_788916 : sel_788913;
  assign add_788920 = sel_788917 + 8'h01;
  assign sel_788921 = array_index_788748 == array_index_772894 ? add_788920 : sel_788917;
  assign add_788924 = sel_788921 + 8'h01;
  assign sel_788925 = array_index_788748 == array_index_772900 ? add_788924 : sel_788921;
  assign add_788928 = sel_788925 + 8'h01;
  assign sel_788929 = array_index_788748 == array_index_772906 ? add_788928 : sel_788925;
  assign add_788932 = sel_788929 + 8'h01;
  assign sel_788933 = array_index_788748 == array_index_772912 ? add_788932 : sel_788929;
  assign add_788936 = sel_788933 + 8'h01;
  assign sel_788937 = array_index_788748 == array_index_772918 ? add_788936 : sel_788933;
  assign add_788940 = sel_788937 + 8'h01;
  assign sel_788941 = array_index_788748 == array_index_772924 ? add_788940 : sel_788937;
  assign add_788944 = sel_788941 + 8'h01;
  assign sel_788945 = array_index_788748 == array_index_772930 ? add_788944 : sel_788941;
  assign add_788948 = sel_788945 + 8'h01;
  assign sel_788949 = array_index_788748 == array_index_772936 ? add_788948 : sel_788945;
  assign add_788952 = sel_788949 + 8'h01;
  assign sel_788953 = array_index_788748 == array_index_772942 ? add_788952 : sel_788949;
  assign add_788956 = sel_788953 + 8'h01;
  assign sel_788957 = array_index_788748 == array_index_772948 ? add_788956 : sel_788953;
  assign add_788960 = sel_788957 + 8'h01;
  assign sel_788961 = array_index_788748 == array_index_772954 ? add_788960 : sel_788957;
  assign add_788964 = sel_788961 + 8'h01;
  assign sel_788965 = array_index_788748 == array_index_772960 ? add_788964 : sel_788961;
  assign add_788968 = sel_788965 + 8'h01;
  assign sel_788969 = array_index_788748 == array_index_772966 ? add_788968 : sel_788965;
  assign add_788972 = sel_788969 + 8'h01;
  assign sel_788973 = array_index_788748 == array_index_772972 ? add_788972 : sel_788969;
  assign add_788976 = sel_788973 + 8'h01;
  assign sel_788977 = array_index_788748 == array_index_772978 ? add_788976 : sel_788973;
  assign add_788980 = sel_788977 + 8'h01;
  assign sel_788981 = array_index_788748 == array_index_772984 ? add_788980 : sel_788977;
  assign add_788984 = sel_788981 + 8'h01;
  assign sel_788985 = array_index_788748 == array_index_772990 ? add_788984 : sel_788981;
  assign add_788988 = sel_788985 + 8'h01;
  assign sel_788989 = array_index_788748 == array_index_772996 ? add_788988 : sel_788985;
  assign add_788992 = sel_788989 + 8'h01;
  assign sel_788993 = array_index_788748 == array_index_773002 ? add_788992 : sel_788989;
  assign add_788996 = sel_788993 + 8'h01;
  assign sel_788997 = array_index_788748 == array_index_773008 ? add_788996 : sel_788993;
  assign add_789000 = sel_788997 + 8'h01;
  assign sel_789001 = array_index_788748 == array_index_773014 ? add_789000 : sel_788997;
  assign add_789004 = sel_789001 + 8'h01;
  assign sel_789005 = array_index_788748 == array_index_773020 ? add_789004 : sel_789001;
  assign add_789008 = sel_789005 + 8'h01;
  assign sel_789009 = array_index_788748 == array_index_773026 ? add_789008 : sel_789005;
  assign add_789012 = sel_789009 + 8'h01;
  assign sel_789013 = array_index_788748 == array_index_773032 ? add_789012 : sel_789009;
  assign add_789016 = sel_789013 + 8'h01;
  assign sel_789017 = array_index_788748 == array_index_773038 ? add_789016 : sel_789013;
  assign add_789020 = sel_789017 + 8'h01;
  assign sel_789021 = array_index_788748 == array_index_773044 ? add_789020 : sel_789017;
  assign add_789024 = sel_789021 + 8'h01;
  assign sel_789025 = array_index_788748 == array_index_773050 ? add_789024 : sel_789021;
  assign add_789028 = sel_789025 + 8'h01;
  assign sel_789029 = array_index_788748 == array_index_773056 ? add_789028 : sel_789025;
  assign add_789032 = sel_789029 + 8'h01;
  assign sel_789033 = array_index_788748 == array_index_773062 ? add_789032 : sel_789029;
  assign add_789036 = sel_789033 + 8'h01;
  assign sel_789037 = array_index_788748 == array_index_773068 ? add_789036 : sel_789033;
  assign add_789040 = sel_789037 + 8'h01;
  assign sel_789041 = array_index_788748 == array_index_773074 ? add_789040 : sel_789037;
  assign add_789044 = sel_789041 + 8'h01;
  assign sel_789045 = array_index_788748 == array_index_773080 ? add_789044 : sel_789041;
  assign add_789048 = sel_789045 + 8'h01;
  assign sel_789049 = array_index_788748 == array_index_773086 ? add_789048 : sel_789045;
  assign add_789052 = sel_789049 + 8'h01;
  assign sel_789053 = array_index_788748 == array_index_773092 ? add_789052 : sel_789049;
  assign add_789056 = sel_789053 + 8'h01;
  assign sel_789057 = array_index_788748 == array_index_773098 ? add_789056 : sel_789053;
  assign add_789060 = sel_789057 + 8'h01;
  assign sel_789061 = array_index_788748 == array_index_773104 ? add_789060 : sel_789057;
  assign add_789064 = sel_789061 + 8'h01;
  assign sel_789065 = array_index_788748 == array_index_773110 ? add_789064 : sel_789061;
  assign add_789068 = sel_789065 + 8'h01;
  assign sel_789069 = array_index_788748 == array_index_773116 ? add_789068 : sel_789065;
  assign add_789072 = sel_789069 + 8'h01;
  assign sel_789073 = array_index_788748 == array_index_773122 ? add_789072 : sel_789069;
  assign add_789076 = sel_789073 + 8'h01;
  assign sel_789077 = array_index_788748 == array_index_773128 ? add_789076 : sel_789073;
  assign add_789080 = sel_789077 + 8'h01;
  assign sel_789081 = array_index_788748 == array_index_773134 ? add_789080 : sel_789077;
  assign add_789084 = sel_789081 + 8'h01;
  assign sel_789085 = array_index_788748 == array_index_773140 ? add_789084 : sel_789081;
  assign add_789088 = sel_789085 + 8'h01;
  assign sel_789089 = array_index_788748 == array_index_773146 ? add_789088 : sel_789085;
  assign add_789092 = sel_789089 + 8'h01;
  assign sel_789093 = array_index_788748 == array_index_773152 ? add_789092 : sel_789089;
  assign add_789096 = sel_789093 + 8'h01;
  assign sel_789097 = array_index_788748 == array_index_773158 ? add_789096 : sel_789093;
  assign add_789100 = sel_789097 + 8'h01;
  assign sel_789101 = array_index_788748 == array_index_773164 ? add_789100 : sel_789097;
  assign add_789104 = sel_789101 + 8'h01;
  assign sel_789105 = array_index_788748 == array_index_773170 ? add_789104 : sel_789101;
  assign add_789109 = sel_789105 + 8'h01;
  assign array_index_789110 = set1_unflattened[7'h2d];
  assign sel_789111 = array_index_788748 == array_index_773176 ? add_789109 : sel_789105;
  assign add_789114 = sel_789111 + 8'h01;
  assign sel_789115 = array_index_789110 == array_index_772632 ? add_789114 : sel_789111;
  assign add_789118 = sel_789115 + 8'h01;
  assign sel_789119 = array_index_789110 == array_index_772636 ? add_789118 : sel_789115;
  assign add_789122 = sel_789119 + 8'h01;
  assign sel_789123 = array_index_789110 == array_index_772644 ? add_789122 : sel_789119;
  assign add_789126 = sel_789123 + 8'h01;
  assign sel_789127 = array_index_789110 == array_index_772652 ? add_789126 : sel_789123;
  assign add_789130 = sel_789127 + 8'h01;
  assign sel_789131 = array_index_789110 == array_index_772660 ? add_789130 : sel_789127;
  assign add_789134 = sel_789131 + 8'h01;
  assign sel_789135 = array_index_789110 == array_index_772668 ? add_789134 : sel_789131;
  assign add_789138 = sel_789135 + 8'h01;
  assign sel_789139 = array_index_789110 == array_index_772676 ? add_789138 : sel_789135;
  assign add_789142 = sel_789139 + 8'h01;
  assign sel_789143 = array_index_789110 == array_index_772684 ? add_789142 : sel_789139;
  assign add_789146 = sel_789143 + 8'h01;
  assign sel_789147 = array_index_789110 == array_index_772690 ? add_789146 : sel_789143;
  assign add_789150 = sel_789147 + 8'h01;
  assign sel_789151 = array_index_789110 == array_index_772696 ? add_789150 : sel_789147;
  assign add_789154 = sel_789151 + 8'h01;
  assign sel_789155 = array_index_789110 == array_index_772702 ? add_789154 : sel_789151;
  assign add_789158 = sel_789155 + 8'h01;
  assign sel_789159 = array_index_789110 == array_index_772708 ? add_789158 : sel_789155;
  assign add_789162 = sel_789159 + 8'h01;
  assign sel_789163 = array_index_789110 == array_index_772714 ? add_789162 : sel_789159;
  assign add_789166 = sel_789163 + 8'h01;
  assign sel_789167 = array_index_789110 == array_index_772720 ? add_789166 : sel_789163;
  assign add_789170 = sel_789167 + 8'h01;
  assign sel_789171 = array_index_789110 == array_index_772726 ? add_789170 : sel_789167;
  assign add_789174 = sel_789171 + 8'h01;
  assign sel_789175 = array_index_789110 == array_index_772732 ? add_789174 : sel_789171;
  assign add_789178 = sel_789175 + 8'h01;
  assign sel_789179 = array_index_789110 == array_index_772738 ? add_789178 : sel_789175;
  assign add_789182 = sel_789179 + 8'h01;
  assign sel_789183 = array_index_789110 == array_index_772744 ? add_789182 : sel_789179;
  assign add_789186 = sel_789183 + 8'h01;
  assign sel_789187 = array_index_789110 == array_index_772750 ? add_789186 : sel_789183;
  assign add_789190 = sel_789187 + 8'h01;
  assign sel_789191 = array_index_789110 == array_index_772756 ? add_789190 : sel_789187;
  assign add_789194 = sel_789191 + 8'h01;
  assign sel_789195 = array_index_789110 == array_index_772762 ? add_789194 : sel_789191;
  assign add_789198 = sel_789195 + 8'h01;
  assign sel_789199 = array_index_789110 == array_index_772768 ? add_789198 : sel_789195;
  assign add_789202 = sel_789199 + 8'h01;
  assign sel_789203 = array_index_789110 == array_index_772774 ? add_789202 : sel_789199;
  assign add_789206 = sel_789203 + 8'h01;
  assign sel_789207 = array_index_789110 == array_index_772780 ? add_789206 : sel_789203;
  assign add_789210 = sel_789207 + 8'h01;
  assign sel_789211 = array_index_789110 == array_index_772786 ? add_789210 : sel_789207;
  assign add_789214 = sel_789211 + 8'h01;
  assign sel_789215 = array_index_789110 == array_index_772792 ? add_789214 : sel_789211;
  assign add_789218 = sel_789215 + 8'h01;
  assign sel_789219 = array_index_789110 == array_index_772798 ? add_789218 : sel_789215;
  assign add_789222 = sel_789219 + 8'h01;
  assign sel_789223 = array_index_789110 == array_index_772804 ? add_789222 : sel_789219;
  assign add_789226 = sel_789223 + 8'h01;
  assign sel_789227 = array_index_789110 == array_index_772810 ? add_789226 : sel_789223;
  assign add_789230 = sel_789227 + 8'h01;
  assign sel_789231 = array_index_789110 == array_index_772816 ? add_789230 : sel_789227;
  assign add_789234 = sel_789231 + 8'h01;
  assign sel_789235 = array_index_789110 == array_index_772822 ? add_789234 : sel_789231;
  assign add_789238 = sel_789235 + 8'h01;
  assign sel_789239 = array_index_789110 == array_index_772828 ? add_789238 : sel_789235;
  assign add_789242 = sel_789239 + 8'h01;
  assign sel_789243 = array_index_789110 == array_index_772834 ? add_789242 : sel_789239;
  assign add_789246 = sel_789243 + 8'h01;
  assign sel_789247 = array_index_789110 == array_index_772840 ? add_789246 : sel_789243;
  assign add_789250 = sel_789247 + 8'h01;
  assign sel_789251 = array_index_789110 == array_index_772846 ? add_789250 : sel_789247;
  assign add_789254 = sel_789251 + 8'h01;
  assign sel_789255 = array_index_789110 == array_index_772852 ? add_789254 : sel_789251;
  assign add_789258 = sel_789255 + 8'h01;
  assign sel_789259 = array_index_789110 == array_index_772858 ? add_789258 : sel_789255;
  assign add_789262 = sel_789259 + 8'h01;
  assign sel_789263 = array_index_789110 == array_index_772864 ? add_789262 : sel_789259;
  assign add_789266 = sel_789263 + 8'h01;
  assign sel_789267 = array_index_789110 == array_index_772870 ? add_789266 : sel_789263;
  assign add_789270 = sel_789267 + 8'h01;
  assign sel_789271 = array_index_789110 == array_index_772876 ? add_789270 : sel_789267;
  assign add_789274 = sel_789271 + 8'h01;
  assign sel_789275 = array_index_789110 == array_index_772882 ? add_789274 : sel_789271;
  assign add_789278 = sel_789275 + 8'h01;
  assign sel_789279 = array_index_789110 == array_index_772888 ? add_789278 : sel_789275;
  assign add_789282 = sel_789279 + 8'h01;
  assign sel_789283 = array_index_789110 == array_index_772894 ? add_789282 : sel_789279;
  assign add_789286 = sel_789283 + 8'h01;
  assign sel_789287 = array_index_789110 == array_index_772900 ? add_789286 : sel_789283;
  assign add_789290 = sel_789287 + 8'h01;
  assign sel_789291 = array_index_789110 == array_index_772906 ? add_789290 : sel_789287;
  assign add_789294 = sel_789291 + 8'h01;
  assign sel_789295 = array_index_789110 == array_index_772912 ? add_789294 : sel_789291;
  assign add_789298 = sel_789295 + 8'h01;
  assign sel_789299 = array_index_789110 == array_index_772918 ? add_789298 : sel_789295;
  assign add_789302 = sel_789299 + 8'h01;
  assign sel_789303 = array_index_789110 == array_index_772924 ? add_789302 : sel_789299;
  assign add_789306 = sel_789303 + 8'h01;
  assign sel_789307 = array_index_789110 == array_index_772930 ? add_789306 : sel_789303;
  assign add_789310 = sel_789307 + 8'h01;
  assign sel_789311 = array_index_789110 == array_index_772936 ? add_789310 : sel_789307;
  assign add_789314 = sel_789311 + 8'h01;
  assign sel_789315 = array_index_789110 == array_index_772942 ? add_789314 : sel_789311;
  assign add_789318 = sel_789315 + 8'h01;
  assign sel_789319 = array_index_789110 == array_index_772948 ? add_789318 : sel_789315;
  assign add_789322 = sel_789319 + 8'h01;
  assign sel_789323 = array_index_789110 == array_index_772954 ? add_789322 : sel_789319;
  assign add_789326 = sel_789323 + 8'h01;
  assign sel_789327 = array_index_789110 == array_index_772960 ? add_789326 : sel_789323;
  assign add_789330 = sel_789327 + 8'h01;
  assign sel_789331 = array_index_789110 == array_index_772966 ? add_789330 : sel_789327;
  assign add_789334 = sel_789331 + 8'h01;
  assign sel_789335 = array_index_789110 == array_index_772972 ? add_789334 : sel_789331;
  assign add_789338 = sel_789335 + 8'h01;
  assign sel_789339 = array_index_789110 == array_index_772978 ? add_789338 : sel_789335;
  assign add_789342 = sel_789339 + 8'h01;
  assign sel_789343 = array_index_789110 == array_index_772984 ? add_789342 : sel_789339;
  assign add_789346 = sel_789343 + 8'h01;
  assign sel_789347 = array_index_789110 == array_index_772990 ? add_789346 : sel_789343;
  assign add_789350 = sel_789347 + 8'h01;
  assign sel_789351 = array_index_789110 == array_index_772996 ? add_789350 : sel_789347;
  assign add_789354 = sel_789351 + 8'h01;
  assign sel_789355 = array_index_789110 == array_index_773002 ? add_789354 : sel_789351;
  assign add_789358 = sel_789355 + 8'h01;
  assign sel_789359 = array_index_789110 == array_index_773008 ? add_789358 : sel_789355;
  assign add_789362 = sel_789359 + 8'h01;
  assign sel_789363 = array_index_789110 == array_index_773014 ? add_789362 : sel_789359;
  assign add_789366 = sel_789363 + 8'h01;
  assign sel_789367 = array_index_789110 == array_index_773020 ? add_789366 : sel_789363;
  assign add_789370 = sel_789367 + 8'h01;
  assign sel_789371 = array_index_789110 == array_index_773026 ? add_789370 : sel_789367;
  assign add_789374 = sel_789371 + 8'h01;
  assign sel_789375 = array_index_789110 == array_index_773032 ? add_789374 : sel_789371;
  assign add_789378 = sel_789375 + 8'h01;
  assign sel_789379 = array_index_789110 == array_index_773038 ? add_789378 : sel_789375;
  assign add_789382 = sel_789379 + 8'h01;
  assign sel_789383 = array_index_789110 == array_index_773044 ? add_789382 : sel_789379;
  assign add_789386 = sel_789383 + 8'h01;
  assign sel_789387 = array_index_789110 == array_index_773050 ? add_789386 : sel_789383;
  assign add_789390 = sel_789387 + 8'h01;
  assign sel_789391 = array_index_789110 == array_index_773056 ? add_789390 : sel_789387;
  assign add_789394 = sel_789391 + 8'h01;
  assign sel_789395 = array_index_789110 == array_index_773062 ? add_789394 : sel_789391;
  assign add_789398 = sel_789395 + 8'h01;
  assign sel_789399 = array_index_789110 == array_index_773068 ? add_789398 : sel_789395;
  assign add_789402 = sel_789399 + 8'h01;
  assign sel_789403 = array_index_789110 == array_index_773074 ? add_789402 : sel_789399;
  assign add_789406 = sel_789403 + 8'h01;
  assign sel_789407 = array_index_789110 == array_index_773080 ? add_789406 : sel_789403;
  assign add_789410 = sel_789407 + 8'h01;
  assign sel_789411 = array_index_789110 == array_index_773086 ? add_789410 : sel_789407;
  assign add_789414 = sel_789411 + 8'h01;
  assign sel_789415 = array_index_789110 == array_index_773092 ? add_789414 : sel_789411;
  assign add_789418 = sel_789415 + 8'h01;
  assign sel_789419 = array_index_789110 == array_index_773098 ? add_789418 : sel_789415;
  assign add_789422 = sel_789419 + 8'h01;
  assign sel_789423 = array_index_789110 == array_index_773104 ? add_789422 : sel_789419;
  assign add_789426 = sel_789423 + 8'h01;
  assign sel_789427 = array_index_789110 == array_index_773110 ? add_789426 : sel_789423;
  assign add_789430 = sel_789427 + 8'h01;
  assign sel_789431 = array_index_789110 == array_index_773116 ? add_789430 : sel_789427;
  assign add_789434 = sel_789431 + 8'h01;
  assign sel_789435 = array_index_789110 == array_index_773122 ? add_789434 : sel_789431;
  assign add_789438 = sel_789435 + 8'h01;
  assign sel_789439 = array_index_789110 == array_index_773128 ? add_789438 : sel_789435;
  assign add_789442 = sel_789439 + 8'h01;
  assign sel_789443 = array_index_789110 == array_index_773134 ? add_789442 : sel_789439;
  assign add_789446 = sel_789443 + 8'h01;
  assign sel_789447 = array_index_789110 == array_index_773140 ? add_789446 : sel_789443;
  assign add_789450 = sel_789447 + 8'h01;
  assign sel_789451 = array_index_789110 == array_index_773146 ? add_789450 : sel_789447;
  assign add_789454 = sel_789451 + 8'h01;
  assign sel_789455 = array_index_789110 == array_index_773152 ? add_789454 : sel_789451;
  assign add_789458 = sel_789455 + 8'h01;
  assign sel_789459 = array_index_789110 == array_index_773158 ? add_789458 : sel_789455;
  assign add_789462 = sel_789459 + 8'h01;
  assign sel_789463 = array_index_789110 == array_index_773164 ? add_789462 : sel_789459;
  assign add_789466 = sel_789463 + 8'h01;
  assign sel_789467 = array_index_789110 == array_index_773170 ? add_789466 : sel_789463;
  assign add_789471 = sel_789467 + 8'h01;
  assign array_index_789472 = set1_unflattened[7'h2e];
  assign sel_789473 = array_index_789110 == array_index_773176 ? add_789471 : sel_789467;
  assign add_789476 = sel_789473 + 8'h01;
  assign sel_789477 = array_index_789472 == array_index_772632 ? add_789476 : sel_789473;
  assign add_789480 = sel_789477 + 8'h01;
  assign sel_789481 = array_index_789472 == array_index_772636 ? add_789480 : sel_789477;
  assign add_789484 = sel_789481 + 8'h01;
  assign sel_789485 = array_index_789472 == array_index_772644 ? add_789484 : sel_789481;
  assign add_789488 = sel_789485 + 8'h01;
  assign sel_789489 = array_index_789472 == array_index_772652 ? add_789488 : sel_789485;
  assign add_789492 = sel_789489 + 8'h01;
  assign sel_789493 = array_index_789472 == array_index_772660 ? add_789492 : sel_789489;
  assign add_789496 = sel_789493 + 8'h01;
  assign sel_789497 = array_index_789472 == array_index_772668 ? add_789496 : sel_789493;
  assign add_789500 = sel_789497 + 8'h01;
  assign sel_789501 = array_index_789472 == array_index_772676 ? add_789500 : sel_789497;
  assign add_789504 = sel_789501 + 8'h01;
  assign sel_789505 = array_index_789472 == array_index_772684 ? add_789504 : sel_789501;
  assign add_789508 = sel_789505 + 8'h01;
  assign sel_789509 = array_index_789472 == array_index_772690 ? add_789508 : sel_789505;
  assign add_789512 = sel_789509 + 8'h01;
  assign sel_789513 = array_index_789472 == array_index_772696 ? add_789512 : sel_789509;
  assign add_789516 = sel_789513 + 8'h01;
  assign sel_789517 = array_index_789472 == array_index_772702 ? add_789516 : sel_789513;
  assign add_789520 = sel_789517 + 8'h01;
  assign sel_789521 = array_index_789472 == array_index_772708 ? add_789520 : sel_789517;
  assign add_789524 = sel_789521 + 8'h01;
  assign sel_789525 = array_index_789472 == array_index_772714 ? add_789524 : sel_789521;
  assign add_789528 = sel_789525 + 8'h01;
  assign sel_789529 = array_index_789472 == array_index_772720 ? add_789528 : sel_789525;
  assign add_789532 = sel_789529 + 8'h01;
  assign sel_789533 = array_index_789472 == array_index_772726 ? add_789532 : sel_789529;
  assign add_789536 = sel_789533 + 8'h01;
  assign sel_789537 = array_index_789472 == array_index_772732 ? add_789536 : sel_789533;
  assign add_789540 = sel_789537 + 8'h01;
  assign sel_789541 = array_index_789472 == array_index_772738 ? add_789540 : sel_789537;
  assign add_789544 = sel_789541 + 8'h01;
  assign sel_789545 = array_index_789472 == array_index_772744 ? add_789544 : sel_789541;
  assign add_789548 = sel_789545 + 8'h01;
  assign sel_789549 = array_index_789472 == array_index_772750 ? add_789548 : sel_789545;
  assign add_789552 = sel_789549 + 8'h01;
  assign sel_789553 = array_index_789472 == array_index_772756 ? add_789552 : sel_789549;
  assign add_789556 = sel_789553 + 8'h01;
  assign sel_789557 = array_index_789472 == array_index_772762 ? add_789556 : sel_789553;
  assign add_789560 = sel_789557 + 8'h01;
  assign sel_789561 = array_index_789472 == array_index_772768 ? add_789560 : sel_789557;
  assign add_789564 = sel_789561 + 8'h01;
  assign sel_789565 = array_index_789472 == array_index_772774 ? add_789564 : sel_789561;
  assign add_789568 = sel_789565 + 8'h01;
  assign sel_789569 = array_index_789472 == array_index_772780 ? add_789568 : sel_789565;
  assign add_789572 = sel_789569 + 8'h01;
  assign sel_789573 = array_index_789472 == array_index_772786 ? add_789572 : sel_789569;
  assign add_789576 = sel_789573 + 8'h01;
  assign sel_789577 = array_index_789472 == array_index_772792 ? add_789576 : sel_789573;
  assign add_789580 = sel_789577 + 8'h01;
  assign sel_789581 = array_index_789472 == array_index_772798 ? add_789580 : sel_789577;
  assign add_789584 = sel_789581 + 8'h01;
  assign sel_789585 = array_index_789472 == array_index_772804 ? add_789584 : sel_789581;
  assign add_789588 = sel_789585 + 8'h01;
  assign sel_789589 = array_index_789472 == array_index_772810 ? add_789588 : sel_789585;
  assign add_789592 = sel_789589 + 8'h01;
  assign sel_789593 = array_index_789472 == array_index_772816 ? add_789592 : sel_789589;
  assign add_789596 = sel_789593 + 8'h01;
  assign sel_789597 = array_index_789472 == array_index_772822 ? add_789596 : sel_789593;
  assign add_789600 = sel_789597 + 8'h01;
  assign sel_789601 = array_index_789472 == array_index_772828 ? add_789600 : sel_789597;
  assign add_789604 = sel_789601 + 8'h01;
  assign sel_789605 = array_index_789472 == array_index_772834 ? add_789604 : sel_789601;
  assign add_789608 = sel_789605 + 8'h01;
  assign sel_789609 = array_index_789472 == array_index_772840 ? add_789608 : sel_789605;
  assign add_789612 = sel_789609 + 8'h01;
  assign sel_789613 = array_index_789472 == array_index_772846 ? add_789612 : sel_789609;
  assign add_789616 = sel_789613 + 8'h01;
  assign sel_789617 = array_index_789472 == array_index_772852 ? add_789616 : sel_789613;
  assign add_789620 = sel_789617 + 8'h01;
  assign sel_789621 = array_index_789472 == array_index_772858 ? add_789620 : sel_789617;
  assign add_789624 = sel_789621 + 8'h01;
  assign sel_789625 = array_index_789472 == array_index_772864 ? add_789624 : sel_789621;
  assign add_789628 = sel_789625 + 8'h01;
  assign sel_789629 = array_index_789472 == array_index_772870 ? add_789628 : sel_789625;
  assign add_789632 = sel_789629 + 8'h01;
  assign sel_789633 = array_index_789472 == array_index_772876 ? add_789632 : sel_789629;
  assign add_789636 = sel_789633 + 8'h01;
  assign sel_789637 = array_index_789472 == array_index_772882 ? add_789636 : sel_789633;
  assign add_789640 = sel_789637 + 8'h01;
  assign sel_789641 = array_index_789472 == array_index_772888 ? add_789640 : sel_789637;
  assign add_789644 = sel_789641 + 8'h01;
  assign sel_789645 = array_index_789472 == array_index_772894 ? add_789644 : sel_789641;
  assign add_789648 = sel_789645 + 8'h01;
  assign sel_789649 = array_index_789472 == array_index_772900 ? add_789648 : sel_789645;
  assign add_789652 = sel_789649 + 8'h01;
  assign sel_789653 = array_index_789472 == array_index_772906 ? add_789652 : sel_789649;
  assign add_789656 = sel_789653 + 8'h01;
  assign sel_789657 = array_index_789472 == array_index_772912 ? add_789656 : sel_789653;
  assign add_789660 = sel_789657 + 8'h01;
  assign sel_789661 = array_index_789472 == array_index_772918 ? add_789660 : sel_789657;
  assign add_789664 = sel_789661 + 8'h01;
  assign sel_789665 = array_index_789472 == array_index_772924 ? add_789664 : sel_789661;
  assign add_789668 = sel_789665 + 8'h01;
  assign sel_789669 = array_index_789472 == array_index_772930 ? add_789668 : sel_789665;
  assign add_789672 = sel_789669 + 8'h01;
  assign sel_789673 = array_index_789472 == array_index_772936 ? add_789672 : sel_789669;
  assign add_789676 = sel_789673 + 8'h01;
  assign sel_789677 = array_index_789472 == array_index_772942 ? add_789676 : sel_789673;
  assign add_789680 = sel_789677 + 8'h01;
  assign sel_789681 = array_index_789472 == array_index_772948 ? add_789680 : sel_789677;
  assign add_789684 = sel_789681 + 8'h01;
  assign sel_789685 = array_index_789472 == array_index_772954 ? add_789684 : sel_789681;
  assign add_789688 = sel_789685 + 8'h01;
  assign sel_789689 = array_index_789472 == array_index_772960 ? add_789688 : sel_789685;
  assign add_789692 = sel_789689 + 8'h01;
  assign sel_789693 = array_index_789472 == array_index_772966 ? add_789692 : sel_789689;
  assign add_789696 = sel_789693 + 8'h01;
  assign sel_789697 = array_index_789472 == array_index_772972 ? add_789696 : sel_789693;
  assign add_789700 = sel_789697 + 8'h01;
  assign sel_789701 = array_index_789472 == array_index_772978 ? add_789700 : sel_789697;
  assign add_789704 = sel_789701 + 8'h01;
  assign sel_789705 = array_index_789472 == array_index_772984 ? add_789704 : sel_789701;
  assign add_789708 = sel_789705 + 8'h01;
  assign sel_789709 = array_index_789472 == array_index_772990 ? add_789708 : sel_789705;
  assign add_789712 = sel_789709 + 8'h01;
  assign sel_789713 = array_index_789472 == array_index_772996 ? add_789712 : sel_789709;
  assign add_789716 = sel_789713 + 8'h01;
  assign sel_789717 = array_index_789472 == array_index_773002 ? add_789716 : sel_789713;
  assign add_789720 = sel_789717 + 8'h01;
  assign sel_789721 = array_index_789472 == array_index_773008 ? add_789720 : sel_789717;
  assign add_789724 = sel_789721 + 8'h01;
  assign sel_789725 = array_index_789472 == array_index_773014 ? add_789724 : sel_789721;
  assign add_789728 = sel_789725 + 8'h01;
  assign sel_789729 = array_index_789472 == array_index_773020 ? add_789728 : sel_789725;
  assign add_789732 = sel_789729 + 8'h01;
  assign sel_789733 = array_index_789472 == array_index_773026 ? add_789732 : sel_789729;
  assign add_789736 = sel_789733 + 8'h01;
  assign sel_789737 = array_index_789472 == array_index_773032 ? add_789736 : sel_789733;
  assign add_789740 = sel_789737 + 8'h01;
  assign sel_789741 = array_index_789472 == array_index_773038 ? add_789740 : sel_789737;
  assign add_789744 = sel_789741 + 8'h01;
  assign sel_789745 = array_index_789472 == array_index_773044 ? add_789744 : sel_789741;
  assign add_789748 = sel_789745 + 8'h01;
  assign sel_789749 = array_index_789472 == array_index_773050 ? add_789748 : sel_789745;
  assign add_789752 = sel_789749 + 8'h01;
  assign sel_789753 = array_index_789472 == array_index_773056 ? add_789752 : sel_789749;
  assign add_789756 = sel_789753 + 8'h01;
  assign sel_789757 = array_index_789472 == array_index_773062 ? add_789756 : sel_789753;
  assign add_789760 = sel_789757 + 8'h01;
  assign sel_789761 = array_index_789472 == array_index_773068 ? add_789760 : sel_789757;
  assign add_789764 = sel_789761 + 8'h01;
  assign sel_789765 = array_index_789472 == array_index_773074 ? add_789764 : sel_789761;
  assign add_789768 = sel_789765 + 8'h01;
  assign sel_789769 = array_index_789472 == array_index_773080 ? add_789768 : sel_789765;
  assign add_789772 = sel_789769 + 8'h01;
  assign sel_789773 = array_index_789472 == array_index_773086 ? add_789772 : sel_789769;
  assign add_789776 = sel_789773 + 8'h01;
  assign sel_789777 = array_index_789472 == array_index_773092 ? add_789776 : sel_789773;
  assign add_789780 = sel_789777 + 8'h01;
  assign sel_789781 = array_index_789472 == array_index_773098 ? add_789780 : sel_789777;
  assign add_789784 = sel_789781 + 8'h01;
  assign sel_789785 = array_index_789472 == array_index_773104 ? add_789784 : sel_789781;
  assign add_789788 = sel_789785 + 8'h01;
  assign sel_789789 = array_index_789472 == array_index_773110 ? add_789788 : sel_789785;
  assign add_789792 = sel_789789 + 8'h01;
  assign sel_789793 = array_index_789472 == array_index_773116 ? add_789792 : sel_789789;
  assign add_789796 = sel_789793 + 8'h01;
  assign sel_789797 = array_index_789472 == array_index_773122 ? add_789796 : sel_789793;
  assign add_789800 = sel_789797 + 8'h01;
  assign sel_789801 = array_index_789472 == array_index_773128 ? add_789800 : sel_789797;
  assign add_789804 = sel_789801 + 8'h01;
  assign sel_789805 = array_index_789472 == array_index_773134 ? add_789804 : sel_789801;
  assign add_789808 = sel_789805 + 8'h01;
  assign sel_789809 = array_index_789472 == array_index_773140 ? add_789808 : sel_789805;
  assign add_789812 = sel_789809 + 8'h01;
  assign sel_789813 = array_index_789472 == array_index_773146 ? add_789812 : sel_789809;
  assign add_789816 = sel_789813 + 8'h01;
  assign sel_789817 = array_index_789472 == array_index_773152 ? add_789816 : sel_789813;
  assign add_789820 = sel_789817 + 8'h01;
  assign sel_789821 = array_index_789472 == array_index_773158 ? add_789820 : sel_789817;
  assign add_789824 = sel_789821 + 8'h01;
  assign sel_789825 = array_index_789472 == array_index_773164 ? add_789824 : sel_789821;
  assign add_789828 = sel_789825 + 8'h01;
  assign sel_789829 = array_index_789472 == array_index_773170 ? add_789828 : sel_789825;
  assign add_789833 = sel_789829 + 8'h01;
  assign array_index_789834 = set1_unflattened[7'h2f];
  assign sel_789835 = array_index_789472 == array_index_773176 ? add_789833 : sel_789829;
  assign add_789838 = sel_789835 + 8'h01;
  assign sel_789839 = array_index_789834 == array_index_772632 ? add_789838 : sel_789835;
  assign add_789842 = sel_789839 + 8'h01;
  assign sel_789843 = array_index_789834 == array_index_772636 ? add_789842 : sel_789839;
  assign add_789846 = sel_789843 + 8'h01;
  assign sel_789847 = array_index_789834 == array_index_772644 ? add_789846 : sel_789843;
  assign add_789850 = sel_789847 + 8'h01;
  assign sel_789851 = array_index_789834 == array_index_772652 ? add_789850 : sel_789847;
  assign add_789854 = sel_789851 + 8'h01;
  assign sel_789855 = array_index_789834 == array_index_772660 ? add_789854 : sel_789851;
  assign add_789858 = sel_789855 + 8'h01;
  assign sel_789859 = array_index_789834 == array_index_772668 ? add_789858 : sel_789855;
  assign add_789862 = sel_789859 + 8'h01;
  assign sel_789863 = array_index_789834 == array_index_772676 ? add_789862 : sel_789859;
  assign add_789866 = sel_789863 + 8'h01;
  assign sel_789867 = array_index_789834 == array_index_772684 ? add_789866 : sel_789863;
  assign add_789870 = sel_789867 + 8'h01;
  assign sel_789871 = array_index_789834 == array_index_772690 ? add_789870 : sel_789867;
  assign add_789874 = sel_789871 + 8'h01;
  assign sel_789875 = array_index_789834 == array_index_772696 ? add_789874 : sel_789871;
  assign add_789878 = sel_789875 + 8'h01;
  assign sel_789879 = array_index_789834 == array_index_772702 ? add_789878 : sel_789875;
  assign add_789882 = sel_789879 + 8'h01;
  assign sel_789883 = array_index_789834 == array_index_772708 ? add_789882 : sel_789879;
  assign add_789886 = sel_789883 + 8'h01;
  assign sel_789887 = array_index_789834 == array_index_772714 ? add_789886 : sel_789883;
  assign add_789890 = sel_789887 + 8'h01;
  assign sel_789891 = array_index_789834 == array_index_772720 ? add_789890 : sel_789887;
  assign add_789894 = sel_789891 + 8'h01;
  assign sel_789895 = array_index_789834 == array_index_772726 ? add_789894 : sel_789891;
  assign add_789898 = sel_789895 + 8'h01;
  assign sel_789899 = array_index_789834 == array_index_772732 ? add_789898 : sel_789895;
  assign add_789902 = sel_789899 + 8'h01;
  assign sel_789903 = array_index_789834 == array_index_772738 ? add_789902 : sel_789899;
  assign add_789906 = sel_789903 + 8'h01;
  assign sel_789907 = array_index_789834 == array_index_772744 ? add_789906 : sel_789903;
  assign add_789910 = sel_789907 + 8'h01;
  assign sel_789911 = array_index_789834 == array_index_772750 ? add_789910 : sel_789907;
  assign add_789914 = sel_789911 + 8'h01;
  assign sel_789915 = array_index_789834 == array_index_772756 ? add_789914 : sel_789911;
  assign add_789918 = sel_789915 + 8'h01;
  assign sel_789919 = array_index_789834 == array_index_772762 ? add_789918 : sel_789915;
  assign add_789922 = sel_789919 + 8'h01;
  assign sel_789923 = array_index_789834 == array_index_772768 ? add_789922 : sel_789919;
  assign add_789926 = sel_789923 + 8'h01;
  assign sel_789927 = array_index_789834 == array_index_772774 ? add_789926 : sel_789923;
  assign add_789930 = sel_789927 + 8'h01;
  assign sel_789931 = array_index_789834 == array_index_772780 ? add_789930 : sel_789927;
  assign add_789934 = sel_789931 + 8'h01;
  assign sel_789935 = array_index_789834 == array_index_772786 ? add_789934 : sel_789931;
  assign add_789938 = sel_789935 + 8'h01;
  assign sel_789939 = array_index_789834 == array_index_772792 ? add_789938 : sel_789935;
  assign add_789942 = sel_789939 + 8'h01;
  assign sel_789943 = array_index_789834 == array_index_772798 ? add_789942 : sel_789939;
  assign add_789946 = sel_789943 + 8'h01;
  assign sel_789947 = array_index_789834 == array_index_772804 ? add_789946 : sel_789943;
  assign add_789950 = sel_789947 + 8'h01;
  assign sel_789951 = array_index_789834 == array_index_772810 ? add_789950 : sel_789947;
  assign add_789954 = sel_789951 + 8'h01;
  assign sel_789955 = array_index_789834 == array_index_772816 ? add_789954 : sel_789951;
  assign add_789958 = sel_789955 + 8'h01;
  assign sel_789959 = array_index_789834 == array_index_772822 ? add_789958 : sel_789955;
  assign add_789962 = sel_789959 + 8'h01;
  assign sel_789963 = array_index_789834 == array_index_772828 ? add_789962 : sel_789959;
  assign add_789966 = sel_789963 + 8'h01;
  assign sel_789967 = array_index_789834 == array_index_772834 ? add_789966 : sel_789963;
  assign add_789970 = sel_789967 + 8'h01;
  assign sel_789971 = array_index_789834 == array_index_772840 ? add_789970 : sel_789967;
  assign add_789974 = sel_789971 + 8'h01;
  assign sel_789975 = array_index_789834 == array_index_772846 ? add_789974 : sel_789971;
  assign add_789978 = sel_789975 + 8'h01;
  assign sel_789979 = array_index_789834 == array_index_772852 ? add_789978 : sel_789975;
  assign add_789982 = sel_789979 + 8'h01;
  assign sel_789983 = array_index_789834 == array_index_772858 ? add_789982 : sel_789979;
  assign add_789986 = sel_789983 + 8'h01;
  assign sel_789987 = array_index_789834 == array_index_772864 ? add_789986 : sel_789983;
  assign add_789990 = sel_789987 + 8'h01;
  assign sel_789991 = array_index_789834 == array_index_772870 ? add_789990 : sel_789987;
  assign add_789994 = sel_789991 + 8'h01;
  assign sel_789995 = array_index_789834 == array_index_772876 ? add_789994 : sel_789991;
  assign add_789998 = sel_789995 + 8'h01;
  assign sel_789999 = array_index_789834 == array_index_772882 ? add_789998 : sel_789995;
  assign add_790002 = sel_789999 + 8'h01;
  assign sel_790003 = array_index_789834 == array_index_772888 ? add_790002 : sel_789999;
  assign add_790006 = sel_790003 + 8'h01;
  assign sel_790007 = array_index_789834 == array_index_772894 ? add_790006 : sel_790003;
  assign add_790010 = sel_790007 + 8'h01;
  assign sel_790011 = array_index_789834 == array_index_772900 ? add_790010 : sel_790007;
  assign add_790014 = sel_790011 + 8'h01;
  assign sel_790015 = array_index_789834 == array_index_772906 ? add_790014 : sel_790011;
  assign add_790018 = sel_790015 + 8'h01;
  assign sel_790019 = array_index_789834 == array_index_772912 ? add_790018 : sel_790015;
  assign add_790022 = sel_790019 + 8'h01;
  assign sel_790023 = array_index_789834 == array_index_772918 ? add_790022 : sel_790019;
  assign add_790026 = sel_790023 + 8'h01;
  assign sel_790027 = array_index_789834 == array_index_772924 ? add_790026 : sel_790023;
  assign add_790030 = sel_790027 + 8'h01;
  assign sel_790031 = array_index_789834 == array_index_772930 ? add_790030 : sel_790027;
  assign add_790034 = sel_790031 + 8'h01;
  assign sel_790035 = array_index_789834 == array_index_772936 ? add_790034 : sel_790031;
  assign add_790038 = sel_790035 + 8'h01;
  assign sel_790039 = array_index_789834 == array_index_772942 ? add_790038 : sel_790035;
  assign add_790042 = sel_790039 + 8'h01;
  assign sel_790043 = array_index_789834 == array_index_772948 ? add_790042 : sel_790039;
  assign add_790046 = sel_790043 + 8'h01;
  assign sel_790047 = array_index_789834 == array_index_772954 ? add_790046 : sel_790043;
  assign add_790050 = sel_790047 + 8'h01;
  assign sel_790051 = array_index_789834 == array_index_772960 ? add_790050 : sel_790047;
  assign add_790054 = sel_790051 + 8'h01;
  assign sel_790055 = array_index_789834 == array_index_772966 ? add_790054 : sel_790051;
  assign add_790058 = sel_790055 + 8'h01;
  assign sel_790059 = array_index_789834 == array_index_772972 ? add_790058 : sel_790055;
  assign add_790062 = sel_790059 + 8'h01;
  assign sel_790063 = array_index_789834 == array_index_772978 ? add_790062 : sel_790059;
  assign add_790066 = sel_790063 + 8'h01;
  assign sel_790067 = array_index_789834 == array_index_772984 ? add_790066 : sel_790063;
  assign add_790070 = sel_790067 + 8'h01;
  assign sel_790071 = array_index_789834 == array_index_772990 ? add_790070 : sel_790067;
  assign add_790074 = sel_790071 + 8'h01;
  assign sel_790075 = array_index_789834 == array_index_772996 ? add_790074 : sel_790071;
  assign add_790078 = sel_790075 + 8'h01;
  assign sel_790079 = array_index_789834 == array_index_773002 ? add_790078 : sel_790075;
  assign add_790082 = sel_790079 + 8'h01;
  assign sel_790083 = array_index_789834 == array_index_773008 ? add_790082 : sel_790079;
  assign add_790086 = sel_790083 + 8'h01;
  assign sel_790087 = array_index_789834 == array_index_773014 ? add_790086 : sel_790083;
  assign add_790090 = sel_790087 + 8'h01;
  assign sel_790091 = array_index_789834 == array_index_773020 ? add_790090 : sel_790087;
  assign add_790094 = sel_790091 + 8'h01;
  assign sel_790095 = array_index_789834 == array_index_773026 ? add_790094 : sel_790091;
  assign add_790098 = sel_790095 + 8'h01;
  assign sel_790099 = array_index_789834 == array_index_773032 ? add_790098 : sel_790095;
  assign add_790102 = sel_790099 + 8'h01;
  assign sel_790103 = array_index_789834 == array_index_773038 ? add_790102 : sel_790099;
  assign add_790106 = sel_790103 + 8'h01;
  assign sel_790107 = array_index_789834 == array_index_773044 ? add_790106 : sel_790103;
  assign add_790110 = sel_790107 + 8'h01;
  assign sel_790111 = array_index_789834 == array_index_773050 ? add_790110 : sel_790107;
  assign add_790114 = sel_790111 + 8'h01;
  assign sel_790115 = array_index_789834 == array_index_773056 ? add_790114 : sel_790111;
  assign add_790118 = sel_790115 + 8'h01;
  assign sel_790119 = array_index_789834 == array_index_773062 ? add_790118 : sel_790115;
  assign add_790122 = sel_790119 + 8'h01;
  assign sel_790123 = array_index_789834 == array_index_773068 ? add_790122 : sel_790119;
  assign add_790126 = sel_790123 + 8'h01;
  assign sel_790127 = array_index_789834 == array_index_773074 ? add_790126 : sel_790123;
  assign add_790130 = sel_790127 + 8'h01;
  assign sel_790131 = array_index_789834 == array_index_773080 ? add_790130 : sel_790127;
  assign add_790134 = sel_790131 + 8'h01;
  assign sel_790135 = array_index_789834 == array_index_773086 ? add_790134 : sel_790131;
  assign add_790138 = sel_790135 + 8'h01;
  assign sel_790139 = array_index_789834 == array_index_773092 ? add_790138 : sel_790135;
  assign add_790142 = sel_790139 + 8'h01;
  assign sel_790143 = array_index_789834 == array_index_773098 ? add_790142 : sel_790139;
  assign add_790146 = sel_790143 + 8'h01;
  assign sel_790147 = array_index_789834 == array_index_773104 ? add_790146 : sel_790143;
  assign add_790150 = sel_790147 + 8'h01;
  assign sel_790151 = array_index_789834 == array_index_773110 ? add_790150 : sel_790147;
  assign add_790154 = sel_790151 + 8'h01;
  assign sel_790155 = array_index_789834 == array_index_773116 ? add_790154 : sel_790151;
  assign add_790158 = sel_790155 + 8'h01;
  assign sel_790159 = array_index_789834 == array_index_773122 ? add_790158 : sel_790155;
  assign add_790162 = sel_790159 + 8'h01;
  assign sel_790163 = array_index_789834 == array_index_773128 ? add_790162 : sel_790159;
  assign add_790166 = sel_790163 + 8'h01;
  assign sel_790167 = array_index_789834 == array_index_773134 ? add_790166 : sel_790163;
  assign add_790170 = sel_790167 + 8'h01;
  assign sel_790171 = array_index_789834 == array_index_773140 ? add_790170 : sel_790167;
  assign add_790174 = sel_790171 + 8'h01;
  assign sel_790175 = array_index_789834 == array_index_773146 ? add_790174 : sel_790171;
  assign add_790178 = sel_790175 + 8'h01;
  assign sel_790179 = array_index_789834 == array_index_773152 ? add_790178 : sel_790175;
  assign add_790182 = sel_790179 + 8'h01;
  assign sel_790183 = array_index_789834 == array_index_773158 ? add_790182 : sel_790179;
  assign add_790186 = sel_790183 + 8'h01;
  assign sel_790187 = array_index_789834 == array_index_773164 ? add_790186 : sel_790183;
  assign add_790190 = sel_790187 + 8'h01;
  assign sel_790191 = array_index_789834 == array_index_773170 ? add_790190 : sel_790187;
  assign add_790195 = sel_790191 + 8'h01;
  assign array_index_790196 = set1_unflattened[7'h30];
  assign sel_790197 = array_index_789834 == array_index_773176 ? add_790195 : sel_790191;
  assign add_790200 = sel_790197 + 8'h01;
  assign sel_790201 = array_index_790196 == array_index_772632 ? add_790200 : sel_790197;
  assign add_790204 = sel_790201 + 8'h01;
  assign sel_790205 = array_index_790196 == array_index_772636 ? add_790204 : sel_790201;
  assign add_790208 = sel_790205 + 8'h01;
  assign sel_790209 = array_index_790196 == array_index_772644 ? add_790208 : sel_790205;
  assign add_790212 = sel_790209 + 8'h01;
  assign sel_790213 = array_index_790196 == array_index_772652 ? add_790212 : sel_790209;
  assign add_790216 = sel_790213 + 8'h01;
  assign sel_790217 = array_index_790196 == array_index_772660 ? add_790216 : sel_790213;
  assign add_790220 = sel_790217 + 8'h01;
  assign sel_790221 = array_index_790196 == array_index_772668 ? add_790220 : sel_790217;
  assign add_790224 = sel_790221 + 8'h01;
  assign sel_790225 = array_index_790196 == array_index_772676 ? add_790224 : sel_790221;
  assign add_790228 = sel_790225 + 8'h01;
  assign sel_790229 = array_index_790196 == array_index_772684 ? add_790228 : sel_790225;
  assign add_790232 = sel_790229 + 8'h01;
  assign sel_790233 = array_index_790196 == array_index_772690 ? add_790232 : sel_790229;
  assign add_790236 = sel_790233 + 8'h01;
  assign sel_790237 = array_index_790196 == array_index_772696 ? add_790236 : sel_790233;
  assign add_790240 = sel_790237 + 8'h01;
  assign sel_790241 = array_index_790196 == array_index_772702 ? add_790240 : sel_790237;
  assign add_790244 = sel_790241 + 8'h01;
  assign sel_790245 = array_index_790196 == array_index_772708 ? add_790244 : sel_790241;
  assign add_790248 = sel_790245 + 8'h01;
  assign sel_790249 = array_index_790196 == array_index_772714 ? add_790248 : sel_790245;
  assign add_790252 = sel_790249 + 8'h01;
  assign sel_790253 = array_index_790196 == array_index_772720 ? add_790252 : sel_790249;
  assign add_790256 = sel_790253 + 8'h01;
  assign sel_790257 = array_index_790196 == array_index_772726 ? add_790256 : sel_790253;
  assign add_790260 = sel_790257 + 8'h01;
  assign sel_790261 = array_index_790196 == array_index_772732 ? add_790260 : sel_790257;
  assign add_790264 = sel_790261 + 8'h01;
  assign sel_790265 = array_index_790196 == array_index_772738 ? add_790264 : sel_790261;
  assign add_790268 = sel_790265 + 8'h01;
  assign sel_790269 = array_index_790196 == array_index_772744 ? add_790268 : sel_790265;
  assign add_790272 = sel_790269 + 8'h01;
  assign sel_790273 = array_index_790196 == array_index_772750 ? add_790272 : sel_790269;
  assign add_790276 = sel_790273 + 8'h01;
  assign sel_790277 = array_index_790196 == array_index_772756 ? add_790276 : sel_790273;
  assign add_790280 = sel_790277 + 8'h01;
  assign sel_790281 = array_index_790196 == array_index_772762 ? add_790280 : sel_790277;
  assign add_790284 = sel_790281 + 8'h01;
  assign sel_790285 = array_index_790196 == array_index_772768 ? add_790284 : sel_790281;
  assign add_790288 = sel_790285 + 8'h01;
  assign sel_790289 = array_index_790196 == array_index_772774 ? add_790288 : sel_790285;
  assign add_790292 = sel_790289 + 8'h01;
  assign sel_790293 = array_index_790196 == array_index_772780 ? add_790292 : sel_790289;
  assign add_790296 = sel_790293 + 8'h01;
  assign sel_790297 = array_index_790196 == array_index_772786 ? add_790296 : sel_790293;
  assign add_790300 = sel_790297 + 8'h01;
  assign sel_790301 = array_index_790196 == array_index_772792 ? add_790300 : sel_790297;
  assign add_790304 = sel_790301 + 8'h01;
  assign sel_790305 = array_index_790196 == array_index_772798 ? add_790304 : sel_790301;
  assign add_790308 = sel_790305 + 8'h01;
  assign sel_790309 = array_index_790196 == array_index_772804 ? add_790308 : sel_790305;
  assign add_790312 = sel_790309 + 8'h01;
  assign sel_790313 = array_index_790196 == array_index_772810 ? add_790312 : sel_790309;
  assign add_790316 = sel_790313 + 8'h01;
  assign sel_790317 = array_index_790196 == array_index_772816 ? add_790316 : sel_790313;
  assign add_790320 = sel_790317 + 8'h01;
  assign sel_790321 = array_index_790196 == array_index_772822 ? add_790320 : sel_790317;
  assign add_790324 = sel_790321 + 8'h01;
  assign sel_790325 = array_index_790196 == array_index_772828 ? add_790324 : sel_790321;
  assign add_790328 = sel_790325 + 8'h01;
  assign sel_790329 = array_index_790196 == array_index_772834 ? add_790328 : sel_790325;
  assign add_790332 = sel_790329 + 8'h01;
  assign sel_790333 = array_index_790196 == array_index_772840 ? add_790332 : sel_790329;
  assign add_790336 = sel_790333 + 8'h01;
  assign sel_790337 = array_index_790196 == array_index_772846 ? add_790336 : sel_790333;
  assign add_790340 = sel_790337 + 8'h01;
  assign sel_790341 = array_index_790196 == array_index_772852 ? add_790340 : sel_790337;
  assign add_790344 = sel_790341 + 8'h01;
  assign sel_790345 = array_index_790196 == array_index_772858 ? add_790344 : sel_790341;
  assign add_790348 = sel_790345 + 8'h01;
  assign sel_790349 = array_index_790196 == array_index_772864 ? add_790348 : sel_790345;
  assign add_790352 = sel_790349 + 8'h01;
  assign sel_790353 = array_index_790196 == array_index_772870 ? add_790352 : sel_790349;
  assign add_790356 = sel_790353 + 8'h01;
  assign sel_790357 = array_index_790196 == array_index_772876 ? add_790356 : sel_790353;
  assign add_790360 = sel_790357 + 8'h01;
  assign sel_790361 = array_index_790196 == array_index_772882 ? add_790360 : sel_790357;
  assign add_790364 = sel_790361 + 8'h01;
  assign sel_790365 = array_index_790196 == array_index_772888 ? add_790364 : sel_790361;
  assign add_790368 = sel_790365 + 8'h01;
  assign sel_790369 = array_index_790196 == array_index_772894 ? add_790368 : sel_790365;
  assign add_790372 = sel_790369 + 8'h01;
  assign sel_790373 = array_index_790196 == array_index_772900 ? add_790372 : sel_790369;
  assign add_790376 = sel_790373 + 8'h01;
  assign sel_790377 = array_index_790196 == array_index_772906 ? add_790376 : sel_790373;
  assign add_790380 = sel_790377 + 8'h01;
  assign sel_790381 = array_index_790196 == array_index_772912 ? add_790380 : sel_790377;
  assign add_790384 = sel_790381 + 8'h01;
  assign sel_790385 = array_index_790196 == array_index_772918 ? add_790384 : sel_790381;
  assign add_790388 = sel_790385 + 8'h01;
  assign sel_790389 = array_index_790196 == array_index_772924 ? add_790388 : sel_790385;
  assign add_790392 = sel_790389 + 8'h01;
  assign sel_790393 = array_index_790196 == array_index_772930 ? add_790392 : sel_790389;
  assign add_790396 = sel_790393 + 8'h01;
  assign sel_790397 = array_index_790196 == array_index_772936 ? add_790396 : sel_790393;
  assign add_790400 = sel_790397 + 8'h01;
  assign sel_790401 = array_index_790196 == array_index_772942 ? add_790400 : sel_790397;
  assign add_790404 = sel_790401 + 8'h01;
  assign sel_790405 = array_index_790196 == array_index_772948 ? add_790404 : sel_790401;
  assign add_790408 = sel_790405 + 8'h01;
  assign sel_790409 = array_index_790196 == array_index_772954 ? add_790408 : sel_790405;
  assign add_790412 = sel_790409 + 8'h01;
  assign sel_790413 = array_index_790196 == array_index_772960 ? add_790412 : sel_790409;
  assign add_790416 = sel_790413 + 8'h01;
  assign sel_790417 = array_index_790196 == array_index_772966 ? add_790416 : sel_790413;
  assign add_790420 = sel_790417 + 8'h01;
  assign sel_790421 = array_index_790196 == array_index_772972 ? add_790420 : sel_790417;
  assign add_790424 = sel_790421 + 8'h01;
  assign sel_790425 = array_index_790196 == array_index_772978 ? add_790424 : sel_790421;
  assign add_790428 = sel_790425 + 8'h01;
  assign sel_790429 = array_index_790196 == array_index_772984 ? add_790428 : sel_790425;
  assign add_790432 = sel_790429 + 8'h01;
  assign sel_790433 = array_index_790196 == array_index_772990 ? add_790432 : sel_790429;
  assign add_790436 = sel_790433 + 8'h01;
  assign sel_790437 = array_index_790196 == array_index_772996 ? add_790436 : sel_790433;
  assign add_790440 = sel_790437 + 8'h01;
  assign sel_790441 = array_index_790196 == array_index_773002 ? add_790440 : sel_790437;
  assign add_790444 = sel_790441 + 8'h01;
  assign sel_790445 = array_index_790196 == array_index_773008 ? add_790444 : sel_790441;
  assign add_790448 = sel_790445 + 8'h01;
  assign sel_790449 = array_index_790196 == array_index_773014 ? add_790448 : sel_790445;
  assign add_790452 = sel_790449 + 8'h01;
  assign sel_790453 = array_index_790196 == array_index_773020 ? add_790452 : sel_790449;
  assign add_790456 = sel_790453 + 8'h01;
  assign sel_790457 = array_index_790196 == array_index_773026 ? add_790456 : sel_790453;
  assign add_790460 = sel_790457 + 8'h01;
  assign sel_790461 = array_index_790196 == array_index_773032 ? add_790460 : sel_790457;
  assign add_790464 = sel_790461 + 8'h01;
  assign sel_790465 = array_index_790196 == array_index_773038 ? add_790464 : sel_790461;
  assign add_790468 = sel_790465 + 8'h01;
  assign sel_790469 = array_index_790196 == array_index_773044 ? add_790468 : sel_790465;
  assign add_790472 = sel_790469 + 8'h01;
  assign sel_790473 = array_index_790196 == array_index_773050 ? add_790472 : sel_790469;
  assign add_790476 = sel_790473 + 8'h01;
  assign sel_790477 = array_index_790196 == array_index_773056 ? add_790476 : sel_790473;
  assign add_790480 = sel_790477 + 8'h01;
  assign sel_790481 = array_index_790196 == array_index_773062 ? add_790480 : sel_790477;
  assign add_790484 = sel_790481 + 8'h01;
  assign sel_790485 = array_index_790196 == array_index_773068 ? add_790484 : sel_790481;
  assign add_790488 = sel_790485 + 8'h01;
  assign sel_790489 = array_index_790196 == array_index_773074 ? add_790488 : sel_790485;
  assign add_790492 = sel_790489 + 8'h01;
  assign sel_790493 = array_index_790196 == array_index_773080 ? add_790492 : sel_790489;
  assign add_790496 = sel_790493 + 8'h01;
  assign sel_790497 = array_index_790196 == array_index_773086 ? add_790496 : sel_790493;
  assign add_790500 = sel_790497 + 8'h01;
  assign sel_790501 = array_index_790196 == array_index_773092 ? add_790500 : sel_790497;
  assign add_790504 = sel_790501 + 8'h01;
  assign sel_790505 = array_index_790196 == array_index_773098 ? add_790504 : sel_790501;
  assign add_790508 = sel_790505 + 8'h01;
  assign sel_790509 = array_index_790196 == array_index_773104 ? add_790508 : sel_790505;
  assign add_790512 = sel_790509 + 8'h01;
  assign sel_790513 = array_index_790196 == array_index_773110 ? add_790512 : sel_790509;
  assign add_790516 = sel_790513 + 8'h01;
  assign sel_790517 = array_index_790196 == array_index_773116 ? add_790516 : sel_790513;
  assign add_790520 = sel_790517 + 8'h01;
  assign sel_790521 = array_index_790196 == array_index_773122 ? add_790520 : sel_790517;
  assign add_790524 = sel_790521 + 8'h01;
  assign sel_790525 = array_index_790196 == array_index_773128 ? add_790524 : sel_790521;
  assign add_790528 = sel_790525 + 8'h01;
  assign sel_790529 = array_index_790196 == array_index_773134 ? add_790528 : sel_790525;
  assign add_790532 = sel_790529 + 8'h01;
  assign sel_790533 = array_index_790196 == array_index_773140 ? add_790532 : sel_790529;
  assign add_790536 = sel_790533 + 8'h01;
  assign sel_790537 = array_index_790196 == array_index_773146 ? add_790536 : sel_790533;
  assign add_790540 = sel_790537 + 8'h01;
  assign sel_790541 = array_index_790196 == array_index_773152 ? add_790540 : sel_790537;
  assign add_790544 = sel_790541 + 8'h01;
  assign sel_790545 = array_index_790196 == array_index_773158 ? add_790544 : sel_790541;
  assign add_790548 = sel_790545 + 8'h01;
  assign sel_790549 = array_index_790196 == array_index_773164 ? add_790548 : sel_790545;
  assign add_790552 = sel_790549 + 8'h01;
  assign sel_790553 = array_index_790196 == array_index_773170 ? add_790552 : sel_790549;
  assign add_790557 = sel_790553 + 8'h01;
  assign array_index_790558 = set1_unflattened[7'h31];
  assign sel_790559 = array_index_790196 == array_index_773176 ? add_790557 : sel_790553;
  assign add_790562 = sel_790559 + 8'h01;
  assign sel_790563 = array_index_790558 == array_index_772632 ? add_790562 : sel_790559;
  assign add_790566 = sel_790563 + 8'h01;
  assign sel_790567 = array_index_790558 == array_index_772636 ? add_790566 : sel_790563;
  assign add_790570 = sel_790567 + 8'h01;
  assign sel_790571 = array_index_790558 == array_index_772644 ? add_790570 : sel_790567;
  assign add_790574 = sel_790571 + 8'h01;
  assign sel_790575 = array_index_790558 == array_index_772652 ? add_790574 : sel_790571;
  assign add_790578 = sel_790575 + 8'h01;
  assign sel_790579 = array_index_790558 == array_index_772660 ? add_790578 : sel_790575;
  assign add_790582 = sel_790579 + 8'h01;
  assign sel_790583 = array_index_790558 == array_index_772668 ? add_790582 : sel_790579;
  assign add_790586 = sel_790583 + 8'h01;
  assign sel_790587 = array_index_790558 == array_index_772676 ? add_790586 : sel_790583;
  assign add_790590 = sel_790587 + 8'h01;
  assign sel_790591 = array_index_790558 == array_index_772684 ? add_790590 : sel_790587;
  assign add_790594 = sel_790591 + 8'h01;
  assign sel_790595 = array_index_790558 == array_index_772690 ? add_790594 : sel_790591;
  assign add_790598 = sel_790595 + 8'h01;
  assign sel_790599 = array_index_790558 == array_index_772696 ? add_790598 : sel_790595;
  assign add_790602 = sel_790599 + 8'h01;
  assign sel_790603 = array_index_790558 == array_index_772702 ? add_790602 : sel_790599;
  assign add_790606 = sel_790603 + 8'h01;
  assign sel_790607 = array_index_790558 == array_index_772708 ? add_790606 : sel_790603;
  assign add_790610 = sel_790607 + 8'h01;
  assign sel_790611 = array_index_790558 == array_index_772714 ? add_790610 : sel_790607;
  assign add_790614 = sel_790611 + 8'h01;
  assign sel_790615 = array_index_790558 == array_index_772720 ? add_790614 : sel_790611;
  assign add_790618 = sel_790615 + 8'h01;
  assign sel_790619 = array_index_790558 == array_index_772726 ? add_790618 : sel_790615;
  assign add_790622 = sel_790619 + 8'h01;
  assign sel_790623 = array_index_790558 == array_index_772732 ? add_790622 : sel_790619;
  assign add_790626 = sel_790623 + 8'h01;
  assign sel_790627 = array_index_790558 == array_index_772738 ? add_790626 : sel_790623;
  assign add_790630 = sel_790627 + 8'h01;
  assign sel_790631 = array_index_790558 == array_index_772744 ? add_790630 : sel_790627;
  assign add_790634 = sel_790631 + 8'h01;
  assign sel_790635 = array_index_790558 == array_index_772750 ? add_790634 : sel_790631;
  assign add_790638 = sel_790635 + 8'h01;
  assign sel_790639 = array_index_790558 == array_index_772756 ? add_790638 : sel_790635;
  assign add_790642 = sel_790639 + 8'h01;
  assign sel_790643 = array_index_790558 == array_index_772762 ? add_790642 : sel_790639;
  assign add_790646 = sel_790643 + 8'h01;
  assign sel_790647 = array_index_790558 == array_index_772768 ? add_790646 : sel_790643;
  assign add_790650 = sel_790647 + 8'h01;
  assign sel_790651 = array_index_790558 == array_index_772774 ? add_790650 : sel_790647;
  assign add_790654 = sel_790651 + 8'h01;
  assign sel_790655 = array_index_790558 == array_index_772780 ? add_790654 : sel_790651;
  assign add_790658 = sel_790655 + 8'h01;
  assign sel_790659 = array_index_790558 == array_index_772786 ? add_790658 : sel_790655;
  assign add_790662 = sel_790659 + 8'h01;
  assign sel_790663 = array_index_790558 == array_index_772792 ? add_790662 : sel_790659;
  assign add_790666 = sel_790663 + 8'h01;
  assign sel_790667 = array_index_790558 == array_index_772798 ? add_790666 : sel_790663;
  assign add_790670 = sel_790667 + 8'h01;
  assign sel_790671 = array_index_790558 == array_index_772804 ? add_790670 : sel_790667;
  assign add_790674 = sel_790671 + 8'h01;
  assign sel_790675 = array_index_790558 == array_index_772810 ? add_790674 : sel_790671;
  assign add_790678 = sel_790675 + 8'h01;
  assign sel_790679 = array_index_790558 == array_index_772816 ? add_790678 : sel_790675;
  assign add_790682 = sel_790679 + 8'h01;
  assign sel_790683 = array_index_790558 == array_index_772822 ? add_790682 : sel_790679;
  assign add_790686 = sel_790683 + 8'h01;
  assign sel_790687 = array_index_790558 == array_index_772828 ? add_790686 : sel_790683;
  assign add_790690 = sel_790687 + 8'h01;
  assign sel_790691 = array_index_790558 == array_index_772834 ? add_790690 : sel_790687;
  assign add_790694 = sel_790691 + 8'h01;
  assign sel_790695 = array_index_790558 == array_index_772840 ? add_790694 : sel_790691;
  assign add_790698 = sel_790695 + 8'h01;
  assign sel_790699 = array_index_790558 == array_index_772846 ? add_790698 : sel_790695;
  assign add_790702 = sel_790699 + 8'h01;
  assign sel_790703 = array_index_790558 == array_index_772852 ? add_790702 : sel_790699;
  assign add_790706 = sel_790703 + 8'h01;
  assign sel_790707 = array_index_790558 == array_index_772858 ? add_790706 : sel_790703;
  assign add_790710 = sel_790707 + 8'h01;
  assign sel_790711 = array_index_790558 == array_index_772864 ? add_790710 : sel_790707;
  assign add_790714 = sel_790711 + 8'h01;
  assign sel_790715 = array_index_790558 == array_index_772870 ? add_790714 : sel_790711;
  assign add_790718 = sel_790715 + 8'h01;
  assign sel_790719 = array_index_790558 == array_index_772876 ? add_790718 : sel_790715;
  assign add_790722 = sel_790719 + 8'h01;
  assign sel_790723 = array_index_790558 == array_index_772882 ? add_790722 : sel_790719;
  assign add_790726 = sel_790723 + 8'h01;
  assign sel_790727 = array_index_790558 == array_index_772888 ? add_790726 : sel_790723;
  assign add_790730 = sel_790727 + 8'h01;
  assign sel_790731 = array_index_790558 == array_index_772894 ? add_790730 : sel_790727;
  assign add_790734 = sel_790731 + 8'h01;
  assign sel_790735 = array_index_790558 == array_index_772900 ? add_790734 : sel_790731;
  assign add_790738 = sel_790735 + 8'h01;
  assign sel_790739 = array_index_790558 == array_index_772906 ? add_790738 : sel_790735;
  assign add_790742 = sel_790739 + 8'h01;
  assign sel_790743 = array_index_790558 == array_index_772912 ? add_790742 : sel_790739;
  assign add_790746 = sel_790743 + 8'h01;
  assign sel_790747 = array_index_790558 == array_index_772918 ? add_790746 : sel_790743;
  assign add_790750 = sel_790747 + 8'h01;
  assign sel_790751 = array_index_790558 == array_index_772924 ? add_790750 : sel_790747;
  assign add_790754 = sel_790751 + 8'h01;
  assign sel_790755 = array_index_790558 == array_index_772930 ? add_790754 : sel_790751;
  assign add_790758 = sel_790755 + 8'h01;
  assign sel_790759 = array_index_790558 == array_index_772936 ? add_790758 : sel_790755;
  assign add_790762 = sel_790759 + 8'h01;
  assign sel_790763 = array_index_790558 == array_index_772942 ? add_790762 : sel_790759;
  assign add_790766 = sel_790763 + 8'h01;
  assign sel_790767 = array_index_790558 == array_index_772948 ? add_790766 : sel_790763;
  assign add_790770 = sel_790767 + 8'h01;
  assign sel_790771 = array_index_790558 == array_index_772954 ? add_790770 : sel_790767;
  assign add_790774 = sel_790771 + 8'h01;
  assign sel_790775 = array_index_790558 == array_index_772960 ? add_790774 : sel_790771;
  assign add_790778 = sel_790775 + 8'h01;
  assign sel_790779 = array_index_790558 == array_index_772966 ? add_790778 : sel_790775;
  assign add_790782 = sel_790779 + 8'h01;
  assign sel_790783 = array_index_790558 == array_index_772972 ? add_790782 : sel_790779;
  assign add_790786 = sel_790783 + 8'h01;
  assign sel_790787 = array_index_790558 == array_index_772978 ? add_790786 : sel_790783;
  assign add_790790 = sel_790787 + 8'h01;
  assign sel_790791 = array_index_790558 == array_index_772984 ? add_790790 : sel_790787;
  assign add_790794 = sel_790791 + 8'h01;
  assign sel_790795 = array_index_790558 == array_index_772990 ? add_790794 : sel_790791;
  assign add_790798 = sel_790795 + 8'h01;
  assign sel_790799 = array_index_790558 == array_index_772996 ? add_790798 : sel_790795;
  assign add_790802 = sel_790799 + 8'h01;
  assign sel_790803 = array_index_790558 == array_index_773002 ? add_790802 : sel_790799;
  assign add_790806 = sel_790803 + 8'h01;
  assign sel_790807 = array_index_790558 == array_index_773008 ? add_790806 : sel_790803;
  assign add_790810 = sel_790807 + 8'h01;
  assign sel_790811 = array_index_790558 == array_index_773014 ? add_790810 : sel_790807;
  assign add_790814 = sel_790811 + 8'h01;
  assign sel_790815 = array_index_790558 == array_index_773020 ? add_790814 : sel_790811;
  assign add_790818 = sel_790815 + 8'h01;
  assign sel_790819 = array_index_790558 == array_index_773026 ? add_790818 : sel_790815;
  assign add_790822 = sel_790819 + 8'h01;
  assign sel_790823 = array_index_790558 == array_index_773032 ? add_790822 : sel_790819;
  assign add_790826 = sel_790823 + 8'h01;
  assign sel_790827 = array_index_790558 == array_index_773038 ? add_790826 : sel_790823;
  assign add_790830 = sel_790827 + 8'h01;
  assign sel_790831 = array_index_790558 == array_index_773044 ? add_790830 : sel_790827;
  assign add_790834 = sel_790831 + 8'h01;
  assign sel_790835 = array_index_790558 == array_index_773050 ? add_790834 : sel_790831;
  assign add_790838 = sel_790835 + 8'h01;
  assign sel_790839 = array_index_790558 == array_index_773056 ? add_790838 : sel_790835;
  assign add_790842 = sel_790839 + 8'h01;
  assign sel_790843 = array_index_790558 == array_index_773062 ? add_790842 : sel_790839;
  assign add_790846 = sel_790843 + 8'h01;
  assign sel_790847 = array_index_790558 == array_index_773068 ? add_790846 : sel_790843;
  assign add_790850 = sel_790847 + 8'h01;
  assign sel_790851 = array_index_790558 == array_index_773074 ? add_790850 : sel_790847;
  assign add_790854 = sel_790851 + 8'h01;
  assign sel_790855 = array_index_790558 == array_index_773080 ? add_790854 : sel_790851;
  assign add_790858 = sel_790855 + 8'h01;
  assign sel_790859 = array_index_790558 == array_index_773086 ? add_790858 : sel_790855;
  assign add_790862 = sel_790859 + 8'h01;
  assign sel_790863 = array_index_790558 == array_index_773092 ? add_790862 : sel_790859;
  assign add_790866 = sel_790863 + 8'h01;
  assign sel_790867 = array_index_790558 == array_index_773098 ? add_790866 : sel_790863;
  assign add_790870 = sel_790867 + 8'h01;
  assign sel_790871 = array_index_790558 == array_index_773104 ? add_790870 : sel_790867;
  assign add_790874 = sel_790871 + 8'h01;
  assign sel_790875 = array_index_790558 == array_index_773110 ? add_790874 : sel_790871;
  assign add_790878 = sel_790875 + 8'h01;
  assign sel_790879 = array_index_790558 == array_index_773116 ? add_790878 : sel_790875;
  assign add_790882 = sel_790879 + 8'h01;
  assign sel_790883 = array_index_790558 == array_index_773122 ? add_790882 : sel_790879;
  assign add_790886 = sel_790883 + 8'h01;
  assign sel_790887 = array_index_790558 == array_index_773128 ? add_790886 : sel_790883;
  assign add_790890 = sel_790887 + 8'h01;
  assign sel_790891 = array_index_790558 == array_index_773134 ? add_790890 : sel_790887;
  assign add_790894 = sel_790891 + 8'h01;
  assign sel_790895 = array_index_790558 == array_index_773140 ? add_790894 : sel_790891;
  assign add_790898 = sel_790895 + 8'h01;
  assign sel_790899 = array_index_790558 == array_index_773146 ? add_790898 : sel_790895;
  assign add_790902 = sel_790899 + 8'h01;
  assign sel_790903 = array_index_790558 == array_index_773152 ? add_790902 : sel_790899;
  assign add_790906 = sel_790903 + 8'h01;
  assign sel_790907 = array_index_790558 == array_index_773158 ? add_790906 : sel_790903;
  assign add_790910 = sel_790907 + 8'h01;
  assign sel_790911 = array_index_790558 == array_index_773164 ? add_790910 : sel_790907;
  assign add_790914 = sel_790911 + 8'h01;
  assign sel_790915 = array_index_790558 == array_index_773170 ? add_790914 : sel_790911;
  assign add_790919 = sel_790915 + 8'h01;
  assign array_index_790920 = set1_unflattened[7'h32];
  assign sel_790921 = array_index_790558 == array_index_773176 ? add_790919 : sel_790915;
  assign add_790924 = sel_790921 + 8'h01;
  assign sel_790925 = array_index_790920 == array_index_772632 ? add_790924 : sel_790921;
  assign add_790928 = sel_790925 + 8'h01;
  assign sel_790929 = array_index_790920 == array_index_772636 ? add_790928 : sel_790925;
  assign add_790932 = sel_790929 + 8'h01;
  assign sel_790933 = array_index_790920 == array_index_772644 ? add_790932 : sel_790929;
  assign add_790936 = sel_790933 + 8'h01;
  assign sel_790937 = array_index_790920 == array_index_772652 ? add_790936 : sel_790933;
  assign add_790940 = sel_790937 + 8'h01;
  assign sel_790941 = array_index_790920 == array_index_772660 ? add_790940 : sel_790937;
  assign add_790944 = sel_790941 + 8'h01;
  assign sel_790945 = array_index_790920 == array_index_772668 ? add_790944 : sel_790941;
  assign add_790948 = sel_790945 + 8'h01;
  assign sel_790949 = array_index_790920 == array_index_772676 ? add_790948 : sel_790945;
  assign add_790952 = sel_790949 + 8'h01;
  assign sel_790953 = array_index_790920 == array_index_772684 ? add_790952 : sel_790949;
  assign add_790956 = sel_790953 + 8'h01;
  assign sel_790957 = array_index_790920 == array_index_772690 ? add_790956 : sel_790953;
  assign add_790960 = sel_790957 + 8'h01;
  assign sel_790961 = array_index_790920 == array_index_772696 ? add_790960 : sel_790957;
  assign add_790964 = sel_790961 + 8'h01;
  assign sel_790965 = array_index_790920 == array_index_772702 ? add_790964 : sel_790961;
  assign add_790968 = sel_790965 + 8'h01;
  assign sel_790969 = array_index_790920 == array_index_772708 ? add_790968 : sel_790965;
  assign add_790972 = sel_790969 + 8'h01;
  assign sel_790973 = array_index_790920 == array_index_772714 ? add_790972 : sel_790969;
  assign add_790976 = sel_790973 + 8'h01;
  assign sel_790977 = array_index_790920 == array_index_772720 ? add_790976 : sel_790973;
  assign add_790980 = sel_790977 + 8'h01;
  assign sel_790981 = array_index_790920 == array_index_772726 ? add_790980 : sel_790977;
  assign add_790984 = sel_790981 + 8'h01;
  assign sel_790985 = array_index_790920 == array_index_772732 ? add_790984 : sel_790981;
  assign add_790988 = sel_790985 + 8'h01;
  assign sel_790989 = array_index_790920 == array_index_772738 ? add_790988 : sel_790985;
  assign add_790992 = sel_790989 + 8'h01;
  assign sel_790993 = array_index_790920 == array_index_772744 ? add_790992 : sel_790989;
  assign add_790996 = sel_790993 + 8'h01;
  assign sel_790997 = array_index_790920 == array_index_772750 ? add_790996 : sel_790993;
  assign add_791000 = sel_790997 + 8'h01;
  assign sel_791001 = array_index_790920 == array_index_772756 ? add_791000 : sel_790997;
  assign add_791004 = sel_791001 + 8'h01;
  assign sel_791005 = array_index_790920 == array_index_772762 ? add_791004 : sel_791001;
  assign add_791008 = sel_791005 + 8'h01;
  assign sel_791009 = array_index_790920 == array_index_772768 ? add_791008 : sel_791005;
  assign add_791012 = sel_791009 + 8'h01;
  assign sel_791013 = array_index_790920 == array_index_772774 ? add_791012 : sel_791009;
  assign add_791016 = sel_791013 + 8'h01;
  assign sel_791017 = array_index_790920 == array_index_772780 ? add_791016 : sel_791013;
  assign add_791020 = sel_791017 + 8'h01;
  assign sel_791021 = array_index_790920 == array_index_772786 ? add_791020 : sel_791017;
  assign add_791024 = sel_791021 + 8'h01;
  assign sel_791025 = array_index_790920 == array_index_772792 ? add_791024 : sel_791021;
  assign add_791028 = sel_791025 + 8'h01;
  assign sel_791029 = array_index_790920 == array_index_772798 ? add_791028 : sel_791025;
  assign add_791032 = sel_791029 + 8'h01;
  assign sel_791033 = array_index_790920 == array_index_772804 ? add_791032 : sel_791029;
  assign add_791036 = sel_791033 + 8'h01;
  assign sel_791037 = array_index_790920 == array_index_772810 ? add_791036 : sel_791033;
  assign add_791040 = sel_791037 + 8'h01;
  assign sel_791041 = array_index_790920 == array_index_772816 ? add_791040 : sel_791037;
  assign add_791044 = sel_791041 + 8'h01;
  assign sel_791045 = array_index_790920 == array_index_772822 ? add_791044 : sel_791041;
  assign add_791048 = sel_791045 + 8'h01;
  assign sel_791049 = array_index_790920 == array_index_772828 ? add_791048 : sel_791045;
  assign add_791052 = sel_791049 + 8'h01;
  assign sel_791053 = array_index_790920 == array_index_772834 ? add_791052 : sel_791049;
  assign add_791056 = sel_791053 + 8'h01;
  assign sel_791057 = array_index_790920 == array_index_772840 ? add_791056 : sel_791053;
  assign add_791060 = sel_791057 + 8'h01;
  assign sel_791061 = array_index_790920 == array_index_772846 ? add_791060 : sel_791057;
  assign add_791064 = sel_791061 + 8'h01;
  assign sel_791065 = array_index_790920 == array_index_772852 ? add_791064 : sel_791061;
  assign add_791068 = sel_791065 + 8'h01;
  assign sel_791069 = array_index_790920 == array_index_772858 ? add_791068 : sel_791065;
  assign add_791072 = sel_791069 + 8'h01;
  assign sel_791073 = array_index_790920 == array_index_772864 ? add_791072 : sel_791069;
  assign add_791076 = sel_791073 + 8'h01;
  assign sel_791077 = array_index_790920 == array_index_772870 ? add_791076 : sel_791073;
  assign add_791080 = sel_791077 + 8'h01;
  assign sel_791081 = array_index_790920 == array_index_772876 ? add_791080 : sel_791077;
  assign add_791084 = sel_791081 + 8'h01;
  assign sel_791085 = array_index_790920 == array_index_772882 ? add_791084 : sel_791081;
  assign add_791088 = sel_791085 + 8'h01;
  assign sel_791089 = array_index_790920 == array_index_772888 ? add_791088 : sel_791085;
  assign add_791092 = sel_791089 + 8'h01;
  assign sel_791093 = array_index_790920 == array_index_772894 ? add_791092 : sel_791089;
  assign add_791096 = sel_791093 + 8'h01;
  assign sel_791097 = array_index_790920 == array_index_772900 ? add_791096 : sel_791093;
  assign add_791100 = sel_791097 + 8'h01;
  assign sel_791101 = array_index_790920 == array_index_772906 ? add_791100 : sel_791097;
  assign add_791104 = sel_791101 + 8'h01;
  assign sel_791105 = array_index_790920 == array_index_772912 ? add_791104 : sel_791101;
  assign add_791108 = sel_791105 + 8'h01;
  assign sel_791109 = array_index_790920 == array_index_772918 ? add_791108 : sel_791105;
  assign add_791112 = sel_791109 + 8'h01;
  assign sel_791113 = array_index_790920 == array_index_772924 ? add_791112 : sel_791109;
  assign add_791116 = sel_791113 + 8'h01;
  assign sel_791117 = array_index_790920 == array_index_772930 ? add_791116 : sel_791113;
  assign add_791120 = sel_791117 + 8'h01;
  assign sel_791121 = array_index_790920 == array_index_772936 ? add_791120 : sel_791117;
  assign add_791124 = sel_791121 + 8'h01;
  assign sel_791125 = array_index_790920 == array_index_772942 ? add_791124 : sel_791121;
  assign add_791128 = sel_791125 + 8'h01;
  assign sel_791129 = array_index_790920 == array_index_772948 ? add_791128 : sel_791125;
  assign add_791132 = sel_791129 + 8'h01;
  assign sel_791133 = array_index_790920 == array_index_772954 ? add_791132 : sel_791129;
  assign add_791136 = sel_791133 + 8'h01;
  assign sel_791137 = array_index_790920 == array_index_772960 ? add_791136 : sel_791133;
  assign add_791140 = sel_791137 + 8'h01;
  assign sel_791141 = array_index_790920 == array_index_772966 ? add_791140 : sel_791137;
  assign add_791144 = sel_791141 + 8'h01;
  assign sel_791145 = array_index_790920 == array_index_772972 ? add_791144 : sel_791141;
  assign add_791148 = sel_791145 + 8'h01;
  assign sel_791149 = array_index_790920 == array_index_772978 ? add_791148 : sel_791145;
  assign add_791152 = sel_791149 + 8'h01;
  assign sel_791153 = array_index_790920 == array_index_772984 ? add_791152 : sel_791149;
  assign add_791156 = sel_791153 + 8'h01;
  assign sel_791157 = array_index_790920 == array_index_772990 ? add_791156 : sel_791153;
  assign add_791160 = sel_791157 + 8'h01;
  assign sel_791161 = array_index_790920 == array_index_772996 ? add_791160 : sel_791157;
  assign add_791164 = sel_791161 + 8'h01;
  assign sel_791165 = array_index_790920 == array_index_773002 ? add_791164 : sel_791161;
  assign add_791168 = sel_791165 + 8'h01;
  assign sel_791169 = array_index_790920 == array_index_773008 ? add_791168 : sel_791165;
  assign add_791172 = sel_791169 + 8'h01;
  assign sel_791173 = array_index_790920 == array_index_773014 ? add_791172 : sel_791169;
  assign add_791176 = sel_791173 + 8'h01;
  assign sel_791177 = array_index_790920 == array_index_773020 ? add_791176 : sel_791173;
  assign add_791180 = sel_791177 + 8'h01;
  assign sel_791181 = array_index_790920 == array_index_773026 ? add_791180 : sel_791177;
  assign add_791184 = sel_791181 + 8'h01;
  assign sel_791185 = array_index_790920 == array_index_773032 ? add_791184 : sel_791181;
  assign add_791188 = sel_791185 + 8'h01;
  assign sel_791189 = array_index_790920 == array_index_773038 ? add_791188 : sel_791185;
  assign add_791192 = sel_791189 + 8'h01;
  assign sel_791193 = array_index_790920 == array_index_773044 ? add_791192 : sel_791189;
  assign add_791196 = sel_791193 + 8'h01;
  assign sel_791197 = array_index_790920 == array_index_773050 ? add_791196 : sel_791193;
  assign add_791200 = sel_791197 + 8'h01;
  assign sel_791201 = array_index_790920 == array_index_773056 ? add_791200 : sel_791197;
  assign add_791204 = sel_791201 + 8'h01;
  assign sel_791205 = array_index_790920 == array_index_773062 ? add_791204 : sel_791201;
  assign add_791208 = sel_791205 + 8'h01;
  assign sel_791209 = array_index_790920 == array_index_773068 ? add_791208 : sel_791205;
  assign add_791212 = sel_791209 + 8'h01;
  assign sel_791213 = array_index_790920 == array_index_773074 ? add_791212 : sel_791209;
  assign add_791216 = sel_791213 + 8'h01;
  assign sel_791217 = array_index_790920 == array_index_773080 ? add_791216 : sel_791213;
  assign add_791220 = sel_791217 + 8'h01;
  assign sel_791221 = array_index_790920 == array_index_773086 ? add_791220 : sel_791217;
  assign add_791224 = sel_791221 + 8'h01;
  assign sel_791225 = array_index_790920 == array_index_773092 ? add_791224 : sel_791221;
  assign add_791228 = sel_791225 + 8'h01;
  assign sel_791229 = array_index_790920 == array_index_773098 ? add_791228 : sel_791225;
  assign add_791232 = sel_791229 + 8'h01;
  assign sel_791233 = array_index_790920 == array_index_773104 ? add_791232 : sel_791229;
  assign add_791236 = sel_791233 + 8'h01;
  assign sel_791237 = array_index_790920 == array_index_773110 ? add_791236 : sel_791233;
  assign add_791240 = sel_791237 + 8'h01;
  assign sel_791241 = array_index_790920 == array_index_773116 ? add_791240 : sel_791237;
  assign add_791244 = sel_791241 + 8'h01;
  assign sel_791245 = array_index_790920 == array_index_773122 ? add_791244 : sel_791241;
  assign add_791248 = sel_791245 + 8'h01;
  assign sel_791249 = array_index_790920 == array_index_773128 ? add_791248 : sel_791245;
  assign add_791252 = sel_791249 + 8'h01;
  assign sel_791253 = array_index_790920 == array_index_773134 ? add_791252 : sel_791249;
  assign add_791256 = sel_791253 + 8'h01;
  assign sel_791257 = array_index_790920 == array_index_773140 ? add_791256 : sel_791253;
  assign add_791260 = sel_791257 + 8'h01;
  assign sel_791261 = array_index_790920 == array_index_773146 ? add_791260 : sel_791257;
  assign add_791264 = sel_791261 + 8'h01;
  assign sel_791265 = array_index_790920 == array_index_773152 ? add_791264 : sel_791261;
  assign add_791268 = sel_791265 + 8'h01;
  assign sel_791269 = array_index_790920 == array_index_773158 ? add_791268 : sel_791265;
  assign add_791272 = sel_791269 + 8'h01;
  assign sel_791273 = array_index_790920 == array_index_773164 ? add_791272 : sel_791269;
  assign add_791276 = sel_791273 + 8'h01;
  assign sel_791277 = array_index_790920 == array_index_773170 ? add_791276 : sel_791273;
  assign add_791281 = sel_791277 + 8'h01;
  assign array_index_791282 = set1_unflattened[7'h33];
  assign sel_791283 = array_index_790920 == array_index_773176 ? add_791281 : sel_791277;
  assign add_791286 = sel_791283 + 8'h01;
  assign sel_791287 = array_index_791282 == array_index_772632 ? add_791286 : sel_791283;
  assign add_791290 = sel_791287 + 8'h01;
  assign sel_791291 = array_index_791282 == array_index_772636 ? add_791290 : sel_791287;
  assign add_791294 = sel_791291 + 8'h01;
  assign sel_791295 = array_index_791282 == array_index_772644 ? add_791294 : sel_791291;
  assign add_791298 = sel_791295 + 8'h01;
  assign sel_791299 = array_index_791282 == array_index_772652 ? add_791298 : sel_791295;
  assign add_791302 = sel_791299 + 8'h01;
  assign sel_791303 = array_index_791282 == array_index_772660 ? add_791302 : sel_791299;
  assign add_791306 = sel_791303 + 8'h01;
  assign sel_791307 = array_index_791282 == array_index_772668 ? add_791306 : sel_791303;
  assign add_791310 = sel_791307 + 8'h01;
  assign sel_791311 = array_index_791282 == array_index_772676 ? add_791310 : sel_791307;
  assign add_791314 = sel_791311 + 8'h01;
  assign sel_791315 = array_index_791282 == array_index_772684 ? add_791314 : sel_791311;
  assign add_791318 = sel_791315 + 8'h01;
  assign sel_791319 = array_index_791282 == array_index_772690 ? add_791318 : sel_791315;
  assign add_791322 = sel_791319 + 8'h01;
  assign sel_791323 = array_index_791282 == array_index_772696 ? add_791322 : sel_791319;
  assign add_791326 = sel_791323 + 8'h01;
  assign sel_791327 = array_index_791282 == array_index_772702 ? add_791326 : sel_791323;
  assign add_791330 = sel_791327 + 8'h01;
  assign sel_791331 = array_index_791282 == array_index_772708 ? add_791330 : sel_791327;
  assign add_791334 = sel_791331 + 8'h01;
  assign sel_791335 = array_index_791282 == array_index_772714 ? add_791334 : sel_791331;
  assign add_791338 = sel_791335 + 8'h01;
  assign sel_791339 = array_index_791282 == array_index_772720 ? add_791338 : sel_791335;
  assign add_791342 = sel_791339 + 8'h01;
  assign sel_791343 = array_index_791282 == array_index_772726 ? add_791342 : sel_791339;
  assign add_791346 = sel_791343 + 8'h01;
  assign sel_791347 = array_index_791282 == array_index_772732 ? add_791346 : sel_791343;
  assign add_791350 = sel_791347 + 8'h01;
  assign sel_791351 = array_index_791282 == array_index_772738 ? add_791350 : sel_791347;
  assign add_791354 = sel_791351 + 8'h01;
  assign sel_791355 = array_index_791282 == array_index_772744 ? add_791354 : sel_791351;
  assign add_791358 = sel_791355 + 8'h01;
  assign sel_791359 = array_index_791282 == array_index_772750 ? add_791358 : sel_791355;
  assign add_791362 = sel_791359 + 8'h01;
  assign sel_791363 = array_index_791282 == array_index_772756 ? add_791362 : sel_791359;
  assign add_791366 = sel_791363 + 8'h01;
  assign sel_791367 = array_index_791282 == array_index_772762 ? add_791366 : sel_791363;
  assign add_791370 = sel_791367 + 8'h01;
  assign sel_791371 = array_index_791282 == array_index_772768 ? add_791370 : sel_791367;
  assign add_791374 = sel_791371 + 8'h01;
  assign sel_791375 = array_index_791282 == array_index_772774 ? add_791374 : sel_791371;
  assign add_791378 = sel_791375 + 8'h01;
  assign sel_791379 = array_index_791282 == array_index_772780 ? add_791378 : sel_791375;
  assign add_791382 = sel_791379 + 8'h01;
  assign sel_791383 = array_index_791282 == array_index_772786 ? add_791382 : sel_791379;
  assign add_791386 = sel_791383 + 8'h01;
  assign sel_791387 = array_index_791282 == array_index_772792 ? add_791386 : sel_791383;
  assign add_791390 = sel_791387 + 8'h01;
  assign sel_791391 = array_index_791282 == array_index_772798 ? add_791390 : sel_791387;
  assign add_791394 = sel_791391 + 8'h01;
  assign sel_791395 = array_index_791282 == array_index_772804 ? add_791394 : sel_791391;
  assign add_791398 = sel_791395 + 8'h01;
  assign sel_791399 = array_index_791282 == array_index_772810 ? add_791398 : sel_791395;
  assign add_791402 = sel_791399 + 8'h01;
  assign sel_791403 = array_index_791282 == array_index_772816 ? add_791402 : sel_791399;
  assign add_791406 = sel_791403 + 8'h01;
  assign sel_791407 = array_index_791282 == array_index_772822 ? add_791406 : sel_791403;
  assign add_791410 = sel_791407 + 8'h01;
  assign sel_791411 = array_index_791282 == array_index_772828 ? add_791410 : sel_791407;
  assign add_791414 = sel_791411 + 8'h01;
  assign sel_791415 = array_index_791282 == array_index_772834 ? add_791414 : sel_791411;
  assign add_791418 = sel_791415 + 8'h01;
  assign sel_791419 = array_index_791282 == array_index_772840 ? add_791418 : sel_791415;
  assign add_791422 = sel_791419 + 8'h01;
  assign sel_791423 = array_index_791282 == array_index_772846 ? add_791422 : sel_791419;
  assign add_791426 = sel_791423 + 8'h01;
  assign sel_791427 = array_index_791282 == array_index_772852 ? add_791426 : sel_791423;
  assign add_791430 = sel_791427 + 8'h01;
  assign sel_791431 = array_index_791282 == array_index_772858 ? add_791430 : sel_791427;
  assign add_791434 = sel_791431 + 8'h01;
  assign sel_791435 = array_index_791282 == array_index_772864 ? add_791434 : sel_791431;
  assign add_791438 = sel_791435 + 8'h01;
  assign sel_791439 = array_index_791282 == array_index_772870 ? add_791438 : sel_791435;
  assign add_791442 = sel_791439 + 8'h01;
  assign sel_791443 = array_index_791282 == array_index_772876 ? add_791442 : sel_791439;
  assign add_791446 = sel_791443 + 8'h01;
  assign sel_791447 = array_index_791282 == array_index_772882 ? add_791446 : sel_791443;
  assign add_791450 = sel_791447 + 8'h01;
  assign sel_791451 = array_index_791282 == array_index_772888 ? add_791450 : sel_791447;
  assign add_791454 = sel_791451 + 8'h01;
  assign sel_791455 = array_index_791282 == array_index_772894 ? add_791454 : sel_791451;
  assign add_791458 = sel_791455 + 8'h01;
  assign sel_791459 = array_index_791282 == array_index_772900 ? add_791458 : sel_791455;
  assign add_791462 = sel_791459 + 8'h01;
  assign sel_791463 = array_index_791282 == array_index_772906 ? add_791462 : sel_791459;
  assign add_791466 = sel_791463 + 8'h01;
  assign sel_791467 = array_index_791282 == array_index_772912 ? add_791466 : sel_791463;
  assign add_791470 = sel_791467 + 8'h01;
  assign sel_791471 = array_index_791282 == array_index_772918 ? add_791470 : sel_791467;
  assign add_791474 = sel_791471 + 8'h01;
  assign sel_791475 = array_index_791282 == array_index_772924 ? add_791474 : sel_791471;
  assign add_791478 = sel_791475 + 8'h01;
  assign sel_791479 = array_index_791282 == array_index_772930 ? add_791478 : sel_791475;
  assign add_791482 = sel_791479 + 8'h01;
  assign sel_791483 = array_index_791282 == array_index_772936 ? add_791482 : sel_791479;
  assign add_791486 = sel_791483 + 8'h01;
  assign sel_791487 = array_index_791282 == array_index_772942 ? add_791486 : sel_791483;
  assign add_791490 = sel_791487 + 8'h01;
  assign sel_791491 = array_index_791282 == array_index_772948 ? add_791490 : sel_791487;
  assign add_791494 = sel_791491 + 8'h01;
  assign sel_791495 = array_index_791282 == array_index_772954 ? add_791494 : sel_791491;
  assign add_791498 = sel_791495 + 8'h01;
  assign sel_791499 = array_index_791282 == array_index_772960 ? add_791498 : sel_791495;
  assign add_791502 = sel_791499 + 8'h01;
  assign sel_791503 = array_index_791282 == array_index_772966 ? add_791502 : sel_791499;
  assign add_791506 = sel_791503 + 8'h01;
  assign sel_791507 = array_index_791282 == array_index_772972 ? add_791506 : sel_791503;
  assign add_791510 = sel_791507 + 8'h01;
  assign sel_791511 = array_index_791282 == array_index_772978 ? add_791510 : sel_791507;
  assign add_791514 = sel_791511 + 8'h01;
  assign sel_791515 = array_index_791282 == array_index_772984 ? add_791514 : sel_791511;
  assign add_791518 = sel_791515 + 8'h01;
  assign sel_791519 = array_index_791282 == array_index_772990 ? add_791518 : sel_791515;
  assign add_791522 = sel_791519 + 8'h01;
  assign sel_791523 = array_index_791282 == array_index_772996 ? add_791522 : sel_791519;
  assign add_791526 = sel_791523 + 8'h01;
  assign sel_791527 = array_index_791282 == array_index_773002 ? add_791526 : sel_791523;
  assign add_791530 = sel_791527 + 8'h01;
  assign sel_791531 = array_index_791282 == array_index_773008 ? add_791530 : sel_791527;
  assign add_791534 = sel_791531 + 8'h01;
  assign sel_791535 = array_index_791282 == array_index_773014 ? add_791534 : sel_791531;
  assign add_791538 = sel_791535 + 8'h01;
  assign sel_791539 = array_index_791282 == array_index_773020 ? add_791538 : sel_791535;
  assign add_791542 = sel_791539 + 8'h01;
  assign sel_791543 = array_index_791282 == array_index_773026 ? add_791542 : sel_791539;
  assign add_791546 = sel_791543 + 8'h01;
  assign sel_791547 = array_index_791282 == array_index_773032 ? add_791546 : sel_791543;
  assign add_791550 = sel_791547 + 8'h01;
  assign sel_791551 = array_index_791282 == array_index_773038 ? add_791550 : sel_791547;
  assign add_791554 = sel_791551 + 8'h01;
  assign sel_791555 = array_index_791282 == array_index_773044 ? add_791554 : sel_791551;
  assign add_791558 = sel_791555 + 8'h01;
  assign sel_791559 = array_index_791282 == array_index_773050 ? add_791558 : sel_791555;
  assign add_791562 = sel_791559 + 8'h01;
  assign sel_791563 = array_index_791282 == array_index_773056 ? add_791562 : sel_791559;
  assign add_791566 = sel_791563 + 8'h01;
  assign sel_791567 = array_index_791282 == array_index_773062 ? add_791566 : sel_791563;
  assign add_791570 = sel_791567 + 8'h01;
  assign sel_791571 = array_index_791282 == array_index_773068 ? add_791570 : sel_791567;
  assign add_791574 = sel_791571 + 8'h01;
  assign sel_791575 = array_index_791282 == array_index_773074 ? add_791574 : sel_791571;
  assign add_791578 = sel_791575 + 8'h01;
  assign sel_791579 = array_index_791282 == array_index_773080 ? add_791578 : sel_791575;
  assign add_791582 = sel_791579 + 8'h01;
  assign sel_791583 = array_index_791282 == array_index_773086 ? add_791582 : sel_791579;
  assign add_791586 = sel_791583 + 8'h01;
  assign sel_791587 = array_index_791282 == array_index_773092 ? add_791586 : sel_791583;
  assign add_791590 = sel_791587 + 8'h01;
  assign sel_791591 = array_index_791282 == array_index_773098 ? add_791590 : sel_791587;
  assign add_791594 = sel_791591 + 8'h01;
  assign sel_791595 = array_index_791282 == array_index_773104 ? add_791594 : sel_791591;
  assign add_791598 = sel_791595 + 8'h01;
  assign sel_791599 = array_index_791282 == array_index_773110 ? add_791598 : sel_791595;
  assign add_791602 = sel_791599 + 8'h01;
  assign sel_791603 = array_index_791282 == array_index_773116 ? add_791602 : sel_791599;
  assign add_791606 = sel_791603 + 8'h01;
  assign sel_791607 = array_index_791282 == array_index_773122 ? add_791606 : sel_791603;
  assign add_791610 = sel_791607 + 8'h01;
  assign sel_791611 = array_index_791282 == array_index_773128 ? add_791610 : sel_791607;
  assign add_791614 = sel_791611 + 8'h01;
  assign sel_791615 = array_index_791282 == array_index_773134 ? add_791614 : sel_791611;
  assign add_791618 = sel_791615 + 8'h01;
  assign sel_791619 = array_index_791282 == array_index_773140 ? add_791618 : sel_791615;
  assign add_791622 = sel_791619 + 8'h01;
  assign sel_791623 = array_index_791282 == array_index_773146 ? add_791622 : sel_791619;
  assign add_791626 = sel_791623 + 8'h01;
  assign sel_791627 = array_index_791282 == array_index_773152 ? add_791626 : sel_791623;
  assign add_791630 = sel_791627 + 8'h01;
  assign sel_791631 = array_index_791282 == array_index_773158 ? add_791630 : sel_791627;
  assign add_791634 = sel_791631 + 8'h01;
  assign sel_791635 = array_index_791282 == array_index_773164 ? add_791634 : sel_791631;
  assign add_791638 = sel_791635 + 8'h01;
  assign sel_791639 = array_index_791282 == array_index_773170 ? add_791638 : sel_791635;
  assign add_791643 = sel_791639 + 8'h01;
  assign array_index_791644 = set1_unflattened[7'h34];
  assign sel_791645 = array_index_791282 == array_index_773176 ? add_791643 : sel_791639;
  assign add_791648 = sel_791645 + 8'h01;
  assign sel_791649 = array_index_791644 == array_index_772632 ? add_791648 : sel_791645;
  assign add_791652 = sel_791649 + 8'h01;
  assign sel_791653 = array_index_791644 == array_index_772636 ? add_791652 : sel_791649;
  assign add_791656 = sel_791653 + 8'h01;
  assign sel_791657 = array_index_791644 == array_index_772644 ? add_791656 : sel_791653;
  assign add_791660 = sel_791657 + 8'h01;
  assign sel_791661 = array_index_791644 == array_index_772652 ? add_791660 : sel_791657;
  assign add_791664 = sel_791661 + 8'h01;
  assign sel_791665 = array_index_791644 == array_index_772660 ? add_791664 : sel_791661;
  assign add_791668 = sel_791665 + 8'h01;
  assign sel_791669 = array_index_791644 == array_index_772668 ? add_791668 : sel_791665;
  assign add_791672 = sel_791669 + 8'h01;
  assign sel_791673 = array_index_791644 == array_index_772676 ? add_791672 : sel_791669;
  assign add_791676 = sel_791673 + 8'h01;
  assign sel_791677 = array_index_791644 == array_index_772684 ? add_791676 : sel_791673;
  assign add_791680 = sel_791677 + 8'h01;
  assign sel_791681 = array_index_791644 == array_index_772690 ? add_791680 : sel_791677;
  assign add_791684 = sel_791681 + 8'h01;
  assign sel_791685 = array_index_791644 == array_index_772696 ? add_791684 : sel_791681;
  assign add_791688 = sel_791685 + 8'h01;
  assign sel_791689 = array_index_791644 == array_index_772702 ? add_791688 : sel_791685;
  assign add_791692 = sel_791689 + 8'h01;
  assign sel_791693 = array_index_791644 == array_index_772708 ? add_791692 : sel_791689;
  assign add_791696 = sel_791693 + 8'h01;
  assign sel_791697 = array_index_791644 == array_index_772714 ? add_791696 : sel_791693;
  assign add_791700 = sel_791697 + 8'h01;
  assign sel_791701 = array_index_791644 == array_index_772720 ? add_791700 : sel_791697;
  assign add_791704 = sel_791701 + 8'h01;
  assign sel_791705 = array_index_791644 == array_index_772726 ? add_791704 : sel_791701;
  assign add_791708 = sel_791705 + 8'h01;
  assign sel_791709 = array_index_791644 == array_index_772732 ? add_791708 : sel_791705;
  assign add_791712 = sel_791709 + 8'h01;
  assign sel_791713 = array_index_791644 == array_index_772738 ? add_791712 : sel_791709;
  assign add_791716 = sel_791713 + 8'h01;
  assign sel_791717 = array_index_791644 == array_index_772744 ? add_791716 : sel_791713;
  assign add_791720 = sel_791717 + 8'h01;
  assign sel_791721 = array_index_791644 == array_index_772750 ? add_791720 : sel_791717;
  assign add_791724 = sel_791721 + 8'h01;
  assign sel_791725 = array_index_791644 == array_index_772756 ? add_791724 : sel_791721;
  assign add_791728 = sel_791725 + 8'h01;
  assign sel_791729 = array_index_791644 == array_index_772762 ? add_791728 : sel_791725;
  assign add_791732 = sel_791729 + 8'h01;
  assign sel_791733 = array_index_791644 == array_index_772768 ? add_791732 : sel_791729;
  assign add_791736 = sel_791733 + 8'h01;
  assign sel_791737 = array_index_791644 == array_index_772774 ? add_791736 : sel_791733;
  assign add_791740 = sel_791737 + 8'h01;
  assign sel_791741 = array_index_791644 == array_index_772780 ? add_791740 : sel_791737;
  assign add_791744 = sel_791741 + 8'h01;
  assign sel_791745 = array_index_791644 == array_index_772786 ? add_791744 : sel_791741;
  assign add_791748 = sel_791745 + 8'h01;
  assign sel_791749 = array_index_791644 == array_index_772792 ? add_791748 : sel_791745;
  assign add_791752 = sel_791749 + 8'h01;
  assign sel_791753 = array_index_791644 == array_index_772798 ? add_791752 : sel_791749;
  assign add_791756 = sel_791753 + 8'h01;
  assign sel_791757 = array_index_791644 == array_index_772804 ? add_791756 : sel_791753;
  assign add_791760 = sel_791757 + 8'h01;
  assign sel_791761 = array_index_791644 == array_index_772810 ? add_791760 : sel_791757;
  assign add_791764 = sel_791761 + 8'h01;
  assign sel_791765 = array_index_791644 == array_index_772816 ? add_791764 : sel_791761;
  assign add_791768 = sel_791765 + 8'h01;
  assign sel_791769 = array_index_791644 == array_index_772822 ? add_791768 : sel_791765;
  assign add_791772 = sel_791769 + 8'h01;
  assign sel_791773 = array_index_791644 == array_index_772828 ? add_791772 : sel_791769;
  assign add_791776 = sel_791773 + 8'h01;
  assign sel_791777 = array_index_791644 == array_index_772834 ? add_791776 : sel_791773;
  assign add_791780 = sel_791777 + 8'h01;
  assign sel_791781 = array_index_791644 == array_index_772840 ? add_791780 : sel_791777;
  assign add_791784 = sel_791781 + 8'h01;
  assign sel_791785 = array_index_791644 == array_index_772846 ? add_791784 : sel_791781;
  assign add_791788 = sel_791785 + 8'h01;
  assign sel_791789 = array_index_791644 == array_index_772852 ? add_791788 : sel_791785;
  assign add_791792 = sel_791789 + 8'h01;
  assign sel_791793 = array_index_791644 == array_index_772858 ? add_791792 : sel_791789;
  assign add_791796 = sel_791793 + 8'h01;
  assign sel_791797 = array_index_791644 == array_index_772864 ? add_791796 : sel_791793;
  assign add_791800 = sel_791797 + 8'h01;
  assign sel_791801 = array_index_791644 == array_index_772870 ? add_791800 : sel_791797;
  assign add_791804 = sel_791801 + 8'h01;
  assign sel_791805 = array_index_791644 == array_index_772876 ? add_791804 : sel_791801;
  assign add_791808 = sel_791805 + 8'h01;
  assign sel_791809 = array_index_791644 == array_index_772882 ? add_791808 : sel_791805;
  assign add_791812 = sel_791809 + 8'h01;
  assign sel_791813 = array_index_791644 == array_index_772888 ? add_791812 : sel_791809;
  assign add_791816 = sel_791813 + 8'h01;
  assign sel_791817 = array_index_791644 == array_index_772894 ? add_791816 : sel_791813;
  assign add_791820 = sel_791817 + 8'h01;
  assign sel_791821 = array_index_791644 == array_index_772900 ? add_791820 : sel_791817;
  assign add_791824 = sel_791821 + 8'h01;
  assign sel_791825 = array_index_791644 == array_index_772906 ? add_791824 : sel_791821;
  assign add_791828 = sel_791825 + 8'h01;
  assign sel_791829 = array_index_791644 == array_index_772912 ? add_791828 : sel_791825;
  assign add_791832 = sel_791829 + 8'h01;
  assign sel_791833 = array_index_791644 == array_index_772918 ? add_791832 : sel_791829;
  assign add_791836 = sel_791833 + 8'h01;
  assign sel_791837 = array_index_791644 == array_index_772924 ? add_791836 : sel_791833;
  assign add_791840 = sel_791837 + 8'h01;
  assign sel_791841 = array_index_791644 == array_index_772930 ? add_791840 : sel_791837;
  assign add_791844 = sel_791841 + 8'h01;
  assign sel_791845 = array_index_791644 == array_index_772936 ? add_791844 : sel_791841;
  assign add_791848 = sel_791845 + 8'h01;
  assign sel_791849 = array_index_791644 == array_index_772942 ? add_791848 : sel_791845;
  assign add_791852 = sel_791849 + 8'h01;
  assign sel_791853 = array_index_791644 == array_index_772948 ? add_791852 : sel_791849;
  assign add_791856 = sel_791853 + 8'h01;
  assign sel_791857 = array_index_791644 == array_index_772954 ? add_791856 : sel_791853;
  assign add_791860 = sel_791857 + 8'h01;
  assign sel_791861 = array_index_791644 == array_index_772960 ? add_791860 : sel_791857;
  assign add_791864 = sel_791861 + 8'h01;
  assign sel_791865 = array_index_791644 == array_index_772966 ? add_791864 : sel_791861;
  assign add_791868 = sel_791865 + 8'h01;
  assign sel_791869 = array_index_791644 == array_index_772972 ? add_791868 : sel_791865;
  assign add_791872 = sel_791869 + 8'h01;
  assign sel_791873 = array_index_791644 == array_index_772978 ? add_791872 : sel_791869;
  assign add_791876 = sel_791873 + 8'h01;
  assign sel_791877 = array_index_791644 == array_index_772984 ? add_791876 : sel_791873;
  assign add_791880 = sel_791877 + 8'h01;
  assign sel_791881 = array_index_791644 == array_index_772990 ? add_791880 : sel_791877;
  assign add_791884 = sel_791881 + 8'h01;
  assign sel_791885 = array_index_791644 == array_index_772996 ? add_791884 : sel_791881;
  assign add_791888 = sel_791885 + 8'h01;
  assign sel_791889 = array_index_791644 == array_index_773002 ? add_791888 : sel_791885;
  assign add_791892 = sel_791889 + 8'h01;
  assign sel_791893 = array_index_791644 == array_index_773008 ? add_791892 : sel_791889;
  assign add_791896 = sel_791893 + 8'h01;
  assign sel_791897 = array_index_791644 == array_index_773014 ? add_791896 : sel_791893;
  assign add_791900 = sel_791897 + 8'h01;
  assign sel_791901 = array_index_791644 == array_index_773020 ? add_791900 : sel_791897;
  assign add_791904 = sel_791901 + 8'h01;
  assign sel_791905 = array_index_791644 == array_index_773026 ? add_791904 : sel_791901;
  assign add_791908 = sel_791905 + 8'h01;
  assign sel_791909 = array_index_791644 == array_index_773032 ? add_791908 : sel_791905;
  assign add_791912 = sel_791909 + 8'h01;
  assign sel_791913 = array_index_791644 == array_index_773038 ? add_791912 : sel_791909;
  assign add_791916 = sel_791913 + 8'h01;
  assign sel_791917 = array_index_791644 == array_index_773044 ? add_791916 : sel_791913;
  assign add_791920 = sel_791917 + 8'h01;
  assign sel_791921 = array_index_791644 == array_index_773050 ? add_791920 : sel_791917;
  assign add_791924 = sel_791921 + 8'h01;
  assign sel_791925 = array_index_791644 == array_index_773056 ? add_791924 : sel_791921;
  assign add_791928 = sel_791925 + 8'h01;
  assign sel_791929 = array_index_791644 == array_index_773062 ? add_791928 : sel_791925;
  assign add_791932 = sel_791929 + 8'h01;
  assign sel_791933 = array_index_791644 == array_index_773068 ? add_791932 : sel_791929;
  assign add_791936 = sel_791933 + 8'h01;
  assign sel_791937 = array_index_791644 == array_index_773074 ? add_791936 : sel_791933;
  assign add_791940 = sel_791937 + 8'h01;
  assign sel_791941 = array_index_791644 == array_index_773080 ? add_791940 : sel_791937;
  assign add_791944 = sel_791941 + 8'h01;
  assign sel_791945 = array_index_791644 == array_index_773086 ? add_791944 : sel_791941;
  assign add_791948 = sel_791945 + 8'h01;
  assign sel_791949 = array_index_791644 == array_index_773092 ? add_791948 : sel_791945;
  assign add_791952 = sel_791949 + 8'h01;
  assign sel_791953 = array_index_791644 == array_index_773098 ? add_791952 : sel_791949;
  assign add_791956 = sel_791953 + 8'h01;
  assign sel_791957 = array_index_791644 == array_index_773104 ? add_791956 : sel_791953;
  assign add_791960 = sel_791957 + 8'h01;
  assign sel_791961 = array_index_791644 == array_index_773110 ? add_791960 : sel_791957;
  assign add_791964 = sel_791961 + 8'h01;
  assign sel_791965 = array_index_791644 == array_index_773116 ? add_791964 : sel_791961;
  assign add_791968 = sel_791965 + 8'h01;
  assign sel_791969 = array_index_791644 == array_index_773122 ? add_791968 : sel_791965;
  assign add_791972 = sel_791969 + 8'h01;
  assign sel_791973 = array_index_791644 == array_index_773128 ? add_791972 : sel_791969;
  assign add_791976 = sel_791973 + 8'h01;
  assign sel_791977 = array_index_791644 == array_index_773134 ? add_791976 : sel_791973;
  assign add_791980 = sel_791977 + 8'h01;
  assign sel_791981 = array_index_791644 == array_index_773140 ? add_791980 : sel_791977;
  assign add_791984 = sel_791981 + 8'h01;
  assign sel_791985 = array_index_791644 == array_index_773146 ? add_791984 : sel_791981;
  assign add_791988 = sel_791985 + 8'h01;
  assign sel_791989 = array_index_791644 == array_index_773152 ? add_791988 : sel_791985;
  assign add_791992 = sel_791989 + 8'h01;
  assign sel_791993 = array_index_791644 == array_index_773158 ? add_791992 : sel_791989;
  assign add_791996 = sel_791993 + 8'h01;
  assign sel_791997 = array_index_791644 == array_index_773164 ? add_791996 : sel_791993;
  assign add_792000 = sel_791997 + 8'h01;
  assign sel_792001 = array_index_791644 == array_index_773170 ? add_792000 : sel_791997;
  assign add_792005 = sel_792001 + 8'h01;
  assign array_index_792006 = set1_unflattened[7'h35];
  assign sel_792007 = array_index_791644 == array_index_773176 ? add_792005 : sel_792001;
  assign add_792010 = sel_792007 + 8'h01;
  assign sel_792011 = array_index_792006 == array_index_772632 ? add_792010 : sel_792007;
  assign add_792014 = sel_792011 + 8'h01;
  assign sel_792015 = array_index_792006 == array_index_772636 ? add_792014 : sel_792011;
  assign add_792018 = sel_792015 + 8'h01;
  assign sel_792019 = array_index_792006 == array_index_772644 ? add_792018 : sel_792015;
  assign add_792022 = sel_792019 + 8'h01;
  assign sel_792023 = array_index_792006 == array_index_772652 ? add_792022 : sel_792019;
  assign add_792026 = sel_792023 + 8'h01;
  assign sel_792027 = array_index_792006 == array_index_772660 ? add_792026 : sel_792023;
  assign add_792030 = sel_792027 + 8'h01;
  assign sel_792031 = array_index_792006 == array_index_772668 ? add_792030 : sel_792027;
  assign add_792034 = sel_792031 + 8'h01;
  assign sel_792035 = array_index_792006 == array_index_772676 ? add_792034 : sel_792031;
  assign add_792038 = sel_792035 + 8'h01;
  assign sel_792039 = array_index_792006 == array_index_772684 ? add_792038 : sel_792035;
  assign add_792042 = sel_792039 + 8'h01;
  assign sel_792043 = array_index_792006 == array_index_772690 ? add_792042 : sel_792039;
  assign add_792046 = sel_792043 + 8'h01;
  assign sel_792047 = array_index_792006 == array_index_772696 ? add_792046 : sel_792043;
  assign add_792050 = sel_792047 + 8'h01;
  assign sel_792051 = array_index_792006 == array_index_772702 ? add_792050 : sel_792047;
  assign add_792054 = sel_792051 + 8'h01;
  assign sel_792055 = array_index_792006 == array_index_772708 ? add_792054 : sel_792051;
  assign add_792058 = sel_792055 + 8'h01;
  assign sel_792059 = array_index_792006 == array_index_772714 ? add_792058 : sel_792055;
  assign add_792062 = sel_792059 + 8'h01;
  assign sel_792063 = array_index_792006 == array_index_772720 ? add_792062 : sel_792059;
  assign add_792066 = sel_792063 + 8'h01;
  assign sel_792067 = array_index_792006 == array_index_772726 ? add_792066 : sel_792063;
  assign add_792070 = sel_792067 + 8'h01;
  assign sel_792071 = array_index_792006 == array_index_772732 ? add_792070 : sel_792067;
  assign add_792074 = sel_792071 + 8'h01;
  assign sel_792075 = array_index_792006 == array_index_772738 ? add_792074 : sel_792071;
  assign add_792078 = sel_792075 + 8'h01;
  assign sel_792079 = array_index_792006 == array_index_772744 ? add_792078 : sel_792075;
  assign add_792082 = sel_792079 + 8'h01;
  assign sel_792083 = array_index_792006 == array_index_772750 ? add_792082 : sel_792079;
  assign add_792086 = sel_792083 + 8'h01;
  assign sel_792087 = array_index_792006 == array_index_772756 ? add_792086 : sel_792083;
  assign add_792090 = sel_792087 + 8'h01;
  assign sel_792091 = array_index_792006 == array_index_772762 ? add_792090 : sel_792087;
  assign add_792094 = sel_792091 + 8'h01;
  assign sel_792095 = array_index_792006 == array_index_772768 ? add_792094 : sel_792091;
  assign add_792098 = sel_792095 + 8'h01;
  assign sel_792099 = array_index_792006 == array_index_772774 ? add_792098 : sel_792095;
  assign add_792102 = sel_792099 + 8'h01;
  assign sel_792103 = array_index_792006 == array_index_772780 ? add_792102 : sel_792099;
  assign add_792106 = sel_792103 + 8'h01;
  assign sel_792107 = array_index_792006 == array_index_772786 ? add_792106 : sel_792103;
  assign add_792110 = sel_792107 + 8'h01;
  assign sel_792111 = array_index_792006 == array_index_772792 ? add_792110 : sel_792107;
  assign add_792114 = sel_792111 + 8'h01;
  assign sel_792115 = array_index_792006 == array_index_772798 ? add_792114 : sel_792111;
  assign add_792118 = sel_792115 + 8'h01;
  assign sel_792119 = array_index_792006 == array_index_772804 ? add_792118 : sel_792115;
  assign add_792122 = sel_792119 + 8'h01;
  assign sel_792123 = array_index_792006 == array_index_772810 ? add_792122 : sel_792119;
  assign add_792126 = sel_792123 + 8'h01;
  assign sel_792127 = array_index_792006 == array_index_772816 ? add_792126 : sel_792123;
  assign add_792130 = sel_792127 + 8'h01;
  assign sel_792131 = array_index_792006 == array_index_772822 ? add_792130 : sel_792127;
  assign add_792134 = sel_792131 + 8'h01;
  assign sel_792135 = array_index_792006 == array_index_772828 ? add_792134 : sel_792131;
  assign add_792138 = sel_792135 + 8'h01;
  assign sel_792139 = array_index_792006 == array_index_772834 ? add_792138 : sel_792135;
  assign add_792142 = sel_792139 + 8'h01;
  assign sel_792143 = array_index_792006 == array_index_772840 ? add_792142 : sel_792139;
  assign add_792146 = sel_792143 + 8'h01;
  assign sel_792147 = array_index_792006 == array_index_772846 ? add_792146 : sel_792143;
  assign add_792150 = sel_792147 + 8'h01;
  assign sel_792151 = array_index_792006 == array_index_772852 ? add_792150 : sel_792147;
  assign add_792154 = sel_792151 + 8'h01;
  assign sel_792155 = array_index_792006 == array_index_772858 ? add_792154 : sel_792151;
  assign add_792158 = sel_792155 + 8'h01;
  assign sel_792159 = array_index_792006 == array_index_772864 ? add_792158 : sel_792155;
  assign add_792162 = sel_792159 + 8'h01;
  assign sel_792163 = array_index_792006 == array_index_772870 ? add_792162 : sel_792159;
  assign add_792166 = sel_792163 + 8'h01;
  assign sel_792167 = array_index_792006 == array_index_772876 ? add_792166 : sel_792163;
  assign add_792170 = sel_792167 + 8'h01;
  assign sel_792171 = array_index_792006 == array_index_772882 ? add_792170 : sel_792167;
  assign add_792174 = sel_792171 + 8'h01;
  assign sel_792175 = array_index_792006 == array_index_772888 ? add_792174 : sel_792171;
  assign add_792178 = sel_792175 + 8'h01;
  assign sel_792179 = array_index_792006 == array_index_772894 ? add_792178 : sel_792175;
  assign add_792182 = sel_792179 + 8'h01;
  assign sel_792183 = array_index_792006 == array_index_772900 ? add_792182 : sel_792179;
  assign add_792186 = sel_792183 + 8'h01;
  assign sel_792187 = array_index_792006 == array_index_772906 ? add_792186 : sel_792183;
  assign add_792190 = sel_792187 + 8'h01;
  assign sel_792191 = array_index_792006 == array_index_772912 ? add_792190 : sel_792187;
  assign add_792194 = sel_792191 + 8'h01;
  assign sel_792195 = array_index_792006 == array_index_772918 ? add_792194 : sel_792191;
  assign add_792198 = sel_792195 + 8'h01;
  assign sel_792199 = array_index_792006 == array_index_772924 ? add_792198 : sel_792195;
  assign add_792202 = sel_792199 + 8'h01;
  assign sel_792203 = array_index_792006 == array_index_772930 ? add_792202 : sel_792199;
  assign add_792206 = sel_792203 + 8'h01;
  assign sel_792207 = array_index_792006 == array_index_772936 ? add_792206 : sel_792203;
  assign add_792210 = sel_792207 + 8'h01;
  assign sel_792211 = array_index_792006 == array_index_772942 ? add_792210 : sel_792207;
  assign add_792214 = sel_792211 + 8'h01;
  assign sel_792215 = array_index_792006 == array_index_772948 ? add_792214 : sel_792211;
  assign add_792218 = sel_792215 + 8'h01;
  assign sel_792219 = array_index_792006 == array_index_772954 ? add_792218 : sel_792215;
  assign add_792222 = sel_792219 + 8'h01;
  assign sel_792223 = array_index_792006 == array_index_772960 ? add_792222 : sel_792219;
  assign add_792226 = sel_792223 + 8'h01;
  assign sel_792227 = array_index_792006 == array_index_772966 ? add_792226 : sel_792223;
  assign add_792230 = sel_792227 + 8'h01;
  assign sel_792231 = array_index_792006 == array_index_772972 ? add_792230 : sel_792227;
  assign add_792234 = sel_792231 + 8'h01;
  assign sel_792235 = array_index_792006 == array_index_772978 ? add_792234 : sel_792231;
  assign add_792238 = sel_792235 + 8'h01;
  assign sel_792239 = array_index_792006 == array_index_772984 ? add_792238 : sel_792235;
  assign add_792242 = sel_792239 + 8'h01;
  assign sel_792243 = array_index_792006 == array_index_772990 ? add_792242 : sel_792239;
  assign add_792246 = sel_792243 + 8'h01;
  assign sel_792247 = array_index_792006 == array_index_772996 ? add_792246 : sel_792243;
  assign add_792250 = sel_792247 + 8'h01;
  assign sel_792251 = array_index_792006 == array_index_773002 ? add_792250 : sel_792247;
  assign add_792254 = sel_792251 + 8'h01;
  assign sel_792255 = array_index_792006 == array_index_773008 ? add_792254 : sel_792251;
  assign add_792258 = sel_792255 + 8'h01;
  assign sel_792259 = array_index_792006 == array_index_773014 ? add_792258 : sel_792255;
  assign add_792262 = sel_792259 + 8'h01;
  assign sel_792263 = array_index_792006 == array_index_773020 ? add_792262 : sel_792259;
  assign add_792266 = sel_792263 + 8'h01;
  assign sel_792267 = array_index_792006 == array_index_773026 ? add_792266 : sel_792263;
  assign add_792270 = sel_792267 + 8'h01;
  assign sel_792271 = array_index_792006 == array_index_773032 ? add_792270 : sel_792267;
  assign add_792274 = sel_792271 + 8'h01;
  assign sel_792275 = array_index_792006 == array_index_773038 ? add_792274 : sel_792271;
  assign add_792278 = sel_792275 + 8'h01;
  assign sel_792279 = array_index_792006 == array_index_773044 ? add_792278 : sel_792275;
  assign add_792282 = sel_792279 + 8'h01;
  assign sel_792283 = array_index_792006 == array_index_773050 ? add_792282 : sel_792279;
  assign add_792286 = sel_792283 + 8'h01;
  assign sel_792287 = array_index_792006 == array_index_773056 ? add_792286 : sel_792283;
  assign add_792290 = sel_792287 + 8'h01;
  assign sel_792291 = array_index_792006 == array_index_773062 ? add_792290 : sel_792287;
  assign add_792294 = sel_792291 + 8'h01;
  assign sel_792295 = array_index_792006 == array_index_773068 ? add_792294 : sel_792291;
  assign add_792298 = sel_792295 + 8'h01;
  assign sel_792299 = array_index_792006 == array_index_773074 ? add_792298 : sel_792295;
  assign add_792302 = sel_792299 + 8'h01;
  assign sel_792303 = array_index_792006 == array_index_773080 ? add_792302 : sel_792299;
  assign add_792306 = sel_792303 + 8'h01;
  assign sel_792307 = array_index_792006 == array_index_773086 ? add_792306 : sel_792303;
  assign add_792310 = sel_792307 + 8'h01;
  assign sel_792311 = array_index_792006 == array_index_773092 ? add_792310 : sel_792307;
  assign add_792314 = sel_792311 + 8'h01;
  assign sel_792315 = array_index_792006 == array_index_773098 ? add_792314 : sel_792311;
  assign add_792318 = sel_792315 + 8'h01;
  assign sel_792319 = array_index_792006 == array_index_773104 ? add_792318 : sel_792315;
  assign add_792322 = sel_792319 + 8'h01;
  assign sel_792323 = array_index_792006 == array_index_773110 ? add_792322 : sel_792319;
  assign add_792326 = sel_792323 + 8'h01;
  assign sel_792327 = array_index_792006 == array_index_773116 ? add_792326 : sel_792323;
  assign add_792330 = sel_792327 + 8'h01;
  assign sel_792331 = array_index_792006 == array_index_773122 ? add_792330 : sel_792327;
  assign add_792334 = sel_792331 + 8'h01;
  assign sel_792335 = array_index_792006 == array_index_773128 ? add_792334 : sel_792331;
  assign add_792338 = sel_792335 + 8'h01;
  assign sel_792339 = array_index_792006 == array_index_773134 ? add_792338 : sel_792335;
  assign add_792342 = sel_792339 + 8'h01;
  assign sel_792343 = array_index_792006 == array_index_773140 ? add_792342 : sel_792339;
  assign add_792346 = sel_792343 + 8'h01;
  assign sel_792347 = array_index_792006 == array_index_773146 ? add_792346 : sel_792343;
  assign add_792350 = sel_792347 + 8'h01;
  assign sel_792351 = array_index_792006 == array_index_773152 ? add_792350 : sel_792347;
  assign add_792354 = sel_792351 + 8'h01;
  assign sel_792355 = array_index_792006 == array_index_773158 ? add_792354 : sel_792351;
  assign add_792358 = sel_792355 + 8'h01;
  assign sel_792359 = array_index_792006 == array_index_773164 ? add_792358 : sel_792355;
  assign add_792362 = sel_792359 + 8'h01;
  assign sel_792363 = array_index_792006 == array_index_773170 ? add_792362 : sel_792359;
  assign add_792367 = sel_792363 + 8'h01;
  assign array_index_792368 = set1_unflattened[7'h36];
  assign sel_792369 = array_index_792006 == array_index_773176 ? add_792367 : sel_792363;
  assign add_792372 = sel_792369 + 8'h01;
  assign sel_792373 = array_index_792368 == array_index_772632 ? add_792372 : sel_792369;
  assign add_792376 = sel_792373 + 8'h01;
  assign sel_792377 = array_index_792368 == array_index_772636 ? add_792376 : sel_792373;
  assign add_792380 = sel_792377 + 8'h01;
  assign sel_792381 = array_index_792368 == array_index_772644 ? add_792380 : sel_792377;
  assign add_792384 = sel_792381 + 8'h01;
  assign sel_792385 = array_index_792368 == array_index_772652 ? add_792384 : sel_792381;
  assign add_792388 = sel_792385 + 8'h01;
  assign sel_792389 = array_index_792368 == array_index_772660 ? add_792388 : sel_792385;
  assign add_792392 = sel_792389 + 8'h01;
  assign sel_792393 = array_index_792368 == array_index_772668 ? add_792392 : sel_792389;
  assign add_792396 = sel_792393 + 8'h01;
  assign sel_792397 = array_index_792368 == array_index_772676 ? add_792396 : sel_792393;
  assign add_792400 = sel_792397 + 8'h01;
  assign sel_792401 = array_index_792368 == array_index_772684 ? add_792400 : sel_792397;
  assign add_792404 = sel_792401 + 8'h01;
  assign sel_792405 = array_index_792368 == array_index_772690 ? add_792404 : sel_792401;
  assign add_792408 = sel_792405 + 8'h01;
  assign sel_792409 = array_index_792368 == array_index_772696 ? add_792408 : sel_792405;
  assign add_792412 = sel_792409 + 8'h01;
  assign sel_792413 = array_index_792368 == array_index_772702 ? add_792412 : sel_792409;
  assign add_792416 = sel_792413 + 8'h01;
  assign sel_792417 = array_index_792368 == array_index_772708 ? add_792416 : sel_792413;
  assign add_792420 = sel_792417 + 8'h01;
  assign sel_792421 = array_index_792368 == array_index_772714 ? add_792420 : sel_792417;
  assign add_792424 = sel_792421 + 8'h01;
  assign sel_792425 = array_index_792368 == array_index_772720 ? add_792424 : sel_792421;
  assign add_792428 = sel_792425 + 8'h01;
  assign sel_792429 = array_index_792368 == array_index_772726 ? add_792428 : sel_792425;
  assign add_792432 = sel_792429 + 8'h01;
  assign sel_792433 = array_index_792368 == array_index_772732 ? add_792432 : sel_792429;
  assign add_792436 = sel_792433 + 8'h01;
  assign sel_792437 = array_index_792368 == array_index_772738 ? add_792436 : sel_792433;
  assign add_792440 = sel_792437 + 8'h01;
  assign sel_792441 = array_index_792368 == array_index_772744 ? add_792440 : sel_792437;
  assign add_792444 = sel_792441 + 8'h01;
  assign sel_792445 = array_index_792368 == array_index_772750 ? add_792444 : sel_792441;
  assign add_792448 = sel_792445 + 8'h01;
  assign sel_792449 = array_index_792368 == array_index_772756 ? add_792448 : sel_792445;
  assign add_792452 = sel_792449 + 8'h01;
  assign sel_792453 = array_index_792368 == array_index_772762 ? add_792452 : sel_792449;
  assign add_792456 = sel_792453 + 8'h01;
  assign sel_792457 = array_index_792368 == array_index_772768 ? add_792456 : sel_792453;
  assign add_792460 = sel_792457 + 8'h01;
  assign sel_792461 = array_index_792368 == array_index_772774 ? add_792460 : sel_792457;
  assign add_792464 = sel_792461 + 8'h01;
  assign sel_792465 = array_index_792368 == array_index_772780 ? add_792464 : sel_792461;
  assign add_792468 = sel_792465 + 8'h01;
  assign sel_792469 = array_index_792368 == array_index_772786 ? add_792468 : sel_792465;
  assign add_792472 = sel_792469 + 8'h01;
  assign sel_792473 = array_index_792368 == array_index_772792 ? add_792472 : sel_792469;
  assign add_792476 = sel_792473 + 8'h01;
  assign sel_792477 = array_index_792368 == array_index_772798 ? add_792476 : sel_792473;
  assign add_792480 = sel_792477 + 8'h01;
  assign sel_792481 = array_index_792368 == array_index_772804 ? add_792480 : sel_792477;
  assign add_792484 = sel_792481 + 8'h01;
  assign sel_792485 = array_index_792368 == array_index_772810 ? add_792484 : sel_792481;
  assign add_792488 = sel_792485 + 8'h01;
  assign sel_792489 = array_index_792368 == array_index_772816 ? add_792488 : sel_792485;
  assign add_792492 = sel_792489 + 8'h01;
  assign sel_792493 = array_index_792368 == array_index_772822 ? add_792492 : sel_792489;
  assign add_792496 = sel_792493 + 8'h01;
  assign sel_792497 = array_index_792368 == array_index_772828 ? add_792496 : sel_792493;
  assign add_792500 = sel_792497 + 8'h01;
  assign sel_792501 = array_index_792368 == array_index_772834 ? add_792500 : sel_792497;
  assign add_792504 = sel_792501 + 8'h01;
  assign sel_792505 = array_index_792368 == array_index_772840 ? add_792504 : sel_792501;
  assign add_792508 = sel_792505 + 8'h01;
  assign sel_792509 = array_index_792368 == array_index_772846 ? add_792508 : sel_792505;
  assign add_792512 = sel_792509 + 8'h01;
  assign sel_792513 = array_index_792368 == array_index_772852 ? add_792512 : sel_792509;
  assign add_792516 = sel_792513 + 8'h01;
  assign sel_792517 = array_index_792368 == array_index_772858 ? add_792516 : sel_792513;
  assign add_792520 = sel_792517 + 8'h01;
  assign sel_792521 = array_index_792368 == array_index_772864 ? add_792520 : sel_792517;
  assign add_792524 = sel_792521 + 8'h01;
  assign sel_792525 = array_index_792368 == array_index_772870 ? add_792524 : sel_792521;
  assign add_792528 = sel_792525 + 8'h01;
  assign sel_792529 = array_index_792368 == array_index_772876 ? add_792528 : sel_792525;
  assign add_792532 = sel_792529 + 8'h01;
  assign sel_792533 = array_index_792368 == array_index_772882 ? add_792532 : sel_792529;
  assign add_792536 = sel_792533 + 8'h01;
  assign sel_792537 = array_index_792368 == array_index_772888 ? add_792536 : sel_792533;
  assign add_792540 = sel_792537 + 8'h01;
  assign sel_792541 = array_index_792368 == array_index_772894 ? add_792540 : sel_792537;
  assign add_792544 = sel_792541 + 8'h01;
  assign sel_792545 = array_index_792368 == array_index_772900 ? add_792544 : sel_792541;
  assign add_792548 = sel_792545 + 8'h01;
  assign sel_792549 = array_index_792368 == array_index_772906 ? add_792548 : sel_792545;
  assign add_792552 = sel_792549 + 8'h01;
  assign sel_792553 = array_index_792368 == array_index_772912 ? add_792552 : sel_792549;
  assign add_792556 = sel_792553 + 8'h01;
  assign sel_792557 = array_index_792368 == array_index_772918 ? add_792556 : sel_792553;
  assign add_792560 = sel_792557 + 8'h01;
  assign sel_792561 = array_index_792368 == array_index_772924 ? add_792560 : sel_792557;
  assign add_792564 = sel_792561 + 8'h01;
  assign sel_792565 = array_index_792368 == array_index_772930 ? add_792564 : sel_792561;
  assign add_792568 = sel_792565 + 8'h01;
  assign sel_792569 = array_index_792368 == array_index_772936 ? add_792568 : sel_792565;
  assign add_792572 = sel_792569 + 8'h01;
  assign sel_792573 = array_index_792368 == array_index_772942 ? add_792572 : sel_792569;
  assign add_792576 = sel_792573 + 8'h01;
  assign sel_792577 = array_index_792368 == array_index_772948 ? add_792576 : sel_792573;
  assign add_792580 = sel_792577 + 8'h01;
  assign sel_792581 = array_index_792368 == array_index_772954 ? add_792580 : sel_792577;
  assign add_792584 = sel_792581 + 8'h01;
  assign sel_792585 = array_index_792368 == array_index_772960 ? add_792584 : sel_792581;
  assign add_792588 = sel_792585 + 8'h01;
  assign sel_792589 = array_index_792368 == array_index_772966 ? add_792588 : sel_792585;
  assign add_792592 = sel_792589 + 8'h01;
  assign sel_792593 = array_index_792368 == array_index_772972 ? add_792592 : sel_792589;
  assign add_792596 = sel_792593 + 8'h01;
  assign sel_792597 = array_index_792368 == array_index_772978 ? add_792596 : sel_792593;
  assign add_792600 = sel_792597 + 8'h01;
  assign sel_792601 = array_index_792368 == array_index_772984 ? add_792600 : sel_792597;
  assign add_792604 = sel_792601 + 8'h01;
  assign sel_792605 = array_index_792368 == array_index_772990 ? add_792604 : sel_792601;
  assign add_792608 = sel_792605 + 8'h01;
  assign sel_792609 = array_index_792368 == array_index_772996 ? add_792608 : sel_792605;
  assign add_792612 = sel_792609 + 8'h01;
  assign sel_792613 = array_index_792368 == array_index_773002 ? add_792612 : sel_792609;
  assign add_792616 = sel_792613 + 8'h01;
  assign sel_792617 = array_index_792368 == array_index_773008 ? add_792616 : sel_792613;
  assign add_792620 = sel_792617 + 8'h01;
  assign sel_792621 = array_index_792368 == array_index_773014 ? add_792620 : sel_792617;
  assign add_792624 = sel_792621 + 8'h01;
  assign sel_792625 = array_index_792368 == array_index_773020 ? add_792624 : sel_792621;
  assign add_792628 = sel_792625 + 8'h01;
  assign sel_792629 = array_index_792368 == array_index_773026 ? add_792628 : sel_792625;
  assign add_792632 = sel_792629 + 8'h01;
  assign sel_792633 = array_index_792368 == array_index_773032 ? add_792632 : sel_792629;
  assign add_792636 = sel_792633 + 8'h01;
  assign sel_792637 = array_index_792368 == array_index_773038 ? add_792636 : sel_792633;
  assign add_792640 = sel_792637 + 8'h01;
  assign sel_792641 = array_index_792368 == array_index_773044 ? add_792640 : sel_792637;
  assign add_792644 = sel_792641 + 8'h01;
  assign sel_792645 = array_index_792368 == array_index_773050 ? add_792644 : sel_792641;
  assign add_792648 = sel_792645 + 8'h01;
  assign sel_792649 = array_index_792368 == array_index_773056 ? add_792648 : sel_792645;
  assign add_792652 = sel_792649 + 8'h01;
  assign sel_792653 = array_index_792368 == array_index_773062 ? add_792652 : sel_792649;
  assign add_792656 = sel_792653 + 8'h01;
  assign sel_792657 = array_index_792368 == array_index_773068 ? add_792656 : sel_792653;
  assign add_792660 = sel_792657 + 8'h01;
  assign sel_792661 = array_index_792368 == array_index_773074 ? add_792660 : sel_792657;
  assign add_792664 = sel_792661 + 8'h01;
  assign sel_792665 = array_index_792368 == array_index_773080 ? add_792664 : sel_792661;
  assign add_792668 = sel_792665 + 8'h01;
  assign sel_792669 = array_index_792368 == array_index_773086 ? add_792668 : sel_792665;
  assign add_792672 = sel_792669 + 8'h01;
  assign sel_792673 = array_index_792368 == array_index_773092 ? add_792672 : sel_792669;
  assign add_792676 = sel_792673 + 8'h01;
  assign sel_792677 = array_index_792368 == array_index_773098 ? add_792676 : sel_792673;
  assign add_792680 = sel_792677 + 8'h01;
  assign sel_792681 = array_index_792368 == array_index_773104 ? add_792680 : sel_792677;
  assign add_792684 = sel_792681 + 8'h01;
  assign sel_792685 = array_index_792368 == array_index_773110 ? add_792684 : sel_792681;
  assign add_792688 = sel_792685 + 8'h01;
  assign sel_792689 = array_index_792368 == array_index_773116 ? add_792688 : sel_792685;
  assign add_792692 = sel_792689 + 8'h01;
  assign sel_792693 = array_index_792368 == array_index_773122 ? add_792692 : sel_792689;
  assign add_792696 = sel_792693 + 8'h01;
  assign sel_792697 = array_index_792368 == array_index_773128 ? add_792696 : sel_792693;
  assign add_792700 = sel_792697 + 8'h01;
  assign sel_792701 = array_index_792368 == array_index_773134 ? add_792700 : sel_792697;
  assign add_792704 = sel_792701 + 8'h01;
  assign sel_792705 = array_index_792368 == array_index_773140 ? add_792704 : sel_792701;
  assign add_792708 = sel_792705 + 8'h01;
  assign sel_792709 = array_index_792368 == array_index_773146 ? add_792708 : sel_792705;
  assign add_792712 = sel_792709 + 8'h01;
  assign sel_792713 = array_index_792368 == array_index_773152 ? add_792712 : sel_792709;
  assign add_792716 = sel_792713 + 8'h01;
  assign sel_792717 = array_index_792368 == array_index_773158 ? add_792716 : sel_792713;
  assign add_792720 = sel_792717 + 8'h01;
  assign sel_792721 = array_index_792368 == array_index_773164 ? add_792720 : sel_792717;
  assign add_792724 = sel_792721 + 8'h01;
  assign sel_792725 = array_index_792368 == array_index_773170 ? add_792724 : sel_792721;
  assign add_792729 = sel_792725 + 8'h01;
  assign array_index_792730 = set1_unflattened[7'h37];
  assign sel_792731 = array_index_792368 == array_index_773176 ? add_792729 : sel_792725;
  assign add_792734 = sel_792731 + 8'h01;
  assign sel_792735 = array_index_792730 == array_index_772632 ? add_792734 : sel_792731;
  assign add_792738 = sel_792735 + 8'h01;
  assign sel_792739 = array_index_792730 == array_index_772636 ? add_792738 : sel_792735;
  assign add_792742 = sel_792739 + 8'h01;
  assign sel_792743 = array_index_792730 == array_index_772644 ? add_792742 : sel_792739;
  assign add_792746 = sel_792743 + 8'h01;
  assign sel_792747 = array_index_792730 == array_index_772652 ? add_792746 : sel_792743;
  assign add_792750 = sel_792747 + 8'h01;
  assign sel_792751 = array_index_792730 == array_index_772660 ? add_792750 : sel_792747;
  assign add_792754 = sel_792751 + 8'h01;
  assign sel_792755 = array_index_792730 == array_index_772668 ? add_792754 : sel_792751;
  assign add_792758 = sel_792755 + 8'h01;
  assign sel_792759 = array_index_792730 == array_index_772676 ? add_792758 : sel_792755;
  assign add_792762 = sel_792759 + 8'h01;
  assign sel_792763 = array_index_792730 == array_index_772684 ? add_792762 : sel_792759;
  assign add_792766 = sel_792763 + 8'h01;
  assign sel_792767 = array_index_792730 == array_index_772690 ? add_792766 : sel_792763;
  assign add_792770 = sel_792767 + 8'h01;
  assign sel_792771 = array_index_792730 == array_index_772696 ? add_792770 : sel_792767;
  assign add_792774 = sel_792771 + 8'h01;
  assign sel_792775 = array_index_792730 == array_index_772702 ? add_792774 : sel_792771;
  assign add_792778 = sel_792775 + 8'h01;
  assign sel_792779 = array_index_792730 == array_index_772708 ? add_792778 : sel_792775;
  assign add_792782 = sel_792779 + 8'h01;
  assign sel_792783 = array_index_792730 == array_index_772714 ? add_792782 : sel_792779;
  assign add_792786 = sel_792783 + 8'h01;
  assign sel_792787 = array_index_792730 == array_index_772720 ? add_792786 : sel_792783;
  assign add_792790 = sel_792787 + 8'h01;
  assign sel_792791 = array_index_792730 == array_index_772726 ? add_792790 : sel_792787;
  assign add_792794 = sel_792791 + 8'h01;
  assign sel_792795 = array_index_792730 == array_index_772732 ? add_792794 : sel_792791;
  assign add_792798 = sel_792795 + 8'h01;
  assign sel_792799 = array_index_792730 == array_index_772738 ? add_792798 : sel_792795;
  assign add_792802 = sel_792799 + 8'h01;
  assign sel_792803 = array_index_792730 == array_index_772744 ? add_792802 : sel_792799;
  assign add_792806 = sel_792803 + 8'h01;
  assign sel_792807 = array_index_792730 == array_index_772750 ? add_792806 : sel_792803;
  assign add_792810 = sel_792807 + 8'h01;
  assign sel_792811 = array_index_792730 == array_index_772756 ? add_792810 : sel_792807;
  assign add_792814 = sel_792811 + 8'h01;
  assign sel_792815 = array_index_792730 == array_index_772762 ? add_792814 : sel_792811;
  assign add_792818 = sel_792815 + 8'h01;
  assign sel_792819 = array_index_792730 == array_index_772768 ? add_792818 : sel_792815;
  assign add_792822 = sel_792819 + 8'h01;
  assign sel_792823 = array_index_792730 == array_index_772774 ? add_792822 : sel_792819;
  assign add_792826 = sel_792823 + 8'h01;
  assign sel_792827 = array_index_792730 == array_index_772780 ? add_792826 : sel_792823;
  assign add_792830 = sel_792827 + 8'h01;
  assign sel_792831 = array_index_792730 == array_index_772786 ? add_792830 : sel_792827;
  assign add_792834 = sel_792831 + 8'h01;
  assign sel_792835 = array_index_792730 == array_index_772792 ? add_792834 : sel_792831;
  assign add_792838 = sel_792835 + 8'h01;
  assign sel_792839 = array_index_792730 == array_index_772798 ? add_792838 : sel_792835;
  assign add_792842 = sel_792839 + 8'h01;
  assign sel_792843 = array_index_792730 == array_index_772804 ? add_792842 : sel_792839;
  assign add_792846 = sel_792843 + 8'h01;
  assign sel_792847 = array_index_792730 == array_index_772810 ? add_792846 : sel_792843;
  assign add_792850 = sel_792847 + 8'h01;
  assign sel_792851 = array_index_792730 == array_index_772816 ? add_792850 : sel_792847;
  assign add_792854 = sel_792851 + 8'h01;
  assign sel_792855 = array_index_792730 == array_index_772822 ? add_792854 : sel_792851;
  assign add_792858 = sel_792855 + 8'h01;
  assign sel_792859 = array_index_792730 == array_index_772828 ? add_792858 : sel_792855;
  assign add_792862 = sel_792859 + 8'h01;
  assign sel_792863 = array_index_792730 == array_index_772834 ? add_792862 : sel_792859;
  assign add_792866 = sel_792863 + 8'h01;
  assign sel_792867 = array_index_792730 == array_index_772840 ? add_792866 : sel_792863;
  assign add_792870 = sel_792867 + 8'h01;
  assign sel_792871 = array_index_792730 == array_index_772846 ? add_792870 : sel_792867;
  assign add_792874 = sel_792871 + 8'h01;
  assign sel_792875 = array_index_792730 == array_index_772852 ? add_792874 : sel_792871;
  assign add_792878 = sel_792875 + 8'h01;
  assign sel_792879 = array_index_792730 == array_index_772858 ? add_792878 : sel_792875;
  assign add_792882 = sel_792879 + 8'h01;
  assign sel_792883 = array_index_792730 == array_index_772864 ? add_792882 : sel_792879;
  assign add_792886 = sel_792883 + 8'h01;
  assign sel_792887 = array_index_792730 == array_index_772870 ? add_792886 : sel_792883;
  assign add_792890 = sel_792887 + 8'h01;
  assign sel_792891 = array_index_792730 == array_index_772876 ? add_792890 : sel_792887;
  assign add_792894 = sel_792891 + 8'h01;
  assign sel_792895 = array_index_792730 == array_index_772882 ? add_792894 : sel_792891;
  assign add_792898 = sel_792895 + 8'h01;
  assign sel_792899 = array_index_792730 == array_index_772888 ? add_792898 : sel_792895;
  assign add_792902 = sel_792899 + 8'h01;
  assign sel_792903 = array_index_792730 == array_index_772894 ? add_792902 : sel_792899;
  assign add_792906 = sel_792903 + 8'h01;
  assign sel_792907 = array_index_792730 == array_index_772900 ? add_792906 : sel_792903;
  assign add_792910 = sel_792907 + 8'h01;
  assign sel_792911 = array_index_792730 == array_index_772906 ? add_792910 : sel_792907;
  assign add_792914 = sel_792911 + 8'h01;
  assign sel_792915 = array_index_792730 == array_index_772912 ? add_792914 : sel_792911;
  assign add_792918 = sel_792915 + 8'h01;
  assign sel_792919 = array_index_792730 == array_index_772918 ? add_792918 : sel_792915;
  assign add_792922 = sel_792919 + 8'h01;
  assign sel_792923 = array_index_792730 == array_index_772924 ? add_792922 : sel_792919;
  assign add_792926 = sel_792923 + 8'h01;
  assign sel_792927 = array_index_792730 == array_index_772930 ? add_792926 : sel_792923;
  assign add_792930 = sel_792927 + 8'h01;
  assign sel_792931 = array_index_792730 == array_index_772936 ? add_792930 : sel_792927;
  assign add_792934 = sel_792931 + 8'h01;
  assign sel_792935 = array_index_792730 == array_index_772942 ? add_792934 : sel_792931;
  assign add_792938 = sel_792935 + 8'h01;
  assign sel_792939 = array_index_792730 == array_index_772948 ? add_792938 : sel_792935;
  assign add_792942 = sel_792939 + 8'h01;
  assign sel_792943 = array_index_792730 == array_index_772954 ? add_792942 : sel_792939;
  assign add_792946 = sel_792943 + 8'h01;
  assign sel_792947 = array_index_792730 == array_index_772960 ? add_792946 : sel_792943;
  assign add_792950 = sel_792947 + 8'h01;
  assign sel_792951 = array_index_792730 == array_index_772966 ? add_792950 : sel_792947;
  assign add_792954 = sel_792951 + 8'h01;
  assign sel_792955 = array_index_792730 == array_index_772972 ? add_792954 : sel_792951;
  assign add_792958 = sel_792955 + 8'h01;
  assign sel_792959 = array_index_792730 == array_index_772978 ? add_792958 : sel_792955;
  assign add_792962 = sel_792959 + 8'h01;
  assign sel_792963 = array_index_792730 == array_index_772984 ? add_792962 : sel_792959;
  assign add_792966 = sel_792963 + 8'h01;
  assign sel_792967 = array_index_792730 == array_index_772990 ? add_792966 : sel_792963;
  assign add_792970 = sel_792967 + 8'h01;
  assign sel_792971 = array_index_792730 == array_index_772996 ? add_792970 : sel_792967;
  assign add_792974 = sel_792971 + 8'h01;
  assign sel_792975 = array_index_792730 == array_index_773002 ? add_792974 : sel_792971;
  assign add_792978 = sel_792975 + 8'h01;
  assign sel_792979 = array_index_792730 == array_index_773008 ? add_792978 : sel_792975;
  assign add_792982 = sel_792979 + 8'h01;
  assign sel_792983 = array_index_792730 == array_index_773014 ? add_792982 : sel_792979;
  assign add_792986 = sel_792983 + 8'h01;
  assign sel_792987 = array_index_792730 == array_index_773020 ? add_792986 : sel_792983;
  assign add_792990 = sel_792987 + 8'h01;
  assign sel_792991 = array_index_792730 == array_index_773026 ? add_792990 : sel_792987;
  assign add_792994 = sel_792991 + 8'h01;
  assign sel_792995 = array_index_792730 == array_index_773032 ? add_792994 : sel_792991;
  assign add_792998 = sel_792995 + 8'h01;
  assign sel_792999 = array_index_792730 == array_index_773038 ? add_792998 : sel_792995;
  assign add_793002 = sel_792999 + 8'h01;
  assign sel_793003 = array_index_792730 == array_index_773044 ? add_793002 : sel_792999;
  assign add_793006 = sel_793003 + 8'h01;
  assign sel_793007 = array_index_792730 == array_index_773050 ? add_793006 : sel_793003;
  assign add_793010 = sel_793007 + 8'h01;
  assign sel_793011 = array_index_792730 == array_index_773056 ? add_793010 : sel_793007;
  assign add_793014 = sel_793011 + 8'h01;
  assign sel_793015 = array_index_792730 == array_index_773062 ? add_793014 : sel_793011;
  assign add_793018 = sel_793015 + 8'h01;
  assign sel_793019 = array_index_792730 == array_index_773068 ? add_793018 : sel_793015;
  assign add_793022 = sel_793019 + 8'h01;
  assign sel_793023 = array_index_792730 == array_index_773074 ? add_793022 : sel_793019;
  assign add_793026 = sel_793023 + 8'h01;
  assign sel_793027 = array_index_792730 == array_index_773080 ? add_793026 : sel_793023;
  assign add_793030 = sel_793027 + 8'h01;
  assign sel_793031 = array_index_792730 == array_index_773086 ? add_793030 : sel_793027;
  assign add_793034 = sel_793031 + 8'h01;
  assign sel_793035 = array_index_792730 == array_index_773092 ? add_793034 : sel_793031;
  assign add_793038 = sel_793035 + 8'h01;
  assign sel_793039 = array_index_792730 == array_index_773098 ? add_793038 : sel_793035;
  assign add_793042 = sel_793039 + 8'h01;
  assign sel_793043 = array_index_792730 == array_index_773104 ? add_793042 : sel_793039;
  assign add_793046 = sel_793043 + 8'h01;
  assign sel_793047 = array_index_792730 == array_index_773110 ? add_793046 : sel_793043;
  assign add_793050 = sel_793047 + 8'h01;
  assign sel_793051 = array_index_792730 == array_index_773116 ? add_793050 : sel_793047;
  assign add_793054 = sel_793051 + 8'h01;
  assign sel_793055 = array_index_792730 == array_index_773122 ? add_793054 : sel_793051;
  assign add_793058 = sel_793055 + 8'h01;
  assign sel_793059 = array_index_792730 == array_index_773128 ? add_793058 : sel_793055;
  assign add_793062 = sel_793059 + 8'h01;
  assign sel_793063 = array_index_792730 == array_index_773134 ? add_793062 : sel_793059;
  assign add_793066 = sel_793063 + 8'h01;
  assign sel_793067 = array_index_792730 == array_index_773140 ? add_793066 : sel_793063;
  assign add_793070 = sel_793067 + 8'h01;
  assign sel_793071 = array_index_792730 == array_index_773146 ? add_793070 : sel_793067;
  assign add_793074 = sel_793071 + 8'h01;
  assign sel_793075 = array_index_792730 == array_index_773152 ? add_793074 : sel_793071;
  assign add_793078 = sel_793075 + 8'h01;
  assign sel_793079 = array_index_792730 == array_index_773158 ? add_793078 : sel_793075;
  assign add_793082 = sel_793079 + 8'h01;
  assign sel_793083 = array_index_792730 == array_index_773164 ? add_793082 : sel_793079;
  assign add_793086 = sel_793083 + 8'h01;
  assign sel_793087 = array_index_792730 == array_index_773170 ? add_793086 : sel_793083;
  assign add_793091 = sel_793087 + 8'h01;
  assign array_index_793092 = set1_unflattened[7'h38];
  assign sel_793093 = array_index_792730 == array_index_773176 ? add_793091 : sel_793087;
  assign add_793096 = sel_793093 + 8'h01;
  assign sel_793097 = array_index_793092 == array_index_772632 ? add_793096 : sel_793093;
  assign add_793100 = sel_793097 + 8'h01;
  assign sel_793101 = array_index_793092 == array_index_772636 ? add_793100 : sel_793097;
  assign add_793104 = sel_793101 + 8'h01;
  assign sel_793105 = array_index_793092 == array_index_772644 ? add_793104 : sel_793101;
  assign add_793108 = sel_793105 + 8'h01;
  assign sel_793109 = array_index_793092 == array_index_772652 ? add_793108 : sel_793105;
  assign add_793112 = sel_793109 + 8'h01;
  assign sel_793113 = array_index_793092 == array_index_772660 ? add_793112 : sel_793109;
  assign add_793116 = sel_793113 + 8'h01;
  assign sel_793117 = array_index_793092 == array_index_772668 ? add_793116 : sel_793113;
  assign add_793120 = sel_793117 + 8'h01;
  assign sel_793121 = array_index_793092 == array_index_772676 ? add_793120 : sel_793117;
  assign add_793124 = sel_793121 + 8'h01;
  assign sel_793125 = array_index_793092 == array_index_772684 ? add_793124 : sel_793121;
  assign add_793128 = sel_793125 + 8'h01;
  assign sel_793129 = array_index_793092 == array_index_772690 ? add_793128 : sel_793125;
  assign add_793132 = sel_793129 + 8'h01;
  assign sel_793133 = array_index_793092 == array_index_772696 ? add_793132 : sel_793129;
  assign add_793136 = sel_793133 + 8'h01;
  assign sel_793137 = array_index_793092 == array_index_772702 ? add_793136 : sel_793133;
  assign add_793140 = sel_793137 + 8'h01;
  assign sel_793141 = array_index_793092 == array_index_772708 ? add_793140 : sel_793137;
  assign add_793144 = sel_793141 + 8'h01;
  assign sel_793145 = array_index_793092 == array_index_772714 ? add_793144 : sel_793141;
  assign add_793148 = sel_793145 + 8'h01;
  assign sel_793149 = array_index_793092 == array_index_772720 ? add_793148 : sel_793145;
  assign add_793152 = sel_793149 + 8'h01;
  assign sel_793153 = array_index_793092 == array_index_772726 ? add_793152 : sel_793149;
  assign add_793156 = sel_793153 + 8'h01;
  assign sel_793157 = array_index_793092 == array_index_772732 ? add_793156 : sel_793153;
  assign add_793160 = sel_793157 + 8'h01;
  assign sel_793161 = array_index_793092 == array_index_772738 ? add_793160 : sel_793157;
  assign add_793164 = sel_793161 + 8'h01;
  assign sel_793165 = array_index_793092 == array_index_772744 ? add_793164 : sel_793161;
  assign add_793168 = sel_793165 + 8'h01;
  assign sel_793169 = array_index_793092 == array_index_772750 ? add_793168 : sel_793165;
  assign add_793172 = sel_793169 + 8'h01;
  assign sel_793173 = array_index_793092 == array_index_772756 ? add_793172 : sel_793169;
  assign add_793176 = sel_793173 + 8'h01;
  assign sel_793177 = array_index_793092 == array_index_772762 ? add_793176 : sel_793173;
  assign add_793180 = sel_793177 + 8'h01;
  assign sel_793181 = array_index_793092 == array_index_772768 ? add_793180 : sel_793177;
  assign add_793184 = sel_793181 + 8'h01;
  assign sel_793185 = array_index_793092 == array_index_772774 ? add_793184 : sel_793181;
  assign add_793188 = sel_793185 + 8'h01;
  assign sel_793189 = array_index_793092 == array_index_772780 ? add_793188 : sel_793185;
  assign add_793192 = sel_793189 + 8'h01;
  assign sel_793193 = array_index_793092 == array_index_772786 ? add_793192 : sel_793189;
  assign add_793196 = sel_793193 + 8'h01;
  assign sel_793197 = array_index_793092 == array_index_772792 ? add_793196 : sel_793193;
  assign add_793200 = sel_793197 + 8'h01;
  assign sel_793201 = array_index_793092 == array_index_772798 ? add_793200 : sel_793197;
  assign add_793204 = sel_793201 + 8'h01;
  assign sel_793205 = array_index_793092 == array_index_772804 ? add_793204 : sel_793201;
  assign add_793208 = sel_793205 + 8'h01;
  assign sel_793209 = array_index_793092 == array_index_772810 ? add_793208 : sel_793205;
  assign add_793212 = sel_793209 + 8'h01;
  assign sel_793213 = array_index_793092 == array_index_772816 ? add_793212 : sel_793209;
  assign add_793216 = sel_793213 + 8'h01;
  assign sel_793217 = array_index_793092 == array_index_772822 ? add_793216 : sel_793213;
  assign add_793220 = sel_793217 + 8'h01;
  assign sel_793221 = array_index_793092 == array_index_772828 ? add_793220 : sel_793217;
  assign add_793224 = sel_793221 + 8'h01;
  assign sel_793225 = array_index_793092 == array_index_772834 ? add_793224 : sel_793221;
  assign add_793228 = sel_793225 + 8'h01;
  assign sel_793229 = array_index_793092 == array_index_772840 ? add_793228 : sel_793225;
  assign add_793232 = sel_793229 + 8'h01;
  assign sel_793233 = array_index_793092 == array_index_772846 ? add_793232 : sel_793229;
  assign add_793236 = sel_793233 + 8'h01;
  assign sel_793237 = array_index_793092 == array_index_772852 ? add_793236 : sel_793233;
  assign add_793240 = sel_793237 + 8'h01;
  assign sel_793241 = array_index_793092 == array_index_772858 ? add_793240 : sel_793237;
  assign add_793244 = sel_793241 + 8'h01;
  assign sel_793245 = array_index_793092 == array_index_772864 ? add_793244 : sel_793241;
  assign add_793248 = sel_793245 + 8'h01;
  assign sel_793249 = array_index_793092 == array_index_772870 ? add_793248 : sel_793245;
  assign add_793252 = sel_793249 + 8'h01;
  assign sel_793253 = array_index_793092 == array_index_772876 ? add_793252 : sel_793249;
  assign add_793256 = sel_793253 + 8'h01;
  assign sel_793257 = array_index_793092 == array_index_772882 ? add_793256 : sel_793253;
  assign add_793260 = sel_793257 + 8'h01;
  assign sel_793261 = array_index_793092 == array_index_772888 ? add_793260 : sel_793257;
  assign add_793264 = sel_793261 + 8'h01;
  assign sel_793265 = array_index_793092 == array_index_772894 ? add_793264 : sel_793261;
  assign add_793268 = sel_793265 + 8'h01;
  assign sel_793269 = array_index_793092 == array_index_772900 ? add_793268 : sel_793265;
  assign add_793272 = sel_793269 + 8'h01;
  assign sel_793273 = array_index_793092 == array_index_772906 ? add_793272 : sel_793269;
  assign add_793276 = sel_793273 + 8'h01;
  assign sel_793277 = array_index_793092 == array_index_772912 ? add_793276 : sel_793273;
  assign add_793280 = sel_793277 + 8'h01;
  assign sel_793281 = array_index_793092 == array_index_772918 ? add_793280 : sel_793277;
  assign add_793284 = sel_793281 + 8'h01;
  assign sel_793285 = array_index_793092 == array_index_772924 ? add_793284 : sel_793281;
  assign add_793288 = sel_793285 + 8'h01;
  assign sel_793289 = array_index_793092 == array_index_772930 ? add_793288 : sel_793285;
  assign add_793292 = sel_793289 + 8'h01;
  assign sel_793293 = array_index_793092 == array_index_772936 ? add_793292 : sel_793289;
  assign add_793296 = sel_793293 + 8'h01;
  assign sel_793297 = array_index_793092 == array_index_772942 ? add_793296 : sel_793293;
  assign add_793300 = sel_793297 + 8'h01;
  assign sel_793301 = array_index_793092 == array_index_772948 ? add_793300 : sel_793297;
  assign add_793304 = sel_793301 + 8'h01;
  assign sel_793305 = array_index_793092 == array_index_772954 ? add_793304 : sel_793301;
  assign add_793308 = sel_793305 + 8'h01;
  assign sel_793309 = array_index_793092 == array_index_772960 ? add_793308 : sel_793305;
  assign add_793312 = sel_793309 + 8'h01;
  assign sel_793313 = array_index_793092 == array_index_772966 ? add_793312 : sel_793309;
  assign add_793316 = sel_793313 + 8'h01;
  assign sel_793317 = array_index_793092 == array_index_772972 ? add_793316 : sel_793313;
  assign add_793320 = sel_793317 + 8'h01;
  assign sel_793321 = array_index_793092 == array_index_772978 ? add_793320 : sel_793317;
  assign add_793324 = sel_793321 + 8'h01;
  assign sel_793325 = array_index_793092 == array_index_772984 ? add_793324 : sel_793321;
  assign add_793328 = sel_793325 + 8'h01;
  assign sel_793329 = array_index_793092 == array_index_772990 ? add_793328 : sel_793325;
  assign add_793332 = sel_793329 + 8'h01;
  assign sel_793333 = array_index_793092 == array_index_772996 ? add_793332 : sel_793329;
  assign add_793336 = sel_793333 + 8'h01;
  assign sel_793337 = array_index_793092 == array_index_773002 ? add_793336 : sel_793333;
  assign add_793340 = sel_793337 + 8'h01;
  assign sel_793341 = array_index_793092 == array_index_773008 ? add_793340 : sel_793337;
  assign add_793344 = sel_793341 + 8'h01;
  assign sel_793345 = array_index_793092 == array_index_773014 ? add_793344 : sel_793341;
  assign add_793348 = sel_793345 + 8'h01;
  assign sel_793349 = array_index_793092 == array_index_773020 ? add_793348 : sel_793345;
  assign add_793352 = sel_793349 + 8'h01;
  assign sel_793353 = array_index_793092 == array_index_773026 ? add_793352 : sel_793349;
  assign add_793356 = sel_793353 + 8'h01;
  assign sel_793357 = array_index_793092 == array_index_773032 ? add_793356 : sel_793353;
  assign add_793360 = sel_793357 + 8'h01;
  assign sel_793361 = array_index_793092 == array_index_773038 ? add_793360 : sel_793357;
  assign add_793364 = sel_793361 + 8'h01;
  assign sel_793365 = array_index_793092 == array_index_773044 ? add_793364 : sel_793361;
  assign add_793368 = sel_793365 + 8'h01;
  assign sel_793369 = array_index_793092 == array_index_773050 ? add_793368 : sel_793365;
  assign add_793372 = sel_793369 + 8'h01;
  assign sel_793373 = array_index_793092 == array_index_773056 ? add_793372 : sel_793369;
  assign add_793376 = sel_793373 + 8'h01;
  assign sel_793377 = array_index_793092 == array_index_773062 ? add_793376 : sel_793373;
  assign add_793380 = sel_793377 + 8'h01;
  assign sel_793381 = array_index_793092 == array_index_773068 ? add_793380 : sel_793377;
  assign add_793384 = sel_793381 + 8'h01;
  assign sel_793385 = array_index_793092 == array_index_773074 ? add_793384 : sel_793381;
  assign add_793388 = sel_793385 + 8'h01;
  assign sel_793389 = array_index_793092 == array_index_773080 ? add_793388 : sel_793385;
  assign add_793392 = sel_793389 + 8'h01;
  assign sel_793393 = array_index_793092 == array_index_773086 ? add_793392 : sel_793389;
  assign add_793396 = sel_793393 + 8'h01;
  assign sel_793397 = array_index_793092 == array_index_773092 ? add_793396 : sel_793393;
  assign add_793400 = sel_793397 + 8'h01;
  assign sel_793401 = array_index_793092 == array_index_773098 ? add_793400 : sel_793397;
  assign add_793404 = sel_793401 + 8'h01;
  assign sel_793405 = array_index_793092 == array_index_773104 ? add_793404 : sel_793401;
  assign add_793408 = sel_793405 + 8'h01;
  assign sel_793409 = array_index_793092 == array_index_773110 ? add_793408 : sel_793405;
  assign add_793412 = sel_793409 + 8'h01;
  assign sel_793413 = array_index_793092 == array_index_773116 ? add_793412 : sel_793409;
  assign add_793416 = sel_793413 + 8'h01;
  assign sel_793417 = array_index_793092 == array_index_773122 ? add_793416 : sel_793413;
  assign add_793420 = sel_793417 + 8'h01;
  assign sel_793421 = array_index_793092 == array_index_773128 ? add_793420 : sel_793417;
  assign add_793424 = sel_793421 + 8'h01;
  assign sel_793425 = array_index_793092 == array_index_773134 ? add_793424 : sel_793421;
  assign add_793428 = sel_793425 + 8'h01;
  assign sel_793429 = array_index_793092 == array_index_773140 ? add_793428 : sel_793425;
  assign add_793432 = sel_793429 + 8'h01;
  assign sel_793433 = array_index_793092 == array_index_773146 ? add_793432 : sel_793429;
  assign add_793436 = sel_793433 + 8'h01;
  assign sel_793437 = array_index_793092 == array_index_773152 ? add_793436 : sel_793433;
  assign add_793440 = sel_793437 + 8'h01;
  assign sel_793441 = array_index_793092 == array_index_773158 ? add_793440 : sel_793437;
  assign add_793444 = sel_793441 + 8'h01;
  assign sel_793445 = array_index_793092 == array_index_773164 ? add_793444 : sel_793441;
  assign add_793448 = sel_793445 + 8'h01;
  assign sel_793449 = array_index_793092 == array_index_773170 ? add_793448 : sel_793445;
  assign add_793453 = sel_793449 + 8'h01;
  assign array_index_793454 = set1_unflattened[7'h39];
  assign sel_793455 = array_index_793092 == array_index_773176 ? add_793453 : sel_793449;
  assign add_793458 = sel_793455 + 8'h01;
  assign sel_793459 = array_index_793454 == array_index_772632 ? add_793458 : sel_793455;
  assign add_793462 = sel_793459 + 8'h01;
  assign sel_793463 = array_index_793454 == array_index_772636 ? add_793462 : sel_793459;
  assign add_793466 = sel_793463 + 8'h01;
  assign sel_793467 = array_index_793454 == array_index_772644 ? add_793466 : sel_793463;
  assign add_793470 = sel_793467 + 8'h01;
  assign sel_793471 = array_index_793454 == array_index_772652 ? add_793470 : sel_793467;
  assign add_793474 = sel_793471 + 8'h01;
  assign sel_793475 = array_index_793454 == array_index_772660 ? add_793474 : sel_793471;
  assign add_793478 = sel_793475 + 8'h01;
  assign sel_793479 = array_index_793454 == array_index_772668 ? add_793478 : sel_793475;
  assign add_793482 = sel_793479 + 8'h01;
  assign sel_793483 = array_index_793454 == array_index_772676 ? add_793482 : sel_793479;
  assign add_793486 = sel_793483 + 8'h01;
  assign sel_793487 = array_index_793454 == array_index_772684 ? add_793486 : sel_793483;
  assign add_793490 = sel_793487 + 8'h01;
  assign sel_793491 = array_index_793454 == array_index_772690 ? add_793490 : sel_793487;
  assign add_793494 = sel_793491 + 8'h01;
  assign sel_793495 = array_index_793454 == array_index_772696 ? add_793494 : sel_793491;
  assign add_793498 = sel_793495 + 8'h01;
  assign sel_793499 = array_index_793454 == array_index_772702 ? add_793498 : sel_793495;
  assign add_793502 = sel_793499 + 8'h01;
  assign sel_793503 = array_index_793454 == array_index_772708 ? add_793502 : sel_793499;
  assign add_793506 = sel_793503 + 8'h01;
  assign sel_793507 = array_index_793454 == array_index_772714 ? add_793506 : sel_793503;
  assign add_793510 = sel_793507 + 8'h01;
  assign sel_793511 = array_index_793454 == array_index_772720 ? add_793510 : sel_793507;
  assign add_793514 = sel_793511 + 8'h01;
  assign sel_793515 = array_index_793454 == array_index_772726 ? add_793514 : sel_793511;
  assign add_793518 = sel_793515 + 8'h01;
  assign sel_793519 = array_index_793454 == array_index_772732 ? add_793518 : sel_793515;
  assign add_793522 = sel_793519 + 8'h01;
  assign sel_793523 = array_index_793454 == array_index_772738 ? add_793522 : sel_793519;
  assign add_793526 = sel_793523 + 8'h01;
  assign sel_793527 = array_index_793454 == array_index_772744 ? add_793526 : sel_793523;
  assign add_793530 = sel_793527 + 8'h01;
  assign sel_793531 = array_index_793454 == array_index_772750 ? add_793530 : sel_793527;
  assign add_793534 = sel_793531 + 8'h01;
  assign sel_793535 = array_index_793454 == array_index_772756 ? add_793534 : sel_793531;
  assign add_793538 = sel_793535 + 8'h01;
  assign sel_793539 = array_index_793454 == array_index_772762 ? add_793538 : sel_793535;
  assign add_793542 = sel_793539 + 8'h01;
  assign sel_793543 = array_index_793454 == array_index_772768 ? add_793542 : sel_793539;
  assign add_793546 = sel_793543 + 8'h01;
  assign sel_793547 = array_index_793454 == array_index_772774 ? add_793546 : sel_793543;
  assign add_793550 = sel_793547 + 8'h01;
  assign sel_793551 = array_index_793454 == array_index_772780 ? add_793550 : sel_793547;
  assign add_793554 = sel_793551 + 8'h01;
  assign sel_793555 = array_index_793454 == array_index_772786 ? add_793554 : sel_793551;
  assign add_793558 = sel_793555 + 8'h01;
  assign sel_793559 = array_index_793454 == array_index_772792 ? add_793558 : sel_793555;
  assign add_793562 = sel_793559 + 8'h01;
  assign sel_793563 = array_index_793454 == array_index_772798 ? add_793562 : sel_793559;
  assign add_793566 = sel_793563 + 8'h01;
  assign sel_793567 = array_index_793454 == array_index_772804 ? add_793566 : sel_793563;
  assign add_793570 = sel_793567 + 8'h01;
  assign sel_793571 = array_index_793454 == array_index_772810 ? add_793570 : sel_793567;
  assign add_793574 = sel_793571 + 8'h01;
  assign sel_793575 = array_index_793454 == array_index_772816 ? add_793574 : sel_793571;
  assign add_793578 = sel_793575 + 8'h01;
  assign sel_793579 = array_index_793454 == array_index_772822 ? add_793578 : sel_793575;
  assign add_793582 = sel_793579 + 8'h01;
  assign sel_793583 = array_index_793454 == array_index_772828 ? add_793582 : sel_793579;
  assign add_793586 = sel_793583 + 8'h01;
  assign sel_793587 = array_index_793454 == array_index_772834 ? add_793586 : sel_793583;
  assign add_793590 = sel_793587 + 8'h01;
  assign sel_793591 = array_index_793454 == array_index_772840 ? add_793590 : sel_793587;
  assign add_793594 = sel_793591 + 8'h01;
  assign sel_793595 = array_index_793454 == array_index_772846 ? add_793594 : sel_793591;
  assign add_793598 = sel_793595 + 8'h01;
  assign sel_793599 = array_index_793454 == array_index_772852 ? add_793598 : sel_793595;
  assign add_793602 = sel_793599 + 8'h01;
  assign sel_793603 = array_index_793454 == array_index_772858 ? add_793602 : sel_793599;
  assign add_793606 = sel_793603 + 8'h01;
  assign sel_793607 = array_index_793454 == array_index_772864 ? add_793606 : sel_793603;
  assign add_793610 = sel_793607 + 8'h01;
  assign sel_793611 = array_index_793454 == array_index_772870 ? add_793610 : sel_793607;
  assign add_793614 = sel_793611 + 8'h01;
  assign sel_793615 = array_index_793454 == array_index_772876 ? add_793614 : sel_793611;
  assign add_793618 = sel_793615 + 8'h01;
  assign sel_793619 = array_index_793454 == array_index_772882 ? add_793618 : sel_793615;
  assign add_793622 = sel_793619 + 8'h01;
  assign sel_793623 = array_index_793454 == array_index_772888 ? add_793622 : sel_793619;
  assign add_793626 = sel_793623 + 8'h01;
  assign sel_793627 = array_index_793454 == array_index_772894 ? add_793626 : sel_793623;
  assign add_793630 = sel_793627 + 8'h01;
  assign sel_793631 = array_index_793454 == array_index_772900 ? add_793630 : sel_793627;
  assign add_793634 = sel_793631 + 8'h01;
  assign sel_793635 = array_index_793454 == array_index_772906 ? add_793634 : sel_793631;
  assign add_793638 = sel_793635 + 8'h01;
  assign sel_793639 = array_index_793454 == array_index_772912 ? add_793638 : sel_793635;
  assign add_793642 = sel_793639 + 8'h01;
  assign sel_793643 = array_index_793454 == array_index_772918 ? add_793642 : sel_793639;
  assign add_793646 = sel_793643 + 8'h01;
  assign sel_793647 = array_index_793454 == array_index_772924 ? add_793646 : sel_793643;
  assign add_793650 = sel_793647 + 8'h01;
  assign sel_793651 = array_index_793454 == array_index_772930 ? add_793650 : sel_793647;
  assign add_793654 = sel_793651 + 8'h01;
  assign sel_793655 = array_index_793454 == array_index_772936 ? add_793654 : sel_793651;
  assign add_793658 = sel_793655 + 8'h01;
  assign sel_793659 = array_index_793454 == array_index_772942 ? add_793658 : sel_793655;
  assign add_793662 = sel_793659 + 8'h01;
  assign sel_793663 = array_index_793454 == array_index_772948 ? add_793662 : sel_793659;
  assign add_793666 = sel_793663 + 8'h01;
  assign sel_793667 = array_index_793454 == array_index_772954 ? add_793666 : sel_793663;
  assign add_793670 = sel_793667 + 8'h01;
  assign sel_793671 = array_index_793454 == array_index_772960 ? add_793670 : sel_793667;
  assign add_793674 = sel_793671 + 8'h01;
  assign sel_793675 = array_index_793454 == array_index_772966 ? add_793674 : sel_793671;
  assign add_793678 = sel_793675 + 8'h01;
  assign sel_793679 = array_index_793454 == array_index_772972 ? add_793678 : sel_793675;
  assign add_793682 = sel_793679 + 8'h01;
  assign sel_793683 = array_index_793454 == array_index_772978 ? add_793682 : sel_793679;
  assign add_793686 = sel_793683 + 8'h01;
  assign sel_793687 = array_index_793454 == array_index_772984 ? add_793686 : sel_793683;
  assign add_793690 = sel_793687 + 8'h01;
  assign sel_793691 = array_index_793454 == array_index_772990 ? add_793690 : sel_793687;
  assign add_793694 = sel_793691 + 8'h01;
  assign sel_793695 = array_index_793454 == array_index_772996 ? add_793694 : sel_793691;
  assign add_793698 = sel_793695 + 8'h01;
  assign sel_793699 = array_index_793454 == array_index_773002 ? add_793698 : sel_793695;
  assign add_793702 = sel_793699 + 8'h01;
  assign sel_793703 = array_index_793454 == array_index_773008 ? add_793702 : sel_793699;
  assign add_793706 = sel_793703 + 8'h01;
  assign sel_793707 = array_index_793454 == array_index_773014 ? add_793706 : sel_793703;
  assign add_793710 = sel_793707 + 8'h01;
  assign sel_793711 = array_index_793454 == array_index_773020 ? add_793710 : sel_793707;
  assign add_793714 = sel_793711 + 8'h01;
  assign sel_793715 = array_index_793454 == array_index_773026 ? add_793714 : sel_793711;
  assign add_793718 = sel_793715 + 8'h01;
  assign sel_793719 = array_index_793454 == array_index_773032 ? add_793718 : sel_793715;
  assign add_793722 = sel_793719 + 8'h01;
  assign sel_793723 = array_index_793454 == array_index_773038 ? add_793722 : sel_793719;
  assign add_793726 = sel_793723 + 8'h01;
  assign sel_793727 = array_index_793454 == array_index_773044 ? add_793726 : sel_793723;
  assign add_793730 = sel_793727 + 8'h01;
  assign sel_793731 = array_index_793454 == array_index_773050 ? add_793730 : sel_793727;
  assign add_793734 = sel_793731 + 8'h01;
  assign sel_793735 = array_index_793454 == array_index_773056 ? add_793734 : sel_793731;
  assign add_793738 = sel_793735 + 8'h01;
  assign sel_793739 = array_index_793454 == array_index_773062 ? add_793738 : sel_793735;
  assign add_793742 = sel_793739 + 8'h01;
  assign sel_793743 = array_index_793454 == array_index_773068 ? add_793742 : sel_793739;
  assign add_793746 = sel_793743 + 8'h01;
  assign sel_793747 = array_index_793454 == array_index_773074 ? add_793746 : sel_793743;
  assign add_793750 = sel_793747 + 8'h01;
  assign sel_793751 = array_index_793454 == array_index_773080 ? add_793750 : sel_793747;
  assign add_793754 = sel_793751 + 8'h01;
  assign sel_793755 = array_index_793454 == array_index_773086 ? add_793754 : sel_793751;
  assign add_793758 = sel_793755 + 8'h01;
  assign sel_793759 = array_index_793454 == array_index_773092 ? add_793758 : sel_793755;
  assign add_793762 = sel_793759 + 8'h01;
  assign sel_793763 = array_index_793454 == array_index_773098 ? add_793762 : sel_793759;
  assign add_793766 = sel_793763 + 8'h01;
  assign sel_793767 = array_index_793454 == array_index_773104 ? add_793766 : sel_793763;
  assign add_793770 = sel_793767 + 8'h01;
  assign sel_793771 = array_index_793454 == array_index_773110 ? add_793770 : sel_793767;
  assign add_793774 = sel_793771 + 8'h01;
  assign sel_793775 = array_index_793454 == array_index_773116 ? add_793774 : sel_793771;
  assign add_793778 = sel_793775 + 8'h01;
  assign sel_793779 = array_index_793454 == array_index_773122 ? add_793778 : sel_793775;
  assign add_793782 = sel_793779 + 8'h01;
  assign sel_793783 = array_index_793454 == array_index_773128 ? add_793782 : sel_793779;
  assign add_793786 = sel_793783 + 8'h01;
  assign sel_793787 = array_index_793454 == array_index_773134 ? add_793786 : sel_793783;
  assign add_793790 = sel_793787 + 8'h01;
  assign sel_793791 = array_index_793454 == array_index_773140 ? add_793790 : sel_793787;
  assign add_793794 = sel_793791 + 8'h01;
  assign sel_793795 = array_index_793454 == array_index_773146 ? add_793794 : sel_793791;
  assign add_793798 = sel_793795 + 8'h01;
  assign sel_793799 = array_index_793454 == array_index_773152 ? add_793798 : sel_793795;
  assign add_793802 = sel_793799 + 8'h01;
  assign sel_793803 = array_index_793454 == array_index_773158 ? add_793802 : sel_793799;
  assign add_793806 = sel_793803 + 8'h01;
  assign sel_793807 = array_index_793454 == array_index_773164 ? add_793806 : sel_793803;
  assign add_793810 = sel_793807 + 8'h01;
  assign sel_793811 = array_index_793454 == array_index_773170 ? add_793810 : sel_793807;
  assign add_793815 = sel_793811 + 8'h01;
  assign array_index_793816 = set1_unflattened[7'h3a];
  assign sel_793817 = array_index_793454 == array_index_773176 ? add_793815 : sel_793811;
  assign add_793820 = sel_793817 + 8'h01;
  assign sel_793821 = array_index_793816 == array_index_772632 ? add_793820 : sel_793817;
  assign add_793824 = sel_793821 + 8'h01;
  assign sel_793825 = array_index_793816 == array_index_772636 ? add_793824 : sel_793821;
  assign add_793828 = sel_793825 + 8'h01;
  assign sel_793829 = array_index_793816 == array_index_772644 ? add_793828 : sel_793825;
  assign add_793832 = sel_793829 + 8'h01;
  assign sel_793833 = array_index_793816 == array_index_772652 ? add_793832 : sel_793829;
  assign add_793836 = sel_793833 + 8'h01;
  assign sel_793837 = array_index_793816 == array_index_772660 ? add_793836 : sel_793833;
  assign add_793840 = sel_793837 + 8'h01;
  assign sel_793841 = array_index_793816 == array_index_772668 ? add_793840 : sel_793837;
  assign add_793844 = sel_793841 + 8'h01;
  assign sel_793845 = array_index_793816 == array_index_772676 ? add_793844 : sel_793841;
  assign add_793848 = sel_793845 + 8'h01;
  assign sel_793849 = array_index_793816 == array_index_772684 ? add_793848 : sel_793845;
  assign add_793852 = sel_793849 + 8'h01;
  assign sel_793853 = array_index_793816 == array_index_772690 ? add_793852 : sel_793849;
  assign add_793856 = sel_793853 + 8'h01;
  assign sel_793857 = array_index_793816 == array_index_772696 ? add_793856 : sel_793853;
  assign add_793860 = sel_793857 + 8'h01;
  assign sel_793861 = array_index_793816 == array_index_772702 ? add_793860 : sel_793857;
  assign add_793864 = sel_793861 + 8'h01;
  assign sel_793865 = array_index_793816 == array_index_772708 ? add_793864 : sel_793861;
  assign add_793868 = sel_793865 + 8'h01;
  assign sel_793869 = array_index_793816 == array_index_772714 ? add_793868 : sel_793865;
  assign add_793872 = sel_793869 + 8'h01;
  assign sel_793873 = array_index_793816 == array_index_772720 ? add_793872 : sel_793869;
  assign add_793876 = sel_793873 + 8'h01;
  assign sel_793877 = array_index_793816 == array_index_772726 ? add_793876 : sel_793873;
  assign add_793880 = sel_793877 + 8'h01;
  assign sel_793881 = array_index_793816 == array_index_772732 ? add_793880 : sel_793877;
  assign add_793884 = sel_793881 + 8'h01;
  assign sel_793885 = array_index_793816 == array_index_772738 ? add_793884 : sel_793881;
  assign add_793888 = sel_793885 + 8'h01;
  assign sel_793889 = array_index_793816 == array_index_772744 ? add_793888 : sel_793885;
  assign add_793892 = sel_793889 + 8'h01;
  assign sel_793893 = array_index_793816 == array_index_772750 ? add_793892 : sel_793889;
  assign add_793896 = sel_793893 + 8'h01;
  assign sel_793897 = array_index_793816 == array_index_772756 ? add_793896 : sel_793893;
  assign add_793900 = sel_793897 + 8'h01;
  assign sel_793901 = array_index_793816 == array_index_772762 ? add_793900 : sel_793897;
  assign add_793904 = sel_793901 + 8'h01;
  assign sel_793905 = array_index_793816 == array_index_772768 ? add_793904 : sel_793901;
  assign add_793908 = sel_793905 + 8'h01;
  assign sel_793909 = array_index_793816 == array_index_772774 ? add_793908 : sel_793905;
  assign add_793912 = sel_793909 + 8'h01;
  assign sel_793913 = array_index_793816 == array_index_772780 ? add_793912 : sel_793909;
  assign add_793916 = sel_793913 + 8'h01;
  assign sel_793917 = array_index_793816 == array_index_772786 ? add_793916 : sel_793913;
  assign add_793920 = sel_793917 + 8'h01;
  assign sel_793921 = array_index_793816 == array_index_772792 ? add_793920 : sel_793917;
  assign add_793924 = sel_793921 + 8'h01;
  assign sel_793925 = array_index_793816 == array_index_772798 ? add_793924 : sel_793921;
  assign add_793928 = sel_793925 + 8'h01;
  assign sel_793929 = array_index_793816 == array_index_772804 ? add_793928 : sel_793925;
  assign add_793932 = sel_793929 + 8'h01;
  assign sel_793933 = array_index_793816 == array_index_772810 ? add_793932 : sel_793929;
  assign add_793936 = sel_793933 + 8'h01;
  assign sel_793937 = array_index_793816 == array_index_772816 ? add_793936 : sel_793933;
  assign add_793940 = sel_793937 + 8'h01;
  assign sel_793941 = array_index_793816 == array_index_772822 ? add_793940 : sel_793937;
  assign add_793944 = sel_793941 + 8'h01;
  assign sel_793945 = array_index_793816 == array_index_772828 ? add_793944 : sel_793941;
  assign add_793948 = sel_793945 + 8'h01;
  assign sel_793949 = array_index_793816 == array_index_772834 ? add_793948 : sel_793945;
  assign add_793952 = sel_793949 + 8'h01;
  assign sel_793953 = array_index_793816 == array_index_772840 ? add_793952 : sel_793949;
  assign add_793956 = sel_793953 + 8'h01;
  assign sel_793957 = array_index_793816 == array_index_772846 ? add_793956 : sel_793953;
  assign add_793960 = sel_793957 + 8'h01;
  assign sel_793961 = array_index_793816 == array_index_772852 ? add_793960 : sel_793957;
  assign add_793964 = sel_793961 + 8'h01;
  assign sel_793965 = array_index_793816 == array_index_772858 ? add_793964 : sel_793961;
  assign add_793968 = sel_793965 + 8'h01;
  assign sel_793969 = array_index_793816 == array_index_772864 ? add_793968 : sel_793965;
  assign add_793972 = sel_793969 + 8'h01;
  assign sel_793973 = array_index_793816 == array_index_772870 ? add_793972 : sel_793969;
  assign add_793976 = sel_793973 + 8'h01;
  assign sel_793977 = array_index_793816 == array_index_772876 ? add_793976 : sel_793973;
  assign add_793980 = sel_793977 + 8'h01;
  assign sel_793981 = array_index_793816 == array_index_772882 ? add_793980 : sel_793977;
  assign add_793984 = sel_793981 + 8'h01;
  assign sel_793985 = array_index_793816 == array_index_772888 ? add_793984 : sel_793981;
  assign add_793988 = sel_793985 + 8'h01;
  assign sel_793989 = array_index_793816 == array_index_772894 ? add_793988 : sel_793985;
  assign add_793992 = sel_793989 + 8'h01;
  assign sel_793993 = array_index_793816 == array_index_772900 ? add_793992 : sel_793989;
  assign add_793996 = sel_793993 + 8'h01;
  assign sel_793997 = array_index_793816 == array_index_772906 ? add_793996 : sel_793993;
  assign add_794000 = sel_793997 + 8'h01;
  assign sel_794001 = array_index_793816 == array_index_772912 ? add_794000 : sel_793997;
  assign add_794004 = sel_794001 + 8'h01;
  assign sel_794005 = array_index_793816 == array_index_772918 ? add_794004 : sel_794001;
  assign add_794008 = sel_794005 + 8'h01;
  assign sel_794009 = array_index_793816 == array_index_772924 ? add_794008 : sel_794005;
  assign add_794012 = sel_794009 + 8'h01;
  assign sel_794013 = array_index_793816 == array_index_772930 ? add_794012 : sel_794009;
  assign add_794016 = sel_794013 + 8'h01;
  assign sel_794017 = array_index_793816 == array_index_772936 ? add_794016 : sel_794013;
  assign add_794020 = sel_794017 + 8'h01;
  assign sel_794021 = array_index_793816 == array_index_772942 ? add_794020 : sel_794017;
  assign add_794024 = sel_794021 + 8'h01;
  assign sel_794025 = array_index_793816 == array_index_772948 ? add_794024 : sel_794021;
  assign add_794028 = sel_794025 + 8'h01;
  assign sel_794029 = array_index_793816 == array_index_772954 ? add_794028 : sel_794025;
  assign add_794032 = sel_794029 + 8'h01;
  assign sel_794033 = array_index_793816 == array_index_772960 ? add_794032 : sel_794029;
  assign add_794036 = sel_794033 + 8'h01;
  assign sel_794037 = array_index_793816 == array_index_772966 ? add_794036 : sel_794033;
  assign add_794040 = sel_794037 + 8'h01;
  assign sel_794041 = array_index_793816 == array_index_772972 ? add_794040 : sel_794037;
  assign add_794044 = sel_794041 + 8'h01;
  assign sel_794045 = array_index_793816 == array_index_772978 ? add_794044 : sel_794041;
  assign add_794048 = sel_794045 + 8'h01;
  assign sel_794049 = array_index_793816 == array_index_772984 ? add_794048 : sel_794045;
  assign add_794052 = sel_794049 + 8'h01;
  assign sel_794053 = array_index_793816 == array_index_772990 ? add_794052 : sel_794049;
  assign add_794056 = sel_794053 + 8'h01;
  assign sel_794057 = array_index_793816 == array_index_772996 ? add_794056 : sel_794053;
  assign add_794060 = sel_794057 + 8'h01;
  assign sel_794061 = array_index_793816 == array_index_773002 ? add_794060 : sel_794057;
  assign add_794064 = sel_794061 + 8'h01;
  assign sel_794065 = array_index_793816 == array_index_773008 ? add_794064 : sel_794061;
  assign add_794068 = sel_794065 + 8'h01;
  assign sel_794069 = array_index_793816 == array_index_773014 ? add_794068 : sel_794065;
  assign add_794072 = sel_794069 + 8'h01;
  assign sel_794073 = array_index_793816 == array_index_773020 ? add_794072 : sel_794069;
  assign add_794076 = sel_794073 + 8'h01;
  assign sel_794077 = array_index_793816 == array_index_773026 ? add_794076 : sel_794073;
  assign add_794080 = sel_794077 + 8'h01;
  assign sel_794081 = array_index_793816 == array_index_773032 ? add_794080 : sel_794077;
  assign add_794084 = sel_794081 + 8'h01;
  assign sel_794085 = array_index_793816 == array_index_773038 ? add_794084 : sel_794081;
  assign add_794088 = sel_794085 + 8'h01;
  assign sel_794089 = array_index_793816 == array_index_773044 ? add_794088 : sel_794085;
  assign add_794092 = sel_794089 + 8'h01;
  assign sel_794093 = array_index_793816 == array_index_773050 ? add_794092 : sel_794089;
  assign add_794096 = sel_794093 + 8'h01;
  assign sel_794097 = array_index_793816 == array_index_773056 ? add_794096 : sel_794093;
  assign add_794100 = sel_794097 + 8'h01;
  assign sel_794101 = array_index_793816 == array_index_773062 ? add_794100 : sel_794097;
  assign add_794104 = sel_794101 + 8'h01;
  assign sel_794105 = array_index_793816 == array_index_773068 ? add_794104 : sel_794101;
  assign add_794108 = sel_794105 + 8'h01;
  assign sel_794109 = array_index_793816 == array_index_773074 ? add_794108 : sel_794105;
  assign add_794112 = sel_794109 + 8'h01;
  assign sel_794113 = array_index_793816 == array_index_773080 ? add_794112 : sel_794109;
  assign add_794116 = sel_794113 + 8'h01;
  assign sel_794117 = array_index_793816 == array_index_773086 ? add_794116 : sel_794113;
  assign add_794120 = sel_794117 + 8'h01;
  assign sel_794121 = array_index_793816 == array_index_773092 ? add_794120 : sel_794117;
  assign add_794124 = sel_794121 + 8'h01;
  assign sel_794125 = array_index_793816 == array_index_773098 ? add_794124 : sel_794121;
  assign add_794128 = sel_794125 + 8'h01;
  assign sel_794129 = array_index_793816 == array_index_773104 ? add_794128 : sel_794125;
  assign add_794132 = sel_794129 + 8'h01;
  assign sel_794133 = array_index_793816 == array_index_773110 ? add_794132 : sel_794129;
  assign add_794136 = sel_794133 + 8'h01;
  assign sel_794137 = array_index_793816 == array_index_773116 ? add_794136 : sel_794133;
  assign add_794140 = sel_794137 + 8'h01;
  assign sel_794141 = array_index_793816 == array_index_773122 ? add_794140 : sel_794137;
  assign add_794144 = sel_794141 + 8'h01;
  assign sel_794145 = array_index_793816 == array_index_773128 ? add_794144 : sel_794141;
  assign add_794148 = sel_794145 + 8'h01;
  assign sel_794149 = array_index_793816 == array_index_773134 ? add_794148 : sel_794145;
  assign add_794152 = sel_794149 + 8'h01;
  assign sel_794153 = array_index_793816 == array_index_773140 ? add_794152 : sel_794149;
  assign add_794156 = sel_794153 + 8'h01;
  assign sel_794157 = array_index_793816 == array_index_773146 ? add_794156 : sel_794153;
  assign add_794160 = sel_794157 + 8'h01;
  assign sel_794161 = array_index_793816 == array_index_773152 ? add_794160 : sel_794157;
  assign add_794164 = sel_794161 + 8'h01;
  assign sel_794165 = array_index_793816 == array_index_773158 ? add_794164 : sel_794161;
  assign add_794168 = sel_794165 + 8'h01;
  assign sel_794169 = array_index_793816 == array_index_773164 ? add_794168 : sel_794165;
  assign add_794172 = sel_794169 + 8'h01;
  assign sel_794173 = array_index_793816 == array_index_773170 ? add_794172 : sel_794169;
  assign add_794177 = sel_794173 + 8'h01;
  assign array_index_794178 = set1_unflattened[7'h3b];
  assign sel_794179 = array_index_793816 == array_index_773176 ? add_794177 : sel_794173;
  assign add_794182 = sel_794179 + 8'h01;
  assign sel_794183 = array_index_794178 == array_index_772632 ? add_794182 : sel_794179;
  assign add_794186 = sel_794183 + 8'h01;
  assign sel_794187 = array_index_794178 == array_index_772636 ? add_794186 : sel_794183;
  assign add_794190 = sel_794187 + 8'h01;
  assign sel_794191 = array_index_794178 == array_index_772644 ? add_794190 : sel_794187;
  assign add_794194 = sel_794191 + 8'h01;
  assign sel_794195 = array_index_794178 == array_index_772652 ? add_794194 : sel_794191;
  assign add_794198 = sel_794195 + 8'h01;
  assign sel_794199 = array_index_794178 == array_index_772660 ? add_794198 : sel_794195;
  assign add_794202 = sel_794199 + 8'h01;
  assign sel_794203 = array_index_794178 == array_index_772668 ? add_794202 : sel_794199;
  assign add_794206 = sel_794203 + 8'h01;
  assign sel_794207 = array_index_794178 == array_index_772676 ? add_794206 : sel_794203;
  assign add_794210 = sel_794207 + 8'h01;
  assign sel_794211 = array_index_794178 == array_index_772684 ? add_794210 : sel_794207;
  assign add_794214 = sel_794211 + 8'h01;
  assign sel_794215 = array_index_794178 == array_index_772690 ? add_794214 : sel_794211;
  assign add_794218 = sel_794215 + 8'h01;
  assign sel_794219 = array_index_794178 == array_index_772696 ? add_794218 : sel_794215;
  assign add_794222 = sel_794219 + 8'h01;
  assign sel_794223 = array_index_794178 == array_index_772702 ? add_794222 : sel_794219;
  assign add_794226 = sel_794223 + 8'h01;
  assign sel_794227 = array_index_794178 == array_index_772708 ? add_794226 : sel_794223;
  assign add_794230 = sel_794227 + 8'h01;
  assign sel_794231 = array_index_794178 == array_index_772714 ? add_794230 : sel_794227;
  assign add_794234 = sel_794231 + 8'h01;
  assign sel_794235 = array_index_794178 == array_index_772720 ? add_794234 : sel_794231;
  assign add_794238 = sel_794235 + 8'h01;
  assign sel_794239 = array_index_794178 == array_index_772726 ? add_794238 : sel_794235;
  assign add_794242 = sel_794239 + 8'h01;
  assign sel_794243 = array_index_794178 == array_index_772732 ? add_794242 : sel_794239;
  assign add_794246 = sel_794243 + 8'h01;
  assign sel_794247 = array_index_794178 == array_index_772738 ? add_794246 : sel_794243;
  assign add_794250 = sel_794247 + 8'h01;
  assign sel_794251 = array_index_794178 == array_index_772744 ? add_794250 : sel_794247;
  assign add_794254 = sel_794251 + 8'h01;
  assign sel_794255 = array_index_794178 == array_index_772750 ? add_794254 : sel_794251;
  assign add_794258 = sel_794255 + 8'h01;
  assign sel_794259 = array_index_794178 == array_index_772756 ? add_794258 : sel_794255;
  assign add_794262 = sel_794259 + 8'h01;
  assign sel_794263 = array_index_794178 == array_index_772762 ? add_794262 : sel_794259;
  assign add_794266 = sel_794263 + 8'h01;
  assign sel_794267 = array_index_794178 == array_index_772768 ? add_794266 : sel_794263;
  assign add_794270 = sel_794267 + 8'h01;
  assign sel_794271 = array_index_794178 == array_index_772774 ? add_794270 : sel_794267;
  assign add_794274 = sel_794271 + 8'h01;
  assign sel_794275 = array_index_794178 == array_index_772780 ? add_794274 : sel_794271;
  assign add_794278 = sel_794275 + 8'h01;
  assign sel_794279 = array_index_794178 == array_index_772786 ? add_794278 : sel_794275;
  assign add_794282 = sel_794279 + 8'h01;
  assign sel_794283 = array_index_794178 == array_index_772792 ? add_794282 : sel_794279;
  assign add_794286 = sel_794283 + 8'h01;
  assign sel_794287 = array_index_794178 == array_index_772798 ? add_794286 : sel_794283;
  assign add_794290 = sel_794287 + 8'h01;
  assign sel_794291 = array_index_794178 == array_index_772804 ? add_794290 : sel_794287;
  assign add_794294 = sel_794291 + 8'h01;
  assign sel_794295 = array_index_794178 == array_index_772810 ? add_794294 : sel_794291;
  assign add_794298 = sel_794295 + 8'h01;
  assign sel_794299 = array_index_794178 == array_index_772816 ? add_794298 : sel_794295;
  assign add_794302 = sel_794299 + 8'h01;
  assign sel_794303 = array_index_794178 == array_index_772822 ? add_794302 : sel_794299;
  assign add_794306 = sel_794303 + 8'h01;
  assign sel_794307 = array_index_794178 == array_index_772828 ? add_794306 : sel_794303;
  assign add_794310 = sel_794307 + 8'h01;
  assign sel_794311 = array_index_794178 == array_index_772834 ? add_794310 : sel_794307;
  assign add_794314 = sel_794311 + 8'h01;
  assign sel_794315 = array_index_794178 == array_index_772840 ? add_794314 : sel_794311;
  assign add_794318 = sel_794315 + 8'h01;
  assign sel_794319 = array_index_794178 == array_index_772846 ? add_794318 : sel_794315;
  assign add_794322 = sel_794319 + 8'h01;
  assign sel_794323 = array_index_794178 == array_index_772852 ? add_794322 : sel_794319;
  assign add_794326 = sel_794323 + 8'h01;
  assign sel_794327 = array_index_794178 == array_index_772858 ? add_794326 : sel_794323;
  assign add_794330 = sel_794327 + 8'h01;
  assign sel_794331 = array_index_794178 == array_index_772864 ? add_794330 : sel_794327;
  assign add_794334 = sel_794331 + 8'h01;
  assign sel_794335 = array_index_794178 == array_index_772870 ? add_794334 : sel_794331;
  assign add_794338 = sel_794335 + 8'h01;
  assign sel_794339 = array_index_794178 == array_index_772876 ? add_794338 : sel_794335;
  assign add_794342 = sel_794339 + 8'h01;
  assign sel_794343 = array_index_794178 == array_index_772882 ? add_794342 : sel_794339;
  assign add_794346 = sel_794343 + 8'h01;
  assign sel_794347 = array_index_794178 == array_index_772888 ? add_794346 : sel_794343;
  assign add_794350 = sel_794347 + 8'h01;
  assign sel_794351 = array_index_794178 == array_index_772894 ? add_794350 : sel_794347;
  assign add_794354 = sel_794351 + 8'h01;
  assign sel_794355 = array_index_794178 == array_index_772900 ? add_794354 : sel_794351;
  assign add_794358 = sel_794355 + 8'h01;
  assign sel_794359 = array_index_794178 == array_index_772906 ? add_794358 : sel_794355;
  assign add_794362 = sel_794359 + 8'h01;
  assign sel_794363 = array_index_794178 == array_index_772912 ? add_794362 : sel_794359;
  assign add_794366 = sel_794363 + 8'h01;
  assign sel_794367 = array_index_794178 == array_index_772918 ? add_794366 : sel_794363;
  assign add_794370 = sel_794367 + 8'h01;
  assign sel_794371 = array_index_794178 == array_index_772924 ? add_794370 : sel_794367;
  assign add_794374 = sel_794371 + 8'h01;
  assign sel_794375 = array_index_794178 == array_index_772930 ? add_794374 : sel_794371;
  assign add_794378 = sel_794375 + 8'h01;
  assign sel_794379 = array_index_794178 == array_index_772936 ? add_794378 : sel_794375;
  assign add_794382 = sel_794379 + 8'h01;
  assign sel_794383 = array_index_794178 == array_index_772942 ? add_794382 : sel_794379;
  assign add_794386 = sel_794383 + 8'h01;
  assign sel_794387 = array_index_794178 == array_index_772948 ? add_794386 : sel_794383;
  assign add_794390 = sel_794387 + 8'h01;
  assign sel_794391 = array_index_794178 == array_index_772954 ? add_794390 : sel_794387;
  assign add_794394 = sel_794391 + 8'h01;
  assign sel_794395 = array_index_794178 == array_index_772960 ? add_794394 : sel_794391;
  assign add_794398 = sel_794395 + 8'h01;
  assign sel_794399 = array_index_794178 == array_index_772966 ? add_794398 : sel_794395;
  assign add_794402 = sel_794399 + 8'h01;
  assign sel_794403 = array_index_794178 == array_index_772972 ? add_794402 : sel_794399;
  assign add_794406 = sel_794403 + 8'h01;
  assign sel_794407 = array_index_794178 == array_index_772978 ? add_794406 : sel_794403;
  assign add_794410 = sel_794407 + 8'h01;
  assign sel_794411 = array_index_794178 == array_index_772984 ? add_794410 : sel_794407;
  assign add_794414 = sel_794411 + 8'h01;
  assign sel_794415 = array_index_794178 == array_index_772990 ? add_794414 : sel_794411;
  assign add_794418 = sel_794415 + 8'h01;
  assign sel_794419 = array_index_794178 == array_index_772996 ? add_794418 : sel_794415;
  assign add_794422 = sel_794419 + 8'h01;
  assign sel_794423 = array_index_794178 == array_index_773002 ? add_794422 : sel_794419;
  assign add_794426 = sel_794423 + 8'h01;
  assign sel_794427 = array_index_794178 == array_index_773008 ? add_794426 : sel_794423;
  assign add_794430 = sel_794427 + 8'h01;
  assign sel_794431 = array_index_794178 == array_index_773014 ? add_794430 : sel_794427;
  assign add_794434 = sel_794431 + 8'h01;
  assign sel_794435 = array_index_794178 == array_index_773020 ? add_794434 : sel_794431;
  assign add_794438 = sel_794435 + 8'h01;
  assign sel_794439 = array_index_794178 == array_index_773026 ? add_794438 : sel_794435;
  assign add_794442 = sel_794439 + 8'h01;
  assign sel_794443 = array_index_794178 == array_index_773032 ? add_794442 : sel_794439;
  assign add_794446 = sel_794443 + 8'h01;
  assign sel_794447 = array_index_794178 == array_index_773038 ? add_794446 : sel_794443;
  assign add_794450 = sel_794447 + 8'h01;
  assign sel_794451 = array_index_794178 == array_index_773044 ? add_794450 : sel_794447;
  assign add_794454 = sel_794451 + 8'h01;
  assign sel_794455 = array_index_794178 == array_index_773050 ? add_794454 : sel_794451;
  assign add_794458 = sel_794455 + 8'h01;
  assign sel_794459 = array_index_794178 == array_index_773056 ? add_794458 : sel_794455;
  assign add_794462 = sel_794459 + 8'h01;
  assign sel_794463 = array_index_794178 == array_index_773062 ? add_794462 : sel_794459;
  assign add_794466 = sel_794463 + 8'h01;
  assign sel_794467 = array_index_794178 == array_index_773068 ? add_794466 : sel_794463;
  assign add_794470 = sel_794467 + 8'h01;
  assign sel_794471 = array_index_794178 == array_index_773074 ? add_794470 : sel_794467;
  assign add_794474 = sel_794471 + 8'h01;
  assign sel_794475 = array_index_794178 == array_index_773080 ? add_794474 : sel_794471;
  assign add_794478 = sel_794475 + 8'h01;
  assign sel_794479 = array_index_794178 == array_index_773086 ? add_794478 : sel_794475;
  assign add_794482 = sel_794479 + 8'h01;
  assign sel_794483 = array_index_794178 == array_index_773092 ? add_794482 : sel_794479;
  assign add_794486 = sel_794483 + 8'h01;
  assign sel_794487 = array_index_794178 == array_index_773098 ? add_794486 : sel_794483;
  assign add_794490 = sel_794487 + 8'h01;
  assign sel_794491 = array_index_794178 == array_index_773104 ? add_794490 : sel_794487;
  assign add_794494 = sel_794491 + 8'h01;
  assign sel_794495 = array_index_794178 == array_index_773110 ? add_794494 : sel_794491;
  assign add_794498 = sel_794495 + 8'h01;
  assign sel_794499 = array_index_794178 == array_index_773116 ? add_794498 : sel_794495;
  assign add_794502 = sel_794499 + 8'h01;
  assign sel_794503 = array_index_794178 == array_index_773122 ? add_794502 : sel_794499;
  assign add_794506 = sel_794503 + 8'h01;
  assign sel_794507 = array_index_794178 == array_index_773128 ? add_794506 : sel_794503;
  assign add_794510 = sel_794507 + 8'h01;
  assign sel_794511 = array_index_794178 == array_index_773134 ? add_794510 : sel_794507;
  assign add_794514 = sel_794511 + 8'h01;
  assign sel_794515 = array_index_794178 == array_index_773140 ? add_794514 : sel_794511;
  assign add_794518 = sel_794515 + 8'h01;
  assign sel_794519 = array_index_794178 == array_index_773146 ? add_794518 : sel_794515;
  assign add_794522 = sel_794519 + 8'h01;
  assign sel_794523 = array_index_794178 == array_index_773152 ? add_794522 : sel_794519;
  assign add_794526 = sel_794523 + 8'h01;
  assign sel_794527 = array_index_794178 == array_index_773158 ? add_794526 : sel_794523;
  assign add_794530 = sel_794527 + 8'h01;
  assign sel_794531 = array_index_794178 == array_index_773164 ? add_794530 : sel_794527;
  assign add_794534 = sel_794531 + 8'h01;
  assign sel_794535 = array_index_794178 == array_index_773170 ? add_794534 : sel_794531;
  assign add_794539 = sel_794535 + 8'h01;
  assign array_index_794540 = set1_unflattened[7'h3c];
  assign sel_794541 = array_index_794178 == array_index_773176 ? add_794539 : sel_794535;
  assign add_794544 = sel_794541 + 8'h01;
  assign sel_794545 = array_index_794540 == array_index_772632 ? add_794544 : sel_794541;
  assign add_794548 = sel_794545 + 8'h01;
  assign sel_794549 = array_index_794540 == array_index_772636 ? add_794548 : sel_794545;
  assign add_794552 = sel_794549 + 8'h01;
  assign sel_794553 = array_index_794540 == array_index_772644 ? add_794552 : sel_794549;
  assign add_794556 = sel_794553 + 8'h01;
  assign sel_794557 = array_index_794540 == array_index_772652 ? add_794556 : sel_794553;
  assign add_794560 = sel_794557 + 8'h01;
  assign sel_794561 = array_index_794540 == array_index_772660 ? add_794560 : sel_794557;
  assign add_794564 = sel_794561 + 8'h01;
  assign sel_794565 = array_index_794540 == array_index_772668 ? add_794564 : sel_794561;
  assign add_794568 = sel_794565 + 8'h01;
  assign sel_794569 = array_index_794540 == array_index_772676 ? add_794568 : sel_794565;
  assign add_794572 = sel_794569 + 8'h01;
  assign sel_794573 = array_index_794540 == array_index_772684 ? add_794572 : sel_794569;
  assign add_794576 = sel_794573 + 8'h01;
  assign sel_794577 = array_index_794540 == array_index_772690 ? add_794576 : sel_794573;
  assign add_794580 = sel_794577 + 8'h01;
  assign sel_794581 = array_index_794540 == array_index_772696 ? add_794580 : sel_794577;
  assign add_794584 = sel_794581 + 8'h01;
  assign sel_794585 = array_index_794540 == array_index_772702 ? add_794584 : sel_794581;
  assign add_794588 = sel_794585 + 8'h01;
  assign sel_794589 = array_index_794540 == array_index_772708 ? add_794588 : sel_794585;
  assign add_794592 = sel_794589 + 8'h01;
  assign sel_794593 = array_index_794540 == array_index_772714 ? add_794592 : sel_794589;
  assign add_794596 = sel_794593 + 8'h01;
  assign sel_794597 = array_index_794540 == array_index_772720 ? add_794596 : sel_794593;
  assign add_794600 = sel_794597 + 8'h01;
  assign sel_794601 = array_index_794540 == array_index_772726 ? add_794600 : sel_794597;
  assign add_794604 = sel_794601 + 8'h01;
  assign sel_794605 = array_index_794540 == array_index_772732 ? add_794604 : sel_794601;
  assign add_794608 = sel_794605 + 8'h01;
  assign sel_794609 = array_index_794540 == array_index_772738 ? add_794608 : sel_794605;
  assign add_794612 = sel_794609 + 8'h01;
  assign sel_794613 = array_index_794540 == array_index_772744 ? add_794612 : sel_794609;
  assign add_794616 = sel_794613 + 8'h01;
  assign sel_794617 = array_index_794540 == array_index_772750 ? add_794616 : sel_794613;
  assign add_794620 = sel_794617 + 8'h01;
  assign sel_794621 = array_index_794540 == array_index_772756 ? add_794620 : sel_794617;
  assign add_794624 = sel_794621 + 8'h01;
  assign sel_794625 = array_index_794540 == array_index_772762 ? add_794624 : sel_794621;
  assign add_794628 = sel_794625 + 8'h01;
  assign sel_794629 = array_index_794540 == array_index_772768 ? add_794628 : sel_794625;
  assign add_794632 = sel_794629 + 8'h01;
  assign sel_794633 = array_index_794540 == array_index_772774 ? add_794632 : sel_794629;
  assign add_794636 = sel_794633 + 8'h01;
  assign sel_794637 = array_index_794540 == array_index_772780 ? add_794636 : sel_794633;
  assign add_794640 = sel_794637 + 8'h01;
  assign sel_794641 = array_index_794540 == array_index_772786 ? add_794640 : sel_794637;
  assign add_794644 = sel_794641 + 8'h01;
  assign sel_794645 = array_index_794540 == array_index_772792 ? add_794644 : sel_794641;
  assign add_794648 = sel_794645 + 8'h01;
  assign sel_794649 = array_index_794540 == array_index_772798 ? add_794648 : sel_794645;
  assign add_794652 = sel_794649 + 8'h01;
  assign sel_794653 = array_index_794540 == array_index_772804 ? add_794652 : sel_794649;
  assign add_794656 = sel_794653 + 8'h01;
  assign sel_794657 = array_index_794540 == array_index_772810 ? add_794656 : sel_794653;
  assign add_794660 = sel_794657 + 8'h01;
  assign sel_794661 = array_index_794540 == array_index_772816 ? add_794660 : sel_794657;
  assign add_794664 = sel_794661 + 8'h01;
  assign sel_794665 = array_index_794540 == array_index_772822 ? add_794664 : sel_794661;
  assign add_794668 = sel_794665 + 8'h01;
  assign sel_794669 = array_index_794540 == array_index_772828 ? add_794668 : sel_794665;
  assign add_794672 = sel_794669 + 8'h01;
  assign sel_794673 = array_index_794540 == array_index_772834 ? add_794672 : sel_794669;
  assign add_794676 = sel_794673 + 8'h01;
  assign sel_794677 = array_index_794540 == array_index_772840 ? add_794676 : sel_794673;
  assign add_794680 = sel_794677 + 8'h01;
  assign sel_794681 = array_index_794540 == array_index_772846 ? add_794680 : sel_794677;
  assign add_794684 = sel_794681 + 8'h01;
  assign sel_794685 = array_index_794540 == array_index_772852 ? add_794684 : sel_794681;
  assign add_794688 = sel_794685 + 8'h01;
  assign sel_794689 = array_index_794540 == array_index_772858 ? add_794688 : sel_794685;
  assign add_794692 = sel_794689 + 8'h01;
  assign sel_794693 = array_index_794540 == array_index_772864 ? add_794692 : sel_794689;
  assign add_794696 = sel_794693 + 8'h01;
  assign sel_794697 = array_index_794540 == array_index_772870 ? add_794696 : sel_794693;
  assign add_794700 = sel_794697 + 8'h01;
  assign sel_794701 = array_index_794540 == array_index_772876 ? add_794700 : sel_794697;
  assign add_794704 = sel_794701 + 8'h01;
  assign sel_794705 = array_index_794540 == array_index_772882 ? add_794704 : sel_794701;
  assign add_794708 = sel_794705 + 8'h01;
  assign sel_794709 = array_index_794540 == array_index_772888 ? add_794708 : sel_794705;
  assign add_794712 = sel_794709 + 8'h01;
  assign sel_794713 = array_index_794540 == array_index_772894 ? add_794712 : sel_794709;
  assign add_794716 = sel_794713 + 8'h01;
  assign sel_794717 = array_index_794540 == array_index_772900 ? add_794716 : sel_794713;
  assign add_794720 = sel_794717 + 8'h01;
  assign sel_794721 = array_index_794540 == array_index_772906 ? add_794720 : sel_794717;
  assign add_794724 = sel_794721 + 8'h01;
  assign sel_794725 = array_index_794540 == array_index_772912 ? add_794724 : sel_794721;
  assign add_794728 = sel_794725 + 8'h01;
  assign sel_794729 = array_index_794540 == array_index_772918 ? add_794728 : sel_794725;
  assign add_794732 = sel_794729 + 8'h01;
  assign sel_794733 = array_index_794540 == array_index_772924 ? add_794732 : sel_794729;
  assign add_794736 = sel_794733 + 8'h01;
  assign sel_794737 = array_index_794540 == array_index_772930 ? add_794736 : sel_794733;
  assign add_794740 = sel_794737 + 8'h01;
  assign sel_794741 = array_index_794540 == array_index_772936 ? add_794740 : sel_794737;
  assign add_794744 = sel_794741 + 8'h01;
  assign sel_794745 = array_index_794540 == array_index_772942 ? add_794744 : sel_794741;
  assign add_794748 = sel_794745 + 8'h01;
  assign sel_794749 = array_index_794540 == array_index_772948 ? add_794748 : sel_794745;
  assign add_794752 = sel_794749 + 8'h01;
  assign sel_794753 = array_index_794540 == array_index_772954 ? add_794752 : sel_794749;
  assign add_794756 = sel_794753 + 8'h01;
  assign sel_794757 = array_index_794540 == array_index_772960 ? add_794756 : sel_794753;
  assign add_794760 = sel_794757 + 8'h01;
  assign sel_794761 = array_index_794540 == array_index_772966 ? add_794760 : sel_794757;
  assign add_794764 = sel_794761 + 8'h01;
  assign sel_794765 = array_index_794540 == array_index_772972 ? add_794764 : sel_794761;
  assign add_794768 = sel_794765 + 8'h01;
  assign sel_794769 = array_index_794540 == array_index_772978 ? add_794768 : sel_794765;
  assign add_794772 = sel_794769 + 8'h01;
  assign sel_794773 = array_index_794540 == array_index_772984 ? add_794772 : sel_794769;
  assign add_794776 = sel_794773 + 8'h01;
  assign sel_794777 = array_index_794540 == array_index_772990 ? add_794776 : sel_794773;
  assign add_794780 = sel_794777 + 8'h01;
  assign sel_794781 = array_index_794540 == array_index_772996 ? add_794780 : sel_794777;
  assign add_794784 = sel_794781 + 8'h01;
  assign sel_794785 = array_index_794540 == array_index_773002 ? add_794784 : sel_794781;
  assign add_794788 = sel_794785 + 8'h01;
  assign sel_794789 = array_index_794540 == array_index_773008 ? add_794788 : sel_794785;
  assign add_794792 = sel_794789 + 8'h01;
  assign sel_794793 = array_index_794540 == array_index_773014 ? add_794792 : sel_794789;
  assign add_794796 = sel_794793 + 8'h01;
  assign sel_794797 = array_index_794540 == array_index_773020 ? add_794796 : sel_794793;
  assign add_794800 = sel_794797 + 8'h01;
  assign sel_794801 = array_index_794540 == array_index_773026 ? add_794800 : sel_794797;
  assign add_794804 = sel_794801 + 8'h01;
  assign sel_794805 = array_index_794540 == array_index_773032 ? add_794804 : sel_794801;
  assign add_794808 = sel_794805 + 8'h01;
  assign sel_794809 = array_index_794540 == array_index_773038 ? add_794808 : sel_794805;
  assign add_794812 = sel_794809 + 8'h01;
  assign sel_794813 = array_index_794540 == array_index_773044 ? add_794812 : sel_794809;
  assign add_794816 = sel_794813 + 8'h01;
  assign sel_794817 = array_index_794540 == array_index_773050 ? add_794816 : sel_794813;
  assign add_794820 = sel_794817 + 8'h01;
  assign sel_794821 = array_index_794540 == array_index_773056 ? add_794820 : sel_794817;
  assign add_794824 = sel_794821 + 8'h01;
  assign sel_794825 = array_index_794540 == array_index_773062 ? add_794824 : sel_794821;
  assign add_794828 = sel_794825 + 8'h01;
  assign sel_794829 = array_index_794540 == array_index_773068 ? add_794828 : sel_794825;
  assign add_794832 = sel_794829 + 8'h01;
  assign sel_794833 = array_index_794540 == array_index_773074 ? add_794832 : sel_794829;
  assign add_794836 = sel_794833 + 8'h01;
  assign sel_794837 = array_index_794540 == array_index_773080 ? add_794836 : sel_794833;
  assign add_794840 = sel_794837 + 8'h01;
  assign sel_794841 = array_index_794540 == array_index_773086 ? add_794840 : sel_794837;
  assign add_794844 = sel_794841 + 8'h01;
  assign sel_794845 = array_index_794540 == array_index_773092 ? add_794844 : sel_794841;
  assign add_794848 = sel_794845 + 8'h01;
  assign sel_794849 = array_index_794540 == array_index_773098 ? add_794848 : sel_794845;
  assign add_794852 = sel_794849 + 8'h01;
  assign sel_794853 = array_index_794540 == array_index_773104 ? add_794852 : sel_794849;
  assign add_794856 = sel_794853 + 8'h01;
  assign sel_794857 = array_index_794540 == array_index_773110 ? add_794856 : sel_794853;
  assign add_794860 = sel_794857 + 8'h01;
  assign sel_794861 = array_index_794540 == array_index_773116 ? add_794860 : sel_794857;
  assign add_794864 = sel_794861 + 8'h01;
  assign sel_794865 = array_index_794540 == array_index_773122 ? add_794864 : sel_794861;
  assign add_794868 = sel_794865 + 8'h01;
  assign sel_794869 = array_index_794540 == array_index_773128 ? add_794868 : sel_794865;
  assign add_794872 = sel_794869 + 8'h01;
  assign sel_794873 = array_index_794540 == array_index_773134 ? add_794872 : sel_794869;
  assign add_794876 = sel_794873 + 8'h01;
  assign sel_794877 = array_index_794540 == array_index_773140 ? add_794876 : sel_794873;
  assign add_794880 = sel_794877 + 8'h01;
  assign sel_794881 = array_index_794540 == array_index_773146 ? add_794880 : sel_794877;
  assign add_794884 = sel_794881 + 8'h01;
  assign sel_794885 = array_index_794540 == array_index_773152 ? add_794884 : sel_794881;
  assign add_794888 = sel_794885 + 8'h01;
  assign sel_794889 = array_index_794540 == array_index_773158 ? add_794888 : sel_794885;
  assign add_794892 = sel_794889 + 8'h01;
  assign sel_794893 = array_index_794540 == array_index_773164 ? add_794892 : sel_794889;
  assign add_794896 = sel_794893 + 8'h01;
  assign sel_794897 = array_index_794540 == array_index_773170 ? add_794896 : sel_794893;
  assign add_794901 = sel_794897 + 8'h01;
  assign array_index_794902 = set1_unflattened[7'h3d];
  assign sel_794903 = array_index_794540 == array_index_773176 ? add_794901 : sel_794897;
  assign add_794906 = sel_794903 + 8'h01;
  assign sel_794907 = array_index_794902 == array_index_772632 ? add_794906 : sel_794903;
  assign add_794910 = sel_794907 + 8'h01;
  assign sel_794911 = array_index_794902 == array_index_772636 ? add_794910 : sel_794907;
  assign add_794914 = sel_794911 + 8'h01;
  assign sel_794915 = array_index_794902 == array_index_772644 ? add_794914 : sel_794911;
  assign add_794918 = sel_794915 + 8'h01;
  assign sel_794919 = array_index_794902 == array_index_772652 ? add_794918 : sel_794915;
  assign add_794922 = sel_794919 + 8'h01;
  assign sel_794923 = array_index_794902 == array_index_772660 ? add_794922 : sel_794919;
  assign add_794926 = sel_794923 + 8'h01;
  assign sel_794927 = array_index_794902 == array_index_772668 ? add_794926 : sel_794923;
  assign add_794930 = sel_794927 + 8'h01;
  assign sel_794931 = array_index_794902 == array_index_772676 ? add_794930 : sel_794927;
  assign add_794934 = sel_794931 + 8'h01;
  assign sel_794935 = array_index_794902 == array_index_772684 ? add_794934 : sel_794931;
  assign add_794938 = sel_794935 + 8'h01;
  assign sel_794939 = array_index_794902 == array_index_772690 ? add_794938 : sel_794935;
  assign add_794942 = sel_794939 + 8'h01;
  assign sel_794943 = array_index_794902 == array_index_772696 ? add_794942 : sel_794939;
  assign add_794946 = sel_794943 + 8'h01;
  assign sel_794947 = array_index_794902 == array_index_772702 ? add_794946 : sel_794943;
  assign add_794950 = sel_794947 + 8'h01;
  assign sel_794951 = array_index_794902 == array_index_772708 ? add_794950 : sel_794947;
  assign add_794954 = sel_794951 + 8'h01;
  assign sel_794955 = array_index_794902 == array_index_772714 ? add_794954 : sel_794951;
  assign add_794958 = sel_794955 + 8'h01;
  assign sel_794959 = array_index_794902 == array_index_772720 ? add_794958 : sel_794955;
  assign add_794962 = sel_794959 + 8'h01;
  assign sel_794963 = array_index_794902 == array_index_772726 ? add_794962 : sel_794959;
  assign add_794966 = sel_794963 + 8'h01;
  assign sel_794967 = array_index_794902 == array_index_772732 ? add_794966 : sel_794963;
  assign add_794970 = sel_794967 + 8'h01;
  assign sel_794971 = array_index_794902 == array_index_772738 ? add_794970 : sel_794967;
  assign add_794974 = sel_794971 + 8'h01;
  assign sel_794975 = array_index_794902 == array_index_772744 ? add_794974 : sel_794971;
  assign add_794978 = sel_794975 + 8'h01;
  assign sel_794979 = array_index_794902 == array_index_772750 ? add_794978 : sel_794975;
  assign add_794982 = sel_794979 + 8'h01;
  assign sel_794983 = array_index_794902 == array_index_772756 ? add_794982 : sel_794979;
  assign add_794986 = sel_794983 + 8'h01;
  assign sel_794987 = array_index_794902 == array_index_772762 ? add_794986 : sel_794983;
  assign add_794990 = sel_794987 + 8'h01;
  assign sel_794991 = array_index_794902 == array_index_772768 ? add_794990 : sel_794987;
  assign add_794994 = sel_794991 + 8'h01;
  assign sel_794995 = array_index_794902 == array_index_772774 ? add_794994 : sel_794991;
  assign add_794998 = sel_794995 + 8'h01;
  assign sel_794999 = array_index_794902 == array_index_772780 ? add_794998 : sel_794995;
  assign add_795002 = sel_794999 + 8'h01;
  assign sel_795003 = array_index_794902 == array_index_772786 ? add_795002 : sel_794999;
  assign add_795006 = sel_795003 + 8'h01;
  assign sel_795007 = array_index_794902 == array_index_772792 ? add_795006 : sel_795003;
  assign add_795010 = sel_795007 + 8'h01;
  assign sel_795011 = array_index_794902 == array_index_772798 ? add_795010 : sel_795007;
  assign add_795014 = sel_795011 + 8'h01;
  assign sel_795015 = array_index_794902 == array_index_772804 ? add_795014 : sel_795011;
  assign add_795018 = sel_795015 + 8'h01;
  assign sel_795019 = array_index_794902 == array_index_772810 ? add_795018 : sel_795015;
  assign add_795022 = sel_795019 + 8'h01;
  assign sel_795023 = array_index_794902 == array_index_772816 ? add_795022 : sel_795019;
  assign add_795026 = sel_795023 + 8'h01;
  assign sel_795027 = array_index_794902 == array_index_772822 ? add_795026 : sel_795023;
  assign add_795030 = sel_795027 + 8'h01;
  assign sel_795031 = array_index_794902 == array_index_772828 ? add_795030 : sel_795027;
  assign add_795034 = sel_795031 + 8'h01;
  assign sel_795035 = array_index_794902 == array_index_772834 ? add_795034 : sel_795031;
  assign add_795038 = sel_795035 + 8'h01;
  assign sel_795039 = array_index_794902 == array_index_772840 ? add_795038 : sel_795035;
  assign add_795042 = sel_795039 + 8'h01;
  assign sel_795043 = array_index_794902 == array_index_772846 ? add_795042 : sel_795039;
  assign add_795046 = sel_795043 + 8'h01;
  assign sel_795047 = array_index_794902 == array_index_772852 ? add_795046 : sel_795043;
  assign add_795050 = sel_795047 + 8'h01;
  assign sel_795051 = array_index_794902 == array_index_772858 ? add_795050 : sel_795047;
  assign add_795054 = sel_795051 + 8'h01;
  assign sel_795055 = array_index_794902 == array_index_772864 ? add_795054 : sel_795051;
  assign add_795058 = sel_795055 + 8'h01;
  assign sel_795059 = array_index_794902 == array_index_772870 ? add_795058 : sel_795055;
  assign add_795062 = sel_795059 + 8'h01;
  assign sel_795063 = array_index_794902 == array_index_772876 ? add_795062 : sel_795059;
  assign add_795066 = sel_795063 + 8'h01;
  assign sel_795067 = array_index_794902 == array_index_772882 ? add_795066 : sel_795063;
  assign add_795070 = sel_795067 + 8'h01;
  assign sel_795071 = array_index_794902 == array_index_772888 ? add_795070 : sel_795067;
  assign add_795074 = sel_795071 + 8'h01;
  assign sel_795075 = array_index_794902 == array_index_772894 ? add_795074 : sel_795071;
  assign add_795078 = sel_795075 + 8'h01;
  assign sel_795079 = array_index_794902 == array_index_772900 ? add_795078 : sel_795075;
  assign add_795082 = sel_795079 + 8'h01;
  assign sel_795083 = array_index_794902 == array_index_772906 ? add_795082 : sel_795079;
  assign add_795086 = sel_795083 + 8'h01;
  assign sel_795087 = array_index_794902 == array_index_772912 ? add_795086 : sel_795083;
  assign add_795090 = sel_795087 + 8'h01;
  assign sel_795091 = array_index_794902 == array_index_772918 ? add_795090 : sel_795087;
  assign add_795094 = sel_795091 + 8'h01;
  assign sel_795095 = array_index_794902 == array_index_772924 ? add_795094 : sel_795091;
  assign add_795098 = sel_795095 + 8'h01;
  assign sel_795099 = array_index_794902 == array_index_772930 ? add_795098 : sel_795095;
  assign add_795102 = sel_795099 + 8'h01;
  assign sel_795103 = array_index_794902 == array_index_772936 ? add_795102 : sel_795099;
  assign add_795106 = sel_795103 + 8'h01;
  assign sel_795107 = array_index_794902 == array_index_772942 ? add_795106 : sel_795103;
  assign add_795110 = sel_795107 + 8'h01;
  assign sel_795111 = array_index_794902 == array_index_772948 ? add_795110 : sel_795107;
  assign add_795114 = sel_795111 + 8'h01;
  assign sel_795115 = array_index_794902 == array_index_772954 ? add_795114 : sel_795111;
  assign add_795118 = sel_795115 + 8'h01;
  assign sel_795119 = array_index_794902 == array_index_772960 ? add_795118 : sel_795115;
  assign add_795122 = sel_795119 + 8'h01;
  assign sel_795123 = array_index_794902 == array_index_772966 ? add_795122 : sel_795119;
  assign add_795126 = sel_795123 + 8'h01;
  assign sel_795127 = array_index_794902 == array_index_772972 ? add_795126 : sel_795123;
  assign add_795130 = sel_795127 + 8'h01;
  assign sel_795131 = array_index_794902 == array_index_772978 ? add_795130 : sel_795127;
  assign add_795134 = sel_795131 + 8'h01;
  assign sel_795135 = array_index_794902 == array_index_772984 ? add_795134 : sel_795131;
  assign add_795138 = sel_795135 + 8'h01;
  assign sel_795139 = array_index_794902 == array_index_772990 ? add_795138 : sel_795135;
  assign add_795142 = sel_795139 + 8'h01;
  assign sel_795143 = array_index_794902 == array_index_772996 ? add_795142 : sel_795139;
  assign add_795146 = sel_795143 + 8'h01;
  assign sel_795147 = array_index_794902 == array_index_773002 ? add_795146 : sel_795143;
  assign add_795150 = sel_795147 + 8'h01;
  assign sel_795151 = array_index_794902 == array_index_773008 ? add_795150 : sel_795147;
  assign add_795154 = sel_795151 + 8'h01;
  assign sel_795155 = array_index_794902 == array_index_773014 ? add_795154 : sel_795151;
  assign add_795158 = sel_795155 + 8'h01;
  assign sel_795159 = array_index_794902 == array_index_773020 ? add_795158 : sel_795155;
  assign add_795162 = sel_795159 + 8'h01;
  assign sel_795163 = array_index_794902 == array_index_773026 ? add_795162 : sel_795159;
  assign add_795166 = sel_795163 + 8'h01;
  assign sel_795167 = array_index_794902 == array_index_773032 ? add_795166 : sel_795163;
  assign add_795170 = sel_795167 + 8'h01;
  assign sel_795171 = array_index_794902 == array_index_773038 ? add_795170 : sel_795167;
  assign add_795174 = sel_795171 + 8'h01;
  assign sel_795175 = array_index_794902 == array_index_773044 ? add_795174 : sel_795171;
  assign add_795178 = sel_795175 + 8'h01;
  assign sel_795179 = array_index_794902 == array_index_773050 ? add_795178 : sel_795175;
  assign add_795182 = sel_795179 + 8'h01;
  assign sel_795183 = array_index_794902 == array_index_773056 ? add_795182 : sel_795179;
  assign add_795186 = sel_795183 + 8'h01;
  assign sel_795187 = array_index_794902 == array_index_773062 ? add_795186 : sel_795183;
  assign add_795190 = sel_795187 + 8'h01;
  assign sel_795191 = array_index_794902 == array_index_773068 ? add_795190 : sel_795187;
  assign add_795194 = sel_795191 + 8'h01;
  assign sel_795195 = array_index_794902 == array_index_773074 ? add_795194 : sel_795191;
  assign add_795198 = sel_795195 + 8'h01;
  assign sel_795199 = array_index_794902 == array_index_773080 ? add_795198 : sel_795195;
  assign add_795202 = sel_795199 + 8'h01;
  assign sel_795203 = array_index_794902 == array_index_773086 ? add_795202 : sel_795199;
  assign add_795206 = sel_795203 + 8'h01;
  assign sel_795207 = array_index_794902 == array_index_773092 ? add_795206 : sel_795203;
  assign add_795210 = sel_795207 + 8'h01;
  assign sel_795211 = array_index_794902 == array_index_773098 ? add_795210 : sel_795207;
  assign add_795214 = sel_795211 + 8'h01;
  assign sel_795215 = array_index_794902 == array_index_773104 ? add_795214 : sel_795211;
  assign add_795218 = sel_795215 + 8'h01;
  assign sel_795219 = array_index_794902 == array_index_773110 ? add_795218 : sel_795215;
  assign add_795222 = sel_795219 + 8'h01;
  assign sel_795223 = array_index_794902 == array_index_773116 ? add_795222 : sel_795219;
  assign add_795226 = sel_795223 + 8'h01;
  assign sel_795227 = array_index_794902 == array_index_773122 ? add_795226 : sel_795223;
  assign add_795230 = sel_795227 + 8'h01;
  assign sel_795231 = array_index_794902 == array_index_773128 ? add_795230 : sel_795227;
  assign add_795234 = sel_795231 + 8'h01;
  assign sel_795235 = array_index_794902 == array_index_773134 ? add_795234 : sel_795231;
  assign add_795238 = sel_795235 + 8'h01;
  assign sel_795239 = array_index_794902 == array_index_773140 ? add_795238 : sel_795235;
  assign add_795242 = sel_795239 + 8'h01;
  assign sel_795243 = array_index_794902 == array_index_773146 ? add_795242 : sel_795239;
  assign add_795246 = sel_795243 + 8'h01;
  assign sel_795247 = array_index_794902 == array_index_773152 ? add_795246 : sel_795243;
  assign add_795250 = sel_795247 + 8'h01;
  assign sel_795251 = array_index_794902 == array_index_773158 ? add_795250 : sel_795247;
  assign add_795254 = sel_795251 + 8'h01;
  assign sel_795255 = array_index_794902 == array_index_773164 ? add_795254 : sel_795251;
  assign add_795258 = sel_795255 + 8'h01;
  assign sel_795259 = array_index_794902 == array_index_773170 ? add_795258 : sel_795255;
  assign add_795263 = sel_795259 + 8'h01;
  assign array_index_795264 = set1_unflattened[7'h3e];
  assign sel_795265 = array_index_794902 == array_index_773176 ? add_795263 : sel_795259;
  assign add_795268 = sel_795265 + 8'h01;
  assign sel_795269 = array_index_795264 == array_index_772632 ? add_795268 : sel_795265;
  assign add_795272 = sel_795269 + 8'h01;
  assign sel_795273 = array_index_795264 == array_index_772636 ? add_795272 : sel_795269;
  assign add_795276 = sel_795273 + 8'h01;
  assign sel_795277 = array_index_795264 == array_index_772644 ? add_795276 : sel_795273;
  assign add_795280 = sel_795277 + 8'h01;
  assign sel_795281 = array_index_795264 == array_index_772652 ? add_795280 : sel_795277;
  assign add_795284 = sel_795281 + 8'h01;
  assign sel_795285 = array_index_795264 == array_index_772660 ? add_795284 : sel_795281;
  assign add_795288 = sel_795285 + 8'h01;
  assign sel_795289 = array_index_795264 == array_index_772668 ? add_795288 : sel_795285;
  assign add_795292 = sel_795289 + 8'h01;
  assign sel_795293 = array_index_795264 == array_index_772676 ? add_795292 : sel_795289;
  assign add_795296 = sel_795293 + 8'h01;
  assign sel_795297 = array_index_795264 == array_index_772684 ? add_795296 : sel_795293;
  assign add_795300 = sel_795297 + 8'h01;
  assign sel_795301 = array_index_795264 == array_index_772690 ? add_795300 : sel_795297;
  assign add_795304 = sel_795301 + 8'h01;
  assign sel_795305 = array_index_795264 == array_index_772696 ? add_795304 : sel_795301;
  assign add_795308 = sel_795305 + 8'h01;
  assign sel_795309 = array_index_795264 == array_index_772702 ? add_795308 : sel_795305;
  assign add_795312 = sel_795309 + 8'h01;
  assign sel_795313 = array_index_795264 == array_index_772708 ? add_795312 : sel_795309;
  assign add_795316 = sel_795313 + 8'h01;
  assign sel_795317 = array_index_795264 == array_index_772714 ? add_795316 : sel_795313;
  assign add_795320 = sel_795317 + 8'h01;
  assign sel_795321 = array_index_795264 == array_index_772720 ? add_795320 : sel_795317;
  assign add_795324 = sel_795321 + 8'h01;
  assign sel_795325 = array_index_795264 == array_index_772726 ? add_795324 : sel_795321;
  assign add_795328 = sel_795325 + 8'h01;
  assign sel_795329 = array_index_795264 == array_index_772732 ? add_795328 : sel_795325;
  assign add_795332 = sel_795329 + 8'h01;
  assign sel_795333 = array_index_795264 == array_index_772738 ? add_795332 : sel_795329;
  assign add_795336 = sel_795333 + 8'h01;
  assign sel_795337 = array_index_795264 == array_index_772744 ? add_795336 : sel_795333;
  assign add_795340 = sel_795337 + 8'h01;
  assign sel_795341 = array_index_795264 == array_index_772750 ? add_795340 : sel_795337;
  assign add_795344 = sel_795341 + 8'h01;
  assign sel_795345 = array_index_795264 == array_index_772756 ? add_795344 : sel_795341;
  assign add_795348 = sel_795345 + 8'h01;
  assign sel_795349 = array_index_795264 == array_index_772762 ? add_795348 : sel_795345;
  assign add_795352 = sel_795349 + 8'h01;
  assign sel_795353 = array_index_795264 == array_index_772768 ? add_795352 : sel_795349;
  assign add_795356 = sel_795353 + 8'h01;
  assign sel_795357 = array_index_795264 == array_index_772774 ? add_795356 : sel_795353;
  assign add_795360 = sel_795357 + 8'h01;
  assign sel_795361 = array_index_795264 == array_index_772780 ? add_795360 : sel_795357;
  assign add_795364 = sel_795361 + 8'h01;
  assign sel_795365 = array_index_795264 == array_index_772786 ? add_795364 : sel_795361;
  assign add_795368 = sel_795365 + 8'h01;
  assign sel_795369 = array_index_795264 == array_index_772792 ? add_795368 : sel_795365;
  assign add_795372 = sel_795369 + 8'h01;
  assign sel_795373 = array_index_795264 == array_index_772798 ? add_795372 : sel_795369;
  assign add_795376 = sel_795373 + 8'h01;
  assign sel_795377 = array_index_795264 == array_index_772804 ? add_795376 : sel_795373;
  assign add_795380 = sel_795377 + 8'h01;
  assign sel_795381 = array_index_795264 == array_index_772810 ? add_795380 : sel_795377;
  assign add_795384 = sel_795381 + 8'h01;
  assign sel_795385 = array_index_795264 == array_index_772816 ? add_795384 : sel_795381;
  assign add_795388 = sel_795385 + 8'h01;
  assign sel_795389 = array_index_795264 == array_index_772822 ? add_795388 : sel_795385;
  assign add_795392 = sel_795389 + 8'h01;
  assign sel_795393 = array_index_795264 == array_index_772828 ? add_795392 : sel_795389;
  assign add_795396 = sel_795393 + 8'h01;
  assign sel_795397 = array_index_795264 == array_index_772834 ? add_795396 : sel_795393;
  assign add_795400 = sel_795397 + 8'h01;
  assign sel_795401 = array_index_795264 == array_index_772840 ? add_795400 : sel_795397;
  assign add_795404 = sel_795401 + 8'h01;
  assign sel_795405 = array_index_795264 == array_index_772846 ? add_795404 : sel_795401;
  assign add_795408 = sel_795405 + 8'h01;
  assign sel_795409 = array_index_795264 == array_index_772852 ? add_795408 : sel_795405;
  assign add_795412 = sel_795409 + 8'h01;
  assign sel_795413 = array_index_795264 == array_index_772858 ? add_795412 : sel_795409;
  assign add_795416 = sel_795413 + 8'h01;
  assign sel_795417 = array_index_795264 == array_index_772864 ? add_795416 : sel_795413;
  assign add_795420 = sel_795417 + 8'h01;
  assign sel_795421 = array_index_795264 == array_index_772870 ? add_795420 : sel_795417;
  assign add_795424 = sel_795421 + 8'h01;
  assign sel_795425 = array_index_795264 == array_index_772876 ? add_795424 : sel_795421;
  assign add_795428 = sel_795425 + 8'h01;
  assign sel_795429 = array_index_795264 == array_index_772882 ? add_795428 : sel_795425;
  assign add_795432 = sel_795429 + 8'h01;
  assign sel_795433 = array_index_795264 == array_index_772888 ? add_795432 : sel_795429;
  assign add_795436 = sel_795433 + 8'h01;
  assign sel_795437 = array_index_795264 == array_index_772894 ? add_795436 : sel_795433;
  assign add_795440 = sel_795437 + 8'h01;
  assign sel_795441 = array_index_795264 == array_index_772900 ? add_795440 : sel_795437;
  assign add_795444 = sel_795441 + 8'h01;
  assign sel_795445 = array_index_795264 == array_index_772906 ? add_795444 : sel_795441;
  assign add_795448 = sel_795445 + 8'h01;
  assign sel_795449 = array_index_795264 == array_index_772912 ? add_795448 : sel_795445;
  assign add_795452 = sel_795449 + 8'h01;
  assign sel_795453 = array_index_795264 == array_index_772918 ? add_795452 : sel_795449;
  assign add_795456 = sel_795453 + 8'h01;
  assign sel_795457 = array_index_795264 == array_index_772924 ? add_795456 : sel_795453;
  assign add_795460 = sel_795457 + 8'h01;
  assign sel_795461 = array_index_795264 == array_index_772930 ? add_795460 : sel_795457;
  assign add_795464 = sel_795461 + 8'h01;
  assign sel_795465 = array_index_795264 == array_index_772936 ? add_795464 : sel_795461;
  assign add_795468 = sel_795465 + 8'h01;
  assign sel_795469 = array_index_795264 == array_index_772942 ? add_795468 : sel_795465;
  assign add_795472 = sel_795469 + 8'h01;
  assign sel_795473 = array_index_795264 == array_index_772948 ? add_795472 : sel_795469;
  assign add_795476 = sel_795473 + 8'h01;
  assign sel_795477 = array_index_795264 == array_index_772954 ? add_795476 : sel_795473;
  assign add_795480 = sel_795477 + 8'h01;
  assign sel_795481 = array_index_795264 == array_index_772960 ? add_795480 : sel_795477;
  assign add_795484 = sel_795481 + 8'h01;
  assign sel_795485 = array_index_795264 == array_index_772966 ? add_795484 : sel_795481;
  assign add_795488 = sel_795485 + 8'h01;
  assign sel_795489 = array_index_795264 == array_index_772972 ? add_795488 : sel_795485;
  assign add_795492 = sel_795489 + 8'h01;
  assign sel_795493 = array_index_795264 == array_index_772978 ? add_795492 : sel_795489;
  assign add_795496 = sel_795493 + 8'h01;
  assign sel_795497 = array_index_795264 == array_index_772984 ? add_795496 : sel_795493;
  assign add_795500 = sel_795497 + 8'h01;
  assign sel_795501 = array_index_795264 == array_index_772990 ? add_795500 : sel_795497;
  assign add_795504 = sel_795501 + 8'h01;
  assign sel_795505 = array_index_795264 == array_index_772996 ? add_795504 : sel_795501;
  assign add_795508 = sel_795505 + 8'h01;
  assign sel_795509 = array_index_795264 == array_index_773002 ? add_795508 : sel_795505;
  assign add_795512 = sel_795509 + 8'h01;
  assign sel_795513 = array_index_795264 == array_index_773008 ? add_795512 : sel_795509;
  assign add_795516 = sel_795513 + 8'h01;
  assign sel_795517 = array_index_795264 == array_index_773014 ? add_795516 : sel_795513;
  assign add_795520 = sel_795517 + 8'h01;
  assign sel_795521 = array_index_795264 == array_index_773020 ? add_795520 : sel_795517;
  assign add_795524 = sel_795521 + 8'h01;
  assign sel_795525 = array_index_795264 == array_index_773026 ? add_795524 : sel_795521;
  assign add_795528 = sel_795525 + 8'h01;
  assign sel_795529 = array_index_795264 == array_index_773032 ? add_795528 : sel_795525;
  assign add_795532 = sel_795529 + 8'h01;
  assign sel_795533 = array_index_795264 == array_index_773038 ? add_795532 : sel_795529;
  assign add_795536 = sel_795533 + 8'h01;
  assign sel_795537 = array_index_795264 == array_index_773044 ? add_795536 : sel_795533;
  assign add_795540 = sel_795537 + 8'h01;
  assign sel_795541 = array_index_795264 == array_index_773050 ? add_795540 : sel_795537;
  assign add_795544 = sel_795541 + 8'h01;
  assign sel_795545 = array_index_795264 == array_index_773056 ? add_795544 : sel_795541;
  assign add_795548 = sel_795545 + 8'h01;
  assign sel_795549 = array_index_795264 == array_index_773062 ? add_795548 : sel_795545;
  assign add_795552 = sel_795549 + 8'h01;
  assign sel_795553 = array_index_795264 == array_index_773068 ? add_795552 : sel_795549;
  assign add_795556 = sel_795553 + 8'h01;
  assign sel_795557 = array_index_795264 == array_index_773074 ? add_795556 : sel_795553;
  assign add_795560 = sel_795557 + 8'h01;
  assign sel_795561 = array_index_795264 == array_index_773080 ? add_795560 : sel_795557;
  assign add_795564 = sel_795561 + 8'h01;
  assign sel_795565 = array_index_795264 == array_index_773086 ? add_795564 : sel_795561;
  assign add_795568 = sel_795565 + 8'h01;
  assign sel_795569 = array_index_795264 == array_index_773092 ? add_795568 : sel_795565;
  assign add_795572 = sel_795569 + 8'h01;
  assign sel_795573 = array_index_795264 == array_index_773098 ? add_795572 : sel_795569;
  assign add_795576 = sel_795573 + 8'h01;
  assign sel_795577 = array_index_795264 == array_index_773104 ? add_795576 : sel_795573;
  assign add_795580 = sel_795577 + 8'h01;
  assign sel_795581 = array_index_795264 == array_index_773110 ? add_795580 : sel_795577;
  assign add_795584 = sel_795581 + 8'h01;
  assign sel_795585 = array_index_795264 == array_index_773116 ? add_795584 : sel_795581;
  assign add_795588 = sel_795585 + 8'h01;
  assign sel_795589 = array_index_795264 == array_index_773122 ? add_795588 : sel_795585;
  assign add_795592 = sel_795589 + 8'h01;
  assign sel_795593 = array_index_795264 == array_index_773128 ? add_795592 : sel_795589;
  assign add_795596 = sel_795593 + 8'h01;
  assign sel_795597 = array_index_795264 == array_index_773134 ? add_795596 : sel_795593;
  assign add_795600 = sel_795597 + 8'h01;
  assign sel_795601 = array_index_795264 == array_index_773140 ? add_795600 : sel_795597;
  assign add_795604 = sel_795601 + 8'h01;
  assign sel_795605 = array_index_795264 == array_index_773146 ? add_795604 : sel_795601;
  assign add_795608 = sel_795605 + 8'h01;
  assign sel_795609 = array_index_795264 == array_index_773152 ? add_795608 : sel_795605;
  assign add_795612 = sel_795609 + 8'h01;
  assign sel_795613 = array_index_795264 == array_index_773158 ? add_795612 : sel_795609;
  assign add_795616 = sel_795613 + 8'h01;
  assign sel_795617 = array_index_795264 == array_index_773164 ? add_795616 : sel_795613;
  assign add_795620 = sel_795617 + 8'h01;
  assign sel_795621 = array_index_795264 == array_index_773170 ? add_795620 : sel_795617;
  assign add_795625 = sel_795621 + 8'h01;
  assign array_index_795626 = set1_unflattened[7'h3f];
  assign sel_795627 = array_index_795264 == array_index_773176 ? add_795625 : sel_795621;
  assign add_795630 = sel_795627 + 8'h01;
  assign sel_795631 = array_index_795626 == array_index_772632 ? add_795630 : sel_795627;
  assign add_795634 = sel_795631 + 8'h01;
  assign sel_795635 = array_index_795626 == array_index_772636 ? add_795634 : sel_795631;
  assign add_795638 = sel_795635 + 8'h01;
  assign sel_795639 = array_index_795626 == array_index_772644 ? add_795638 : sel_795635;
  assign add_795642 = sel_795639 + 8'h01;
  assign sel_795643 = array_index_795626 == array_index_772652 ? add_795642 : sel_795639;
  assign add_795646 = sel_795643 + 8'h01;
  assign sel_795647 = array_index_795626 == array_index_772660 ? add_795646 : sel_795643;
  assign add_795650 = sel_795647 + 8'h01;
  assign sel_795651 = array_index_795626 == array_index_772668 ? add_795650 : sel_795647;
  assign add_795654 = sel_795651 + 8'h01;
  assign sel_795655 = array_index_795626 == array_index_772676 ? add_795654 : sel_795651;
  assign add_795658 = sel_795655 + 8'h01;
  assign sel_795659 = array_index_795626 == array_index_772684 ? add_795658 : sel_795655;
  assign add_795662 = sel_795659 + 8'h01;
  assign sel_795663 = array_index_795626 == array_index_772690 ? add_795662 : sel_795659;
  assign add_795666 = sel_795663 + 8'h01;
  assign sel_795667 = array_index_795626 == array_index_772696 ? add_795666 : sel_795663;
  assign add_795670 = sel_795667 + 8'h01;
  assign sel_795671 = array_index_795626 == array_index_772702 ? add_795670 : sel_795667;
  assign add_795674 = sel_795671 + 8'h01;
  assign sel_795675 = array_index_795626 == array_index_772708 ? add_795674 : sel_795671;
  assign add_795678 = sel_795675 + 8'h01;
  assign sel_795679 = array_index_795626 == array_index_772714 ? add_795678 : sel_795675;
  assign add_795682 = sel_795679 + 8'h01;
  assign sel_795683 = array_index_795626 == array_index_772720 ? add_795682 : sel_795679;
  assign add_795686 = sel_795683 + 8'h01;
  assign sel_795687 = array_index_795626 == array_index_772726 ? add_795686 : sel_795683;
  assign add_795690 = sel_795687 + 8'h01;
  assign sel_795691 = array_index_795626 == array_index_772732 ? add_795690 : sel_795687;
  assign add_795694 = sel_795691 + 8'h01;
  assign sel_795695 = array_index_795626 == array_index_772738 ? add_795694 : sel_795691;
  assign add_795698 = sel_795695 + 8'h01;
  assign sel_795699 = array_index_795626 == array_index_772744 ? add_795698 : sel_795695;
  assign add_795702 = sel_795699 + 8'h01;
  assign sel_795703 = array_index_795626 == array_index_772750 ? add_795702 : sel_795699;
  assign add_795706 = sel_795703 + 8'h01;
  assign sel_795707 = array_index_795626 == array_index_772756 ? add_795706 : sel_795703;
  assign add_795710 = sel_795707 + 8'h01;
  assign sel_795711 = array_index_795626 == array_index_772762 ? add_795710 : sel_795707;
  assign add_795714 = sel_795711 + 8'h01;
  assign sel_795715 = array_index_795626 == array_index_772768 ? add_795714 : sel_795711;
  assign add_795718 = sel_795715 + 8'h01;
  assign sel_795719 = array_index_795626 == array_index_772774 ? add_795718 : sel_795715;
  assign add_795722 = sel_795719 + 8'h01;
  assign sel_795723 = array_index_795626 == array_index_772780 ? add_795722 : sel_795719;
  assign add_795726 = sel_795723 + 8'h01;
  assign sel_795727 = array_index_795626 == array_index_772786 ? add_795726 : sel_795723;
  assign add_795730 = sel_795727 + 8'h01;
  assign sel_795731 = array_index_795626 == array_index_772792 ? add_795730 : sel_795727;
  assign add_795734 = sel_795731 + 8'h01;
  assign sel_795735 = array_index_795626 == array_index_772798 ? add_795734 : sel_795731;
  assign add_795738 = sel_795735 + 8'h01;
  assign sel_795739 = array_index_795626 == array_index_772804 ? add_795738 : sel_795735;
  assign add_795742 = sel_795739 + 8'h01;
  assign sel_795743 = array_index_795626 == array_index_772810 ? add_795742 : sel_795739;
  assign add_795746 = sel_795743 + 8'h01;
  assign sel_795747 = array_index_795626 == array_index_772816 ? add_795746 : sel_795743;
  assign add_795750 = sel_795747 + 8'h01;
  assign sel_795751 = array_index_795626 == array_index_772822 ? add_795750 : sel_795747;
  assign add_795754 = sel_795751 + 8'h01;
  assign sel_795755 = array_index_795626 == array_index_772828 ? add_795754 : sel_795751;
  assign add_795758 = sel_795755 + 8'h01;
  assign sel_795759 = array_index_795626 == array_index_772834 ? add_795758 : sel_795755;
  assign add_795762 = sel_795759 + 8'h01;
  assign sel_795763 = array_index_795626 == array_index_772840 ? add_795762 : sel_795759;
  assign add_795766 = sel_795763 + 8'h01;
  assign sel_795767 = array_index_795626 == array_index_772846 ? add_795766 : sel_795763;
  assign add_795770 = sel_795767 + 8'h01;
  assign sel_795771 = array_index_795626 == array_index_772852 ? add_795770 : sel_795767;
  assign add_795774 = sel_795771 + 8'h01;
  assign sel_795775 = array_index_795626 == array_index_772858 ? add_795774 : sel_795771;
  assign add_795778 = sel_795775 + 8'h01;
  assign sel_795779 = array_index_795626 == array_index_772864 ? add_795778 : sel_795775;
  assign add_795782 = sel_795779 + 8'h01;
  assign sel_795783 = array_index_795626 == array_index_772870 ? add_795782 : sel_795779;
  assign add_795786 = sel_795783 + 8'h01;
  assign sel_795787 = array_index_795626 == array_index_772876 ? add_795786 : sel_795783;
  assign add_795790 = sel_795787 + 8'h01;
  assign sel_795791 = array_index_795626 == array_index_772882 ? add_795790 : sel_795787;
  assign add_795794 = sel_795791 + 8'h01;
  assign sel_795795 = array_index_795626 == array_index_772888 ? add_795794 : sel_795791;
  assign add_795798 = sel_795795 + 8'h01;
  assign sel_795799 = array_index_795626 == array_index_772894 ? add_795798 : sel_795795;
  assign add_795802 = sel_795799 + 8'h01;
  assign sel_795803 = array_index_795626 == array_index_772900 ? add_795802 : sel_795799;
  assign add_795806 = sel_795803 + 8'h01;
  assign sel_795807 = array_index_795626 == array_index_772906 ? add_795806 : sel_795803;
  assign add_795810 = sel_795807 + 8'h01;
  assign sel_795811 = array_index_795626 == array_index_772912 ? add_795810 : sel_795807;
  assign add_795814 = sel_795811 + 8'h01;
  assign sel_795815 = array_index_795626 == array_index_772918 ? add_795814 : sel_795811;
  assign add_795818 = sel_795815 + 8'h01;
  assign sel_795819 = array_index_795626 == array_index_772924 ? add_795818 : sel_795815;
  assign add_795822 = sel_795819 + 8'h01;
  assign sel_795823 = array_index_795626 == array_index_772930 ? add_795822 : sel_795819;
  assign add_795826 = sel_795823 + 8'h01;
  assign sel_795827 = array_index_795626 == array_index_772936 ? add_795826 : sel_795823;
  assign add_795830 = sel_795827 + 8'h01;
  assign sel_795831 = array_index_795626 == array_index_772942 ? add_795830 : sel_795827;
  assign add_795834 = sel_795831 + 8'h01;
  assign sel_795835 = array_index_795626 == array_index_772948 ? add_795834 : sel_795831;
  assign add_795838 = sel_795835 + 8'h01;
  assign sel_795839 = array_index_795626 == array_index_772954 ? add_795838 : sel_795835;
  assign add_795842 = sel_795839 + 8'h01;
  assign sel_795843 = array_index_795626 == array_index_772960 ? add_795842 : sel_795839;
  assign add_795846 = sel_795843 + 8'h01;
  assign sel_795847 = array_index_795626 == array_index_772966 ? add_795846 : sel_795843;
  assign add_795850 = sel_795847 + 8'h01;
  assign sel_795851 = array_index_795626 == array_index_772972 ? add_795850 : sel_795847;
  assign add_795854 = sel_795851 + 8'h01;
  assign sel_795855 = array_index_795626 == array_index_772978 ? add_795854 : sel_795851;
  assign add_795858 = sel_795855 + 8'h01;
  assign sel_795859 = array_index_795626 == array_index_772984 ? add_795858 : sel_795855;
  assign add_795862 = sel_795859 + 8'h01;
  assign sel_795863 = array_index_795626 == array_index_772990 ? add_795862 : sel_795859;
  assign add_795866 = sel_795863 + 8'h01;
  assign sel_795867 = array_index_795626 == array_index_772996 ? add_795866 : sel_795863;
  assign add_795870 = sel_795867 + 8'h01;
  assign sel_795871 = array_index_795626 == array_index_773002 ? add_795870 : sel_795867;
  assign add_795874 = sel_795871 + 8'h01;
  assign sel_795875 = array_index_795626 == array_index_773008 ? add_795874 : sel_795871;
  assign add_795878 = sel_795875 + 8'h01;
  assign sel_795879 = array_index_795626 == array_index_773014 ? add_795878 : sel_795875;
  assign add_795882 = sel_795879 + 8'h01;
  assign sel_795883 = array_index_795626 == array_index_773020 ? add_795882 : sel_795879;
  assign add_795886 = sel_795883 + 8'h01;
  assign sel_795887 = array_index_795626 == array_index_773026 ? add_795886 : sel_795883;
  assign add_795890 = sel_795887 + 8'h01;
  assign sel_795891 = array_index_795626 == array_index_773032 ? add_795890 : sel_795887;
  assign add_795894 = sel_795891 + 8'h01;
  assign sel_795895 = array_index_795626 == array_index_773038 ? add_795894 : sel_795891;
  assign add_795898 = sel_795895 + 8'h01;
  assign sel_795899 = array_index_795626 == array_index_773044 ? add_795898 : sel_795895;
  assign add_795902 = sel_795899 + 8'h01;
  assign sel_795903 = array_index_795626 == array_index_773050 ? add_795902 : sel_795899;
  assign add_795906 = sel_795903 + 8'h01;
  assign sel_795907 = array_index_795626 == array_index_773056 ? add_795906 : sel_795903;
  assign add_795910 = sel_795907 + 8'h01;
  assign sel_795911 = array_index_795626 == array_index_773062 ? add_795910 : sel_795907;
  assign add_795914 = sel_795911 + 8'h01;
  assign sel_795915 = array_index_795626 == array_index_773068 ? add_795914 : sel_795911;
  assign add_795918 = sel_795915 + 8'h01;
  assign sel_795919 = array_index_795626 == array_index_773074 ? add_795918 : sel_795915;
  assign add_795922 = sel_795919 + 8'h01;
  assign sel_795923 = array_index_795626 == array_index_773080 ? add_795922 : sel_795919;
  assign add_795926 = sel_795923 + 8'h01;
  assign sel_795927 = array_index_795626 == array_index_773086 ? add_795926 : sel_795923;
  assign add_795930 = sel_795927 + 8'h01;
  assign sel_795931 = array_index_795626 == array_index_773092 ? add_795930 : sel_795927;
  assign add_795934 = sel_795931 + 8'h01;
  assign sel_795935 = array_index_795626 == array_index_773098 ? add_795934 : sel_795931;
  assign add_795938 = sel_795935 + 8'h01;
  assign sel_795939 = array_index_795626 == array_index_773104 ? add_795938 : sel_795935;
  assign add_795942 = sel_795939 + 8'h01;
  assign sel_795943 = array_index_795626 == array_index_773110 ? add_795942 : sel_795939;
  assign add_795946 = sel_795943 + 8'h01;
  assign sel_795947 = array_index_795626 == array_index_773116 ? add_795946 : sel_795943;
  assign add_795950 = sel_795947 + 8'h01;
  assign sel_795951 = array_index_795626 == array_index_773122 ? add_795950 : sel_795947;
  assign add_795954 = sel_795951 + 8'h01;
  assign sel_795955 = array_index_795626 == array_index_773128 ? add_795954 : sel_795951;
  assign add_795958 = sel_795955 + 8'h01;
  assign sel_795959 = array_index_795626 == array_index_773134 ? add_795958 : sel_795955;
  assign add_795962 = sel_795959 + 8'h01;
  assign sel_795963 = array_index_795626 == array_index_773140 ? add_795962 : sel_795959;
  assign add_795966 = sel_795963 + 8'h01;
  assign sel_795967 = array_index_795626 == array_index_773146 ? add_795966 : sel_795963;
  assign add_795970 = sel_795967 + 8'h01;
  assign sel_795971 = array_index_795626 == array_index_773152 ? add_795970 : sel_795967;
  assign add_795974 = sel_795971 + 8'h01;
  assign sel_795975 = array_index_795626 == array_index_773158 ? add_795974 : sel_795971;
  assign add_795978 = sel_795975 + 8'h01;
  assign sel_795979 = array_index_795626 == array_index_773164 ? add_795978 : sel_795975;
  assign add_795982 = sel_795979 + 8'h01;
  assign sel_795983 = array_index_795626 == array_index_773170 ? add_795982 : sel_795979;
  assign add_795987 = sel_795983 + 8'h01;
  assign array_index_795988 = set1_unflattened[7'h40];
  assign sel_795989 = array_index_795626 == array_index_773176 ? add_795987 : sel_795983;
  assign add_795992 = sel_795989 + 8'h01;
  assign sel_795993 = array_index_795988 == array_index_772632 ? add_795992 : sel_795989;
  assign add_795996 = sel_795993 + 8'h01;
  assign sel_795997 = array_index_795988 == array_index_772636 ? add_795996 : sel_795993;
  assign add_796000 = sel_795997 + 8'h01;
  assign sel_796001 = array_index_795988 == array_index_772644 ? add_796000 : sel_795997;
  assign add_796004 = sel_796001 + 8'h01;
  assign sel_796005 = array_index_795988 == array_index_772652 ? add_796004 : sel_796001;
  assign add_796008 = sel_796005 + 8'h01;
  assign sel_796009 = array_index_795988 == array_index_772660 ? add_796008 : sel_796005;
  assign add_796012 = sel_796009 + 8'h01;
  assign sel_796013 = array_index_795988 == array_index_772668 ? add_796012 : sel_796009;
  assign add_796016 = sel_796013 + 8'h01;
  assign sel_796017 = array_index_795988 == array_index_772676 ? add_796016 : sel_796013;
  assign add_796020 = sel_796017 + 8'h01;
  assign sel_796021 = array_index_795988 == array_index_772684 ? add_796020 : sel_796017;
  assign add_796024 = sel_796021 + 8'h01;
  assign sel_796025 = array_index_795988 == array_index_772690 ? add_796024 : sel_796021;
  assign add_796028 = sel_796025 + 8'h01;
  assign sel_796029 = array_index_795988 == array_index_772696 ? add_796028 : sel_796025;
  assign add_796032 = sel_796029 + 8'h01;
  assign sel_796033 = array_index_795988 == array_index_772702 ? add_796032 : sel_796029;
  assign add_796036 = sel_796033 + 8'h01;
  assign sel_796037 = array_index_795988 == array_index_772708 ? add_796036 : sel_796033;
  assign add_796040 = sel_796037 + 8'h01;
  assign sel_796041 = array_index_795988 == array_index_772714 ? add_796040 : sel_796037;
  assign add_796044 = sel_796041 + 8'h01;
  assign sel_796045 = array_index_795988 == array_index_772720 ? add_796044 : sel_796041;
  assign add_796048 = sel_796045 + 8'h01;
  assign sel_796049 = array_index_795988 == array_index_772726 ? add_796048 : sel_796045;
  assign add_796052 = sel_796049 + 8'h01;
  assign sel_796053 = array_index_795988 == array_index_772732 ? add_796052 : sel_796049;
  assign add_796056 = sel_796053 + 8'h01;
  assign sel_796057 = array_index_795988 == array_index_772738 ? add_796056 : sel_796053;
  assign add_796060 = sel_796057 + 8'h01;
  assign sel_796061 = array_index_795988 == array_index_772744 ? add_796060 : sel_796057;
  assign add_796064 = sel_796061 + 8'h01;
  assign sel_796065 = array_index_795988 == array_index_772750 ? add_796064 : sel_796061;
  assign add_796068 = sel_796065 + 8'h01;
  assign sel_796069 = array_index_795988 == array_index_772756 ? add_796068 : sel_796065;
  assign add_796072 = sel_796069 + 8'h01;
  assign sel_796073 = array_index_795988 == array_index_772762 ? add_796072 : sel_796069;
  assign add_796076 = sel_796073 + 8'h01;
  assign sel_796077 = array_index_795988 == array_index_772768 ? add_796076 : sel_796073;
  assign add_796080 = sel_796077 + 8'h01;
  assign sel_796081 = array_index_795988 == array_index_772774 ? add_796080 : sel_796077;
  assign add_796084 = sel_796081 + 8'h01;
  assign sel_796085 = array_index_795988 == array_index_772780 ? add_796084 : sel_796081;
  assign add_796088 = sel_796085 + 8'h01;
  assign sel_796089 = array_index_795988 == array_index_772786 ? add_796088 : sel_796085;
  assign add_796092 = sel_796089 + 8'h01;
  assign sel_796093 = array_index_795988 == array_index_772792 ? add_796092 : sel_796089;
  assign add_796096 = sel_796093 + 8'h01;
  assign sel_796097 = array_index_795988 == array_index_772798 ? add_796096 : sel_796093;
  assign add_796100 = sel_796097 + 8'h01;
  assign sel_796101 = array_index_795988 == array_index_772804 ? add_796100 : sel_796097;
  assign add_796104 = sel_796101 + 8'h01;
  assign sel_796105 = array_index_795988 == array_index_772810 ? add_796104 : sel_796101;
  assign add_796108 = sel_796105 + 8'h01;
  assign sel_796109 = array_index_795988 == array_index_772816 ? add_796108 : sel_796105;
  assign add_796112 = sel_796109 + 8'h01;
  assign sel_796113 = array_index_795988 == array_index_772822 ? add_796112 : sel_796109;
  assign add_796116 = sel_796113 + 8'h01;
  assign sel_796117 = array_index_795988 == array_index_772828 ? add_796116 : sel_796113;
  assign add_796120 = sel_796117 + 8'h01;
  assign sel_796121 = array_index_795988 == array_index_772834 ? add_796120 : sel_796117;
  assign add_796124 = sel_796121 + 8'h01;
  assign sel_796125 = array_index_795988 == array_index_772840 ? add_796124 : sel_796121;
  assign add_796128 = sel_796125 + 8'h01;
  assign sel_796129 = array_index_795988 == array_index_772846 ? add_796128 : sel_796125;
  assign add_796132 = sel_796129 + 8'h01;
  assign sel_796133 = array_index_795988 == array_index_772852 ? add_796132 : sel_796129;
  assign add_796136 = sel_796133 + 8'h01;
  assign sel_796137 = array_index_795988 == array_index_772858 ? add_796136 : sel_796133;
  assign add_796140 = sel_796137 + 8'h01;
  assign sel_796141 = array_index_795988 == array_index_772864 ? add_796140 : sel_796137;
  assign add_796144 = sel_796141 + 8'h01;
  assign sel_796145 = array_index_795988 == array_index_772870 ? add_796144 : sel_796141;
  assign add_796148 = sel_796145 + 8'h01;
  assign sel_796149 = array_index_795988 == array_index_772876 ? add_796148 : sel_796145;
  assign add_796152 = sel_796149 + 8'h01;
  assign sel_796153 = array_index_795988 == array_index_772882 ? add_796152 : sel_796149;
  assign add_796156 = sel_796153 + 8'h01;
  assign sel_796157 = array_index_795988 == array_index_772888 ? add_796156 : sel_796153;
  assign add_796160 = sel_796157 + 8'h01;
  assign sel_796161 = array_index_795988 == array_index_772894 ? add_796160 : sel_796157;
  assign add_796164 = sel_796161 + 8'h01;
  assign sel_796165 = array_index_795988 == array_index_772900 ? add_796164 : sel_796161;
  assign add_796168 = sel_796165 + 8'h01;
  assign sel_796169 = array_index_795988 == array_index_772906 ? add_796168 : sel_796165;
  assign add_796172 = sel_796169 + 8'h01;
  assign sel_796173 = array_index_795988 == array_index_772912 ? add_796172 : sel_796169;
  assign add_796176 = sel_796173 + 8'h01;
  assign sel_796177 = array_index_795988 == array_index_772918 ? add_796176 : sel_796173;
  assign add_796180 = sel_796177 + 8'h01;
  assign sel_796181 = array_index_795988 == array_index_772924 ? add_796180 : sel_796177;
  assign add_796184 = sel_796181 + 8'h01;
  assign sel_796185 = array_index_795988 == array_index_772930 ? add_796184 : sel_796181;
  assign add_796188 = sel_796185 + 8'h01;
  assign sel_796189 = array_index_795988 == array_index_772936 ? add_796188 : sel_796185;
  assign add_796192 = sel_796189 + 8'h01;
  assign sel_796193 = array_index_795988 == array_index_772942 ? add_796192 : sel_796189;
  assign add_796196 = sel_796193 + 8'h01;
  assign sel_796197 = array_index_795988 == array_index_772948 ? add_796196 : sel_796193;
  assign add_796200 = sel_796197 + 8'h01;
  assign sel_796201 = array_index_795988 == array_index_772954 ? add_796200 : sel_796197;
  assign add_796204 = sel_796201 + 8'h01;
  assign sel_796205 = array_index_795988 == array_index_772960 ? add_796204 : sel_796201;
  assign add_796208 = sel_796205 + 8'h01;
  assign sel_796209 = array_index_795988 == array_index_772966 ? add_796208 : sel_796205;
  assign add_796212 = sel_796209 + 8'h01;
  assign sel_796213 = array_index_795988 == array_index_772972 ? add_796212 : sel_796209;
  assign add_796216 = sel_796213 + 8'h01;
  assign sel_796217 = array_index_795988 == array_index_772978 ? add_796216 : sel_796213;
  assign add_796220 = sel_796217 + 8'h01;
  assign sel_796221 = array_index_795988 == array_index_772984 ? add_796220 : sel_796217;
  assign add_796224 = sel_796221 + 8'h01;
  assign sel_796225 = array_index_795988 == array_index_772990 ? add_796224 : sel_796221;
  assign add_796228 = sel_796225 + 8'h01;
  assign sel_796229 = array_index_795988 == array_index_772996 ? add_796228 : sel_796225;
  assign add_796232 = sel_796229 + 8'h01;
  assign sel_796233 = array_index_795988 == array_index_773002 ? add_796232 : sel_796229;
  assign add_796236 = sel_796233 + 8'h01;
  assign sel_796237 = array_index_795988 == array_index_773008 ? add_796236 : sel_796233;
  assign add_796240 = sel_796237 + 8'h01;
  assign sel_796241 = array_index_795988 == array_index_773014 ? add_796240 : sel_796237;
  assign add_796244 = sel_796241 + 8'h01;
  assign sel_796245 = array_index_795988 == array_index_773020 ? add_796244 : sel_796241;
  assign add_796248 = sel_796245 + 8'h01;
  assign sel_796249 = array_index_795988 == array_index_773026 ? add_796248 : sel_796245;
  assign add_796252 = sel_796249 + 8'h01;
  assign sel_796253 = array_index_795988 == array_index_773032 ? add_796252 : sel_796249;
  assign add_796256 = sel_796253 + 8'h01;
  assign sel_796257 = array_index_795988 == array_index_773038 ? add_796256 : sel_796253;
  assign add_796260 = sel_796257 + 8'h01;
  assign sel_796261 = array_index_795988 == array_index_773044 ? add_796260 : sel_796257;
  assign add_796264 = sel_796261 + 8'h01;
  assign sel_796265 = array_index_795988 == array_index_773050 ? add_796264 : sel_796261;
  assign add_796268 = sel_796265 + 8'h01;
  assign sel_796269 = array_index_795988 == array_index_773056 ? add_796268 : sel_796265;
  assign add_796272 = sel_796269 + 8'h01;
  assign sel_796273 = array_index_795988 == array_index_773062 ? add_796272 : sel_796269;
  assign add_796276 = sel_796273 + 8'h01;
  assign sel_796277 = array_index_795988 == array_index_773068 ? add_796276 : sel_796273;
  assign add_796280 = sel_796277 + 8'h01;
  assign sel_796281 = array_index_795988 == array_index_773074 ? add_796280 : sel_796277;
  assign add_796284 = sel_796281 + 8'h01;
  assign sel_796285 = array_index_795988 == array_index_773080 ? add_796284 : sel_796281;
  assign add_796288 = sel_796285 + 8'h01;
  assign sel_796289 = array_index_795988 == array_index_773086 ? add_796288 : sel_796285;
  assign add_796292 = sel_796289 + 8'h01;
  assign sel_796293 = array_index_795988 == array_index_773092 ? add_796292 : sel_796289;
  assign add_796296 = sel_796293 + 8'h01;
  assign sel_796297 = array_index_795988 == array_index_773098 ? add_796296 : sel_796293;
  assign add_796300 = sel_796297 + 8'h01;
  assign sel_796301 = array_index_795988 == array_index_773104 ? add_796300 : sel_796297;
  assign add_796304 = sel_796301 + 8'h01;
  assign sel_796305 = array_index_795988 == array_index_773110 ? add_796304 : sel_796301;
  assign add_796308 = sel_796305 + 8'h01;
  assign sel_796309 = array_index_795988 == array_index_773116 ? add_796308 : sel_796305;
  assign add_796312 = sel_796309 + 8'h01;
  assign sel_796313 = array_index_795988 == array_index_773122 ? add_796312 : sel_796309;
  assign add_796316 = sel_796313 + 8'h01;
  assign sel_796317 = array_index_795988 == array_index_773128 ? add_796316 : sel_796313;
  assign add_796320 = sel_796317 + 8'h01;
  assign sel_796321 = array_index_795988 == array_index_773134 ? add_796320 : sel_796317;
  assign add_796324 = sel_796321 + 8'h01;
  assign sel_796325 = array_index_795988 == array_index_773140 ? add_796324 : sel_796321;
  assign add_796328 = sel_796325 + 8'h01;
  assign sel_796329 = array_index_795988 == array_index_773146 ? add_796328 : sel_796325;
  assign add_796332 = sel_796329 + 8'h01;
  assign sel_796333 = array_index_795988 == array_index_773152 ? add_796332 : sel_796329;
  assign add_796336 = sel_796333 + 8'h01;
  assign sel_796337 = array_index_795988 == array_index_773158 ? add_796336 : sel_796333;
  assign add_796340 = sel_796337 + 8'h01;
  assign sel_796341 = array_index_795988 == array_index_773164 ? add_796340 : sel_796337;
  assign add_796344 = sel_796341 + 8'h01;
  assign sel_796345 = array_index_795988 == array_index_773170 ? add_796344 : sel_796341;
  assign add_796349 = sel_796345 + 8'h01;
  assign array_index_796350 = set1_unflattened[7'h41];
  assign sel_796351 = array_index_795988 == array_index_773176 ? add_796349 : sel_796345;
  assign add_796354 = sel_796351 + 8'h01;
  assign sel_796355 = array_index_796350 == array_index_772632 ? add_796354 : sel_796351;
  assign add_796358 = sel_796355 + 8'h01;
  assign sel_796359 = array_index_796350 == array_index_772636 ? add_796358 : sel_796355;
  assign add_796362 = sel_796359 + 8'h01;
  assign sel_796363 = array_index_796350 == array_index_772644 ? add_796362 : sel_796359;
  assign add_796366 = sel_796363 + 8'h01;
  assign sel_796367 = array_index_796350 == array_index_772652 ? add_796366 : sel_796363;
  assign add_796370 = sel_796367 + 8'h01;
  assign sel_796371 = array_index_796350 == array_index_772660 ? add_796370 : sel_796367;
  assign add_796374 = sel_796371 + 8'h01;
  assign sel_796375 = array_index_796350 == array_index_772668 ? add_796374 : sel_796371;
  assign add_796378 = sel_796375 + 8'h01;
  assign sel_796379 = array_index_796350 == array_index_772676 ? add_796378 : sel_796375;
  assign add_796382 = sel_796379 + 8'h01;
  assign sel_796383 = array_index_796350 == array_index_772684 ? add_796382 : sel_796379;
  assign add_796386 = sel_796383 + 8'h01;
  assign sel_796387 = array_index_796350 == array_index_772690 ? add_796386 : sel_796383;
  assign add_796390 = sel_796387 + 8'h01;
  assign sel_796391 = array_index_796350 == array_index_772696 ? add_796390 : sel_796387;
  assign add_796394 = sel_796391 + 8'h01;
  assign sel_796395 = array_index_796350 == array_index_772702 ? add_796394 : sel_796391;
  assign add_796398 = sel_796395 + 8'h01;
  assign sel_796399 = array_index_796350 == array_index_772708 ? add_796398 : sel_796395;
  assign add_796402 = sel_796399 + 8'h01;
  assign sel_796403 = array_index_796350 == array_index_772714 ? add_796402 : sel_796399;
  assign add_796406 = sel_796403 + 8'h01;
  assign sel_796407 = array_index_796350 == array_index_772720 ? add_796406 : sel_796403;
  assign add_796410 = sel_796407 + 8'h01;
  assign sel_796411 = array_index_796350 == array_index_772726 ? add_796410 : sel_796407;
  assign add_796414 = sel_796411 + 8'h01;
  assign sel_796415 = array_index_796350 == array_index_772732 ? add_796414 : sel_796411;
  assign add_796418 = sel_796415 + 8'h01;
  assign sel_796419 = array_index_796350 == array_index_772738 ? add_796418 : sel_796415;
  assign add_796422 = sel_796419 + 8'h01;
  assign sel_796423 = array_index_796350 == array_index_772744 ? add_796422 : sel_796419;
  assign add_796426 = sel_796423 + 8'h01;
  assign sel_796427 = array_index_796350 == array_index_772750 ? add_796426 : sel_796423;
  assign add_796430 = sel_796427 + 8'h01;
  assign sel_796431 = array_index_796350 == array_index_772756 ? add_796430 : sel_796427;
  assign add_796434 = sel_796431 + 8'h01;
  assign sel_796435 = array_index_796350 == array_index_772762 ? add_796434 : sel_796431;
  assign add_796438 = sel_796435 + 8'h01;
  assign sel_796439 = array_index_796350 == array_index_772768 ? add_796438 : sel_796435;
  assign add_796442 = sel_796439 + 8'h01;
  assign sel_796443 = array_index_796350 == array_index_772774 ? add_796442 : sel_796439;
  assign add_796446 = sel_796443 + 8'h01;
  assign sel_796447 = array_index_796350 == array_index_772780 ? add_796446 : sel_796443;
  assign add_796450 = sel_796447 + 8'h01;
  assign sel_796451 = array_index_796350 == array_index_772786 ? add_796450 : sel_796447;
  assign add_796454 = sel_796451 + 8'h01;
  assign sel_796455 = array_index_796350 == array_index_772792 ? add_796454 : sel_796451;
  assign add_796458 = sel_796455 + 8'h01;
  assign sel_796459 = array_index_796350 == array_index_772798 ? add_796458 : sel_796455;
  assign add_796462 = sel_796459 + 8'h01;
  assign sel_796463 = array_index_796350 == array_index_772804 ? add_796462 : sel_796459;
  assign add_796466 = sel_796463 + 8'h01;
  assign sel_796467 = array_index_796350 == array_index_772810 ? add_796466 : sel_796463;
  assign add_796470 = sel_796467 + 8'h01;
  assign sel_796471 = array_index_796350 == array_index_772816 ? add_796470 : sel_796467;
  assign add_796474 = sel_796471 + 8'h01;
  assign sel_796475 = array_index_796350 == array_index_772822 ? add_796474 : sel_796471;
  assign add_796478 = sel_796475 + 8'h01;
  assign sel_796479 = array_index_796350 == array_index_772828 ? add_796478 : sel_796475;
  assign add_796482 = sel_796479 + 8'h01;
  assign sel_796483 = array_index_796350 == array_index_772834 ? add_796482 : sel_796479;
  assign add_796486 = sel_796483 + 8'h01;
  assign sel_796487 = array_index_796350 == array_index_772840 ? add_796486 : sel_796483;
  assign add_796490 = sel_796487 + 8'h01;
  assign sel_796491 = array_index_796350 == array_index_772846 ? add_796490 : sel_796487;
  assign add_796494 = sel_796491 + 8'h01;
  assign sel_796495 = array_index_796350 == array_index_772852 ? add_796494 : sel_796491;
  assign add_796498 = sel_796495 + 8'h01;
  assign sel_796499 = array_index_796350 == array_index_772858 ? add_796498 : sel_796495;
  assign add_796502 = sel_796499 + 8'h01;
  assign sel_796503 = array_index_796350 == array_index_772864 ? add_796502 : sel_796499;
  assign add_796506 = sel_796503 + 8'h01;
  assign sel_796507 = array_index_796350 == array_index_772870 ? add_796506 : sel_796503;
  assign add_796510 = sel_796507 + 8'h01;
  assign sel_796511 = array_index_796350 == array_index_772876 ? add_796510 : sel_796507;
  assign add_796514 = sel_796511 + 8'h01;
  assign sel_796515 = array_index_796350 == array_index_772882 ? add_796514 : sel_796511;
  assign add_796518 = sel_796515 + 8'h01;
  assign sel_796519 = array_index_796350 == array_index_772888 ? add_796518 : sel_796515;
  assign add_796522 = sel_796519 + 8'h01;
  assign sel_796523 = array_index_796350 == array_index_772894 ? add_796522 : sel_796519;
  assign add_796526 = sel_796523 + 8'h01;
  assign sel_796527 = array_index_796350 == array_index_772900 ? add_796526 : sel_796523;
  assign add_796530 = sel_796527 + 8'h01;
  assign sel_796531 = array_index_796350 == array_index_772906 ? add_796530 : sel_796527;
  assign add_796534 = sel_796531 + 8'h01;
  assign sel_796535 = array_index_796350 == array_index_772912 ? add_796534 : sel_796531;
  assign add_796538 = sel_796535 + 8'h01;
  assign sel_796539 = array_index_796350 == array_index_772918 ? add_796538 : sel_796535;
  assign add_796542 = sel_796539 + 8'h01;
  assign sel_796543 = array_index_796350 == array_index_772924 ? add_796542 : sel_796539;
  assign add_796546 = sel_796543 + 8'h01;
  assign sel_796547 = array_index_796350 == array_index_772930 ? add_796546 : sel_796543;
  assign add_796550 = sel_796547 + 8'h01;
  assign sel_796551 = array_index_796350 == array_index_772936 ? add_796550 : sel_796547;
  assign add_796554 = sel_796551 + 8'h01;
  assign sel_796555 = array_index_796350 == array_index_772942 ? add_796554 : sel_796551;
  assign add_796558 = sel_796555 + 8'h01;
  assign sel_796559 = array_index_796350 == array_index_772948 ? add_796558 : sel_796555;
  assign add_796562 = sel_796559 + 8'h01;
  assign sel_796563 = array_index_796350 == array_index_772954 ? add_796562 : sel_796559;
  assign add_796566 = sel_796563 + 8'h01;
  assign sel_796567 = array_index_796350 == array_index_772960 ? add_796566 : sel_796563;
  assign add_796570 = sel_796567 + 8'h01;
  assign sel_796571 = array_index_796350 == array_index_772966 ? add_796570 : sel_796567;
  assign add_796574 = sel_796571 + 8'h01;
  assign sel_796575 = array_index_796350 == array_index_772972 ? add_796574 : sel_796571;
  assign add_796578 = sel_796575 + 8'h01;
  assign sel_796579 = array_index_796350 == array_index_772978 ? add_796578 : sel_796575;
  assign add_796582 = sel_796579 + 8'h01;
  assign sel_796583 = array_index_796350 == array_index_772984 ? add_796582 : sel_796579;
  assign add_796586 = sel_796583 + 8'h01;
  assign sel_796587 = array_index_796350 == array_index_772990 ? add_796586 : sel_796583;
  assign add_796590 = sel_796587 + 8'h01;
  assign sel_796591 = array_index_796350 == array_index_772996 ? add_796590 : sel_796587;
  assign add_796594 = sel_796591 + 8'h01;
  assign sel_796595 = array_index_796350 == array_index_773002 ? add_796594 : sel_796591;
  assign add_796598 = sel_796595 + 8'h01;
  assign sel_796599 = array_index_796350 == array_index_773008 ? add_796598 : sel_796595;
  assign add_796602 = sel_796599 + 8'h01;
  assign sel_796603 = array_index_796350 == array_index_773014 ? add_796602 : sel_796599;
  assign add_796606 = sel_796603 + 8'h01;
  assign sel_796607 = array_index_796350 == array_index_773020 ? add_796606 : sel_796603;
  assign add_796610 = sel_796607 + 8'h01;
  assign sel_796611 = array_index_796350 == array_index_773026 ? add_796610 : sel_796607;
  assign add_796614 = sel_796611 + 8'h01;
  assign sel_796615 = array_index_796350 == array_index_773032 ? add_796614 : sel_796611;
  assign add_796618 = sel_796615 + 8'h01;
  assign sel_796619 = array_index_796350 == array_index_773038 ? add_796618 : sel_796615;
  assign add_796622 = sel_796619 + 8'h01;
  assign sel_796623 = array_index_796350 == array_index_773044 ? add_796622 : sel_796619;
  assign add_796626 = sel_796623 + 8'h01;
  assign sel_796627 = array_index_796350 == array_index_773050 ? add_796626 : sel_796623;
  assign add_796630 = sel_796627 + 8'h01;
  assign sel_796631 = array_index_796350 == array_index_773056 ? add_796630 : sel_796627;
  assign add_796634 = sel_796631 + 8'h01;
  assign sel_796635 = array_index_796350 == array_index_773062 ? add_796634 : sel_796631;
  assign add_796638 = sel_796635 + 8'h01;
  assign sel_796639 = array_index_796350 == array_index_773068 ? add_796638 : sel_796635;
  assign add_796642 = sel_796639 + 8'h01;
  assign sel_796643 = array_index_796350 == array_index_773074 ? add_796642 : sel_796639;
  assign add_796646 = sel_796643 + 8'h01;
  assign sel_796647 = array_index_796350 == array_index_773080 ? add_796646 : sel_796643;
  assign add_796650 = sel_796647 + 8'h01;
  assign sel_796651 = array_index_796350 == array_index_773086 ? add_796650 : sel_796647;
  assign add_796654 = sel_796651 + 8'h01;
  assign sel_796655 = array_index_796350 == array_index_773092 ? add_796654 : sel_796651;
  assign add_796658 = sel_796655 + 8'h01;
  assign sel_796659 = array_index_796350 == array_index_773098 ? add_796658 : sel_796655;
  assign add_796662 = sel_796659 + 8'h01;
  assign sel_796663 = array_index_796350 == array_index_773104 ? add_796662 : sel_796659;
  assign add_796666 = sel_796663 + 8'h01;
  assign sel_796667 = array_index_796350 == array_index_773110 ? add_796666 : sel_796663;
  assign add_796670 = sel_796667 + 8'h01;
  assign sel_796671 = array_index_796350 == array_index_773116 ? add_796670 : sel_796667;
  assign add_796674 = sel_796671 + 8'h01;
  assign sel_796675 = array_index_796350 == array_index_773122 ? add_796674 : sel_796671;
  assign add_796678 = sel_796675 + 8'h01;
  assign sel_796679 = array_index_796350 == array_index_773128 ? add_796678 : sel_796675;
  assign add_796682 = sel_796679 + 8'h01;
  assign sel_796683 = array_index_796350 == array_index_773134 ? add_796682 : sel_796679;
  assign add_796686 = sel_796683 + 8'h01;
  assign sel_796687 = array_index_796350 == array_index_773140 ? add_796686 : sel_796683;
  assign add_796690 = sel_796687 + 8'h01;
  assign sel_796691 = array_index_796350 == array_index_773146 ? add_796690 : sel_796687;
  assign add_796694 = sel_796691 + 8'h01;
  assign sel_796695 = array_index_796350 == array_index_773152 ? add_796694 : sel_796691;
  assign add_796698 = sel_796695 + 8'h01;
  assign sel_796699 = array_index_796350 == array_index_773158 ? add_796698 : sel_796695;
  assign add_796702 = sel_796699 + 8'h01;
  assign sel_796703 = array_index_796350 == array_index_773164 ? add_796702 : sel_796699;
  assign add_796706 = sel_796703 + 8'h01;
  assign sel_796707 = array_index_796350 == array_index_773170 ? add_796706 : sel_796703;
  assign add_796711 = sel_796707 + 8'h01;
  assign array_index_796712 = set1_unflattened[7'h42];
  assign sel_796713 = array_index_796350 == array_index_773176 ? add_796711 : sel_796707;
  assign add_796716 = sel_796713 + 8'h01;
  assign sel_796717 = array_index_796712 == array_index_772632 ? add_796716 : sel_796713;
  assign add_796720 = sel_796717 + 8'h01;
  assign sel_796721 = array_index_796712 == array_index_772636 ? add_796720 : sel_796717;
  assign add_796724 = sel_796721 + 8'h01;
  assign sel_796725 = array_index_796712 == array_index_772644 ? add_796724 : sel_796721;
  assign add_796728 = sel_796725 + 8'h01;
  assign sel_796729 = array_index_796712 == array_index_772652 ? add_796728 : sel_796725;
  assign add_796732 = sel_796729 + 8'h01;
  assign sel_796733 = array_index_796712 == array_index_772660 ? add_796732 : sel_796729;
  assign add_796736 = sel_796733 + 8'h01;
  assign sel_796737 = array_index_796712 == array_index_772668 ? add_796736 : sel_796733;
  assign add_796740 = sel_796737 + 8'h01;
  assign sel_796741 = array_index_796712 == array_index_772676 ? add_796740 : sel_796737;
  assign add_796744 = sel_796741 + 8'h01;
  assign sel_796745 = array_index_796712 == array_index_772684 ? add_796744 : sel_796741;
  assign add_796748 = sel_796745 + 8'h01;
  assign sel_796749 = array_index_796712 == array_index_772690 ? add_796748 : sel_796745;
  assign add_796752 = sel_796749 + 8'h01;
  assign sel_796753 = array_index_796712 == array_index_772696 ? add_796752 : sel_796749;
  assign add_796756 = sel_796753 + 8'h01;
  assign sel_796757 = array_index_796712 == array_index_772702 ? add_796756 : sel_796753;
  assign add_796760 = sel_796757 + 8'h01;
  assign sel_796761 = array_index_796712 == array_index_772708 ? add_796760 : sel_796757;
  assign add_796764 = sel_796761 + 8'h01;
  assign sel_796765 = array_index_796712 == array_index_772714 ? add_796764 : sel_796761;
  assign add_796768 = sel_796765 + 8'h01;
  assign sel_796769 = array_index_796712 == array_index_772720 ? add_796768 : sel_796765;
  assign add_796772 = sel_796769 + 8'h01;
  assign sel_796773 = array_index_796712 == array_index_772726 ? add_796772 : sel_796769;
  assign add_796776 = sel_796773 + 8'h01;
  assign sel_796777 = array_index_796712 == array_index_772732 ? add_796776 : sel_796773;
  assign add_796780 = sel_796777 + 8'h01;
  assign sel_796781 = array_index_796712 == array_index_772738 ? add_796780 : sel_796777;
  assign add_796784 = sel_796781 + 8'h01;
  assign sel_796785 = array_index_796712 == array_index_772744 ? add_796784 : sel_796781;
  assign add_796788 = sel_796785 + 8'h01;
  assign sel_796789 = array_index_796712 == array_index_772750 ? add_796788 : sel_796785;
  assign add_796792 = sel_796789 + 8'h01;
  assign sel_796793 = array_index_796712 == array_index_772756 ? add_796792 : sel_796789;
  assign add_796796 = sel_796793 + 8'h01;
  assign sel_796797 = array_index_796712 == array_index_772762 ? add_796796 : sel_796793;
  assign add_796800 = sel_796797 + 8'h01;
  assign sel_796801 = array_index_796712 == array_index_772768 ? add_796800 : sel_796797;
  assign add_796804 = sel_796801 + 8'h01;
  assign sel_796805 = array_index_796712 == array_index_772774 ? add_796804 : sel_796801;
  assign add_796808 = sel_796805 + 8'h01;
  assign sel_796809 = array_index_796712 == array_index_772780 ? add_796808 : sel_796805;
  assign add_796812 = sel_796809 + 8'h01;
  assign sel_796813 = array_index_796712 == array_index_772786 ? add_796812 : sel_796809;
  assign add_796816 = sel_796813 + 8'h01;
  assign sel_796817 = array_index_796712 == array_index_772792 ? add_796816 : sel_796813;
  assign add_796820 = sel_796817 + 8'h01;
  assign sel_796821 = array_index_796712 == array_index_772798 ? add_796820 : sel_796817;
  assign add_796824 = sel_796821 + 8'h01;
  assign sel_796825 = array_index_796712 == array_index_772804 ? add_796824 : sel_796821;
  assign add_796828 = sel_796825 + 8'h01;
  assign sel_796829 = array_index_796712 == array_index_772810 ? add_796828 : sel_796825;
  assign add_796832 = sel_796829 + 8'h01;
  assign sel_796833 = array_index_796712 == array_index_772816 ? add_796832 : sel_796829;
  assign add_796836 = sel_796833 + 8'h01;
  assign sel_796837 = array_index_796712 == array_index_772822 ? add_796836 : sel_796833;
  assign add_796840 = sel_796837 + 8'h01;
  assign sel_796841 = array_index_796712 == array_index_772828 ? add_796840 : sel_796837;
  assign add_796844 = sel_796841 + 8'h01;
  assign sel_796845 = array_index_796712 == array_index_772834 ? add_796844 : sel_796841;
  assign add_796848 = sel_796845 + 8'h01;
  assign sel_796849 = array_index_796712 == array_index_772840 ? add_796848 : sel_796845;
  assign add_796852 = sel_796849 + 8'h01;
  assign sel_796853 = array_index_796712 == array_index_772846 ? add_796852 : sel_796849;
  assign add_796856 = sel_796853 + 8'h01;
  assign sel_796857 = array_index_796712 == array_index_772852 ? add_796856 : sel_796853;
  assign add_796860 = sel_796857 + 8'h01;
  assign sel_796861 = array_index_796712 == array_index_772858 ? add_796860 : sel_796857;
  assign add_796864 = sel_796861 + 8'h01;
  assign sel_796865 = array_index_796712 == array_index_772864 ? add_796864 : sel_796861;
  assign add_796868 = sel_796865 + 8'h01;
  assign sel_796869 = array_index_796712 == array_index_772870 ? add_796868 : sel_796865;
  assign add_796872 = sel_796869 + 8'h01;
  assign sel_796873 = array_index_796712 == array_index_772876 ? add_796872 : sel_796869;
  assign add_796876 = sel_796873 + 8'h01;
  assign sel_796877 = array_index_796712 == array_index_772882 ? add_796876 : sel_796873;
  assign add_796880 = sel_796877 + 8'h01;
  assign sel_796881 = array_index_796712 == array_index_772888 ? add_796880 : sel_796877;
  assign add_796884 = sel_796881 + 8'h01;
  assign sel_796885 = array_index_796712 == array_index_772894 ? add_796884 : sel_796881;
  assign add_796888 = sel_796885 + 8'h01;
  assign sel_796889 = array_index_796712 == array_index_772900 ? add_796888 : sel_796885;
  assign add_796892 = sel_796889 + 8'h01;
  assign sel_796893 = array_index_796712 == array_index_772906 ? add_796892 : sel_796889;
  assign add_796896 = sel_796893 + 8'h01;
  assign sel_796897 = array_index_796712 == array_index_772912 ? add_796896 : sel_796893;
  assign add_796900 = sel_796897 + 8'h01;
  assign sel_796901 = array_index_796712 == array_index_772918 ? add_796900 : sel_796897;
  assign add_796904 = sel_796901 + 8'h01;
  assign sel_796905 = array_index_796712 == array_index_772924 ? add_796904 : sel_796901;
  assign add_796908 = sel_796905 + 8'h01;
  assign sel_796909 = array_index_796712 == array_index_772930 ? add_796908 : sel_796905;
  assign add_796912 = sel_796909 + 8'h01;
  assign sel_796913 = array_index_796712 == array_index_772936 ? add_796912 : sel_796909;
  assign add_796916 = sel_796913 + 8'h01;
  assign sel_796917 = array_index_796712 == array_index_772942 ? add_796916 : sel_796913;
  assign add_796920 = sel_796917 + 8'h01;
  assign sel_796921 = array_index_796712 == array_index_772948 ? add_796920 : sel_796917;
  assign add_796924 = sel_796921 + 8'h01;
  assign sel_796925 = array_index_796712 == array_index_772954 ? add_796924 : sel_796921;
  assign add_796928 = sel_796925 + 8'h01;
  assign sel_796929 = array_index_796712 == array_index_772960 ? add_796928 : sel_796925;
  assign add_796932 = sel_796929 + 8'h01;
  assign sel_796933 = array_index_796712 == array_index_772966 ? add_796932 : sel_796929;
  assign add_796936 = sel_796933 + 8'h01;
  assign sel_796937 = array_index_796712 == array_index_772972 ? add_796936 : sel_796933;
  assign add_796940 = sel_796937 + 8'h01;
  assign sel_796941 = array_index_796712 == array_index_772978 ? add_796940 : sel_796937;
  assign add_796944 = sel_796941 + 8'h01;
  assign sel_796945 = array_index_796712 == array_index_772984 ? add_796944 : sel_796941;
  assign add_796948 = sel_796945 + 8'h01;
  assign sel_796949 = array_index_796712 == array_index_772990 ? add_796948 : sel_796945;
  assign add_796952 = sel_796949 + 8'h01;
  assign sel_796953 = array_index_796712 == array_index_772996 ? add_796952 : sel_796949;
  assign add_796956 = sel_796953 + 8'h01;
  assign sel_796957 = array_index_796712 == array_index_773002 ? add_796956 : sel_796953;
  assign add_796960 = sel_796957 + 8'h01;
  assign sel_796961 = array_index_796712 == array_index_773008 ? add_796960 : sel_796957;
  assign add_796964 = sel_796961 + 8'h01;
  assign sel_796965 = array_index_796712 == array_index_773014 ? add_796964 : sel_796961;
  assign add_796968 = sel_796965 + 8'h01;
  assign sel_796969 = array_index_796712 == array_index_773020 ? add_796968 : sel_796965;
  assign add_796972 = sel_796969 + 8'h01;
  assign sel_796973 = array_index_796712 == array_index_773026 ? add_796972 : sel_796969;
  assign add_796976 = sel_796973 + 8'h01;
  assign sel_796977 = array_index_796712 == array_index_773032 ? add_796976 : sel_796973;
  assign add_796980 = sel_796977 + 8'h01;
  assign sel_796981 = array_index_796712 == array_index_773038 ? add_796980 : sel_796977;
  assign add_796984 = sel_796981 + 8'h01;
  assign sel_796985 = array_index_796712 == array_index_773044 ? add_796984 : sel_796981;
  assign add_796988 = sel_796985 + 8'h01;
  assign sel_796989 = array_index_796712 == array_index_773050 ? add_796988 : sel_796985;
  assign add_796992 = sel_796989 + 8'h01;
  assign sel_796993 = array_index_796712 == array_index_773056 ? add_796992 : sel_796989;
  assign add_796996 = sel_796993 + 8'h01;
  assign sel_796997 = array_index_796712 == array_index_773062 ? add_796996 : sel_796993;
  assign add_797000 = sel_796997 + 8'h01;
  assign sel_797001 = array_index_796712 == array_index_773068 ? add_797000 : sel_796997;
  assign add_797004 = sel_797001 + 8'h01;
  assign sel_797005 = array_index_796712 == array_index_773074 ? add_797004 : sel_797001;
  assign add_797008 = sel_797005 + 8'h01;
  assign sel_797009 = array_index_796712 == array_index_773080 ? add_797008 : sel_797005;
  assign add_797012 = sel_797009 + 8'h01;
  assign sel_797013 = array_index_796712 == array_index_773086 ? add_797012 : sel_797009;
  assign add_797016 = sel_797013 + 8'h01;
  assign sel_797017 = array_index_796712 == array_index_773092 ? add_797016 : sel_797013;
  assign add_797020 = sel_797017 + 8'h01;
  assign sel_797021 = array_index_796712 == array_index_773098 ? add_797020 : sel_797017;
  assign add_797024 = sel_797021 + 8'h01;
  assign sel_797025 = array_index_796712 == array_index_773104 ? add_797024 : sel_797021;
  assign add_797028 = sel_797025 + 8'h01;
  assign sel_797029 = array_index_796712 == array_index_773110 ? add_797028 : sel_797025;
  assign add_797032 = sel_797029 + 8'h01;
  assign sel_797033 = array_index_796712 == array_index_773116 ? add_797032 : sel_797029;
  assign add_797036 = sel_797033 + 8'h01;
  assign sel_797037 = array_index_796712 == array_index_773122 ? add_797036 : sel_797033;
  assign add_797040 = sel_797037 + 8'h01;
  assign sel_797041 = array_index_796712 == array_index_773128 ? add_797040 : sel_797037;
  assign add_797044 = sel_797041 + 8'h01;
  assign sel_797045 = array_index_796712 == array_index_773134 ? add_797044 : sel_797041;
  assign add_797048 = sel_797045 + 8'h01;
  assign sel_797049 = array_index_796712 == array_index_773140 ? add_797048 : sel_797045;
  assign add_797052 = sel_797049 + 8'h01;
  assign sel_797053 = array_index_796712 == array_index_773146 ? add_797052 : sel_797049;
  assign add_797056 = sel_797053 + 8'h01;
  assign sel_797057 = array_index_796712 == array_index_773152 ? add_797056 : sel_797053;
  assign add_797060 = sel_797057 + 8'h01;
  assign sel_797061 = array_index_796712 == array_index_773158 ? add_797060 : sel_797057;
  assign add_797064 = sel_797061 + 8'h01;
  assign sel_797065 = array_index_796712 == array_index_773164 ? add_797064 : sel_797061;
  assign add_797068 = sel_797065 + 8'h01;
  assign sel_797069 = array_index_796712 == array_index_773170 ? add_797068 : sel_797065;
  assign add_797073 = sel_797069 + 8'h01;
  assign array_index_797074 = set1_unflattened[7'h43];
  assign sel_797075 = array_index_796712 == array_index_773176 ? add_797073 : sel_797069;
  assign add_797078 = sel_797075 + 8'h01;
  assign sel_797079 = array_index_797074 == array_index_772632 ? add_797078 : sel_797075;
  assign add_797082 = sel_797079 + 8'h01;
  assign sel_797083 = array_index_797074 == array_index_772636 ? add_797082 : sel_797079;
  assign add_797086 = sel_797083 + 8'h01;
  assign sel_797087 = array_index_797074 == array_index_772644 ? add_797086 : sel_797083;
  assign add_797090 = sel_797087 + 8'h01;
  assign sel_797091 = array_index_797074 == array_index_772652 ? add_797090 : sel_797087;
  assign add_797094 = sel_797091 + 8'h01;
  assign sel_797095 = array_index_797074 == array_index_772660 ? add_797094 : sel_797091;
  assign add_797098 = sel_797095 + 8'h01;
  assign sel_797099 = array_index_797074 == array_index_772668 ? add_797098 : sel_797095;
  assign add_797102 = sel_797099 + 8'h01;
  assign sel_797103 = array_index_797074 == array_index_772676 ? add_797102 : sel_797099;
  assign add_797106 = sel_797103 + 8'h01;
  assign sel_797107 = array_index_797074 == array_index_772684 ? add_797106 : sel_797103;
  assign add_797110 = sel_797107 + 8'h01;
  assign sel_797111 = array_index_797074 == array_index_772690 ? add_797110 : sel_797107;
  assign add_797114 = sel_797111 + 8'h01;
  assign sel_797115 = array_index_797074 == array_index_772696 ? add_797114 : sel_797111;
  assign add_797118 = sel_797115 + 8'h01;
  assign sel_797119 = array_index_797074 == array_index_772702 ? add_797118 : sel_797115;
  assign add_797122 = sel_797119 + 8'h01;
  assign sel_797123 = array_index_797074 == array_index_772708 ? add_797122 : sel_797119;
  assign add_797126 = sel_797123 + 8'h01;
  assign sel_797127 = array_index_797074 == array_index_772714 ? add_797126 : sel_797123;
  assign add_797130 = sel_797127 + 8'h01;
  assign sel_797131 = array_index_797074 == array_index_772720 ? add_797130 : sel_797127;
  assign add_797134 = sel_797131 + 8'h01;
  assign sel_797135 = array_index_797074 == array_index_772726 ? add_797134 : sel_797131;
  assign add_797138 = sel_797135 + 8'h01;
  assign sel_797139 = array_index_797074 == array_index_772732 ? add_797138 : sel_797135;
  assign add_797142 = sel_797139 + 8'h01;
  assign sel_797143 = array_index_797074 == array_index_772738 ? add_797142 : sel_797139;
  assign add_797146 = sel_797143 + 8'h01;
  assign sel_797147 = array_index_797074 == array_index_772744 ? add_797146 : sel_797143;
  assign add_797150 = sel_797147 + 8'h01;
  assign sel_797151 = array_index_797074 == array_index_772750 ? add_797150 : sel_797147;
  assign add_797154 = sel_797151 + 8'h01;
  assign sel_797155 = array_index_797074 == array_index_772756 ? add_797154 : sel_797151;
  assign add_797158 = sel_797155 + 8'h01;
  assign sel_797159 = array_index_797074 == array_index_772762 ? add_797158 : sel_797155;
  assign add_797162 = sel_797159 + 8'h01;
  assign sel_797163 = array_index_797074 == array_index_772768 ? add_797162 : sel_797159;
  assign add_797166 = sel_797163 + 8'h01;
  assign sel_797167 = array_index_797074 == array_index_772774 ? add_797166 : sel_797163;
  assign add_797170 = sel_797167 + 8'h01;
  assign sel_797171 = array_index_797074 == array_index_772780 ? add_797170 : sel_797167;
  assign add_797174 = sel_797171 + 8'h01;
  assign sel_797175 = array_index_797074 == array_index_772786 ? add_797174 : sel_797171;
  assign add_797178 = sel_797175 + 8'h01;
  assign sel_797179 = array_index_797074 == array_index_772792 ? add_797178 : sel_797175;
  assign add_797182 = sel_797179 + 8'h01;
  assign sel_797183 = array_index_797074 == array_index_772798 ? add_797182 : sel_797179;
  assign add_797186 = sel_797183 + 8'h01;
  assign sel_797187 = array_index_797074 == array_index_772804 ? add_797186 : sel_797183;
  assign add_797190 = sel_797187 + 8'h01;
  assign sel_797191 = array_index_797074 == array_index_772810 ? add_797190 : sel_797187;
  assign add_797194 = sel_797191 + 8'h01;
  assign sel_797195 = array_index_797074 == array_index_772816 ? add_797194 : sel_797191;
  assign add_797198 = sel_797195 + 8'h01;
  assign sel_797199 = array_index_797074 == array_index_772822 ? add_797198 : sel_797195;
  assign add_797202 = sel_797199 + 8'h01;
  assign sel_797203 = array_index_797074 == array_index_772828 ? add_797202 : sel_797199;
  assign add_797206 = sel_797203 + 8'h01;
  assign sel_797207 = array_index_797074 == array_index_772834 ? add_797206 : sel_797203;
  assign add_797210 = sel_797207 + 8'h01;
  assign sel_797211 = array_index_797074 == array_index_772840 ? add_797210 : sel_797207;
  assign add_797214 = sel_797211 + 8'h01;
  assign sel_797215 = array_index_797074 == array_index_772846 ? add_797214 : sel_797211;
  assign add_797218 = sel_797215 + 8'h01;
  assign sel_797219 = array_index_797074 == array_index_772852 ? add_797218 : sel_797215;
  assign add_797222 = sel_797219 + 8'h01;
  assign sel_797223 = array_index_797074 == array_index_772858 ? add_797222 : sel_797219;
  assign add_797226 = sel_797223 + 8'h01;
  assign sel_797227 = array_index_797074 == array_index_772864 ? add_797226 : sel_797223;
  assign add_797230 = sel_797227 + 8'h01;
  assign sel_797231 = array_index_797074 == array_index_772870 ? add_797230 : sel_797227;
  assign add_797234 = sel_797231 + 8'h01;
  assign sel_797235 = array_index_797074 == array_index_772876 ? add_797234 : sel_797231;
  assign add_797238 = sel_797235 + 8'h01;
  assign sel_797239 = array_index_797074 == array_index_772882 ? add_797238 : sel_797235;
  assign add_797242 = sel_797239 + 8'h01;
  assign sel_797243 = array_index_797074 == array_index_772888 ? add_797242 : sel_797239;
  assign add_797246 = sel_797243 + 8'h01;
  assign sel_797247 = array_index_797074 == array_index_772894 ? add_797246 : sel_797243;
  assign add_797250 = sel_797247 + 8'h01;
  assign sel_797251 = array_index_797074 == array_index_772900 ? add_797250 : sel_797247;
  assign add_797254 = sel_797251 + 8'h01;
  assign sel_797255 = array_index_797074 == array_index_772906 ? add_797254 : sel_797251;
  assign add_797258 = sel_797255 + 8'h01;
  assign sel_797259 = array_index_797074 == array_index_772912 ? add_797258 : sel_797255;
  assign add_797262 = sel_797259 + 8'h01;
  assign sel_797263 = array_index_797074 == array_index_772918 ? add_797262 : sel_797259;
  assign add_797266 = sel_797263 + 8'h01;
  assign sel_797267 = array_index_797074 == array_index_772924 ? add_797266 : sel_797263;
  assign add_797270 = sel_797267 + 8'h01;
  assign sel_797271 = array_index_797074 == array_index_772930 ? add_797270 : sel_797267;
  assign add_797274 = sel_797271 + 8'h01;
  assign sel_797275 = array_index_797074 == array_index_772936 ? add_797274 : sel_797271;
  assign add_797278 = sel_797275 + 8'h01;
  assign sel_797279 = array_index_797074 == array_index_772942 ? add_797278 : sel_797275;
  assign add_797282 = sel_797279 + 8'h01;
  assign sel_797283 = array_index_797074 == array_index_772948 ? add_797282 : sel_797279;
  assign add_797286 = sel_797283 + 8'h01;
  assign sel_797287 = array_index_797074 == array_index_772954 ? add_797286 : sel_797283;
  assign add_797290 = sel_797287 + 8'h01;
  assign sel_797291 = array_index_797074 == array_index_772960 ? add_797290 : sel_797287;
  assign add_797294 = sel_797291 + 8'h01;
  assign sel_797295 = array_index_797074 == array_index_772966 ? add_797294 : sel_797291;
  assign add_797298 = sel_797295 + 8'h01;
  assign sel_797299 = array_index_797074 == array_index_772972 ? add_797298 : sel_797295;
  assign add_797302 = sel_797299 + 8'h01;
  assign sel_797303 = array_index_797074 == array_index_772978 ? add_797302 : sel_797299;
  assign add_797306 = sel_797303 + 8'h01;
  assign sel_797307 = array_index_797074 == array_index_772984 ? add_797306 : sel_797303;
  assign add_797310 = sel_797307 + 8'h01;
  assign sel_797311 = array_index_797074 == array_index_772990 ? add_797310 : sel_797307;
  assign add_797314 = sel_797311 + 8'h01;
  assign sel_797315 = array_index_797074 == array_index_772996 ? add_797314 : sel_797311;
  assign add_797318 = sel_797315 + 8'h01;
  assign sel_797319 = array_index_797074 == array_index_773002 ? add_797318 : sel_797315;
  assign add_797322 = sel_797319 + 8'h01;
  assign sel_797323 = array_index_797074 == array_index_773008 ? add_797322 : sel_797319;
  assign add_797326 = sel_797323 + 8'h01;
  assign sel_797327 = array_index_797074 == array_index_773014 ? add_797326 : sel_797323;
  assign add_797330 = sel_797327 + 8'h01;
  assign sel_797331 = array_index_797074 == array_index_773020 ? add_797330 : sel_797327;
  assign add_797334 = sel_797331 + 8'h01;
  assign sel_797335 = array_index_797074 == array_index_773026 ? add_797334 : sel_797331;
  assign add_797338 = sel_797335 + 8'h01;
  assign sel_797339 = array_index_797074 == array_index_773032 ? add_797338 : sel_797335;
  assign add_797342 = sel_797339 + 8'h01;
  assign sel_797343 = array_index_797074 == array_index_773038 ? add_797342 : sel_797339;
  assign add_797346 = sel_797343 + 8'h01;
  assign sel_797347 = array_index_797074 == array_index_773044 ? add_797346 : sel_797343;
  assign add_797350 = sel_797347 + 8'h01;
  assign sel_797351 = array_index_797074 == array_index_773050 ? add_797350 : sel_797347;
  assign add_797354 = sel_797351 + 8'h01;
  assign sel_797355 = array_index_797074 == array_index_773056 ? add_797354 : sel_797351;
  assign add_797358 = sel_797355 + 8'h01;
  assign sel_797359 = array_index_797074 == array_index_773062 ? add_797358 : sel_797355;
  assign add_797362 = sel_797359 + 8'h01;
  assign sel_797363 = array_index_797074 == array_index_773068 ? add_797362 : sel_797359;
  assign add_797366 = sel_797363 + 8'h01;
  assign sel_797367 = array_index_797074 == array_index_773074 ? add_797366 : sel_797363;
  assign add_797370 = sel_797367 + 8'h01;
  assign sel_797371 = array_index_797074 == array_index_773080 ? add_797370 : sel_797367;
  assign add_797374 = sel_797371 + 8'h01;
  assign sel_797375 = array_index_797074 == array_index_773086 ? add_797374 : sel_797371;
  assign add_797378 = sel_797375 + 8'h01;
  assign sel_797379 = array_index_797074 == array_index_773092 ? add_797378 : sel_797375;
  assign add_797382 = sel_797379 + 8'h01;
  assign sel_797383 = array_index_797074 == array_index_773098 ? add_797382 : sel_797379;
  assign add_797386 = sel_797383 + 8'h01;
  assign sel_797387 = array_index_797074 == array_index_773104 ? add_797386 : sel_797383;
  assign add_797390 = sel_797387 + 8'h01;
  assign sel_797391 = array_index_797074 == array_index_773110 ? add_797390 : sel_797387;
  assign add_797394 = sel_797391 + 8'h01;
  assign sel_797395 = array_index_797074 == array_index_773116 ? add_797394 : sel_797391;
  assign add_797398 = sel_797395 + 8'h01;
  assign sel_797399 = array_index_797074 == array_index_773122 ? add_797398 : sel_797395;
  assign add_797402 = sel_797399 + 8'h01;
  assign sel_797403 = array_index_797074 == array_index_773128 ? add_797402 : sel_797399;
  assign add_797406 = sel_797403 + 8'h01;
  assign sel_797407 = array_index_797074 == array_index_773134 ? add_797406 : sel_797403;
  assign add_797410 = sel_797407 + 8'h01;
  assign sel_797411 = array_index_797074 == array_index_773140 ? add_797410 : sel_797407;
  assign add_797414 = sel_797411 + 8'h01;
  assign sel_797415 = array_index_797074 == array_index_773146 ? add_797414 : sel_797411;
  assign add_797418 = sel_797415 + 8'h01;
  assign sel_797419 = array_index_797074 == array_index_773152 ? add_797418 : sel_797415;
  assign add_797422 = sel_797419 + 8'h01;
  assign sel_797423 = array_index_797074 == array_index_773158 ? add_797422 : sel_797419;
  assign add_797426 = sel_797423 + 8'h01;
  assign sel_797427 = array_index_797074 == array_index_773164 ? add_797426 : sel_797423;
  assign add_797430 = sel_797427 + 8'h01;
  assign sel_797431 = array_index_797074 == array_index_773170 ? add_797430 : sel_797427;
  assign add_797435 = sel_797431 + 8'h01;
  assign array_index_797436 = set1_unflattened[7'h44];
  assign sel_797437 = array_index_797074 == array_index_773176 ? add_797435 : sel_797431;
  assign add_797440 = sel_797437 + 8'h01;
  assign sel_797441 = array_index_797436 == array_index_772632 ? add_797440 : sel_797437;
  assign add_797444 = sel_797441 + 8'h01;
  assign sel_797445 = array_index_797436 == array_index_772636 ? add_797444 : sel_797441;
  assign add_797448 = sel_797445 + 8'h01;
  assign sel_797449 = array_index_797436 == array_index_772644 ? add_797448 : sel_797445;
  assign add_797452 = sel_797449 + 8'h01;
  assign sel_797453 = array_index_797436 == array_index_772652 ? add_797452 : sel_797449;
  assign add_797456 = sel_797453 + 8'h01;
  assign sel_797457 = array_index_797436 == array_index_772660 ? add_797456 : sel_797453;
  assign add_797460 = sel_797457 + 8'h01;
  assign sel_797461 = array_index_797436 == array_index_772668 ? add_797460 : sel_797457;
  assign add_797464 = sel_797461 + 8'h01;
  assign sel_797465 = array_index_797436 == array_index_772676 ? add_797464 : sel_797461;
  assign add_797468 = sel_797465 + 8'h01;
  assign sel_797469 = array_index_797436 == array_index_772684 ? add_797468 : sel_797465;
  assign add_797472 = sel_797469 + 8'h01;
  assign sel_797473 = array_index_797436 == array_index_772690 ? add_797472 : sel_797469;
  assign add_797476 = sel_797473 + 8'h01;
  assign sel_797477 = array_index_797436 == array_index_772696 ? add_797476 : sel_797473;
  assign add_797480 = sel_797477 + 8'h01;
  assign sel_797481 = array_index_797436 == array_index_772702 ? add_797480 : sel_797477;
  assign add_797484 = sel_797481 + 8'h01;
  assign sel_797485 = array_index_797436 == array_index_772708 ? add_797484 : sel_797481;
  assign add_797488 = sel_797485 + 8'h01;
  assign sel_797489 = array_index_797436 == array_index_772714 ? add_797488 : sel_797485;
  assign add_797492 = sel_797489 + 8'h01;
  assign sel_797493 = array_index_797436 == array_index_772720 ? add_797492 : sel_797489;
  assign add_797496 = sel_797493 + 8'h01;
  assign sel_797497 = array_index_797436 == array_index_772726 ? add_797496 : sel_797493;
  assign add_797500 = sel_797497 + 8'h01;
  assign sel_797501 = array_index_797436 == array_index_772732 ? add_797500 : sel_797497;
  assign add_797504 = sel_797501 + 8'h01;
  assign sel_797505 = array_index_797436 == array_index_772738 ? add_797504 : sel_797501;
  assign add_797508 = sel_797505 + 8'h01;
  assign sel_797509 = array_index_797436 == array_index_772744 ? add_797508 : sel_797505;
  assign add_797512 = sel_797509 + 8'h01;
  assign sel_797513 = array_index_797436 == array_index_772750 ? add_797512 : sel_797509;
  assign add_797516 = sel_797513 + 8'h01;
  assign sel_797517 = array_index_797436 == array_index_772756 ? add_797516 : sel_797513;
  assign add_797520 = sel_797517 + 8'h01;
  assign sel_797521 = array_index_797436 == array_index_772762 ? add_797520 : sel_797517;
  assign add_797524 = sel_797521 + 8'h01;
  assign sel_797525 = array_index_797436 == array_index_772768 ? add_797524 : sel_797521;
  assign add_797528 = sel_797525 + 8'h01;
  assign sel_797529 = array_index_797436 == array_index_772774 ? add_797528 : sel_797525;
  assign add_797532 = sel_797529 + 8'h01;
  assign sel_797533 = array_index_797436 == array_index_772780 ? add_797532 : sel_797529;
  assign add_797536 = sel_797533 + 8'h01;
  assign sel_797537 = array_index_797436 == array_index_772786 ? add_797536 : sel_797533;
  assign add_797540 = sel_797537 + 8'h01;
  assign sel_797541 = array_index_797436 == array_index_772792 ? add_797540 : sel_797537;
  assign add_797544 = sel_797541 + 8'h01;
  assign sel_797545 = array_index_797436 == array_index_772798 ? add_797544 : sel_797541;
  assign add_797548 = sel_797545 + 8'h01;
  assign sel_797549 = array_index_797436 == array_index_772804 ? add_797548 : sel_797545;
  assign add_797552 = sel_797549 + 8'h01;
  assign sel_797553 = array_index_797436 == array_index_772810 ? add_797552 : sel_797549;
  assign add_797556 = sel_797553 + 8'h01;
  assign sel_797557 = array_index_797436 == array_index_772816 ? add_797556 : sel_797553;
  assign add_797560 = sel_797557 + 8'h01;
  assign sel_797561 = array_index_797436 == array_index_772822 ? add_797560 : sel_797557;
  assign add_797564 = sel_797561 + 8'h01;
  assign sel_797565 = array_index_797436 == array_index_772828 ? add_797564 : sel_797561;
  assign add_797568 = sel_797565 + 8'h01;
  assign sel_797569 = array_index_797436 == array_index_772834 ? add_797568 : sel_797565;
  assign add_797572 = sel_797569 + 8'h01;
  assign sel_797573 = array_index_797436 == array_index_772840 ? add_797572 : sel_797569;
  assign add_797576 = sel_797573 + 8'h01;
  assign sel_797577 = array_index_797436 == array_index_772846 ? add_797576 : sel_797573;
  assign add_797580 = sel_797577 + 8'h01;
  assign sel_797581 = array_index_797436 == array_index_772852 ? add_797580 : sel_797577;
  assign add_797584 = sel_797581 + 8'h01;
  assign sel_797585 = array_index_797436 == array_index_772858 ? add_797584 : sel_797581;
  assign add_797588 = sel_797585 + 8'h01;
  assign sel_797589 = array_index_797436 == array_index_772864 ? add_797588 : sel_797585;
  assign add_797592 = sel_797589 + 8'h01;
  assign sel_797593 = array_index_797436 == array_index_772870 ? add_797592 : sel_797589;
  assign add_797596 = sel_797593 + 8'h01;
  assign sel_797597 = array_index_797436 == array_index_772876 ? add_797596 : sel_797593;
  assign add_797600 = sel_797597 + 8'h01;
  assign sel_797601 = array_index_797436 == array_index_772882 ? add_797600 : sel_797597;
  assign add_797604 = sel_797601 + 8'h01;
  assign sel_797605 = array_index_797436 == array_index_772888 ? add_797604 : sel_797601;
  assign add_797608 = sel_797605 + 8'h01;
  assign sel_797609 = array_index_797436 == array_index_772894 ? add_797608 : sel_797605;
  assign add_797612 = sel_797609 + 8'h01;
  assign sel_797613 = array_index_797436 == array_index_772900 ? add_797612 : sel_797609;
  assign add_797616 = sel_797613 + 8'h01;
  assign sel_797617 = array_index_797436 == array_index_772906 ? add_797616 : sel_797613;
  assign add_797620 = sel_797617 + 8'h01;
  assign sel_797621 = array_index_797436 == array_index_772912 ? add_797620 : sel_797617;
  assign add_797624 = sel_797621 + 8'h01;
  assign sel_797625 = array_index_797436 == array_index_772918 ? add_797624 : sel_797621;
  assign add_797628 = sel_797625 + 8'h01;
  assign sel_797629 = array_index_797436 == array_index_772924 ? add_797628 : sel_797625;
  assign add_797632 = sel_797629 + 8'h01;
  assign sel_797633 = array_index_797436 == array_index_772930 ? add_797632 : sel_797629;
  assign add_797636 = sel_797633 + 8'h01;
  assign sel_797637 = array_index_797436 == array_index_772936 ? add_797636 : sel_797633;
  assign add_797640 = sel_797637 + 8'h01;
  assign sel_797641 = array_index_797436 == array_index_772942 ? add_797640 : sel_797637;
  assign add_797644 = sel_797641 + 8'h01;
  assign sel_797645 = array_index_797436 == array_index_772948 ? add_797644 : sel_797641;
  assign add_797648 = sel_797645 + 8'h01;
  assign sel_797649 = array_index_797436 == array_index_772954 ? add_797648 : sel_797645;
  assign add_797652 = sel_797649 + 8'h01;
  assign sel_797653 = array_index_797436 == array_index_772960 ? add_797652 : sel_797649;
  assign add_797656 = sel_797653 + 8'h01;
  assign sel_797657 = array_index_797436 == array_index_772966 ? add_797656 : sel_797653;
  assign add_797660 = sel_797657 + 8'h01;
  assign sel_797661 = array_index_797436 == array_index_772972 ? add_797660 : sel_797657;
  assign add_797664 = sel_797661 + 8'h01;
  assign sel_797665 = array_index_797436 == array_index_772978 ? add_797664 : sel_797661;
  assign add_797668 = sel_797665 + 8'h01;
  assign sel_797669 = array_index_797436 == array_index_772984 ? add_797668 : sel_797665;
  assign add_797672 = sel_797669 + 8'h01;
  assign sel_797673 = array_index_797436 == array_index_772990 ? add_797672 : sel_797669;
  assign add_797676 = sel_797673 + 8'h01;
  assign sel_797677 = array_index_797436 == array_index_772996 ? add_797676 : sel_797673;
  assign add_797680 = sel_797677 + 8'h01;
  assign sel_797681 = array_index_797436 == array_index_773002 ? add_797680 : sel_797677;
  assign add_797684 = sel_797681 + 8'h01;
  assign sel_797685 = array_index_797436 == array_index_773008 ? add_797684 : sel_797681;
  assign add_797688 = sel_797685 + 8'h01;
  assign sel_797689 = array_index_797436 == array_index_773014 ? add_797688 : sel_797685;
  assign add_797692 = sel_797689 + 8'h01;
  assign sel_797693 = array_index_797436 == array_index_773020 ? add_797692 : sel_797689;
  assign add_797696 = sel_797693 + 8'h01;
  assign sel_797697 = array_index_797436 == array_index_773026 ? add_797696 : sel_797693;
  assign add_797700 = sel_797697 + 8'h01;
  assign sel_797701 = array_index_797436 == array_index_773032 ? add_797700 : sel_797697;
  assign add_797704 = sel_797701 + 8'h01;
  assign sel_797705 = array_index_797436 == array_index_773038 ? add_797704 : sel_797701;
  assign add_797708 = sel_797705 + 8'h01;
  assign sel_797709 = array_index_797436 == array_index_773044 ? add_797708 : sel_797705;
  assign add_797712 = sel_797709 + 8'h01;
  assign sel_797713 = array_index_797436 == array_index_773050 ? add_797712 : sel_797709;
  assign add_797716 = sel_797713 + 8'h01;
  assign sel_797717 = array_index_797436 == array_index_773056 ? add_797716 : sel_797713;
  assign add_797720 = sel_797717 + 8'h01;
  assign sel_797721 = array_index_797436 == array_index_773062 ? add_797720 : sel_797717;
  assign add_797724 = sel_797721 + 8'h01;
  assign sel_797725 = array_index_797436 == array_index_773068 ? add_797724 : sel_797721;
  assign add_797728 = sel_797725 + 8'h01;
  assign sel_797729 = array_index_797436 == array_index_773074 ? add_797728 : sel_797725;
  assign add_797732 = sel_797729 + 8'h01;
  assign sel_797733 = array_index_797436 == array_index_773080 ? add_797732 : sel_797729;
  assign add_797736 = sel_797733 + 8'h01;
  assign sel_797737 = array_index_797436 == array_index_773086 ? add_797736 : sel_797733;
  assign add_797740 = sel_797737 + 8'h01;
  assign sel_797741 = array_index_797436 == array_index_773092 ? add_797740 : sel_797737;
  assign add_797744 = sel_797741 + 8'h01;
  assign sel_797745 = array_index_797436 == array_index_773098 ? add_797744 : sel_797741;
  assign add_797748 = sel_797745 + 8'h01;
  assign sel_797749 = array_index_797436 == array_index_773104 ? add_797748 : sel_797745;
  assign add_797752 = sel_797749 + 8'h01;
  assign sel_797753 = array_index_797436 == array_index_773110 ? add_797752 : sel_797749;
  assign add_797756 = sel_797753 + 8'h01;
  assign sel_797757 = array_index_797436 == array_index_773116 ? add_797756 : sel_797753;
  assign add_797760 = sel_797757 + 8'h01;
  assign sel_797761 = array_index_797436 == array_index_773122 ? add_797760 : sel_797757;
  assign add_797764 = sel_797761 + 8'h01;
  assign sel_797765 = array_index_797436 == array_index_773128 ? add_797764 : sel_797761;
  assign add_797768 = sel_797765 + 8'h01;
  assign sel_797769 = array_index_797436 == array_index_773134 ? add_797768 : sel_797765;
  assign add_797772 = sel_797769 + 8'h01;
  assign sel_797773 = array_index_797436 == array_index_773140 ? add_797772 : sel_797769;
  assign add_797776 = sel_797773 + 8'h01;
  assign sel_797777 = array_index_797436 == array_index_773146 ? add_797776 : sel_797773;
  assign add_797780 = sel_797777 + 8'h01;
  assign sel_797781 = array_index_797436 == array_index_773152 ? add_797780 : sel_797777;
  assign add_797784 = sel_797781 + 8'h01;
  assign sel_797785 = array_index_797436 == array_index_773158 ? add_797784 : sel_797781;
  assign add_797788 = sel_797785 + 8'h01;
  assign sel_797789 = array_index_797436 == array_index_773164 ? add_797788 : sel_797785;
  assign add_797792 = sel_797789 + 8'h01;
  assign sel_797793 = array_index_797436 == array_index_773170 ? add_797792 : sel_797789;
  assign add_797797 = sel_797793 + 8'h01;
  assign array_index_797798 = set1_unflattened[7'h45];
  assign sel_797799 = array_index_797436 == array_index_773176 ? add_797797 : sel_797793;
  assign add_797802 = sel_797799 + 8'h01;
  assign sel_797803 = array_index_797798 == array_index_772632 ? add_797802 : sel_797799;
  assign add_797806 = sel_797803 + 8'h01;
  assign sel_797807 = array_index_797798 == array_index_772636 ? add_797806 : sel_797803;
  assign add_797810 = sel_797807 + 8'h01;
  assign sel_797811 = array_index_797798 == array_index_772644 ? add_797810 : sel_797807;
  assign add_797814 = sel_797811 + 8'h01;
  assign sel_797815 = array_index_797798 == array_index_772652 ? add_797814 : sel_797811;
  assign add_797818 = sel_797815 + 8'h01;
  assign sel_797819 = array_index_797798 == array_index_772660 ? add_797818 : sel_797815;
  assign add_797822 = sel_797819 + 8'h01;
  assign sel_797823 = array_index_797798 == array_index_772668 ? add_797822 : sel_797819;
  assign add_797826 = sel_797823 + 8'h01;
  assign sel_797827 = array_index_797798 == array_index_772676 ? add_797826 : sel_797823;
  assign add_797830 = sel_797827 + 8'h01;
  assign sel_797831 = array_index_797798 == array_index_772684 ? add_797830 : sel_797827;
  assign add_797834 = sel_797831 + 8'h01;
  assign sel_797835 = array_index_797798 == array_index_772690 ? add_797834 : sel_797831;
  assign add_797838 = sel_797835 + 8'h01;
  assign sel_797839 = array_index_797798 == array_index_772696 ? add_797838 : sel_797835;
  assign add_797842 = sel_797839 + 8'h01;
  assign sel_797843 = array_index_797798 == array_index_772702 ? add_797842 : sel_797839;
  assign add_797846 = sel_797843 + 8'h01;
  assign sel_797847 = array_index_797798 == array_index_772708 ? add_797846 : sel_797843;
  assign add_797850 = sel_797847 + 8'h01;
  assign sel_797851 = array_index_797798 == array_index_772714 ? add_797850 : sel_797847;
  assign add_797854 = sel_797851 + 8'h01;
  assign sel_797855 = array_index_797798 == array_index_772720 ? add_797854 : sel_797851;
  assign add_797858 = sel_797855 + 8'h01;
  assign sel_797859 = array_index_797798 == array_index_772726 ? add_797858 : sel_797855;
  assign add_797862 = sel_797859 + 8'h01;
  assign sel_797863 = array_index_797798 == array_index_772732 ? add_797862 : sel_797859;
  assign add_797866 = sel_797863 + 8'h01;
  assign sel_797867 = array_index_797798 == array_index_772738 ? add_797866 : sel_797863;
  assign add_797870 = sel_797867 + 8'h01;
  assign sel_797871 = array_index_797798 == array_index_772744 ? add_797870 : sel_797867;
  assign add_797874 = sel_797871 + 8'h01;
  assign sel_797875 = array_index_797798 == array_index_772750 ? add_797874 : sel_797871;
  assign add_797878 = sel_797875 + 8'h01;
  assign sel_797879 = array_index_797798 == array_index_772756 ? add_797878 : sel_797875;
  assign add_797882 = sel_797879 + 8'h01;
  assign sel_797883 = array_index_797798 == array_index_772762 ? add_797882 : sel_797879;
  assign add_797886 = sel_797883 + 8'h01;
  assign sel_797887 = array_index_797798 == array_index_772768 ? add_797886 : sel_797883;
  assign add_797890 = sel_797887 + 8'h01;
  assign sel_797891 = array_index_797798 == array_index_772774 ? add_797890 : sel_797887;
  assign add_797894 = sel_797891 + 8'h01;
  assign sel_797895 = array_index_797798 == array_index_772780 ? add_797894 : sel_797891;
  assign add_797898 = sel_797895 + 8'h01;
  assign sel_797899 = array_index_797798 == array_index_772786 ? add_797898 : sel_797895;
  assign add_797902 = sel_797899 + 8'h01;
  assign sel_797903 = array_index_797798 == array_index_772792 ? add_797902 : sel_797899;
  assign add_797906 = sel_797903 + 8'h01;
  assign sel_797907 = array_index_797798 == array_index_772798 ? add_797906 : sel_797903;
  assign add_797910 = sel_797907 + 8'h01;
  assign sel_797911 = array_index_797798 == array_index_772804 ? add_797910 : sel_797907;
  assign add_797914 = sel_797911 + 8'h01;
  assign sel_797915 = array_index_797798 == array_index_772810 ? add_797914 : sel_797911;
  assign add_797918 = sel_797915 + 8'h01;
  assign sel_797919 = array_index_797798 == array_index_772816 ? add_797918 : sel_797915;
  assign add_797922 = sel_797919 + 8'h01;
  assign sel_797923 = array_index_797798 == array_index_772822 ? add_797922 : sel_797919;
  assign add_797926 = sel_797923 + 8'h01;
  assign sel_797927 = array_index_797798 == array_index_772828 ? add_797926 : sel_797923;
  assign add_797930 = sel_797927 + 8'h01;
  assign sel_797931 = array_index_797798 == array_index_772834 ? add_797930 : sel_797927;
  assign add_797934 = sel_797931 + 8'h01;
  assign sel_797935 = array_index_797798 == array_index_772840 ? add_797934 : sel_797931;
  assign add_797938 = sel_797935 + 8'h01;
  assign sel_797939 = array_index_797798 == array_index_772846 ? add_797938 : sel_797935;
  assign add_797942 = sel_797939 + 8'h01;
  assign sel_797943 = array_index_797798 == array_index_772852 ? add_797942 : sel_797939;
  assign add_797946 = sel_797943 + 8'h01;
  assign sel_797947 = array_index_797798 == array_index_772858 ? add_797946 : sel_797943;
  assign add_797950 = sel_797947 + 8'h01;
  assign sel_797951 = array_index_797798 == array_index_772864 ? add_797950 : sel_797947;
  assign add_797954 = sel_797951 + 8'h01;
  assign sel_797955 = array_index_797798 == array_index_772870 ? add_797954 : sel_797951;
  assign add_797958 = sel_797955 + 8'h01;
  assign sel_797959 = array_index_797798 == array_index_772876 ? add_797958 : sel_797955;
  assign add_797962 = sel_797959 + 8'h01;
  assign sel_797963 = array_index_797798 == array_index_772882 ? add_797962 : sel_797959;
  assign add_797966 = sel_797963 + 8'h01;
  assign sel_797967 = array_index_797798 == array_index_772888 ? add_797966 : sel_797963;
  assign add_797970 = sel_797967 + 8'h01;
  assign sel_797971 = array_index_797798 == array_index_772894 ? add_797970 : sel_797967;
  assign add_797974 = sel_797971 + 8'h01;
  assign sel_797975 = array_index_797798 == array_index_772900 ? add_797974 : sel_797971;
  assign add_797978 = sel_797975 + 8'h01;
  assign sel_797979 = array_index_797798 == array_index_772906 ? add_797978 : sel_797975;
  assign add_797982 = sel_797979 + 8'h01;
  assign sel_797983 = array_index_797798 == array_index_772912 ? add_797982 : sel_797979;
  assign add_797986 = sel_797983 + 8'h01;
  assign sel_797987 = array_index_797798 == array_index_772918 ? add_797986 : sel_797983;
  assign add_797990 = sel_797987 + 8'h01;
  assign sel_797991 = array_index_797798 == array_index_772924 ? add_797990 : sel_797987;
  assign add_797994 = sel_797991 + 8'h01;
  assign sel_797995 = array_index_797798 == array_index_772930 ? add_797994 : sel_797991;
  assign add_797998 = sel_797995 + 8'h01;
  assign sel_797999 = array_index_797798 == array_index_772936 ? add_797998 : sel_797995;
  assign add_798002 = sel_797999 + 8'h01;
  assign sel_798003 = array_index_797798 == array_index_772942 ? add_798002 : sel_797999;
  assign add_798006 = sel_798003 + 8'h01;
  assign sel_798007 = array_index_797798 == array_index_772948 ? add_798006 : sel_798003;
  assign add_798010 = sel_798007 + 8'h01;
  assign sel_798011 = array_index_797798 == array_index_772954 ? add_798010 : sel_798007;
  assign add_798014 = sel_798011 + 8'h01;
  assign sel_798015 = array_index_797798 == array_index_772960 ? add_798014 : sel_798011;
  assign add_798018 = sel_798015 + 8'h01;
  assign sel_798019 = array_index_797798 == array_index_772966 ? add_798018 : sel_798015;
  assign add_798022 = sel_798019 + 8'h01;
  assign sel_798023 = array_index_797798 == array_index_772972 ? add_798022 : sel_798019;
  assign add_798026 = sel_798023 + 8'h01;
  assign sel_798027 = array_index_797798 == array_index_772978 ? add_798026 : sel_798023;
  assign add_798030 = sel_798027 + 8'h01;
  assign sel_798031 = array_index_797798 == array_index_772984 ? add_798030 : sel_798027;
  assign add_798034 = sel_798031 + 8'h01;
  assign sel_798035 = array_index_797798 == array_index_772990 ? add_798034 : sel_798031;
  assign add_798038 = sel_798035 + 8'h01;
  assign sel_798039 = array_index_797798 == array_index_772996 ? add_798038 : sel_798035;
  assign add_798042 = sel_798039 + 8'h01;
  assign sel_798043 = array_index_797798 == array_index_773002 ? add_798042 : sel_798039;
  assign add_798046 = sel_798043 + 8'h01;
  assign sel_798047 = array_index_797798 == array_index_773008 ? add_798046 : sel_798043;
  assign add_798050 = sel_798047 + 8'h01;
  assign sel_798051 = array_index_797798 == array_index_773014 ? add_798050 : sel_798047;
  assign add_798054 = sel_798051 + 8'h01;
  assign sel_798055 = array_index_797798 == array_index_773020 ? add_798054 : sel_798051;
  assign add_798058 = sel_798055 + 8'h01;
  assign sel_798059 = array_index_797798 == array_index_773026 ? add_798058 : sel_798055;
  assign add_798062 = sel_798059 + 8'h01;
  assign sel_798063 = array_index_797798 == array_index_773032 ? add_798062 : sel_798059;
  assign add_798066 = sel_798063 + 8'h01;
  assign sel_798067 = array_index_797798 == array_index_773038 ? add_798066 : sel_798063;
  assign add_798070 = sel_798067 + 8'h01;
  assign sel_798071 = array_index_797798 == array_index_773044 ? add_798070 : sel_798067;
  assign add_798074 = sel_798071 + 8'h01;
  assign sel_798075 = array_index_797798 == array_index_773050 ? add_798074 : sel_798071;
  assign add_798078 = sel_798075 + 8'h01;
  assign sel_798079 = array_index_797798 == array_index_773056 ? add_798078 : sel_798075;
  assign add_798082 = sel_798079 + 8'h01;
  assign sel_798083 = array_index_797798 == array_index_773062 ? add_798082 : sel_798079;
  assign add_798086 = sel_798083 + 8'h01;
  assign sel_798087 = array_index_797798 == array_index_773068 ? add_798086 : sel_798083;
  assign add_798090 = sel_798087 + 8'h01;
  assign sel_798091 = array_index_797798 == array_index_773074 ? add_798090 : sel_798087;
  assign add_798094 = sel_798091 + 8'h01;
  assign sel_798095 = array_index_797798 == array_index_773080 ? add_798094 : sel_798091;
  assign add_798098 = sel_798095 + 8'h01;
  assign sel_798099 = array_index_797798 == array_index_773086 ? add_798098 : sel_798095;
  assign add_798102 = sel_798099 + 8'h01;
  assign sel_798103 = array_index_797798 == array_index_773092 ? add_798102 : sel_798099;
  assign add_798106 = sel_798103 + 8'h01;
  assign sel_798107 = array_index_797798 == array_index_773098 ? add_798106 : sel_798103;
  assign add_798110 = sel_798107 + 8'h01;
  assign sel_798111 = array_index_797798 == array_index_773104 ? add_798110 : sel_798107;
  assign add_798114 = sel_798111 + 8'h01;
  assign sel_798115 = array_index_797798 == array_index_773110 ? add_798114 : sel_798111;
  assign add_798118 = sel_798115 + 8'h01;
  assign sel_798119 = array_index_797798 == array_index_773116 ? add_798118 : sel_798115;
  assign add_798122 = sel_798119 + 8'h01;
  assign sel_798123 = array_index_797798 == array_index_773122 ? add_798122 : sel_798119;
  assign add_798126 = sel_798123 + 8'h01;
  assign sel_798127 = array_index_797798 == array_index_773128 ? add_798126 : sel_798123;
  assign add_798130 = sel_798127 + 8'h01;
  assign sel_798131 = array_index_797798 == array_index_773134 ? add_798130 : sel_798127;
  assign add_798134 = sel_798131 + 8'h01;
  assign sel_798135 = array_index_797798 == array_index_773140 ? add_798134 : sel_798131;
  assign add_798138 = sel_798135 + 8'h01;
  assign sel_798139 = array_index_797798 == array_index_773146 ? add_798138 : sel_798135;
  assign add_798142 = sel_798139 + 8'h01;
  assign sel_798143 = array_index_797798 == array_index_773152 ? add_798142 : sel_798139;
  assign add_798146 = sel_798143 + 8'h01;
  assign sel_798147 = array_index_797798 == array_index_773158 ? add_798146 : sel_798143;
  assign add_798150 = sel_798147 + 8'h01;
  assign sel_798151 = array_index_797798 == array_index_773164 ? add_798150 : sel_798147;
  assign add_798154 = sel_798151 + 8'h01;
  assign sel_798155 = array_index_797798 == array_index_773170 ? add_798154 : sel_798151;
  assign add_798159 = sel_798155 + 8'h01;
  assign array_index_798160 = set1_unflattened[7'h46];
  assign sel_798161 = array_index_797798 == array_index_773176 ? add_798159 : sel_798155;
  assign add_798164 = sel_798161 + 8'h01;
  assign sel_798165 = array_index_798160 == array_index_772632 ? add_798164 : sel_798161;
  assign add_798168 = sel_798165 + 8'h01;
  assign sel_798169 = array_index_798160 == array_index_772636 ? add_798168 : sel_798165;
  assign add_798172 = sel_798169 + 8'h01;
  assign sel_798173 = array_index_798160 == array_index_772644 ? add_798172 : sel_798169;
  assign add_798176 = sel_798173 + 8'h01;
  assign sel_798177 = array_index_798160 == array_index_772652 ? add_798176 : sel_798173;
  assign add_798180 = sel_798177 + 8'h01;
  assign sel_798181 = array_index_798160 == array_index_772660 ? add_798180 : sel_798177;
  assign add_798184 = sel_798181 + 8'h01;
  assign sel_798185 = array_index_798160 == array_index_772668 ? add_798184 : sel_798181;
  assign add_798188 = sel_798185 + 8'h01;
  assign sel_798189 = array_index_798160 == array_index_772676 ? add_798188 : sel_798185;
  assign add_798192 = sel_798189 + 8'h01;
  assign sel_798193 = array_index_798160 == array_index_772684 ? add_798192 : sel_798189;
  assign add_798196 = sel_798193 + 8'h01;
  assign sel_798197 = array_index_798160 == array_index_772690 ? add_798196 : sel_798193;
  assign add_798200 = sel_798197 + 8'h01;
  assign sel_798201 = array_index_798160 == array_index_772696 ? add_798200 : sel_798197;
  assign add_798204 = sel_798201 + 8'h01;
  assign sel_798205 = array_index_798160 == array_index_772702 ? add_798204 : sel_798201;
  assign add_798208 = sel_798205 + 8'h01;
  assign sel_798209 = array_index_798160 == array_index_772708 ? add_798208 : sel_798205;
  assign add_798212 = sel_798209 + 8'h01;
  assign sel_798213 = array_index_798160 == array_index_772714 ? add_798212 : sel_798209;
  assign add_798216 = sel_798213 + 8'h01;
  assign sel_798217 = array_index_798160 == array_index_772720 ? add_798216 : sel_798213;
  assign add_798220 = sel_798217 + 8'h01;
  assign sel_798221 = array_index_798160 == array_index_772726 ? add_798220 : sel_798217;
  assign add_798224 = sel_798221 + 8'h01;
  assign sel_798225 = array_index_798160 == array_index_772732 ? add_798224 : sel_798221;
  assign add_798228 = sel_798225 + 8'h01;
  assign sel_798229 = array_index_798160 == array_index_772738 ? add_798228 : sel_798225;
  assign add_798232 = sel_798229 + 8'h01;
  assign sel_798233 = array_index_798160 == array_index_772744 ? add_798232 : sel_798229;
  assign add_798236 = sel_798233 + 8'h01;
  assign sel_798237 = array_index_798160 == array_index_772750 ? add_798236 : sel_798233;
  assign add_798240 = sel_798237 + 8'h01;
  assign sel_798241 = array_index_798160 == array_index_772756 ? add_798240 : sel_798237;
  assign add_798244 = sel_798241 + 8'h01;
  assign sel_798245 = array_index_798160 == array_index_772762 ? add_798244 : sel_798241;
  assign add_798248 = sel_798245 + 8'h01;
  assign sel_798249 = array_index_798160 == array_index_772768 ? add_798248 : sel_798245;
  assign add_798252 = sel_798249 + 8'h01;
  assign sel_798253 = array_index_798160 == array_index_772774 ? add_798252 : sel_798249;
  assign add_798256 = sel_798253 + 8'h01;
  assign sel_798257 = array_index_798160 == array_index_772780 ? add_798256 : sel_798253;
  assign add_798260 = sel_798257 + 8'h01;
  assign sel_798261 = array_index_798160 == array_index_772786 ? add_798260 : sel_798257;
  assign add_798264 = sel_798261 + 8'h01;
  assign sel_798265 = array_index_798160 == array_index_772792 ? add_798264 : sel_798261;
  assign add_798268 = sel_798265 + 8'h01;
  assign sel_798269 = array_index_798160 == array_index_772798 ? add_798268 : sel_798265;
  assign add_798272 = sel_798269 + 8'h01;
  assign sel_798273 = array_index_798160 == array_index_772804 ? add_798272 : sel_798269;
  assign add_798276 = sel_798273 + 8'h01;
  assign sel_798277 = array_index_798160 == array_index_772810 ? add_798276 : sel_798273;
  assign add_798280 = sel_798277 + 8'h01;
  assign sel_798281 = array_index_798160 == array_index_772816 ? add_798280 : sel_798277;
  assign add_798284 = sel_798281 + 8'h01;
  assign sel_798285 = array_index_798160 == array_index_772822 ? add_798284 : sel_798281;
  assign add_798288 = sel_798285 + 8'h01;
  assign sel_798289 = array_index_798160 == array_index_772828 ? add_798288 : sel_798285;
  assign add_798292 = sel_798289 + 8'h01;
  assign sel_798293 = array_index_798160 == array_index_772834 ? add_798292 : sel_798289;
  assign add_798296 = sel_798293 + 8'h01;
  assign sel_798297 = array_index_798160 == array_index_772840 ? add_798296 : sel_798293;
  assign add_798300 = sel_798297 + 8'h01;
  assign sel_798301 = array_index_798160 == array_index_772846 ? add_798300 : sel_798297;
  assign add_798304 = sel_798301 + 8'h01;
  assign sel_798305 = array_index_798160 == array_index_772852 ? add_798304 : sel_798301;
  assign add_798308 = sel_798305 + 8'h01;
  assign sel_798309 = array_index_798160 == array_index_772858 ? add_798308 : sel_798305;
  assign add_798312 = sel_798309 + 8'h01;
  assign sel_798313 = array_index_798160 == array_index_772864 ? add_798312 : sel_798309;
  assign add_798316 = sel_798313 + 8'h01;
  assign sel_798317 = array_index_798160 == array_index_772870 ? add_798316 : sel_798313;
  assign add_798320 = sel_798317 + 8'h01;
  assign sel_798321 = array_index_798160 == array_index_772876 ? add_798320 : sel_798317;
  assign add_798324 = sel_798321 + 8'h01;
  assign sel_798325 = array_index_798160 == array_index_772882 ? add_798324 : sel_798321;
  assign add_798328 = sel_798325 + 8'h01;
  assign sel_798329 = array_index_798160 == array_index_772888 ? add_798328 : sel_798325;
  assign add_798332 = sel_798329 + 8'h01;
  assign sel_798333 = array_index_798160 == array_index_772894 ? add_798332 : sel_798329;
  assign add_798336 = sel_798333 + 8'h01;
  assign sel_798337 = array_index_798160 == array_index_772900 ? add_798336 : sel_798333;
  assign add_798340 = sel_798337 + 8'h01;
  assign sel_798341 = array_index_798160 == array_index_772906 ? add_798340 : sel_798337;
  assign add_798344 = sel_798341 + 8'h01;
  assign sel_798345 = array_index_798160 == array_index_772912 ? add_798344 : sel_798341;
  assign add_798348 = sel_798345 + 8'h01;
  assign sel_798349 = array_index_798160 == array_index_772918 ? add_798348 : sel_798345;
  assign add_798352 = sel_798349 + 8'h01;
  assign sel_798353 = array_index_798160 == array_index_772924 ? add_798352 : sel_798349;
  assign add_798356 = sel_798353 + 8'h01;
  assign sel_798357 = array_index_798160 == array_index_772930 ? add_798356 : sel_798353;
  assign add_798360 = sel_798357 + 8'h01;
  assign sel_798361 = array_index_798160 == array_index_772936 ? add_798360 : sel_798357;
  assign add_798364 = sel_798361 + 8'h01;
  assign sel_798365 = array_index_798160 == array_index_772942 ? add_798364 : sel_798361;
  assign add_798368 = sel_798365 + 8'h01;
  assign sel_798369 = array_index_798160 == array_index_772948 ? add_798368 : sel_798365;
  assign add_798372 = sel_798369 + 8'h01;
  assign sel_798373 = array_index_798160 == array_index_772954 ? add_798372 : sel_798369;
  assign add_798376 = sel_798373 + 8'h01;
  assign sel_798377 = array_index_798160 == array_index_772960 ? add_798376 : sel_798373;
  assign add_798380 = sel_798377 + 8'h01;
  assign sel_798381 = array_index_798160 == array_index_772966 ? add_798380 : sel_798377;
  assign add_798384 = sel_798381 + 8'h01;
  assign sel_798385 = array_index_798160 == array_index_772972 ? add_798384 : sel_798381;
  assign add_798388 = sel_798385 + 8'h01;
  assign sel_798389 = array_index_798160 == array_index_772978 ? add_798388 : sel_798385;
  assign add_798392 = sel_798389 + 8'h01;
  assign sel_798393 = array_index_798160 == array_index_772984 ? add_798392 : sel_798389;
  assign add_798396 = sel_798393 + 8'h01;
  assign sel_798397 = array_index_798160 == array_index_772990 ? add_798396 : sel_798393;
  assign add_798400 = sel_798397 + 8'h01;
  assign sel_798401 = array_index_798160 == array_index_772996 ? add_798400 : sel_798397;
  assign add_798404 = sel_798401 + 8'h01;
  assign sel_798405 = array_index_798160 == array_index_773002 ? add_798404 : sel_798401;
  assign add_798408 = sel_798405 + 8'h01;
  assign sel_798409 = array_index_798160 == array_index_773008 ? add_798408 : sel_798405;
  assign add_798412 = sel_798409 + 8'h01;
  assign sel_798413 = array_index_798160 == array_index_773014 ? add_798412 : sel_798409;
  assign add_798416 = sel_798413 + 8'h01;
  assign sel_798417 = array_index_798160 == array_index_773020 ? add_798416 : sel_798413;
  assign add_798420 = sel_798417 + 8'h01;
  assign sel_798421 = array_index_798160 == array_index_773026 ? add_798420 : sel_798417;
  assign add_798424 = sel_798421 + 8'h01;
  assign sel_798425 = array_index_798160 == array_index_773032 ? add_798424 : sel_798421;
  assign add_798428 = sel_798425 + 8'h01;
  assign sel_798429 = array_index_798160 == array_index_773038 ? add_798428 : sel_798425;
  assign add_798432 = sel_798429 + 8'h01;
  assign sel_798433 = array_index_798160 == array_index_773044 ? add_798432 : sel_798429;
  assign add_798436 = sel_798433 + 8'h01;
  assign sel_798437 = array_index_798160 == array_index_773050 ? add_798436 : sel_798433;
  assign add_798440 = sel_798437 + 8'h01;
  assign sel_798441 = array_index_798160 == array_index_773056 ? add_798440 : sel_798437;
  assign add_798444 = sel_798441 + 8'h01;
  assign sel_798445 = array_index_798160 == array_index_773062 ? add_798444 : sel_798441;
  assign add_798448 = sel_798445 + 8'h01;
  assign sel_798449 = array_index_798160 == array_index_773068 ? add_798448 : sel_798445;
  assign add_798452 = sel_798449 + 8'h01;
  assign sel_798453 = array_index_798160 == array_index_773074 ? add_798452 : sel_798449;
  assign add_798456 = sel_798453 + 8'h01;
  assign sel_798457 = array_index_798160 == array_index_773080 ? add_798456 : sel_798453;
  assign add_798460 = sel_798457 + 8'h01;
  assign sel_798461 = array_index_798160 == array_index_773086 ? add_798460 : sel_798457;
  assign add_798464 = sel_798461 + 8'h01;
  assign sel_798465 = array_index_798160 == array_index_773092 ? add_798464 : sel_798461;
  assign add_798468 = sel_798465 + 8'h01;
  assign sel_798469 = array_index_798160 == array_index_773098 ? add_798468 : sel_798465;
  assign add_798472 = sel_798469 + 8'h01;
  assign sel_798473 = array_index_798160 == array_index_773104 ? add_798472 : sel_798469;
  assign add_798476 = sel_798473 + 8'h01;
  assign sel_798477 = array_index_798160 == array_index_773110 ? add_798476 : sel_798473;
  assign add_798480 = sel_798477 + 8'h01;
  assign sel_798481 = array_index_798160 == array_index_773116 ? add_798480 : sel_798477;
  assign add_798484 = sel_798481 + 8'h01;
  assign sel_798485 = array_index_798160 == array_index_773122 ? add_798484 : sel_798481;
  assign add_798488 = sel_798485 + 8'h01;
  assign sel_798489 = array_index_798160 == array_index_773128 ? add_798488 : sel_798485;
  assign add_798492 = sel_798489 + 8'h01;
  assign sel_798493 = array_index_798160 == array_index_773134 ? add_798492 : sel_798489;
  assign add_798496 = sel_798493 + 8'h01;
  assign sel_798497 = array_index_798160 == array_index_773140 ? add_798496 : sel_798493;
  assign add_798500 = sel_798497 + 8'h01;
  assign sel_798501 = array_index_798160 == array_index_773146 ? add_798500 : sel_798497;
  assign add_798504 = sel_798501 + 8'h01;
  assign sel_798505 = array_index_798160 == array_index_773152 ? add_798504 : sel_798501;
  assign add_798508 = sel_798505 + 8'h01;
  assign sel_798509 = array_index_798160 == array_index_773158 ? add_798508 : sel_798505;
  assign add_798512 = sel_798509 + 8'h01;
  assign sel_798513 = array_index_798160 == array_index_773164 ? add_798512 : sel_798509;
  assign add_798516 = sel_798513 + 8'h01;
  assign sel_798517 = array_index_798160 == array_index_773170 ? add_798516 : sel_798513;
  assign add_798521 = sel_798517 + 8'h01;
  assign array_index_798522 = set1_unflattened[7'h47];
  assign sel_798523 = array_index_798160 == array_index_773176 ? add_798521 : sel_798517;
  assign add_798526 = sel_798523 + 8'h01;
  assign sel_798527 = array_index_798522 == array_index_772632 ? add_798526 : sel_798523;
  assign add_798530 = sel_798527 + 8'h01;
  assign sel_798531 = array_index_798522 == array_index_772636 ? add_798530 : sel_798527;
  assign add_798534 = sel_798531 + 8'h01;
  assign sel_798535 = array_index_798522 == array_index_772644 ? add_798534 : sel_798531;
  assign add_798538 = sel_798535 + 8'h01;
  assign sel_798539 = array_index_798522 == array_index_772652 ? add_798538 : sel_798535;
  assign add_798542 = sel_798539 + 8'h01;
  assign sel_798543 = array_index_798522 == array_index_772660 ? add_798542 : sel_798539;
  assign add_798546 = sel_798543 + 8'h01;
  assign sel_798547 = array_index_798522 == array_index_772668 ? add_798546 : sel_798543;
  assign add_798550 = sel_798547 + 8'h01;
  assign sel_798551 = array_index_798522 == array_index_772676 ? add_798550 : sel_798547;
  assign add_798554 = sel_798551 + 8'h01;
  assign sel_798555 = array_index_798522 == array_index_772684 ? add_798554 : sel_798551;
  assign add_798558 = sel_798555 + 8'h01;
  assign sel_798559 = array_index_798522 == array_index_772690 ? add_798558 : sel_798555;
  assign add_798562 = sel_798559 + 8'h01;
  assign sel_798563 = array_index_798522 == array_index_772696 ? add_798562 : sel_798559;
  assign add_798566 = sel_798563 + 8'h01;
  assign sel_798567 = array_index_798522 == array_index_772702 ? add_798566 : sel_798563;
  assign add_798570 = sel_798567 + 8'h01;
  assign sel_798571 = array_index_798522 == array_index_772708 ? add_798570 : sel_798567;
  assign add_798574 = sel_798571 + 8'h01;
  assign sel_798575 = array_index_798522 == array_index_772714 ? add_798574 : sel_798571;
  assign add_798578 = sel_798575 + 8'h01;
  assign sel_798579 = array_index_798522 == array_index_772720 ? add_798578 : sel_798575;
  assign add_798582 = sel_798579 + 8'h01;
  assign sel_798583 = array_index_798522 == array_index_772726 ? add_798582 : sel_798579;
  assign add_798586 = sel_798583 + 8'h01;
  assign sel_798587 = array_index_798522 == array_index_772732 ? add_798586 : sel_798583;
  assign add_798590 = sel_798587 + 8'h01;
  assign sel_798591 = array_index_798522 == array_index_772738 ? add_798590 : sel_798587;
  assign add_798594 = sel_798591 + 8'h01;
  assign sel_798595 = array_index_798522 == array_index_772744 ? add_798594 : sel_798591;
  assign add_798598 = sel_798595 + 8'h01;
  assign sel_798599 = array_index_798522 == array_index_772750 ? add_798598 : sel_798595;
  assign add_798602 = sel_798599 + 8'h01;
  assign sel_798603 = array_index_798522 == array_index_772756 ? add_798602 : sel_798599;
  assign add_798606 = sel_798603 + 8'h01;
  assign sel_798607 = array_index_798522 == array_index_772762 ? add_798606 : sel_798603;
  assign add_798610 = sel_798607 + 8'h01;
  assign sel_798611 = array_index_798522 == array_index_772768 ? add_798610 : sel_798607;
  assign add_798614 = sel_798611 + 8'h01;
  assign sel_798615 = array_index_798522 == array_index_772774 ? add_798614 : sel_798611;
  assign add_798618 = sel_798615 + 8'h01;
  assign sel_798619 = array_index_798522 == array_index_772780 ? add_798618 : sel_798615;
  assign add_798622 = sel_798619 + 8'h01;
  assign sel_798623 = array_index_798522 == array_index_772786 ? add_798622 : sel_798619;
  assign add_798626 = sel_798623 + 8'h01;
  assign sel_798627 = array_index_798522 == array_index_772792 ? add_798626 : sel_798623;
  assign add_798630 = sel_798627 + 8'h01;
  assign sel_798631 = array_index_798522 == array_index_772798 ? add_798630 : sel_798627;
  assign add_798634 = sel_798631 + 8'h01;
  assign sel_798635 = array_index_798522 == array_index_772804 ? add_798634 : sel_798631;
  assign add_798638 = sel_798635 + 8'h01;
  assign sel_798639 = array_index_798522 == array_index_772810 ? add_798638 : sel_798635;
  assign add_798642 = sel_798639 + 8'h01;
  assign sel_798643 = array_index_798522 == array_index_772816 ? add_798642 : sel_798639;
  assign add_798646 = sel_798643 + 8'h01;
  assign sel_798647 = array_index_798522 == array_index_772822 ? add_798646 : sel_798643;
  assign add_798650 = sel_798647 + 8'h01;
  assign sel_798651 = array_index_798522 == array_index_772828 ? add_798650 : sel_798647;
  assign add_798654 = sel_798651 + 8'h01;
  assign sel_798655 = array_index_798522 == array_index_772834 ? add_798654 : sel_798651;
  assign add_798658 = sel_798655 + 8'h01;
  assign sel_798659 = array_index_798522 == array_index_772840 ? add_798658 : sel_798655;
  assign add_798662 = sel_798659 + 8'h01;
  assign sel_798663 = array_index_798522 == array_index_772846 ? add_798662 : sel_798659;
  assign add_798666 = sel_798663 + 8'h01;
  assign sel_798667 = array_index_798522 == array_index_772852 ? add_798666 : sel_798663;
  assign add_798670 = sel_798667 + 8'h01;
  assign sel_798671 = array_index_798522 == array_index_772858 ? add_798670 : sel_798667;
  assign add_798674 = sel_798671 + 8'h01;
  assign sel_798675 = array_index_798522 == array_index_772864 ? add_798674 : sel_798671;
  assign add_798678 = sel_798675 + 8'h01;
  assign sel_798679 = array_index_798522 == array_index_772870 ? add_798678 : sel_798675;
  assign add_798682 = sel_798679 + 8'h01;
  assign sel_798683 = array_index_798522 == array_index_772876 ? add_798682 : sel_798679;
  assign add_798686 = sel_798683 + 8'h01;
  assign sel_798687 = array_index_798522 == array_index_772882 ? add_798686 : sel_798683;
  assign add_798690 = sel_798687 + 8'h01;
  assign sel_798691 = array_index_798522 == array_index_772888 ? add_798690 : sel_798687;
  assign add_798694 = sel_798691 + 8'h01;
  assign sel_798695 = array_index_798522 == array_index_772894 ? add_798694 : sel_798691;
  assign add_798698 = sel_798695 + 8'h01;
  assign sel_798699 = array_index_798522 == array_index_772900 ? add_798698 : sel_798695;
  assign add_798702 = sel_798699 + 8'h01;
  assign sel_798703 = array_index_798522 == array_index_772906 ? add_798702 : sel_798699;
  assign add_798706 = sel_798703 + 8'h01;
  assign sel_798707 = array_index_798522 == array_index_772912 ? add_798706 : sel_798703;
  assign add_798710 = sel_798707 + 8'h01;
  assign sel_798711 = array_index_798522 == array_index_772918 ? add_798710 : sel_798707;
  assign add_798714 = sel_798711 + 8'h01;
  assign sel_798715 = array_index_798522 == array_index_772924 ? add_798714 : sel_798711;
  assign add_798718 = sel_798715 + 8'h01;
  assign sel_798719 = array_index_798522 == array_index_772930 ? add_798718 : sel_798715;
  assign add_798722 = sel_798719 + 8'h01;
  assign sel_798723 = array_index_798522 == array_index_772936 ? add_798722 : sel_798719;
  assign add_798726 = sel_798723 + 8'h01;
  assign sel_798727 = array_index_798522 == array_index_772942 ? add_798726 : sel_798723;
  assign add_798730 = sel_798727 + 8'h01;
  assign sel_798731 = array_index_798522 == array_index_772948 ? add_798730 : sel_798727;
  assign add_798734 = sel_798731 + 8'h01;
  assign sel_798735 = array_index_798522 == array_index_772954 ? add_798734 : sel_798731;
  assign add_798738 = sel_798735 + 8'h01;
  assign sel_798739 = array_index_798522 == array_index_772960 ? add_798738 : sel_798735;
  assign add_798742 = sel_798739 + 8'h01;
  assign sel_798743 = array_index_798522 == array_index_772966 ? add_798742 : sel_798739;
  assign add_798746 = sel_798743 + 8'h01;
  assign sel_798747 = array_index_798522 == array_index_772972 ? add_798746 : sel_798743;
  assign add_798750 = sel_798747 + 8'h01;
  assign sel_798751 = array_index_798522 == array_index_772978 ? add_798750 : sel_798747;
  assign add_798754 = sel_798751 + 8'h01;
  assign sel_798755 = array_index_798522 == array_index_772984 ? add_798754 : sel_798751;
  assign add_798758 = sel_798755 + 8'h01;
  assign sel_798759 = array_index_798522 == array_index_772990 ? add_798758 : sel_798755;
  assign add_798762 = sel_798759 + 8'h01;
  assign sel_798763 = array_index_798522 == array_index_772996 ? add_798762 : sel_798759;
  assign add_798766 = sel_798763 + 8'h01;
  assign sel_798767 = array_index_798522 == array_index_773002 ? add_798766 : sel_798763;
  assign add_798770 = sel_798767 + 8'h01;
  assign sel_798771 = array_index_798522 == array_index_773008 ? add_798770 : sel_798767;
  assign add_798774 = sel_798771 + 8'h01;
  assign sel_798775 = array_index_798522 == array_index_773014 ? add_798774 : sel_798771;
  assign add_798778 = sel_798775 + 8'h01;
  assign sel_798779 = array_index_798522 == array_index_773020 ? add_798778 : sel_798775;
  assign add_798782 = sel_798779 + 8'h01;
  assign sel_798783 = array_index_798522 == array_index_773026 ? add_798782 : sel_798779;
  assign add_798786 = sel_798783 + 8'h01;
  assign sel_798787 = array_index_798522 == array_index_773032 ? add_798786 : sel_798783;
  assign add_798790 = sel_798787 + 8'h01;
  assign sel_798791 = array_index_798522 == array_index_773038 ? add_798790 : sel_798787;
  assign add_798794 = sel_798791 + 8'h01;
  assign sel_798795 = array_index_798522 == array_index_773044 ? add_798794 : sel_798791;
  assign add_798798 = sel_798795 + 8'h01;
  assign sel_798799 = array_index_798522 == array_index_773050 ? add_798798 : sel_798795;
  assign add_798802 = sel_798799 + 8'h01;
  assign sel_798803 = array_index_798522 == array_index_773056 ? add_798802 : sel_798799;
  assign add_798806 = sel_798803 + 8'h01;
  assign sel_798807 = array_index_798522 == array_index_773062 ? add_798806 : sel_798803;
  assign add_798810 = sel_798807 + 8'h01;
  assign sel_798811 = array_index_798522 == array_index_773068 ? add_798810 : sel_798807;
  assign add_798814 = sel_798811 + 8'h01;
  assign sel_798815 = array_index_798522 == array_index_773074 ? add_798814 : sel_798811;
  assign add_798818 = sel_798815 + 8'h01;
  assign sel_798819 = array_index_798522 == array_index_773080 ? add_798818 : sel_798815;
  assign add_798822 = sel_798819 + 8'h01;
  assign sel_798823 = array_index_798522 == array_index_773086 ? add_798822 : sel_798819;
  assign add_798826 = sel_798823 + 8'h01;
  assign sel_798827 = array_index_798522 == array_index_773092 ? add_798826 : sel_798823;
  assign add_798830 = sel_798827 + 8'h01;
  assign sel_798831 = array_index_798522 == array_index_773098 ? add_798830 : sel_798827;
  assign add_798834 = sel_798831 + 8'h01;
  assign sel_798835 = array_index_798522 == array_index_773104 ? add_798834 : sel_798831;
  assign add_798838 = sel_798835 + 8'h01;
  assign sel_798839 = array_index_798522 == array_index_773110 ? add_798838 : sel_798835;
  assign add_798842 = sel_798839 + 8'h01;
  assign sel_798843 = array_index_798522 == array_index_773116 ? add_798842 : sel_798839;
  assign add_798846 = sel_798843 + 8'h01;
  assign sel_798847 = array_index_798522 == array_index_773122 ? add_798846 : sel_798843;
  assign add_798850 = sel_798847 + 8'h01;
  assign sel_798851 = array_index_798522 == array_index_773128 ? add_798850 : sel_798847;
  assign add_798854 = sel_798851 + 8'h01;
  assign sel_798855 = array_index_798522 == array_index_773134 ? add_798854 : sel_798851;
  assign add_798858 = sel_798855 + 8'h01;
  assign sel_798859 = array_index_798522 == array_index_773140 ? add_798858 : sel_798855;
  assign add_798862 = sel_798859 + 8'h01;
  assign sel_798863 = array_index_798522 == array_index_773146 ? add_798862 : sel_798859;
  assign add_798866 = sel_798863 + 8'h01;
  assign sel_798867 = array_index_798522 == array_index_773152 ? add_798866 : sel_798863;
  assign add_798870 = sel_798867 + 8'h01;
  assign sel_798871 = array_index_798522 == array_index_773158 ? add_798870 : sel_798867;
  assign add_798874 = sel_798871 + 8'h01;
  assign sel_798875 = array_index_798522 == array_index_773164 ? add_798874 : sel_798871;
  assign add_798878 = sel_798875 + 8'h01;
  assign sel_798879 = array_index_798522 == array_index_773170 ? add_798878 : sel_798875;
  assign add_798883 = sel_798879 + 8'h01;
  assign array_index_798884 = set1_unflattened[7'h48];
  assign sel_798885 = array_index_798522 == array_index_773176 ? add_798883 : sel_798879;
  assign add_798888 = sel_798885 + 8'h01;
  assign sel_798889 = array_index_798884 == array_index_772632 ? add_798888 : sel_798885;
  assign add_798892 = sel_798889 + 8'h01;
  assign sel_798893 = array_index_798884 == array_index_772636 ? add_798892 : sel_798889;
  assign add_798896 = sel_798893 + 8'h01;
  assign sel_798897 = array_index_798884 == array_index_772644 ? add_798896 : sel_798893;
  assign add_798900 = sel_798897 + 8'h01;
  assign sel_798901 = array_index_798884 == array_index_772652 ? add_798900 : sel_798897;
  assign add_798904 = sel_798901 + 8'h01;
  assign sel_798905 = array_index_798884 == array_index_772660 ? add_798904 : sel_798901;
  assign add_798908 = sel_798905 + 8'h01;
  assign sel_798909 = array_index_798884 == array_index_772668 ? add_798908 : sel_798905;
  assign add_798912 = sel_798909 + 8'h01;
  assign sel_798913 = array_index_798884 == array_index_772676 ? add_798912 : sel_798909;
  assign add_798916 = sel_798913 + 8'h01;
  assign sel_798917 = array_index_798884 == array_index_772684 ? add_798916 : sel_798913;
  assign add_798920 = sel_798917 + 8'h01;
  assign sel_798921 = array_index_798884 == array_index_772690 ? add_798920 : sel_798917;
  assign add_798924 = sel_798921 + 8'h01;
  assign sel_798925 = array_index_798884 == array_index_772696 ? add_798924 : sel_798921;
  assign add_798928 = sel_798925 + 8'h01;
  assign sel_798929 = array_index_798884 == array_index_772702 ? add_798928 : sel_798925;
  assign add_798932 = sel_798929 + 8'h01;
  assign sel_798933 = array_index_798884 == array_index_772708 ? add_798932 : sel_798929;
  assign add_798936 = sel_798933 + 8'h01;
  assign sel_798937 = array_index_798884 == array_index_772714 ? add_798936 : sel_798933;
  assign add_798940 = sel_798937 + 8'h01;
  assign sel_798941 = array_index_798884 == array_index_772720 ? add_798940 : sel_798937;
  assign add_798944 = sel_798941 + 8'h01;
  assign sel_798945 = array_index_798884 == array_index_772726 ? add_798944 : sel_798941;
  assign add_798948 = sel_798945 + 8'h01;
  assign sel_798949 = array_index_798884 == array_index_772732 ? add_798948 : sel_798945;
  assign add_798952 = sel_798949 + 8'h01;
  assign sel_798953 = array_index_798884 == array_index_772738 ? add_798952 : sel_798949;
  assign add_798956 = sel_798953 + 8'h01;
  assign sel_798957 = array_index_798884 == array_index_772744 ? add_798956 : sel_798953;
  assign add_798960 = sel_798957 + 8'h01;
  assign sel_798961 = array_index_798884 == array_index_772750 ? add_798960 : sel_798957;
  assign add_798964 = sel_798961 + 8'h01;
  assign sel_798965 = array_index_798884 == array_index_772756 ? add_798964 : sel_798961;
  assign add_798968 = sel_798965 + 8'h01;
  assign sel_798969 = array_index_798884 == array_index_772762 ? add_798968 : sel_798965;
  assign add_798972 = sel_798969 + 8'h01;
  assign sel_798973 = array_index_798884 == array_index_772768 ? add_798972 : sel_798969;
  assign add_798976 = sel_798973 + 8'h01;
  assign sel_798977 = array_index_798884 == array_index_772774 ? add_798976 : sel_798973;
  assign add_798980 = sel_798977 + 8'h01;
  assign sel_798981 = array_index_798884 == array_index_772780 ? add_798980 : sel_798977;
  assign add_798984 = sel_798981 + 8'h01;
  assign sel_798985 = array_index_798884 == array_index_772786 ? add_798984 : sel_798981;
  assign add_798988 = sel_798985 + 8'h01;
  assign sel_798989 = array_index_798884 == array_index_772792 ? add_798988 : sel_798985;
  assign add_798992 = sel_798989 + 8'h01;
  assign sel_798993 = array_index_798884 == array_index_772798 ? add_798992 : sel_798989;
  assign add_798996 = sel_798993 + 8'h01;
  assign sel_798997 = array_index_798884 == array_index_772804 ? add_798996 : sel_798993;
  assign add_799000 = sel_798997 + 8'h01;
  assign sel_799001 = array_index_798884 == array_index_772810 ? add_799000 : sel_798997;
  assign add_799004 = sel_799001 + 8'h01;
  assign sel_799005 = array_index_798884 == array_index_772816 ? add_799004 : sel_799001;
  assign add_799008 = sel_799005 + 8'h01;
  assign sel_799009 = array_index_798884 == array_index_772822 ? add_799008 : sel_799005;
  assign add_799012 = sel_799009 + 8'h01;
  assign sel_799013 = array_index_798884 == array_index_772828 ? add_799012 : sel_799009;
  assign add_799016 = sel_799013 + 8'h01;
  assign sel_799017 = array_index_798884 == array_index_772834 ? add_799016 : sel_799013;
  assign add_799020 = sel_799017 + 8'h01;
  assign sel_799021 = array_index_798884 == array_index_772840 ? add_799020 : sel_799017;
  assign add_799024 = sel_799021 + 8'h01;
  assign sel_799025 = array_index_798884 == array_index_772846 ? add_799024 : sel_799021;
  assign add_799028 = sel_799025 + 8'h01;
  assign sel_799029 = array_index_798884 == array_index_772852 ? add_799028 : sel_799025;
  assign add_799032 = sel_799029 + 8'h01;
  assign sel_799033 = array_index_798884 == array_index_772858 ? add_799032 : sel_799029;
  assign add_799036 = sel_799033 + 8'h01;
  assign sel_799037 = array_index_798884 == array_index_772864 ? add_799036 : sel_799033;
  assign add_799040 = sel_799037 + 8'h01;
  assign sel_799041 = array_index_798884 == array_index_772870 ? add_799040 : sel_799037;
  assign add_799044 = sel_799041 + 8'h01;
  assign sel_799045 = array_index_798884 == array_index_772876 ? add_799044 : sel_799041;
  assign add_799048 = sel_799045 + 8'h01;
  assign sel_799049 = array_index_798884 == array_index_772882 ? add_799048 : sel_799045;
  assign add_799052 = sel_799049 + 8'h01;
  assign sel_799053 = array_index_798884 == array_index_772888 ? add_799052 : sel_799049;
  assign add_799056 = sel_799053 + 8'h01;
  assign sel_799057 = array_index_798884 == array_index_772894 ? add_799056 : sel_799053;
  assign add_799060 = sel_799057 + 8'h01;
  assign sel_799061 = array_index_798884 == array_index_772900 ? add_799060 : sel_799057;
  assign add_799064 = sel_799061 + 8'h01;
  assign sel_799065 = array_index_798884 == array_index_772906 ? add_799064 : sel_799061;
  assign add_799068 = sel_799065 + 8'h01;
  assign sel_799069 = array_index_798884 == array_index_772912 ? add_799068 : sel_799065;
  assign add_799072 = sel_799069 + 8'h01;
  assign sel_799073 = array_index_798884 == array_index_772918 ? add_799072 : sel_799069;
  assign add_799076 = sel_799073 + 8'h01;
  assign sel_799077 = array_index_798884 == array_index_772924 ? add_799076 : sel_799073;
  assign add_799080 = sel_799077 + 8'h01;
  assign sel_799081 = array_index_798884 == array_index_772930 ? add_799080 : sel_799077;
  assign add_799084 = sel_799081 + 8'h01;
  assign sel_799085 = array_index_798884 == array_index_772936 ? add_799084 : sel_799081;
  assign add_799088 = sel_799085 + 8'h01;
  assign sel_799089 = array_index_798884 == array_index_772942 ? add_799088 : sel_799085;
  assign add_799092 = sel_799089 + 8'h01;
  assign sel_799093 = array_index_798884 == array_index_772948 ? add_799092 : sel_799089;
  assign add_799096 = sel_799093 + 8'h01;
  assign sel_799097 = array_index_798884 == array_index_772954 ? add_799096 : sel_799093;
  assign add_799100 = sel_799097 + 8'h01;
  assign sel_799101 = array_index_798884 == array_index_772960 ? add_799100 : sel_799097;
  assign add_799104 = sel_799101 + 8'h01;
  assign sel_799105 = array_index_798884 == array_index_772966 ? add_799104 : sel_799101;
  assign add_799108 = sel_799105 + 8'h01;
  assign sel_799109 = array_index_798884 == array_index_772972 ? add_799108 : sel_799105;
  assign add_799112 = sel_799109 + 8'h01;
  assign sel_799113 = array_index_798884 == array_index_772978 ? add_799112 : sel_799109;
  assign add_799116 = sel_799113 + 8'h01;
  assign sel_799117 = array_index_798884 == array_index_772984 ? add_799116 : sel_799113;
  assign add_799120 = sel_799117 + 8'h01;
  assign sel_799121 = array_index_798884 == array_index_772990 ? add_799120 : sel_799117;
  assign add_799124 = sel_799121 + 8'h01;
  assign sel_799125 = array_index_798884 == array_index_772996 ? add_799124 : sel_799121;
  assign add_799128 = sel_799125 + 8'h01;
  assign sel_799129 = array_index_798884 == array_index_773002 ? add_799128 : sel_799125;
  assign add_799132 = sel_799129 + 8'h01;
  assign sel_799133 = array_index_798884 == array_index_773008 ? add_799132 : sel_799129;
  assign add_799136 = sel_799133 + 8'h01;
  assign sel_799137 = array_index_798884 == array_index_773014 ? add_799136 : sel_799133;
  assign add_799140 = sel_799137 + 8'h01;
  assign sel_799141 = array_index_798884 == array_index_773020 ? add_799140 : sel_799137;
  assign add_799144 = sel_799141 + 8'h01;
  assign sel_799145 = array_index_798884 == array_index_773026 ? add_799144 : sel_799141;
  assign add_799148 = sel_799145 + 8'h01;
  assign sel_799149 = array_index_798884 == array_index_773032 ? add_799148 : sel_799145;
  assign add_799152 = sel_799149 + 8'h01;
  assign sel_799153 = array_index_798884 == array_index_773038 ? add_799152 : sel_799149;
  assign add_799156 = sel_799153 + 8'h01;
  assign sel_799157 = array_index_798884 == array_index_773044 ? add_799156 : sel_799153;
  assign add_799160 = sel_799157 + 8'h01;
  assign sel_799161 = array_index_798884 == array_index_773050 ? add_799160 : sel_799157;
  assign add_799164 = sel_799161 + 8'h01;
  assign sel_799165 = array_index_798884 == array_index_773056 ? add_799164 : sel_799161;
  assign add_799168 = sel_799165 + 8'h01;
  assign sel_799169 = array_index_798884 == array_index_773062 ? add_799168 : sel_799165;
  assign add_799172 = sel_799169 + 8'h01;
  assign sel_799173 = array_index_798884 == array_index_773068 ? add_799172 : sel_799169;
  assign add_799176 = sel_799173 + 8'h01;
  assign sel_799177 = array_index_798884 == array_index_773074 ? add_799176 : sel_799173;
  assign add_799180 = sel_799177 + 8'h01;
  assign sel_799181 = array_index_798884 == array_index_773080 ? add_799180 : sel_799177;
  assign add_799184 = sel_799181 + 8'h01;
  assign sel_799185 = array_index_798884 == array_index_773086 ? add_799184 : sel_799181;
  assign add_799188 = sel_799185 + 8'h01;
  assign sel_799189 = array_index_798884 == array_index_773092 ? add_799188 : sel_799185;
  assign add_799192 = sel_799189 + 8'h01;
  assign sel_799193 = array_index_798884 == array_index_773098 ? add_799192 : sel_799189;
  assign add_799196 = sel_799193 + 8'h01;
  assign sel_799197 = array_index_798884 == array_index_773104 ? add_799196 : sel_799193;
  assign add_799200 = sel_799197 + 8'h01;
  assign sel_799201 = array_index_798884 == array_index_773110 ? add_799200 : sel_799197;
  assign add_799204 = sel_799201 + 8'h01;
  assign sel_799205 = array_index_798884 == array_index_773116 ? add_799204 : sel_799201;
  assign add_799208 = sel_799205 + 8'h01;
  assign sel_799209 = array_index_798884 == array_index_773122 ? add_799208 : sel_799205;
  assign add_799212 = sel_799209 + 8'h01;
  assign sel_799213 = array_index_798884 == array_index_773128 ? add_799212 : sel_799209;
  assign add_799216 = sel_799213 + 8'h01;
  assign sel_799217 = array_index_798884 == array_index_773134 ? add_799216 : sel_799213;
  assign add_799220 = sel_799217 + 8'h01;
  assign sel_799221 = array_index_798884 == array_index_773140 ? add_799220 : sel_799217;
  assign add_799224 = sel_799221 + 8'h01;
  assign sel_799225 = array_index_798884 == array_index_773146 ? add_799224 : sel_799221;
  assign add_799228 = sel_799225 + 8'h01;
  assign sel_799229 = array_index_798884 == array_index_773152 ? add_799228 : sel_799225;
  assign add_799232 = sel_799229 + 8'h01;
  assign sel_799233 = array_index_798884 == array_index_773158 ? add_799232 : sel_799229;
  assign add_799236 = sel_799233 + 8'h01;
  assign sel_799237 = array_index_798884 == array_index_773164 ? add_799236 : sel_799233;
  assign add_799240 = sel_799237 + 8'h01;
  assign sel_799241 = array_index_798884 == array_index_773170 ? add_799240 : sel_799237;
  assign add_799245 = sel_799241 + 8'h01;
  assign array_index_799246 = set1_unflattened[7'h49];
  assign sel_799247 = array_index_798884 == array_index_773176 ? add_799245 : sel_799241;
  assign add_799250 = sel_799247 + 8'h01;
  assign sel_799251 = array_index_799246 == array_index_772632 ? add_799250 : sel_799247;
  assign add_799254 = sel_799251 + 8'h01;
  assign sel_799255 = array_index_799246 == array_index_772636 ? add_799254 : sel_799251;
  assign add_799258 = sel_799255 + 8'h01;
  assign sel_799259 = array_index_799246 == array_index_772644 ? add_799258 : sel_799255;
  assign add_799262 = sel_799259 + 8'h01;
  assign sel_799263 = array_index_799246 == array_index_772652 ? add_799262 : sel_799259;
  assign add_799266 = sel_799263 + 8'h01;
  assign sel_799267 = array_index_799246 == array_index_772660 ? add_799266 : sel_799263;
  assign add_799270 = sel_799267 + 8'h01;
  assign sel_799271 = array_index_799246 == array_index_772668 ? add_799270 : sel_799267;
  assign add_799274 = sel_799271 + 8'h01;
  assign sel_799275 = array_index_799246 == array_index_772676 ? add_799274 : sel_799271;
  assign add_799278 = sel_799275 + 8'h01;
  assign sel_799279 = array_index_799246 == array_index_772684 ? add_799278 : sel_799275;
  assign add_799282 = sel_799279 + 8'h01;
  assign sel_799283 = array_index_799246 == array_index_772690 ? add_799282 : sel_799279;
  assign add_799286 = sel_799283 + 8'h01;
  assign sel_799287 = array_index_799246 == array_index_772696 ? add_799286 : sel_799283;
  assign add_799290 = sel_799287 + 8'h01;
  assign sel_799291 = array_index_799246 == array_index_772702 ? add_799290 : sel_799287;
  assign add_799294 = sel_799291 + 8'h01;
  assign sel_799295 = array_index_799246 == array_index_772708 ? add_799294 : sel_799291;
  assign add_799298 = sel_799295 + 8'h01;
  assign sel_799299 = array_index_799246 == array_index_772714 ? add_799298 : sel_799295;
  assign add_799302 = sel_799299 + 8'h01;
  assign sel_799303 = array_index_799246 == array_index_772720 ? add_799302 : sel_799299;
  assign add_799306 = sel_799303 + 8'h01;
  assign sel_799307 = array_index_799246 == array_index_772726 ? add_799306 : sel_799303;
  assign add_799310 = sel_799307 + 8'h01;
  assign sel_799311 = array_index_799246 == array_index_772732 ? add_799310 : sel_799307;
  assign add_799314 = sel_799311 + 8'h01;
  assign sel_799315 = array_index_799246 == array_index_772738 ? add_799314 : sel_799311;
  assign add_799318 = sel_799315 + 8'h01;
  assign sel_799319 = array_index_799246 == array_index_772744 ? add_799318 : sel_799315;
  assign add_799322 = sel_799319 + 8'h01;
  assign sel_799323 = array_index_799246 == array_index_772750 ? add_799322 : sel_799319;
  assign add_799326 = sel_799323 + 8'h01;
  assign sel_799327 = array_index_799246 == array_index_772756 ? add_799326 : sel_799323;
  assign add_799330 = sel_799327 + 8'h01;
  assign sel_799331 = array_index_799246 == array_index_772762 ? add_799330 : sel_799327;
  assign add_799334 = sel_799331 + 8'h01;
  assign sel_799335 = array_index_799246 == array_index_772768 ? add_799334 : sel_799331;
  assign add_799338 = sel_799335 + 8'h01;
  assign sel_799339 = array_index_799246 == array_index_772774 ? add_799338 : sel_799335;
  assign add_799342 = sel_799339 + 8'h01;
  assign sel_799343 = array_index_799246 == array_index_772780 ? add_799342 : sel_799339;
  assign add_799346 = sel_799343 + 8'h01;
  assign sel_799347 = array_index_799246 == array_index_772786 ? add_799346 : sel_799343;
  assign add_799350 = sel_799347 + 8'h01;
  assign sel_799351 = array_index_799246 == array_index_772792 ? add_799350 : sel_799347;
  assign add_799354 = sel_799351 + 8'h01;
  assign sel_799355 = array_index_799246 == array_index_772798 ? add_799354 : sel_799351;
  assign add_799358 = sel_799355 + 8'h01;
  assign sel_799359 = array_index_799246 == array_index_772804 ? add_799358 : sel_799355;
  assign add_799362 = sel_799359 + 8'h01;
  assign sel_799363 = array_index_799246 == array_index_772810 ? add_799362 : sel_799359;
  assign add_799366 = sel_799363 + 8'h01;
  assign sel_799367 = array_index_799246 == array_index_772816 ? add_799366 : sel_799363;
  assign add_799370 = sel_799367 + 8'h01;
  assign sel_799371 = array_index_799246 == array_index_772822 ? add_799370 : sel_799367;
  assign add_799374 = sel_799371 + 8'h01;
  assign sel_799375 = array_index_799246 == array_index_772828 ? add_799374 : sel_799371;
  assign add_799378 = sel_799375 + 8'h01;
  assign sel_799379 = array_index_799246 == array_index_772834 ? add_799378 : sel_799375;
  assign add_799382 = sel_799379 + 8'h01;
  assign sel_799383 = array_index_799246 == array_index_772840 ? add_799382 : sel_799379;
  assign add_799386 = sel_799383 + 8'h01;
  assign sel_799387 = array_index_799246 == array_index_772846 ? add_799386 : sel_799383;
  assign add_799390 = sel_799387 + 8'h01;
  assign sel_799391 = array_index_799246 == array_index_772852 ? add_799390 : sel_799387;
  assign add_799394 = sel_799391 + 8'h01;
  assign sel_799395 = array_index_799246 == array_index_772858 ? add_799394 : sel_799391;
  assign add_799398 = sel_799395 + 8'h01;
  assign sel_799399 = array_index_799246 == array_index_772864 ? add_799398 : sel_799395;
  assign add_799402 = sel_799399 + 8'h01;
  assign sel_799403 = array_index_799246 == array_index_772870 ? add_799402 : sel_799399;
  assign add_799406 = sel_799403 + 8'h01;
  assign sel_799407 = array_index_799246 == array_index_772876 ? add_799406 : sel_799403;
  assign add_799410 = sel_799407 + 8'h01;
  assign sel_799411 = array_index_799246 == array_index_772882 ? add_799410 : sel_799407;
  assign add_799414 = sel_799411 + 8'h01;
  assign sel_799415 = array_index_799246 == array_index_772888 ? add_799414 : sel_799411;
  assign add_799418 = sel_799415 + 8'h01;
  assign sel_799419 = array_index_799246 == array_index_772894 ? add_799418 : sel_799415;
  assign add_799422 = sel_799419 + 8'h01;
  assign sel_799423 = array_index_799246 == array_index_772900 ? add_799422 : sel_799419;
  assign add_799426 = sel_799423 + 8'h01;
  assign sel_799427 = array_index_799246 == array_index_772906 ? add_799426 : sel_799423;
  assign add_799430 = sel_799427 + 8'h01;
  assign sel_799431 = array_index_799246 == array_index_772912 ? add_799430 : sel_799427;
  assign add_799434 = sel_799431 + 8'h01;
  assign sel_799435 = array_index_799246 == array_index_772918 ? add_799434 : sel_799431;
  assign add_799438 = sel_799435 + 8'h01;
  assign sel_799439 = array_index_799246 == array_index_772924 ? add_799438 : sel_799435;
  assign add_799442 = sel_799439 + 8'h01;
  assign sel_799443 = array_index_799246 == array_index_772930 ? add_799442 : sel_799439;
  assign add_799446 = sel_799443 + 8'h01;
  assign sel_799447 = array_index_799246 == array_index_772936 ? add_799446 : sel_799443;
  assign add_799450 = sel_799447 + 8'h01;
  assign sel_799451 = array_index_799246 == array_index_772942 ? add_799450 : sel_799447;
  assign add_799454 = sel_799451 + 8'h01;
  assign sel_799455 = array_index_799246 == array_index_772948 ? add_799454 : sel_799451;
  assign add_799458 = sel_799455 + 8'h01;
  assign sel_799459 = array_index_799246 == array_index_772954 ? add_799458 : sel_799455;
  assign add_799462 = sel_799459 + 8'h01;
  assign sel_799463 = array_index_799246 == array_index_772960 ? add_799462 : sel_799459;
  assign add_799466 = sel_799463 + 8'h01;
  assign sel_799467 = array_index_799246 == array_index_772966 ? add_799466 : sel_799463;
  assign add_799470 = sel_799467 + 8'h01;
  assign sel_799471 = array_index_799246 == array_index_772972 ? add_799470 : sel_799467;
  assign add_799474 = sel_799471 + 8'h01;
  assign sel_799475 = array_index_799246 == array_index_772978 ? add_799474 : sel_799471;
  assign add_799478 = sel_799475 + 8'h01;
  assign sel_799479 = array_index_799246 == array_index_772984 ? add_799478 : sel_799475;
  assign add_799482 = sel_799479 + 8'h01;
  assign sel_799483 = array_index_799246 == array_index_772990 ? add_799482 : sel_799479;
  assign add_799486 = sel_799483 + 8'h01;
  assign sel_799487 = array_index_799246 == array_index_772996 ? add_799486 : sel_799483;
  assign add_799490 = sel_799487 + 8'h01;
  assign sel_799491 = array_index_799246 == array_index_773002 ? add_799490 : sel_799487;
  assign add_799494 = sel_799491 + 8'h01;
  assign sel_799495 = array_index_799246 == array_index_773008 ? add_799494 : sel_799491;
  assign add_799498 = sel_799495 + 8'h01;
  assign sel_799499 = array_index_799246 == array_index_773014 ? add_799498 : sel_799495;
  assign add_799502 = sel_799499 + 8'h01;
  assign sel_799503 = array_index_799246 == array_index_773020 ? add_799502 : sel_799499;
  assign add_799506 = sel_799503 + 8'h01;
  assign sel_799507 = array_index_799246 == array_index_773026 ? add_799506 : sel_799503;
  assign add_799510 = sel_799507 + 8'h01;
  assign sel_799511 = array_index_799246 == array_index_773032 ? add_799510 : sel_799507;
  assign add_799514 = sel_799511 + 8'h01;
  assign sel_799515 = array_index_799246 == array_index_773038 ? add_799514 : sel_799511;
  assign add_799518 = sel_799515 + 8'h01;
  assign sel_799519 = array_index_799246 == array_index_773044 ? add_799518 : sel_799515;
  assign add_799522 = sel_799519 + 8'h01;
  assign sel_799523 = array_index_799246 == array_index_773050 ? add_799522 : sel_799519;
  assign add_799526 = sel_799523 + 8'h01;
  assign sel_799527 = array_index_799246 == array_index_773056 ? add_799526 : sel_799523;
  assign add_799530 = sel_799527 + 8'h01;
  assign sel_799531 = array_index_799246 == array_index_773062 ? add_799530 : sel_799527;
  assign add_799534 = sel_799531 + 8'h01;
  assign sel_799535 = array_index_799246 == array_index_773068 ? add_799534 : sel_799531;
  assign add_799538 = sel_799535 + 8'h01;
  assign sel_799539 = array_index_799246 == array_index_773074 ? add_799538 : sel_799535;
  assign add_799542 = sel_799539 + 8'h01;
  assign sel_799543 = array_index_799246 == array_index_773080 ? add_799542 : sel_799539;
  assign add_799546 = sel_799543 + 8'h01;
  assign sel_799547 = array_index_799246 == array_index_773086 ? add_799546 : sel_799543;
  assign add_799550 = sel_799547 + 8'h01;
  assign sel_799551 = array_index_799246 == array_index_773092 ? add_799550 : sel_799547;
  assign add_799554 = sel_799551 + 8'h01;
  assign sel_799555 = array_index_799246 == array_index_773098 ? add_799554 : sel_799551;
  assign add_799558 = sel_799555 + 8'h01;
  assign sel_799559 = array_index_799246 == array_index_773104 ? add_799558 : sel_799555;
  assign add_799562 = sel_799559 + 8'h01;
  assign sel_799563 = array_index_799246 == array_index_773110 ? add_799562 : sel_799559;
  assign add_799566 = sel_799563 + 8'h01;
  assign sel_799567 = array_index_799246 == array_index_773116 ? add_799566 : sel_799563;
  assign add_799570 = sel_799567 + 8'h01;
  assign sel_799571 = array_index_799246 == array_index_773122 ? add_799570 : sel_799567;
  assign add_799574 = sel_799571 + 8'h01;
  assign sel_799575 = array_index_799246 == array_index_773128 ? add_799574 : sel_799571;
  assign add_799578 = sel_799575 + 8'h01;
  assign sel_799579 = array_index_799246 == array_index_773134 ? add_799578 : sel_799575;
  assign add_799582 = sel_799579 + 8'h01;
  assign sel_799583 = array_index_799246 == array_index_773140 ? add_799582 : sel_799579;
  assign add_799586 = sel_799583 + 8'h01;
  assign sel_799587 = array_index_799246 == array_index_773146 ? add_799586 : sel_799583;
  assign add_799590 = sel_799587 + 8'h01;
  assign sel_799591 = array_index_799246 == array_index_773152 ? add_799590 : sel_799587;
  assign add_799594 = sel_799591 + 8'h01;
  assign sel_799595 = array_index_799246 == array_index_773158 ? add_799594 : sel_799591;
  assign add_799598 = sel_799595 + 8'h01;
  assign sel_799599 = array_index_799246 == array_index_773164 ? add_799598 : sel_799595;
  assign add_799602 = sel_799599 + 8'h01;
  assign sel_799603 = array_index_799246 == array_index_773170 ? add_799602 : sel_799599;
  assign add_799607 = sel_799603 + 8'h01;
  assign array_index_799608 = set1_unflattened[7'h4a];
  assign sel_799609 = array_index_799246 == array_index_773176 ? add_799607 : sel_799603;
  assign add_799612 = sel_799609 + 8'h01;
  assign sel_799613 = array_index_799608 == array_index_772632 ? add_799612 : sel_799609;
  assign add_799616 = sel_799613 + 8'h01;
  assign sel_799617 = array_index_799608 == array_index_772636 ? add_799616 : sel_799613;
  assign add_799620 = sel_799617 + 8'h01;
  assign sel_799621 = array_index_799608 == array_index_772644 ? add_799620 : sel_799617;
  assign add_799624 = sel_799621 + 8'h01;
  assign sel_799625 = array_index_799608 == array_index_772652 ? add_799624 : sel_799621;
  assign add_799628 = sel_799625 + 8'h01;
  assign sel_799629 = array_index_799608 == array_index_772660 ? add_799628 : sel_799625;
  assign add_799632 = sel_799629 + 8'h01;
  assign sel_799633 = array_index_799608 == array_index_772668 ? add_799632 : sel_799629;
  assign add_799636 = sel_799633 + 8'h01;
  assign sel_799637 = array_index_799608 == array_index_772676 ? add_799636 : sel_799633;
  assign add_799640 = sel_799637 + 8'h01;
  assign sel_799641 = array_index_799608 == array_index_772684 ? add_799640 : sel_799637;
  assign add_799644 = sel_799641 + 8'h01;
  assign sel_799645 = array_index_799608 == array_index_772690 ? add_799644 : sel_799641;
  assign add_799648 = sel_799645 + 8'h01;
  assign sel_799649 = array_index_799608 == array_index_772696 ? add_799648 : sel_799645;
  assign add_799652 = sel_799649 + 8'h01;
  assign sel_799653 = array_index_799608 == array_index_772702 ? add_799652 : sel_799649;
  assign add_799656 = sel_799653 + 8'h01;
  assign sel_799657 = array_index_799608 == array_index_772708 ? add_799656 : sel_799653;
  assign add_799660 = sel_799657 + 8'h01;
  assign sel_799661 = array_index_799608 == array_index_772714 ? add_799660 : sel_799657;
  assign add_799664 = sel_799661 + 8'h01;
  assign sel_799665 = array_index_799608 == array_index_772720 ? add_799664 : sel_799661;
  assign add_799668 = sel_799665 + 8'h01;
  assign sel_799669 = array_index_799608 == array_index_772726 ? add_799668 : sel_799665;
  assign add_799672 = sel_799669 + 8'h01;
  assign sel_799673 = array_index_799608 == array_index_772732 ? add_799672 : sel_799669;
  assign add_799676 = sel_799673 + 8'h01;
  assign sel_799677 = array_index_799608 == array_index_772738 ? add_799676 : sel_799673;
  assign add_799680 = sel_799677 + 8'h01;
  assign sel_799681 = array_index_799608 == array_index_772744 ? add_799680 : sel_799677;
  assign add_799684 = sel_799681 + 8'h01;
  assign sel_799685 = array_index_799608 == array_index_772750 ? add_799684 : sel_799681;
  assign add_799688 = sel_799685 + 8'h01;
  assign sel_799689 = array_index_799608 == array_index_772756 ? add_799688 : sel_799685;
  assign add_799692 = sel_799689 + 8'h01;
  assign sel_799693 = array_index_799608 == array_index_772762 ? add_799692 : sel_799689;
  assign add_799696 = sel_799693 + 8'h01;
  assign sel_799697 = array_index_799608 == array_index_772768 ? add_799696 : sel_799693;
  assign add_799700 = sel_799697 + 8'h01;
  assign sel_799701 = array_index_799608 == array_index_772774 ? add_799700 : sel_799697;
  assign add_799704 = sel_799701 + 8'h01;
  assign sel_799705 = array_index_799608 == array_index_772780 ? add_799704 : sel_799701;
  assign add_799708 = sel_799705 + 8'h01;
  assign sel_799709 = array_index_799608 == array_index_772786 ? add_799708 : sel_799705;
  assign add_799712 = sel_799709 + 8'h01;
  assign sel_799713 = array_index_799608 == array_index_772792 ? add_799712 : sel_799709;
  assign add_799716 = sel_799713 + 8'h01;
  assign sel_799717 = array_index_799608 == array_index_772798 ? add_799716 : sel_799713;
  assign add_799720 = sel_799717 + 8'h01;
  assign sel_799721 = array_index_799608 == array_index_772804 ? add_799720 : sel_799717;
  assign add_799724 = sel_799721 + 8'h01;
  assign sel_799725 = array_index_799608 == array_index_772810 ? add_799724 : sel_799721;
  assign add_799728 = sel_799725 + 8'h01;
  assign sel_799729 = array_index_799608 == array_index_772816 ? add_799728 : sel_799725;
  assign add_799732 = sel_799729 + 8'h01;
  assign sel_799733 = array_index_799608 == array_index_772822 ? add_799732 : sel_799729;
  assign add_799736 = sel_799733 + 8'h01;
  assign sel_799737 = array_index_799608 == array_index_772828 ? add_799736 : sel_799733;
  assign add_799740 = sel_799737 + 8'h01;
  assign sel_799741 = array_index_799608 == array_index_772834 ? add_799740 : sel_799737;
  assign add_799744 = sel_799741 + 8'h01;
  assign sel_799745 = array_index_799608 == array_index_772840 ? add_799744 : sel_799741;
  assign add_799748 = sel_799745 + 8'h01;
  assign sel_799749 = array_index_799608 == array_index_772846 ? add_799748 : sel_799745;
  assign add_799752 = sel_799749 + 8'h01;
  assign sel_799753 = array_index_799608 == array_index_772852 ? add_799752 : sel_799749;
  assign add_799756 = sel_799753 + 8'h01;
  assign sel_799757 = array_index_799608 == array_index_772858 ? add_799756 : sel_799753;
  assign add_799760 = sel_799757 + 8'h01;
  assign sel_799761 = array_index_799608 == array_index_772864 ? add_799760 : sel_799757;
  assign add_799764 = sel_799761 + 8'h01;
  assign sel_799765 = array_index_799608 == array_index_772870 ? add_799764 : sel_799761;
  assign add_799768 = sel_799765 + 8'h01;
  assign sel_799769 = array_index_799608 == array_index_772876 ? add_799768 : sel_799765;
  assign add_799772 = sel_799769 + 8'h01;
  assign sel_799773 = array_index_799608 == array_index_772882 ? add_799772 : sel_799769;
  assign add_799776 = sel_799773 + 8'h01;
  assign sel_799777 = array_index_799608 == array_index_772888 ? add_799776 : sel_799773;
  assign add_799780 = sel_799777 + 8'h01;
  assign sel_799781 = array_index_799608 == array_index_772894 ? add_799780 : sel_799777;
  assign add_799784 = sel_799781 + 8'h01;
  assign sel_799785 = array_index_799608 == array_index_772900 ? add_799784 : sel_799781;
  assign add_799788 = sel_799785 + 8'h01;
  assign sel_799789 = array_index_799608 == array_index_772906 ? add_799788 : sel_799785;
  assign add_799792 = sel_799789 + 8'h01;
  assign sel_799793 = array_index_799608 == array_index_772912 ? add_799792 : sel_799789;
  assign add_799796 = sel_799793 + 8'h01;
  assign sel_799797 = array_index_799608 == array_index_772918 ? add_799796 : sel_799793;
  assign add_799800 = sel_799797 + 8'h01;
  assign sel_799801 = array_index_799608 == array_index_772924 ? add_799800 : sel_799797;
  assign add_799804 = sel_799801 + 8'h01;
  assign sel_799805 = array_index_799608 == array_index_772930 ? add_799804 : sel_799801;
  assign add_799808 = sel_799805 + 8'h01;
  assign sel_799809 = array_index_799608 == array_index_772936 ? add_799808 : sel_799805;
  assign add_799812 = sel_799809 + 8'h01;
  assign sel_799813 = array_index_799608 == array_index_772942 ? add_799812 : sel_799809;
  assign add_799816 = sel_799813 + 8'h01;
  assign sel_799817 = array_index_799608 == array_index_772948 ? add_799816 : sel_799813;
  assign add_799820 = sel_799817 + 8'h01;
  assign sel_799821 = array_index_799608 == array_index_772954 ? add_799820 : sel_799817;
  assign add_799824 = sel_799821 + 8'h01;
  assign sel_799825 = array_index_799608 == array_index_772960 ? add_799824 : sel_799821;
  assign add_799828 = sel_799825 + 8'h01;
  assign sel_799829 = array_index_799608 == array_index_772966 ? add_799828 : sel_799825;
  assign add_799832 = sel_799829 + 8'h01;
  assign sel_799833 = array_index_799608 == array_index_772972 ? add_799832 : sel_799829;
  assign add_799836 = sel_799833 + 8'h01;
  assign sel_799837 = array_index_799608 == array_index_772978 ? add_799836 : sel_799833;
  assign add_799840 = sel_799837 + 8'h01;
  assign sel_799841 = array_index_799608 == array_index_772984 ? add_799840 : sel_799837;
  assign add_799844 = sel_799841 + 8'h01;
  assign sel_799845 = array_index_799608 == array_index_772990 ? add_799844 : sel_799841;
  assign add_799848 = sel_799845 + 8'h01;
  assign sel_799849 = array_index_799608 == array_index_772996 ? add_799848 : sel_799845;
  assign add_799852 = sel_799849 + 8'h01;
  assign sel_799853 = array_index_799608 == array_index_773002 ? add_799852 : sel_799849;
  assign add_799856 = sel_799853 + 8'h01;
  assign sel_799857 = array_index_799608 == array_index_773008 ? add_799856 : sel_799853;
  assign add_799860 = sel_799857 + 8'h01;
  assign sel_799861 = array_index_799608 == array_index_773014 ? add_799860 : sel_799857;
  assign add_799864 = sel_799861 + 8'h01;
  assign sel_799865 = array_index_799608 == array_index_773020 ? add_799864 : sel_799861;
  assign add_799868 = sel_799865 + 8'h01;
  assign sel_799869 = array_index_799608 == array_index_773026 ? add_799868 : sel_799865;
  assign add_799872 = sel_799869 + 8'h01;
  assign sel_799873 = array_index_799608 == array_index_773032 ? add_799872 : sel_799869;
  assign add_799876 = sel_799873 + 8'h01;
  assign sel_799877 = array_index_799608 == array_index_773038 ? add_799876 : sel_799873;
  assign add_799880 = sel_799877 + 8'h01;
  assign sel_799881 = array_index_799608 == array_index_773044 ? add_799880 : sel_799877;
  assign add_799884 = sel_799881 + 8'h01;
  assign sel_799885 = array_index_799608 == array_index_773050 ? add_799884 : sel_799881;
  assign add_799888 = sel_799885 + 8'h01;
  assign sel_799889 = array_index_799608 == array_index_773056 ? add_799888 : sel_799885;
  assign add_799892 = sel_799889 + 8'h01;
  assign sel_799893 = array_index_799608 == array_index_773062 ? add_799892 : sel_799889;
  assign add_799896 = sel_799893 + 8'h01;
  assign sel_799897 = array_index_799608 == array_index_773068 ? add_799896 : sel_799893;
  assign add_799900 = sel_799897 + 8'h01;
  assign sel_799901 = array_index_799608 == array_index_773074 ? add_799900 : sel_799897;
  assign add_799904 = sel_799901 + 8'h01;
  assign sel_799905 = array_index_799608 == array_index_773080 ? add_799904 : sel_799901;
  assign add_799908 = sel_799905 + 8'h01;
  assign sel_799909 = array_index_799608 == array_index_773086 ? add_799908 : sel_799905;
  assign add_799912 = sel_799909 + 8'h01;
  assign sel_799913 = array_index_799608 == array_index_773092 ? add_799912 : sel_799909;
  assign add_799916 = sel_799913 + 8'h01;
  assign sel_799917 = array_index_799608 == array_index_773098 ? add_799916 : sel_799913;
  assign add_799920 = sel_799917 + 8'h01;
  assign sel_799921 = array_index_799608 == array_index_773104 ? add_799920 : sel_799917;
  assign add_799924 = sel_799921 + 8'h01;
  assign sel_799925 = array_index_799608 == array_index_773110 ? add_799924 : sel_799921;
  assign add_799928 = sel_799925 + 8'h01;
  assign sel_799929 = array_index_799608 == array_index_773116 ? add_799928 : sel_799925;
  assign add_799932 = sel_799929 + 8'h01;
  assign sel_799933 = array_index_799608 == array_index_773122 ? add_799932 : sel_799929;
  assign add_799936 = sel_799933 + 8'h01;
  assign sel_799937 = array_index_799608 == array_index_773128 ? add_799936 : sel_799933;
  assign add_799940 = sel_799937 + 8'h01;
  assign sel_799941 = array_index_799608 == array_index_773134 ? add_799940 : sel_799937;
  assign add_799944 = sel_799941 + 8'h01;
  assign sel_799945 = array_index_799608 == array_index_773140 ? add_799944 : sel_799941;
  assign add_799948 = sel_799945 + 8'h01;
  assign sel_799949 = array_index_799608 == array_index_773146 ? add_799948 : sel_799945;
  assign add_799952 = sel_799949 + 8'h01;
  assign sel_799953 = array_index_799608 == array_index_773152 ? add_799952 : sel_799949;
  assign add_799956 = sel_799953 + 8'h01;
  assign sel_799957 = array_index_799608 == array_index_773158 ? add_799956 : sel_799953;
  assign add_799960 = sel_799957 + 8'h01;
  assign sel_799961 = array_index_799608 == array_index_773164 ? add_799960 : sel_799957;
  assign add_799964 = sel_799961 + 8'h01;
  assign sel_799965 = array_index_799608 == array_index_773170 ? add_799964 : sel_799961;
  assign add_799969 = sel_799965 + 8'h01;
  assign array_index_799970 = set1_unflattened[7'h4b];
  assign sel_799971 = array_index_799608 == array_index_773176 ? add_799969 : sel_799965;
  assign add_799974 = sel_799971 + 8'h01;
  assign sel_799975 = array_index_799970 == array_index_772632 ? add_799974 : sel_799971;
  assign add_799978 = sel_799975 + 8'h01;
  assign sel_799979 = array_index_799970 == array_index_772636 ? add_799978 : sel_799975;
  assign add_799982 = sel_799979 + 8'h01;
  assign sel_799983 = array_index_799970 == array_index_772644 ? add_799982 : sel_799979;
  assign add_799986 = sel_799983 + 8'h01;
  assign sel_799987 = array_index_799970 == array_index_772652 ? add_799986 : sel_799983;
  assign add_799990 = sel_799987 + 8'h01;
  assign sel_799991 = array_index_799970 == array_index_772660 ? add_799990 : sel_799987;
  assign add_799994 = sel_799991 + 8'h01;
  assign sel_799995 = array_index_799970 == array_index_772668 ? add_799994 : sel_799991;
  assign add_799998 = sel_799995 + 8'h01;
  assign sel_799999 = array_index_799970 == array_index_772676 ? add_799998 : sel_799995;
  assign add_800002 = sel_799999 + 8'h01;
  assign sel_800003 = array_index_799970 == array_index_772684 ? add_800002 : sel_799999;
  assign add_800006 = sel_800003 + 8'h01;
  assign sel_800007 = array_index_799970 == array_index_772690 ? add_800006 : sel_800003;
  assign add_800010 = sel_800007 + 8'h01;
  assign sel_800011 = array_index_799970 == array_index_772696 ? add_800010 : sel_800007;
  assign add_800014 = sel_800011 + 8'h01;
  assign sel_800015 = array_index_799970 == array_index_772702 ? add_800014 : sel_800011;
  assign add_800018 = sel_800015 + 8'h01;
  assign sel_800019 = array_index_799970 == array_index_772708 ? add_800018 : sel_800015;
  assign add_800022 = sel_800019 + 8'h01;
  assign sel_800023 = array_index_799970 == array_index_772714 ? add_800022 : sel_800019;
  assign add_800026 = sel_800023 + 8'h01;
  assign sel_800027 = array_index_799970 == array_index_772720 ? add_800026 : sel_800023;
  assign add_800030 = sel_800027 + 8'h01;
  assign sel_800031 = array_index_799970 == array_index_772726 ? add_800030 : sel_800027;
  assign add_800034 = sel_800031 + 8'h01;
  assign sel_800035 = array_index_799970 == array_index_772732 ? add_800034 : sel_800031;
  assign add_800038 = sel_800035 + 8'h01;
  assign sel_800039 = array_index_799970 == array_index_772738 ? add_800038 : sel_800035;
  assign add_800042 = sel_800039 + 8'h01;
  assign sel_800043 = array_index_799970 == array_index_772744 ? add_800042 : sel_800039;
  assign add_800046 = sel_800043 + 8'h01;
  assign sel_800047 = array_index_799970 == array_index_772750 ? add_800046 : sel_800043;
  assign add_800050 = sel_800047 + 8'h01;
  assign sel_800051 = array_index_799970 == array_index_772756 ? add_800050 : sel_800047;
  assign add_800054 = sel_800051 + 8'h01;
  assign sel_800055 = array_index_799970 == array_index_772762 ? add_800054 : sel_800051;
  assign add_800058 = sel_800055 + 8'h01;
  assign sel_800059 = array_index_799970 == array_index_772768 ? add_800058 : sel_800055;
  assign add_800062 = sel_800059 + 8'h01;
  assign sel_800063 = array_index_799970 == array_index_772774 ? add_800062 : sel_800059;
  assign add_800066 = sel_800063 + 8'h01;
  assign sel_800067 = array_index_799970 == array_index_772780 ? add_800066 : sel_800063;
  assign add_800070 = sel_800067 + 8'h01;
  assign sel_800071 = array_index_799970 == array_index_772786 ? add_800070 : sel_800067;
  assign add_800074 = sel_800071 + 8'h01;
  assign sel_800075 = array_index_799970 == array_index_772792 ? add_800074 : sel_800071;
  assign add_800078 = sel_800075 + 8'h01;
  assign sel_800079 = array_index_799970 == array_index_772798 ? add_800078 : sel_800075;
  assign add_800082 = sel_800079 + 8'h01;
  assign sel_800083 = array_index_799970 == array_index_772804 ? add_800082 : sel_800079;
  assign add_800086 = sel_800083 + 8'h01;
  assign sel_800087 = array_index_799970 == array_index_772810 ? add_800086 : sel_800083;
  assign add_800090 = sel_800087 + 8'h01;
  assign sel_800091 = array_index_799970 == array_index_772816 ? add_800090 : sel_800087;
  assign add_800094 = sel_800091 + 8'h01;
  assign sel_800095 = array_index_799970 == array_index_772822 ? add_800094 : sel_800091;
  assign add_800098 = sel_800095 + 8'h01;
  assign sel_800099 = array_index_799970 == array_index_772828 ? add_800098 : sel_800095;
  assign add_800102 = sel_800099 + 8'h01;
  assign sel_800103 = array_index_799970 == array_index_772834 ? add_800102 : sel_800099;
  assign add_800106 = sel_800103 + 8'h01;
  assign sel_800107 = array_index_799970 == array_index_772840 ? add_800106 : sel_800103;
  assign add_800110 = sel_800107 + 8'h01;
  assign sel_800111 = array_index_799970 == array_index_772846 ? add_800110 : sel_800107;
  assign add_800114 = sel_800111 + 8'h01;
  assign sel_800115 = array_index_799970 == array_index_772852 ? add_800114 : sel_800111;
  assign add_800118 = sel_800115 + 8'h01;
  assign sel_800119 = array_index_799970 == array_index_772858 ? add_800118 : sel_800115;
  assign add_800122 = sel_800119 + 8'h01;
  assign sel_800123 = array_index_799970 == array_index_772864 ? add_800122 : sel_800119;
  assign add_800126 = sel_800123 + 8'h01;
  assign sel_800127 = array_index_799970 == array_index_772870 ? add_800126 : sel_800123;
  assign add_800130 = sel_800127 + 8'h01;
  assign sel_800131 = array_index_799970 == array_index_772876 ? add_800130 : sel_800127;
  assign add_800134 = sel_800131 + 8'h01;
  assign sel_800135 = array_index_799970 == array_index_772882 ? add_800134 : sel_800131;
  assign add_800138 = sel_800135 + 8'h01;
  assign sel_800139 = array_index_799970 == array_index_772888 ? add_800138 : sel_800135;
  assign add_800142 = sel_800139 + 8'h01;
  assign sel_800143 = array_index_799970 == array_index_772894 ? add_800142 : sel_800139;
  assign add_800146 = sel_800143 + 8'h01;
  assign sel_800147 = array_index_799970 == array_index_772900 ? add_800146 : sel_800143;
  assign add_800150 = sel_800147 + 8'h01;
  assign sel_800151 = array_index_799970 == array_index_772906 ? add_800150 : sel_800147;
  assign add_800154 = sel_800151 + 8'h01;
  assign sel_800155 = array_index_799970 == array_index_772912 ? add_800154 : sel_800151;
  assign add_800158 = sel_800155 + 8'h01;
  assign sel_800159 = array_index_799970 == array_index_772918 ? add_800158 : sel_800155;
  assign add_800162 = sel_800159 + 8'h01;
  assign sel_800163 = array_index_799970 == array_index_772924 ? add_800162 : sel_800159;
  assign add_800166 = sel_800163 + 8'h01;
  assign sel_800167 = array_index_799970 == array_index_772930 ? add_800166 : sel_800163;
  assign add_800170 = sel_800167 + 8'h01;
  assign sel_800171 = array_index_799970 == array_index_772936 ? add_800170 : sel_800167;
  assign add_800174 = sel_800171 + 8'h01;
  assign sel_800175 = array_index_799970 == array_index_772942 ? add_800174 : sel_800171;
  assign add_800178 = sel_800175 + 8'h01;
  assign sel_800179 = array_index_799970 == array_index_772948 ? add_800178 : sel_800175;
  assign add_800182 = sel_800179 + 8'h01;
  assign sel_800183 = array_index_799970 == array_index_772954 ? add_800182 : sel_800179;
  assign add_800186 = sel_800183 + 8'h01;
  assign sel_800187 = array_index_799970 == array_index_772960 ? add_800186 : sel_800183;
  assign add_800190 = sel_800187 + 8'h01;
  assign sel_800191 = array_index_799970 == array_index_772966 ? add_800190 : sel_800187;
  assign add_800194 = sel_800191 + 8'h01;
  assign sel_800195 = array_index_799970 == array_index_772972 ? add_800194 : sel_800191;
  assign add_800198 = sel_800195 + 8'h01;
  assign sel_800199 = array_index_799970 == array_index_772978 ? add_800198 : sel_800195;
  assign add_800202 = sel_800199 + 8'h01;
  assign sel_800203 = array_index_799970 == array_index_772984 ? add_800202 : sel_800199;
  assign add_800206 = sel_800203 + 8'h01;
  assign sel_800207 = array_index_799970 == array_index_772990 ? add_800206 : sel_800203;
  assign add_800210 = sel_800207 + 8'h01;
  assign sel_800211 = array_index_799970 == array_index_772996 ? add_800210 : sel_800207;
  assign add_800214 = sel_800211 + 8'h01;
  assign sel_800215 = array_index_799970 == array_index_773002 ? add_800214 : sel_800211;
  assign add_800218 = sel_800215 + 8'h01;
  assign sel_800219 = array_index_799970 == array_index_773008 ? add_800218 : sel_800215;
  assign add_800222 = sel_800219 + 8'h01;
  assign sel_800223 = array_index_799970 == array_index_773014 ? add_800222 : sel_800219;
  assign add_800226 = sel_800223 + 8'h01;
  assign sel_800227 = array_index_799970 == array_index_773020 ? add_800226 : sel_800223;
  assign add_800230 = sel_800227 + 8'h01;
  assign sel_800231 = array_index_799970 == array_index_773026 ? add_800230 : sel_800227;
  assign add_800234 = sel_800231 + 8'h01;
  assign sel_800235 = array_index_799970 == array_index_773032 ? add_800234 : sel_800231;
  assign add_800238 = sel_800235 + 8'h01;
  assign sel_800239 = array_index_799970 == array_index_773038 ? add_800238 : sel_800235;
  assign add_800242 = sel_800239 + 8'h01;
  assign sel_800243 = array_index_799970 == array_index_773044 ? add_800242 : sel_800239;
  assign add_800246 = sel_800243 + 8'h01;
  assign sel_800247 = array_index_799970 == array_index_773050 ? add_800246 : sel_800243;
  assign add_800250 = sel_800247 + 8'h01;
  assign sel_800251 = array_index_799970 == array_index_773056 ? add_800250 : sel_800247;
  assign add_800254 = sel_800251 + 8'h01;
  assign sel_800255 = array_index_799970 == array_index_773062 ? add_800254 : sel_800251;
  assign add_800258 = sel_800255 + 8'h01;
  assign sel_800259 = array_index_799970 == array_index_773068 ? add_800258 : sel_800255;
  assign add_800262 = sel_800259 + 8'h01;
  assign sel_800263 = array_index_799970 == array_index_773074 ? add_800262 : sel_800259;
  assign add_800266 = sel_800263 + 8'h01;
  assign sel_800267 = array_index_799970 == array_index_773080 ? add_800266 : sel_800263;
  assign add_800270 = sel_800267 + 8'h01;
  assign sel_800271 = array_index_799970 == array_index_773086 ? add_800270 : sel_800267;
  assign add_800274 = sel_800271 + 8'h01;
  assign sel_800275 = array_index_799970 == array_index_773092 ? add_800274 : sel_800271;
  assign add_800278 = sel_800275 + 8'h01;
  assign sel_800279 = array_index_799970 == array_index_773098 ? add_800278 : sel_800275;
  assign add_800282 = sel_800279 + 8'h01;
  assign sel_800283 = array_index_799970 == array_index_773104 ? add_800282 : sel_800279;
  assign add_800286 = sel_800283 + 8'h01;
  assign sel_800287 = array_index_799970 == array_index_773110 ? add_800286 : sel_800283;
  assign add_800290 = sel_800287 + 8'h01;
  assign sel_800291 = array_index_799970 == array_index_773116 ? add_800290 : sel_800287;
  assign add_800294 = sel_800291 + 8'h01;
  assign sel_800295 = array_index_799970 == array_index_773122 ? add_800294 : sel_800291;
  assign add_800298 = sel_800295 + 8'h01;
  assign sel_800299 = array_index_799970 == array_index_773128 ? add_800298 : sel_800295;
  assign add_800302 = sel_800299 + 8'h01;
  assign sel_800303 = array_index_799970 == array_index_773134 ? add_800302 : sel_800299;
  assign add_800306 = sel_800303 + 8'h01;
  assign sel_800307 = array_index_799970 == array_index_773140 ? add_800306 : sel_800303;
  assign add_800310 = sel_800307 + 8'h01;
  assign sel_800311 = array_index_799970 == array_index_773146 ? add_800310 : sel_800307;
  assign add_800314 = sel_800311 + 8'h01;
  assign sel_800315 = array_index_799970 == array_index_773152 ? add_800314 : sel_800311;
  assign add_800318 = sel_800315 + 8'h01;
  assign sel_800319 = array_index_799970 == array_index_773158 ? add_800318 : sel_800315;
  assign add_800322 = sel_800319 + 8'h01;
  assign sel_800323 = array_index_799970 == array_index_773164 ? add_800322 : sel_800319;
  assign add_800326 = sel_800323 + 8'h01;
  assign sel_800327 = array_index_799970 == array_index_773170 ? add_800326 : sel_800323;
  assign add_800331 = sel_800327 + 8'h01;
  assign array_index_800332 = set1_unflattened[7'h4c];
  assign sel_800333 = array_index_799970 == array_index_773176 ? add_800331 : sel_800327;
  assign add_800336 = sel_800333 + 8'h01;
  assign sel_800337 = array_index_800332 == array_index_772632 ? add_800336 : sel_800333;
  assign add_800340 = sel_800337 + 8'h01;
  assign sel_800341 = array_index_800332 == array_index_772636 ? add_800340 : sel_800337;
  assign add_800344 = sel_800341 + 8'h01;
  assign sel_800345 = array_index_800332 == array_index_772644 ? add_800344 : sel_800341;
  assign add_800348 = sel_800345 + 8'h01;
  assign sel_800349 = array_index_800332 == array_index_772652 ? add_800348 : sel_800345;
  assign add_800352 = sel_800349 + 8'h01;
  assign sel_800353 = array_index_800332 == array_index_772660 ? add_800352 : sel_800349;
  assign add_800356 = sel_800353 + 8'h01;
  assign sel_800357 = array_index_800332 == array_index_772668 ? add_800356 : sel_800353;
  assign add_800360 = sel_800357 + 8'h01;
  assign sel_800361 = array_index_800332 == array_index_772676 ? add_800360 : sel_800357;
  assign add_800364 = sel_800361 + 8'h01;
  assign sel_800365 = array_index_800332 == array_index_772684 ? add_800364 : sel_800361;
  assign add_800368 = sel_800365 + 8'h01;
  assign sel_800369 = array_index_800332 == array_index_772690 ? add_800368 : sel_800365;
  assign add_800372 = sel_800369 + 8'h01;
  assign sel_800373 = array_index_800332 == array_index_772696 ? add_800372 : sel_800369;
  assign add_800376 = sel_800373 + 8'h01;
  assign sel_800377 = array_index_800332 == array_index_772702 ? add_800376 : sel_800373;
  assign add_800380 = sel_800377 + 8'h01;
  assign sel_800381 = array_index_800332 == array_index_772708 ? add_800380 : sel_800377;
  assign add_800384 = sel_800381 + 8'h01;
  assign sel_800385 = array_index_800332 == array_index_772714 ? add_800384 : sel_800381;
  assign add_800388 = sel_800385 + 8'h01;
  assign sel_800389 = array_index_800332 == array_index_772720 ? add_800388 : sel_800385;
  assign add_800392 = sel_800389 + 8'h01;
  assign sel_800393 = array_index_800332 == array_index_772726 ? add_800392 : sel_800389;
  assign add_800396 = sel_800393 + 8'h01;
  assign sel_800397 = array_index_800332 == array_index_772732 ? add_800396 : sel_800393;
  assign add_800400 = sel_800397 + 8'h01;
  assign sel_800401 = array_index_800332 == array_index_772738 ? add_800400 : sel_800397;
  assign add_800404 = sel_800401 + 8'h01;
  assign sel_800405 = array_index_800332 == array_index_772744 ? add_800404 : sel_800401;
  assign add_800408 = sel_800405 + 8'h01;
  assign sel_800409 = array_index_800332 == array_index_772750 ? add_800408 : sel_800405;
  assign add_800412 = sel_800409 + 8'h01;
  assign sel_800413 = array_index_800332 == array_index_772756 ? add_800412 : sel_800409;
  assign add_800416 = sel_800413 + 8'h01;
  assign sel_800417 = array_index_800332 == array_index_772762 ? add_800416 : sel_800413;
  assign add_800420 = sel_800417 + 8'h01;
  assign sel_800421 = array_index_800332 == array_index_772768 ? add_800420 : sel_800417;
  assign add_800424 = sel_800421 + 8'h01;
  assign sel_800425 = array_index_800332 == array_index_772774 ? add_800424 : sel_800421;
  assign add_800428 = sel_800425 + 8'h01;
  assign sel_800429 = array_index_800332 == array_index_772780 ? add_800428 : sel_800425;
  assign add_800432 = sel_800429 + 8'h01;
  assign sel_800433 = array_index_800332 == array_index_772786 ? add_800432 : sel_800429;
  assign add_800436 = sel_800433 + 8'h01;
  assign sel_800437 = array_index_800332 == array_index_772792 ? add_800436 : sel_800433;
  assign add_800440 = sel_800437 + 8'h01;
  assign sel_800441 = array_index_800332 == array_index_772798 ? add_800440 : sel_800437;
  assign add_800444 = sel_800441 + 8'h01;
  assign sel_800445 = array_index_800332 == array_index_772804 ? add_800444 : sel_800441;
  assign add_800448 = sel_800445 + 8'h01;
  assign sel_800449 = array_index_800332 == array_index_772810 ? add_800448 : sel_800445;
  assign add_800452 = sel_800449 + 8'h01;
  assign sel_800453 = array_index_800332 == array_index_772816 ? add_800452 : sel_800449;
  assign add_800456 = sel_800453 + 8'h01;
  assign sel_800457 = array_index_800332 == array_index_772822 ? add_800456 : sel_800453;
  assign add_800460 = sel_800457 + 8'h01;
  assign sel_800461 = array_index_800332 == array_index_772828 ? add_800460 : sel_800457;
  assign add_800464 = sel_800461 + 8'h01;
  assign sel_800465 = array_index_800332 == array_index_772834 ? add_800464 : sel_800461;
  assign add_800468 = sel_800465 + 8'h01;
  assign sel_800469 = array_index_800332 == array_index_772840 ? add_800468 : sel_800465;
  assign add_800472 = sel_800469 + 8'h01;
  assign sel_800473 = array_index_800332 == array_index_772846 ? add_800472 : sel_800469;
  assign add_800476 = sel_800473 + 8'h01;
  assign sel_800477 = array_index_800332 == array_index_772852 ? add_800476 : sel_800473;
  assign add_800480 = sel_800477 + 8'h01;
  assign sel_800481 = array_index_800332 == array_index_772858 ? add_800480 : sel_800477;
  assign add_800484 = sel_800481 + 8'h01;
  assign sel_800485 = array_index_800332 == array_index_772864 ? add_800484 : sel_800481;
  assign add_800488 = sel_800485 + 8'h01;
  assign sel_800489 = array_index_800332 == array_index_772870 ? add_800488 : sel_800485;
  assign add_800492 = sel_800489 + 8'h01;
  assign sel_800493 = array_index_800332 == array_index_772876 ? add_800492 : sel_800489;
  assign add_800496 = sel_800493 + 8'h01;
  assign sel_800497 = array_index_800332 == array_index_772882 ? add_800496 : sel_800493;
  assign add_800500 = sel_800497 + 8'h01;
  assign sel_800501 = array_index_800332 == array_index_772888 ? add_800500 : sel_800497;
  assign add_800504 = sel_800501 + 8'h01;
  assign sel_800505 = array_index_800332 == array_index_772894 ? add_800504 : sel_800501;
  assign add_800508 = sel_800505 + 8'h01;
  assign sel_800509 = array_index_800332 == array_index_772900 ? add_800508 : sel_800505;
  assign add_800512 = sel_800509 + 8'h01;
  assign sel_800513 = array_index_800332 == array_index_772906 ? add_800512 : sel_800509;
  assign add_800516 = sel_800513 + 8'h01;
  assign sel_800517 = array_index_800332 == array_index_772912 ? add_800516 : sel_800513;
  assign add_800520 = sel_800517 + 8'h01;
  assign sel_800521 = array_index_800332 == array_index_772918 ? add_800520 : sel_800517;
  assign add_800524 = sel_800521 + 8'h01;
  assign sel_800525 = array_index_800332 == array_index_772924 ? add_800524 : sel_800521;
  assign add_800528 = sel_800525 + 8'h01;
  assign sel_800529 = array_index_800332 == array_index_772930 ? add_800528 : sel_800525;
  assign add_800532 = sel_800529 + 8'h01;
  assign sel_800533 = array_index_800332 == array_index_772936 ? add_800532 : sel_800529;
  assign add_800536 = sel_800533 + 8'h01;
  assign sel_800537 = array_index_800332 == array_index_772942 ? add_800536 : sel_800533;
  assign add_800540 = sel_800537 + 8'h01;
  assign sel_800541 = array_index_800332 == array_index_772948 ? add_800540 : sel_800537;
  assign add_800544 = sel_800541 + 8'h01;
  assign sel_800545 = array_index_800332 == array_index_772954 ? add_800544 : sel_800541;
  assign add_800548 = sel_800545 + 8'h01;
  assign sel_800549 = array_index_800332 == array_index_772960 ? add_800548 : sel_800545;
  assign add_800552 = sel_800549 + 8'h01;
  assign sel_800553 = array_index_800332 == array_index_772966 ? add_800552 : sel_800549;
  assign add_800556 = sel_800553 + 8'h01;
  assign sel_800557 = array_index_800332 == array_index_772972 ? add_800556 : sel_800553;
  assign add_800560 = sel_800557 + 8'h01;
  assign sel_800561 = array_index_800332 == array_index_772978 ? add_800560 : sel_800557;
  assign add_800564 = sel_800561 + 8'h01;
  assign sel_800565 = array_index_800332 == array_index_772984 ? add_800564 : sel_800561;
  assign add_800568 = sel_800565 + 8'h01;
  assign sel_800569 = array_index_800332 == array_index_772990 ? add_800568 : sel_800565;
  assign add_800572 = sel_800569 + 8'h01;
  assign sel_800573 = array_index_800332 == array_index_772996 ? add_800572 : sel_800569;
  assign add_800576 = sel_800573 + 8'h01;
  assign sel_800577 = array_index_800332 == array_index_773002 ? add_800576 : sel_800573;
  assign add_800580 = sel_800577 + 8'h01;
  assign sel_800581 = array_index_800332 == array_index_773008 ? add_800580 : sel_800577;
  assign add_800584 = sel_800581 + 8'h01;
  assign sel_800585 = array_index_800332 == array_index_773014 ? add_800584 : sel_800581;
  assign add_800588 = sel_800585 + 8'h01;
  assign sel_800589 = array_index_800332 == array_index_773020 ? add_800588 : sel_800585;
  assign add_800592 = sel_800589 + 8'h01;
  assign sel_800593 = array_index_800332 == array_index_773026 ? add_800592 : sel_800589;
  assign add_800596 = sel_800593 + 8'h01;
  assign sel_800597 = array_index_800332 == array_index_773032 ? add_800596 : sel_800593;
  assign add_800600 = sel_800597 + 8'h01;
  assign sel_800601 = array_index_800332 == array_index_773038 ? add_800600 : sel_800597;
  assign add_800604 = sel_800601 + 8'h01;
  assign sel_800605 = array_index_800332 == array_index_773044 ? add_800604 : sel_800601;
  assign add_800608 = sel_800605 + 8'h01;
  assign sel_800609 = array_index_800332 == array_index_773050 ? add_800608 : sel_800605;
  assign add_800612 = sel_800609 + 8'h01;
  assign sel_800613 = array_index_800332 == array_index_773056 ? add_800612 : sel_800609;
  assign add_800616 = sel_800613 + 8'h01;
  assign sel_800617 = array_index_800332 == array_index_773062 ? add_800616 : sel_800613;
  assign add_800620 = sel_800617 + 8'h01;
  assign sel_800621 = array_index_800332 == array_index_773068 ? add_800620 : sel_800617;
  assign add_800624 = sel_800621 + 8'h01;
  assign sel_800625 = array_index_800332 == array_index_773074 ? add_800624 : sel_800621;
  assign add_800628 = sel_800625 + 8'h01;
  assign sel_800629 = array_index_800332 == array_index_773080 ? add_800628 : sel_800625;
  assign add_800632 = sel_800629 + 8'h01;
  assign sel_800633 = array_index_800332 == array_index_773086 ? add_800632 : sel_800629;
  assign add_800636 = sel_800633 + 8'h01;
  assign sel_800637 = array_index_800332 == array_index_773092 ? add_800636 : sel_800633;
  assign add_800640 = sel_800637 + 8'h01;
  assign sel_800641 = array_index_800332 == array_index_773098 ? add_800640 : sel_800637;
  assign add_800644 = sel_800641 + 8'h01;
  assign sel_800645 = array_index_800332 == array_index_773104 ? add_800644 : sel_800641;
  assign add_800648 = sel_800645 + 8'h01;
  assign sel_800649 = array_index_800332 == array_index_773110 ? add_800648 : sel_800645;
  assign add_800652 = sel_800649 + 8'h01;
  assign sel_800653 = array_index_800332 == array_index_773116 ? add_800652 : sel_800649;
  assign add_800656 = sel_800653 + 8'h01;
  assign sel_800657 = array_index_800332 == array_index_773122 ? add_800656 : sel_800653;
  assign add_800660 = sel_800657 + 8'h01;
  assign sel_800661 = array_index_800332 == array_index_773128 ? add_800660 : sel_800657;
  assign add_800664 = sel_800661 + 8'h01;
  assign sel_800665 = array_index_800332 == array_index_773134 ? add_800664 : sel_800661;
  assign add_800668 = sel_800665 + 8'h01;
  assign sel_800669 = array_index_800332 == array_index_773140 ? add_800668 : sel_800665;
  assign add_800672 = sel_800669 + 8'h01;
  assign sel_800673 = array_index_800332 == array_index_773146 ? add_800672 : sel_800669;
  assign add_800676 = sel_800673 + 8'h01;
  assign sel_800677 = array_index_800332 == array_index_773152 ? add_800676 : sel_800673;
  assign add_800680 = sel_800677 + 8'h01;
  assign sel_800681 = array_index_800332 == array_index_773158 ? add_800680 : sel_800677;
  assign add_800684 = sel_800681 + 8'h01;
  assign sel_800685 = array_index_800332 == array_index_773164 ? add_800684 : sel_800681;
  assign add_800688 = sel_800685 + 8'h01;
  assign sel_800689 = array_index_800332 == array_index_773170 ? add_800688 : sel_800685;
  assign add_800693 = sel_800689 + 8'h01;
  assign array_index_800694 = set1_unflattened[7'h4d];
  assign sel_800695 = array_index_800332 == array_index_773176 ? add_800693 : sel_800689;
  assign add_800698 = sel_800695 + 8'h01;
  assign sel_800699 = array_index_800694 == array_index_772632 ? add_800698 : sel_800695;
  assign add_800702 = sel_800699 + 8'h01;
  assign sel_800703 = array_index_800694 == array_index_772636 ? add_800702 : sel_800699;
  assign add_800706 = sel_800703 + 8'h01;
  assign sel_800707 = array_index_800694 == array_index_772644 ? add_800706 : sel_800703;
  assign add_800710 = sel_800707 + 8'h01;
  assign sel_800711 = array_index_800694 == array_index_772652 ? add_800710 : sel_800707;
  assign add_800714 = sel_800711 + 8'h01;
  assign sel_800715 = array_index_800694 == array_index_772660 ? add_800714 : sel_800711;
  assign add_800718 = sel_800715 + 8'h01;
  assign sel_800719 = array_index_800694 == array_index_772668 ? add_800718 : sel_800715;
  assign add_800722 = sel_800719 + 8'h01;
  assign sel_800723 = array_index_800694 == array_index_772676 ? add_800722 : sel_800719;
  assign add_800726 = sel_800723 + 8'h01;
  assign sel_800727 = array_index_800694 == array_index_772684 ? add_800726 : sel_800723;
  assign add_800730 = sel_800727 + 8'h01;
  assign sel_800731 = array_index_800694 == array_index_772690 ? add_800730 : sel_800727;
  assign add_800734 = sel_800731 + 8'h01;
  assign sel_800735 = array_index_800694 == array_index_772696 ? add_800734 : sel_800731;
  assign add_800738 = sel_800735 + 8'h01;
  assign sel_800739 = array_index_800694 == array_index_772702 ? add_800738 : sel_800735;
  assign add_800742 = sel_800739 + 8'h01;
  assign sel_800743 = array_index_800694 == array_index_772708 ? add_800742 : sel_800739;
  assign add_800746 = sel_800743 + 8'h01;
  assign sel_800747 = array_index_800694 == array_index_772714 ? add_800746 : sel_800743;
  assign add_800750 = sel_800747 + 8'h01;
  assign sel_800751 = array_index_800694 == array_index_772720 ? add_800750 : sel_800747;
  assign add_800754 = sel_800751 + 8'h01;
  assign sel_800755 = array_index_800694 == array_index_772726 ? add_800754 : sel_800751;
  assign add_800758 = sel_800755 + 8'h01;
  assign sel_800759 = array_index_800694 == array_index_772732 ? add_800758 : sel_800755;
  assign add_800762 = sel_800759 + 8'h01;
  assign sel_800763 = array_index_800694 == array_index_772738 ? add_800762 : sel_800759;
  assign add_800766 = sel_800763 + 8'h01;
  assign sel_800767 = array_index_800694 == array_index_772744 ? add_800766 : sel_800763;
  assign add_800770 = sel_800767 + 8'h01;
  assign sel_800771 = array_index_800694 == array_index_772750 ? add_800770 : sel_800767;
  assign add_800774 = sel_800771 + 8'h01;
  assign sel_800775 = array_index_800694 == array_index_772756 ? add_800774 : sel_800771;
  assign add_800778 = sel_800775 + 8'h01;
  assign sel_800779 = array_index_800694 == array_index_772762 ? add_800778 : sel_800775;
  assign add_800782 = sel_800779 + 8'h01;
  assign sel_800783 = array_index_800694 == array_index_772768 ? add_800782 : sel_800779;
  assign add_800786 = sel_800783 + 8'h01;
  assign sel_800787 = array_index_800694 == array_index_772774 ? add_800786 : sel_800783;
  assign add_800790 = sel_800787 + 8'h01;
  assign sel_800791 = array_index_800694 == array_index_772780 ? add_800790 : sel_800787;
  assign add_800794 = sel_800791 + 8'h01;
  assign sel_800795 = array_index_800694 == array_index_772786 ? add_800794 : sel_800791;
  assign add_800798 = sel_800795 + 8'h01;
  assign sel_800799 = array_index_800694 == array_index_772792 ? add_800798 : sel_800795;
  assign add_800802 = sel_800799 + 8'h01;
  assign sel_800803 = array_index_800694 == array_index_772798 ? add_800802 : sel_800799;
  assign add_800806 = sel_800803 + 8'h01;
  assign sel_800807 = array_index_800694 == array_index_772804 ? add_800806 : sel_800803;
  assign add_800810 = sel_800807 + 8'h01;
  assign sel_800811 = array_index_800694 == array_index_772810 ? add_800810 : sel_800807;
  assign add_800814 = sel_800811 + 8'h01;
  assign sel_800815 = array_index_800694 == array_index_772816 ? add_800814 : sel_800811;
  assign add_800818 = sel_800815 + 8'h01;
  assign sel_800819 = array_index_800694 == array_index_772822 ? add_800818 : sel_800815;
  assign add_800822 = sel_800819 + 8'h01;
  assign sel_800823 = array_index_800694 == array_index_772828 ? add_800822 : sel_800819;
  assign add_800826 = sel_800823 + 8'h01;
  assign sel_800827 = array_index_800694 == array_index_772834 ? add_800826 : sel_800823;
  assign add_800830 = sel_800827 + 8'h01;
  assign sel_800831 = array_index_800694 == array_index_772840 ? add_800830 : sel_800827;
  assign add_800834 = sel_800831 + 8'h01;
  assign sel_800835 = array_index_800694 == array_index_772846 ? add_800834 : sel_800831;
  assign add_800838 = sel_800835 + 8'h01;
  assign sel_800839 = array_index_800694 == array_index_772852 ? add_800838 : sel_800835;
  assign add_800842 = sel_800839 + 8'h01;
  assign sel_800843 = array_index_800694 == array_index_772858 ? add_800842 : sel_800839;
  assign add_800846 = sel_800843 + 8'h01;
  assign sel_800847 = array_index_800694 == array_index_772864 ? add_800846 : sel_800843;
  assign add_800850 = sel_800847 + 8'h01;
  assign sel_800851 = array_index_800694 == array_index_772870 ? add_800850 : sel_800847;
  assign add_800854 = sel_800851 + 8'h01;
  assign sel_800855 = array_index_800694 == array_index_772876 ? add_800854 : sel_800851;
  assign add_800858 = sel_800855 + 8'h01;
  assign sel_800859 = array_index_800694 == array_index_772882 ? add_800858 : sel_800855;
  assign add_800862 = sel_800859 + 8'h01;
  assign sel_800863 = array_index_800694 == array_index_772888 ? add_800862 : sel_800859;
  assign add_800866 = sel_800863 + 8'h01;
  assign sel_800867 = array_index_800694 == array_index_772894 ? add_800866 : sel_800863;
  assign add_800870 = sel_800867 + 8'h01;
  assign sel_800871 = array_index_800694 == array_index_772900 ? add_800870 : sel_800867;
  assign add_800874 = sel_800871 + 8'h01;
  assign sel_800875 = array_index_800694 == array_index_772906 ? add_800874 : sel_800871;
  assign add_800878 = sel_800875 + 8'h01;
  assign sel_800879 = array_index_800694 == array_index_772912 ? add_800878 : sel_800875;
  assign add_800882 = sel_800879 + 8'h01;
  assign sel_800883 = array_index_800694 == array_index_772918 ? add_800882 : sel_800879;
  assign add_800886 = sel_800883 + 8'h01;
  assign sel_800887 = array_index_800694 == array_index_772924 ? add_800886 : sel_800883;
  assign add_800890 = sel_800887 + 8'h01;
  assign sel_800891 = array_index_800694 == array_index_772930 ? add_800890 : sel_800887;
  assign add_800894 = sel_800891 + 8'h01;
  assign sel_800895 = array_index_800694 == array_index_772936 ? add_800894 : sel_800891;
  assign add_800898 = sel_800895 + 8'h01;
  assign sel_800899 = array_index_800694 == array_index_772942 ? add_800898 : sel_800895;
  assign add_800902 = sel_800899 + 8'h01;
  assign sel_800903 = array_index_800694 == array_index_772948 ? add_800902 : sel_800899;
  assign add_800906 = sel_800903 + 8'h01;
  assign sel_800907 = array_index_800694 == array_index_772954 ? add_800906 : sel_800903;
  assign add_800910 = sel_800907 + 8'h01;
  assign sel_800911 = array_index_800694 == array_index_772960 ? add_800910 : sel_800907;
  assign add_800914 = sel_800911 + 8'h01;
  assign sel_800915 = array_index_800694 == array_index_772966 ? add_800914 : sel_800911;
  assign add_800918 = sel_800915 + 8'h01;
  assign sel_800919 = array_index_800694 == array_index_772972 ? add_800918 : sel_800915;
  assign add_800922 = sel_800919 + 8'h01;
  assign sel_800923 = array_index_800694 == array_index_772978 ? add_800922 : sel_800919;
  assign add_800926 = sel_800923 + 8'h01;
  assign sel_800927 = array_index_800694 == array_index_772984 ? add_800926 : sel_800923;
  assign add_800930 = sel_800927 + 8'h01;
  assign sel_800931 = array_index_800694 == array_index_772990 ? add_800930 : sel_800927;
  assign add_800934 = sel_800931 + 8'h01;
  assign sel_800935 = array_index_800694 == array_index_772996 ? add_800934 : sel_800931;
  assign add_800938 = sel_800935 + 8'h01;
  assign sel_800939 = array_index_800694 == array_index_773002 ? add_800938 : sel_800935;
  assign add_800942 = sel_800939 + 8'h01;
  assign sel_800943 = array_index_800694 == array_index_773008 ? add_800942 : sel_800939;
  assign add_800946 = sel_800943 + 8'h01;
  assign sel_800947 = array_index_800694 == array_index_773014 ? add_800946 : sel_800943;
  assign add_800950 = sel_800947 + 8'h01;
  assign sel_800951 = array_index_800694 == array_index_773020 ? add_800950 : sel_800947;
  assign add_800954 = sel_800951 + 8'h01;
  assign sel_800955 = array_index_800694 == array_index_773026 ? add_800954 : sel_800951;
  assign add_800958 = sel_800955 + 8'h01;
  assign sel_800959 = array_index_800694 == array_index_773032 ? add_800958 : sel_800955;
  assign add_800962 = sel_800959 + 8'h01;
  assign sel_800963 = array_index_800694 == array_index_773038 ? add_800962 : sel_800959;
  assign add_800966 = sel_800963 + 8'h01;
  assign sel_800967 = array_index_800694 == array_index_773044 ? add_800966 : sel_800963;
  assign add_800970 = sel_800967 + 8'h01;
  assign sel_800971 = array_index_800694 == array_index_773050 ? add_800970 : sel_800967;
  assign add_800974 = sel_800971 + 8'h01;
  assign sel_800975 = array_index_800694 == array_index_773056 ? add_800974 : sel_800971;
  assign add_800978 = sel_800975 + 8'h01;
  assign sel_800979 = array_index_800694 == array_index_773062 ? add_800978 : sel_800975;
  assign add_800982 = sel_800979 + 8'h01;
  assign sel_800983 = array_index_800694 == array_index_773068 ? add_800982 : sel_800979;
  assign add_800986 = sel_800983 + 8'h01;
  assign sel_800987 = array_index_800694 == array_index_773074 ? add_800986 : sel_800983;
  assign add_800990 = sel_800987 + 8'h01;
  assign sel_800991 = array_index_800694 == array_index_773080 ? add_800990 : sel_800987;
  assign add_800994 = sel_800991 + 8'h01;
  assign sel_800995 = array_index_800694 == array_index_773086 ? add_800994 : sel_800991;
  assign add_800998 = sel_800995 + 8'h01;
  assign sel_800999 = array_index_800694 == array_index_773092 ? add_800998 : sel_800995;
  assign add_801002 = sel_800999 + 8'h01;
  assign sel_801003 = array_index_800694 == array_index_773098 ? add_801002 : sel_800999;
  assign add_801006 = sel_801003 + 8'h01;
  assign sel_801007 = array_index_800694 == array_index_773104 ? add_801006 : sel_801003;
  assign add_801010 = sel_801007 + 8'h01;
  assign sel_801011 = array_index_800694 == array_index_773110 ? add_801010 : sel_801007;
  assign add_801014 = sel_801011 + 8'h01;
  assign sel_801015 = array_index_800694 == array_index_773116 ? add_801014 : sel_801011;
  assign add_801018 = sel_801015 + 8'h01;
  assign sel_801019 = array_index_800694 == array_index_773122 ? add_801018 : sel_801015;
  assign add_801022 = sel_801019 + 8'h01;
  assign sel_801023 = array_index_800694 == array_index_773128 ? add_801022 : sel_801019;
  assign add_801026 = sel_801023 + 8'h01;
  assign sel_801027 = array_index_800694 == array_index_773134 ? add_801026 : sel_801023;
  assign add_801030 = sel_801027 + 8'h01;
  assign sel_801031 = array_index_800694 == array_index_773140 ? add_801030 : sel_801027;
  assign add_801034 = sel_801031 + 8'h01;
  assign sel_801035 = array_index_800694 == array_index_773146 ? add_801034 : sel_801031;
  assign add_801038 = sel_801035 + 8'h01;
  assign sel_801039 = array_index_800694 == array_index_773152 ? add_801038 : sel_801035;
  assign add_801042 = sel_801039 + 8'h01;
  assign sel_801043 = array_index_800694 == array_index_773158 ? add_801042 : sel_801039;
  assign add_801046 = sel_801043 + 8'h01;
  assign sel_801047 = array_index_800694 == array_index_773164 ? add_801046 : sel_801043;
  assign add_801050 = sel_801047 + 8'h01;
  assign sel_801051 = array_index_800694 == array_index_773170 ? add_801050 : sel_801047;
  assign add_801055 = sel_801051 + 8'h01;
  assign array_index_801056 = set1_unflattened[7'h4e];
  assign sel_801057 = array_index_800694 == array_index_773176 ? add_801055 : sel_801051;
  assign add_801060 = sel_801057 + 8'h01;
  assign sel_801061 = array_index_801056 == array_index_772632 ? add_801060 : sel_801057;
  assign add_801064 = sel_801061 + 8'h01;
  assign sel_801065 = array_index_801056 == array_index_772636 ? add_801064 : sel_801061;
  assign add_801068 = sel_801065 + 8'h01;
  assign sel_801069 = array_index_801056 == array_index_772644 ? add_801068 : sel_801065;
  assign add_801072 = sel_801069 + 8'h01;
  assign sel_801073 = array_index_801056 == array_index_772652 ? add_801072 : sel_801069;
  assign add_801076 = sel_801073 + 8'h01;
  assign sel_801077 = array_index_801056 == array_index_772660 ? add_801076 : sel_801073;
  assign add_801080 = sel_801077 + 8'h01;
  assign sel_801081 = array_index_801056 == array_index_772668 ? add_801080 : sel_801077;
  assign add_801084 = sel_801081 + 8'h01;
  assign sel_801085 = array_index_801056 == array_index_772676 ? add_801084 : sel_801081;
  assign add_801088 = sel_801085 + 8'h01;
  assign sel_801089 = array_index_801056 == array_index_772684 ? add_801088 : sel_801085;
  assign add_801092 = sel_801089 + 8'h01;
  assign sel_801093 = array_index_801056 == array_index_772690 ? add_801092 : sel_801089;
  assign add_801096 = sel_801093 + 8'h01;
  assign sel_801097 = array_index_801056 == array_index_772696 ? add_801096 : sel_801093;
  assign add_801100 = sel_801097 + 8'h01;
  assign sel_801101 = array_index_801056 == array_index_772702 ? add_801100 : sel_801097;
  assign add_801104 = sel_801101 + 8'h01;
  assign sel_801105 = array_index_801056 == array_index_772708 ? add_801104 : sel_801101;
  assign add_801108 = sel_801105 + 8'h01;
  assign sel_801109 = array_index_801056 == array_index_772714 ? add_801108 : sel_801105;
  assign add_801112 = sel_801109 + 8'h01;
  assign sel_801113 = array_index_801056 == array_index_772720 ? add_801112 : sel_801109;
  assign add_801116 = sel_801113 + 8'h01;
  assign sel_801117 = array_index_801056 == array_index_772726 ? add_801116 : sel_801113;
  assign add_801120 = sel_801117 + 8'h01;
  assign sel_801121 = array_index_801056 == array_index_772732 ? add_801120 : sel_801117;
  assign add_801124 = sel_801121 + 8'h01;
  assign sel_801125 = array_index_801056 == array_index_772738 ? add_801124 : sel_801121;
  assign add_801128 = sel_801125 + 8'h01;
  assign sel_801129 = array_index_801056 == array_index_772744 ? add_801128 : sel_801125;
  assign add_801132 = sel_801129 + 8'h01;
  assign sel_801133 = array_index_801056 == array_index_772750 ? add_801132 : sel_801129;
  assign add_801136 = sel_801133 + 8'h01;
  assign sel_801137 = array_index_801056 == array_index_772756 ? add_801136 : sel_801133;
  assign add_801140 = sel_801137 + 8'h01;
  assign sel_801141 = array_index_801056 == array_index_772762 ? add_801140 : sel_801137;
  assign add_801144 = sel_801141 + 8'h01;
  assign sel_801145 = array_index_801056 == array_index_772768 ? add_801144 : sel_801141;
  assign add_801148 = sel_801145 + 8'h01;
  assign sel_801149 = array_index_801056 == array_index_772774 ? add_801148 : sel_801145;
  assign add_801152 = sel_801149 + 8'h01;
  assign sel_801153 = array_index_801056 == array_index_772780 ? add_801152 : sel_801149;
  assign add_801156 = sel_801153 + 8'h01;
  assign sel_801157 = array_index_801056 == array_index_772786 ? add_801156 : sel_801153;
  assign add_801160 = sel_801157 + 8'h01;
  assign sel_801161 = array_index_801056 == array_index_772792 ? add_801160 : sel_801157;
  assign add_801164 = sel_801161 + 8'h01;
  assign sel_801165 = array_index_801056 == array_index_772798 ? add_801164 : sel_801161;
  assign add_801168 = sel_801165 + 8'h01;
  assign sel_801169 = array_index_801056 == array_index_772804 ? add_801168 : sel_801165;
  assign add_801172 = sel_801169 + 8'h01;
  assign sel_801173 = array_index_801056 == array_index_772810 ? add_801172 : sel_801169;
  assign add_801176 = sel_801173 + 8'h01;
  assign sel_801177 = array_index_801056 == array_index_772816 ? add_801176 : sel_801173;
  assign add_801180 = sel_801177 + 8'h01;
  assign sel_801181 = array_index_801056 == array_index_772822 ? add_801180 : sel_801177;
  assign add_801184 = sel_801181 + 8'h01;
  assign sel_801185 = array_index_801056 == array_index_772828 ? add_801184 : sel_801181;
  assign add_801188 = sel_801185 + 8'h01;
  assign sel_801189 = array_index_801056 == array_index_772834 ? add_801188 : sel_801185;
  assign add_801192 = sel_801189 + 8'h01;
  assign sel_801193 = array_index_801056 == array_index_772840 ? add_801192 : sel_801189;
  assign add_801196 = sel_801193 + 8'h01;
  assign sel_801197 = array_index_801056 == array_index_772846 ? add_801196 : sel_801193;
  assign add_801200 = sel_801197 + 8'h01;
  assign sel_801201 = array_index_801056 == array_index_772852 ? add_801200 : sel_801197;
  assign add_801204 = sel_801201 + 8'h01;
  assign sel_801205 = array_index_801056 == array_index_772858 ? add_801204 : sel_801201;
  assign add_801208 = sel_801205 + 8'h01;
  assign sel_801209 = array_index_801056 == array_index_772864 ? add_801208 : sel_801205;
  assign add_801212 = sel_801209 + 8'h01;
  assign sel_801213 = array_index_801056 == array_index_772870 ? add_801212 : sel_801209;
  assign add_801216 = sel_801213 + 8'h01;
  assign sel_801217 = array_index_801056 == array_index_772876 ? add_801216 : sel_801213;
  assign add_801220 = sel_801217 + 8'h01;
  assign sel_801221 = array_index_801056 == array_index_772882 ? add_801220 : sel_801217;
  assign add_801224 = sel_801221 + 8'h01;
  assign sel_801225 = array_index_801056 == array_index_772888 ? add_801224 : sel_801221;
  assign add_801228 = sel_801225 + 8'h01;
  assign sel_801229 = array_index_801056 == array_index_772894 ? add_801228 : sel_801225;
  assign add_801232 = sel_801229 + 8'h01;
  assign sel_801233 = array_index_801056 == array_index_772900 ? add_801232 : sel_801229;
  assign add_801236 = sel_801233 + 8'h01;
  assign sel_801237 = array_index_801056 == array_index_772906 ? add_801236 : sel_801233;
  assign add_801240 = sel_801237 + 8'h01;
  assign sel_801241 = array_index_801056 == array_index_772912 ? add_801240 : sel_801237;
  assign add_801244 = sel_801241 + 8'h01;
  assign sel_801245 = array_index_801056 == array_index_772918 ? add_801244 : sel_801241;
  assign add_801248 = sel_801245 + 8'h01;
  assign sel_801249 = array_index_801056 == array_index_772924 ? add_801248 : sel_801245;
  assign add_801252 = sel_801249 + 8'h01;
  assign sel_801253 = array_index_801056 == array_index_772930 ? add_801252 : sel_801249;
  assign add_801256 = sel_801253 + 8'h01;
  assign sel_801257 = array_index_801056 == array_index_772936 ? add_801256 : sel_801253;
  assign add_801260 = sel_801257 + 8'h01;
  assign sel_801261 = array_index_801056 == array_index_772942 ? add_801260 : sel_801257;
  assign add_801264 = sel_801261 + 8'h01;
  assign sel_801265 = array_index_801056 == array_index_772948 ? add_801264 : sel_801261;
  assign add_801268 = sel_801265 + 8'h01;
  assign sel_801269 = array_index_801056 == array_index_772954 ? add_801268 : sel_801265;
  assign add_801272 = sel_801269 + 8'h01;
  assign sel_801273 = array_index_801056 == array_index_772960 ? add_801272 : sel_801269;
  assign add_801276 = sel_801273 + 8'h01;
  assign sel_801277 = array_index_801056 == array_index_772966 ? add_801276 : sel_801273;
  assign add_801280 = sel_801277 + 8'h01;
  assign sel_801281 = array_index_801056 == array_index_772972 ? add_801280 : sel_801277;
  assign add_801284 = sel_801281 + 8'h01;
  assign sel_801285 = array_index_801056 == array_index_772978 ? add_801284 : sel_801281;
  assign add_801288 = sel_801285 + 8'h01;
  assign sel_801289 = array_index_801056 == array_index_772984 ? add_801288 : sel_801285;
  assign add_801292 = sel_801289 + 8'h01;
  assign sel_801293 = array_index_801056 == array_index_772990 ? add_801292 : sel_801289;
  assign add_801296 = sel_801293 + 8'h01;
  assign sel_801297 = array_index_801056 == array_index_772996 ? add_801296 : sel_801293;
  assign add_801300 = sel_801297 + 8'h01;
  assign sel_801301 = array_index_801056 == array_index_773002 ? add_801300 : sel_801297;
  assign add_801304 = sel_801301 + 8'h01;
  assign sel_801305 = array_index_801056 == array_index_773008 ? add_801304 : sel_801301;
  assign add_801308 = sel_801305 + 8'h01;
  assign sel_801309 = array_index_801056 == array_index_773014 ? add_801308 : sel_801305;
  assign add_801312 = sel_801309 + 8'h01;
  assign sel_801313 = array_index_801056 == array_index_773020 ? add_801312 : sel_801309;
  assign add_801316 = sel_801313 + 8'h01;
  assign sel_801317 = array_index_801056 == array_index_773026 ? add_801316 : sel_801313;
  assign add_801320 = sel_801317 + 8'h01;
  assign sel_801321 = array_index_801056 == array_index_773032 ? add_801320 : sel_801317;
  assign add_801324 = sel_801321 + 8'h01;
  assign sel_801325 = array_index_801056 == array_index_773038 ? add_801324 : sel_801321;
  assign add_801328 = sel_801325 + 8'h01;
  assign sel_801329 = array_index_801056 == array_index_773044 ? add_801328 : sel_801325;
  assign add_801332 = sel_801329 + 8'h01;
  assign sel_801333 = array_index_801056 == array_index_773050 ? add_801332 : sel_801329;
  assign add_801336 = sel_801333 + 8'h01;
  assign sel_801337 = array_index_801056 == array_index_773056 ? add_801336 : sel_801333;
  assign add_801340 = sel_801337 + 8'h01;
  assign sel_801341 = array_index_801056 == array_index_773062 ? add_801340 : sel_801337;
  assign add_801344 = sel_801341 + 8'h01;
  assign sel_801345 = array_index_801056 == array_index_773068 ? add_801344 : sel_801341;
  assign add_801348 = sel_801345 + 8'h01;
  assign sel_801349 = array_index_801056 == array_index_773074 ? add_801348 : sel_801345;
  assign add_801352 = sel_801349 + 8'h01;
  assign sel_801353 = array_index_801056 == array_index_773080 ? add_801352 : sel_801349;
  assign add_801356 = sel_801353 + 8'h01;
  assign sel_801357 = array_index_801056 == array_index_773086 ? add_801356 : sel_801353;
  assign add_801360 = sel_801357 + 8'h01;
  assign sel_801361 = array_index_801056 == array_index_773092 ? add_801360 : sel_801357;
  assign add_801364 = sel_801361 + 8'h01;
  assign sel_801365 = array_index_801056 == array_index_773098 ? add_801364 : sel_801361;
  assign add_801368 = sel_801365 + 8'h01;
  assign sel_801369 = array_index_801056 == array_index_773104 ? add_801368 : sel_801365;
  assign add_801372 = sel_801369 + 8'h01;
  assign sel_801373 = array_index_801056 == array_index_773110 ? add_801372 : sel_801369;
  assign add_801376 = sel_801373 + 8'h01;
  assign sel_801377 = array_index_801056 == array_index_773116 ? add_801376 : sel_801373;
  assign add_801380 = sel_801377 + 8'h01;
  assign sel_801381 = array_index_801056 == array_index_773122 ? add_801380 : sel_801377;
  assign add_801384 = sel_801381 + 8'h01;
  assign sel_801385 = array_index_801056 == array_index_773128 ? add_801384 : sel_801381;
  assign add_801388 = sel_801385 + 8'h01;
  assign sel_801389 = array_index_801056 == array_index_773134 ? add_801388 : sel_801385;
  assign add_801392 = sel_801389 + 8'h01;
  assign sel_801393 = array_index_801056 == array_index_773140 ? add_801392 : sel_801389;
  assign add_801396 = sel_801393 + 8'h01;
  assign sel_801397 = array_index_801056 == array_index_773146 ? add_801396 : sel_801393;
  assign add_801400 = sel_801397 + 8'h01;
  assign sel_801401 = array_index_801056 == array_index_773152 ? add_801400 : sel_801397;
  assign add_801404 = sel_801401 + 8'h01;
  assign sel_801405 = array_index_801056 == array_index_773158 ? add_801404 : sel_801401;
  assign add_801408 = sel_801405 + 8'h01;
  assign sel_801409 = array_index_801056 == array_index_773164 ? add_801408 : sel_801405;
  assign add_801412 = sel_801409 + 8'h01;
  assign sel_801413 = array_index_801056 == array_index_773170 ? add_801412 : sel_801409;
  assign add_801417 = sel_801413 + 8'h01;
  assign array_index_801418 = set1_unflattened[7'h4f];
  assign sel_801419 = array_index_801056 == array_index_773176 ? add_801417 : sel_801413;
  assign add_801422 = sel_801419 + 8'h01;
  assign sel_801423 = array_index_801418 == array_index_772632 ? add_801422 : sel_801419;
  assign add_801426 = sel_801423 + 8'h01;
  assign sel_801427 = array_index_801418 == array_index_772636 ? add_801426 : sel_801423;
  assign add_801430 = sel_801427 + 8'h01;
  assign sel_801431 = array_index_801418 == array_index_772644 ? add_801430 : sel_801427;
  assign add_801434 = sel_801431 + 8'h01;
  assign sel_801435 = array_index_801418 == array_index_772652 ? add_801434 : sel_801431;
  assign add_801438 = sel_801435 + 8'h01;
  assign sel_801439 = array_index_801418 == array_index_772660 ? add_801438 : sel_801435;
  assign add_801442 = sel_801439 + 8'h01;
  assign sel_801443 = array_index_801418 == array_index_772668 ? add_801442 : sel_801439;
  assign add_801446 = sel_801443 + 8'h01;
  assign sel_801447 = array_index_801418 == array_index_772676 ? add_801446 : sel_801443;
  assign add_801450 = sel_801447 + 8'h01;
  assign sel_801451 = array_index_801418 == array_index_772684 ? add_801450 : sel_801447;
  assign add_801454 = sel_801451 + 8'h01;
  assign sel_801455 = array_index_801418 == array_index_772690 ? add_801454 : sel_801451;
  assign add_801458 = sel_801455 + 8'h01;
  assign sel_801459 = array_index_801418 == array_index_772696 ? add_801458 : sel_801455;
  assign add_801462 = sel_801459 + 8'h01;
  assign sel_801463 = array_index_801418 == array_index_772702 ? add_801462 : sel_801459;
  assign add_801466 = sel_801463 + 8'h01;
  assign sel_801467 = array_index_801418 == array_index_772708 ? add_801466 : sel_801463;
  assign add_801470 = sel_801467 + 8'h01;
  assign sel_801471 = array_index_801418 == array_index_772714 ? add_801470 : sel_801467;
  assign add_801474 = sel_801471 + 8'h01;
  assign sel_801475 = array_index_801418 == array_index_772720 ? add_801474 : sel_801471;
  assign add_801478 = sel_801475 + 8'h01;
  assign sel_801479 = array_index_801418 == array_index_772726 ? add_801478 : sel_801475;
  assign add_801482 = sel_801479 + 8'h01;
  assign sel_801483 = array_index_801418 == array_index_772732 ? add_801482 : sel_801479;
  assign add_801486 = sel_801483 + 8'h01;
  assign sel_801487 = array_index_801418 == array_index_772738 ? add_801486 : sel_801483;
  assign add_801490 = sel_801487 + 8'h01;
  assign sel_801491 = array_index_801418 == array_index_772744 ? add_801490 : sel_801487;
  assign add_801494 = sel_801491 + 8'h01;
  assign sel_801495 = array_index_801418 == array_index_772750 ? add_801494 : sel_801491;
  assign add_801498 = sel_801495 + 8'h01;
  assign sel_801499 = array_index_801418 == array_index_772756 ? add_801498 : sel_801495;
  assign add_801502 = sel_801499 + 8'h01;
  assign sel_801503 = array_index_801418 == array_index_772762 ? add_801502 : sel_801499;
  assign add_801506 = sel_801503 + 8'h01;
  assign sel_801507 = array_index_801418 == array_index_772768 ? add_801506 : sel_801503;
  assign add_801510 = sel_801507 + 8'h01;
  assign sel_801511 = array_index_801418 == array_index_772774 ? add_801510 : sel_801507;
  assign add_801514 = sel_801511 + 8'h01;
  assign sel_801515 = array_index_801418 == array_index_772780 ? add_801514 : sel_801511;
  assign add_801518 = sel_801515 + 8'h01;
  assign sel_801519 = array_index_801418 == array_index_772786 ? add_801518 : sel_801515;
  assign add_801522 = sel_801519 + 8'h01;
  assign sel_801523 = array_index_801418 == array_index_772792 ? add_801522 : sel_801519;
  assign add_801526 = sel_801523 + 8'h01;
  assign sel_801527 = array_index_801418 == array_index_772798 ? add_801526 : sel_801523;
  assign add_801530 = sel_801527 + 8'h01;
  assign sel_801531 = array_index_801418 == array_index_772804 ? add_801530 : sel_801527;
  assign add_801534 = sel_801531 + 8'h01;
  assign sel_801535 = array_index_801418 == array_index_772810 ? add_801534 : sel_801531;
  assign add_801538 = sel_801535 + 8'h01;
  assign sel_801539 = array_index_801418 == array_index_772816 ? add_801538 : sel_801535;
  assign add_801542 = sel_801539 + 8'h01;
  assign sel_801543 = array_index_801418 == array_index_772822 ? add_801542 : sel_801539;
  assign add_801546 = sel_801543 + 8'h01;
  assign sel_801547 = array_index_801418 == array_index_772828 ? add_801546 : sel_801543;
  assign add_801550 = sel_801547 + 8'h01;
  assign sel_801551 = array_index_801418 == array_index_772834 ? add_801550 : sel_801547;
  assign add_801554 = sel_801551 + 8'h01;
  assign sel_801555 = array_index_801418 == array_index_772840 ? add_801554 : sel_801551;
  assign add_801558 = sel_801555 + 8'h01;
  assign sel_801559 = array_index_801418 == array_index_772846 ? add_801558 : sel_801555;
  assign add_801562 = sel_801559 + 8'h01;
  assign sel_801563 = array_index_801418 == array_index_772852 ? add_801562 : sel_801559;
  assign add_801566 = sel_801563 + 8'h01;
  assign sel_801567 = array_index_801418 == array_index_772858 ? add_801566 : sel_801563;
  assign add_801570 = sel_801567 + 8'h01;
  assign sel_801571 = array_index_801418 == array_index_772864 ? add_801570 : sel_801567;
  assign add_801574 = sel_801571 + 8'h01;
  assign sel_801575 = array_index_801418 == array_index_772870 ? add_801574 : sel_801571;
  assign add_801578 = sel_801575 + 8'h01;
  assign sel_801579 = array_index_801418 == array_index_772876 ? add_801578 : sel_801575;
  assign add_801582 = sel_801579 + 8'h01;
  assign sel_801583 = array_index_801418 == array_index_772882 ? add_801582 : sel_801579;
  assign add_801586 = sel_801583 + 8'h01;
  assign sel_801587 = array_index_801418 == array_index_772888 ? add_801586 : sel_801583;
  assign add_801590 = sel_801587 + 8'h01;
  assign sel_801591 = array_index_801418 == array_index_772894 ? add_801590 : sel_801587;
  assign add_801594 = sel_801591 + 8'h01;
  assign sel_801595 = array_index_801418 == array_index_772900 ? add_801594 : sel_801591;
  assign add_801598 = sel_801595 + 8'h01;
  assign sel_801599 = array_index_801418 == array_index_772906 ? add_801598 : sel_801595;
  assign add_801602 = sel_801599 + 8'h01;
  assign sel_801603 = array_index_801418 == array_index_772912 ? add_801602 : sel_801599;
  assign add_801606 = sel_801603 + 8'h01;
  assign sel_801607 = array_index_801418 == array_index_772918 ? add_801606 : sel_801603;
  assign add_801610 = sel_801607 + 8'h01;
  assign sel_801611 = array_index_801418 == array_index_772924 ? add_801610 : sel_801607;
  assign add_801614 = sel_801611 + 8'h01;
  assign sel_801615 = array_index_801418 == array_index_772930 ? add_801614 : sel_801611;
  assign add_801618 = sel_801615 + 8'h01;
  assign sel_801619 = array_index_801418 == array_index_772936 ? add_801618 : sel_801615;
  assign add_801622 = sel_801619 + 8'h01;
  assign sel_801623 = array_index_801418 == array_index_772942 ? add_801622 : sel_801619;
  assign add_801626 = sel_801623 + 8'h01;
  assign sel_801627 = array_index_801418 == array_index_772948 ? add_801626 : sel_801623;
  assign add_801630 = sel_801627 + 8'h01;
  assign sel_801631 = array_index_801418 == array_index_772954 ? add_801630 : sel_801627;
  assign add_801634 = sel_801631 + 8'h01;
  assign sel_801635 = array_index_801418 == array_index_772960 ? add_801634 : sel_801631;
  assign add_801638 = sel_801635 + 8'h01;
  assign sel_801639 = array_index_801418 == array_index_772966 ? add_801638 : sel_801635;
  assign add_801642 = sel_801639 + 8'h01;
  assign sel_801643 = array_index_801418 == array_index_772972 ? add_801642 : sel_801639;
  assign add_801646 = sel_801643 + 8'h01;
  assign sel_801647 = array_index_801418 == array_index_772978 ? add_801646 : sel_801643;
  assign add_801650 = sel_801647 + 8'h01;
  assign sel_801651 = array_index_801418 == array_index_772984 ? add_801650 : sel_801647;
  assign add_801654 = sel_801651 + 8'h01;
  assign sel_801655 = array_index_801418 == array_index_772990 ? add_801654 : sel_801651;
  assign add_801658 = sel_801655 + 8'h01;
  assign sel_801659 = array_index_801418 == array_index_772996 ? add_801658 : sel_801655;
  assign add_801662 = sel_801659 + 8'h01;
  assign sel_801663 = array_index_801418 == array_index_773002 ? add_801662 : sel_801659;
  assign add_801666 = sel_801663 + 8'h01;
  assign sel_801667 = array_index_801418 == array_index_773008 ? add_801666 : sel_801663;
  assign add_801670 = sel_801667 + 8'h01;
  assign sel_801671 = array_index_801418 == array_index_773014 ? add_801670 : sel_801667;
  assign add_801674 = sel_801671 + 8'h01;
  assign sel_801675 = array_index_801418 == array_index_773020 ? add_801674 : sel_801671;
  assign add_801678 = sel_801675 + 8'h01;
  assign sel_801679 = array_index_801418 == array_index_773026 ? add_801678 : sel_801675;
  assign add_801682 = sel_801679 + 8'h01;
  assign sel_801683 = array_index_801418 == array_index_773032 ? add_801682 : sel_801679;
  assign add_801686 = sel_801683 + 8'h01;
  assign sel_801687 = array_index_801418 == array_index_773038 ? add_801686 : sel_801683;
  assign add_801690 = sel_801687 + 8'h01;
  assign sel_801691 = array_index_801418 == array_index_773044 ? add_801690 : sel_801687;
  assign add_801694 = sel_801691 + 8'h01;
  assign sel_801695 = array_index_801418 == array_index_773050 ? add_801694 : sel_801691;
  assign add_801698 = sel_801695 + 8'h01;
  assign sel_801699 = array_index_801418 == array_index_773056 ? add_801698 : sel_801695;
  assign add_801702 = sel_801699 + 8'h01;
  assign sel_801703 = array_index_801418 == array_index_773062 ? add_801702 : sel_801699;
  assign add_801706 = sel_801703 + 8'h01;
  assign sel_801707 = array_index_801418 == array_index_773068 ? add_801706 : sel_801703;
  assign add_801710 = sel_801707 + 8'h01;
  assign sel_801711 = array_index_801418 == array_index_773074 ? add_801710 : sel_801707;
  assign add_801714 = sel_801711 + 8'h01;
  assign sel_801715 = array_index_801418 == array_index_773080 ? add_801714 : sel_801711;
  assign add_801718 = sel_801715 + 8'h01;
  assign sel_801719 = array_index_801418 == array_index_773086 ? add_801718 : sel_801715;
  assign add_801722 = sel_801719 + 8'h01;
  assign sel_801723 = array_index_801418 == array_index_773092 ? add_801722 : sel_801719;
  assign add_801726 = sel_801723 + 8'h01;
  assign sel_801727 = array_index_801418 == array_index_773098 ? add_801726 : sel_801723;
  assign add_801730 = sel_801727 + 8'h01;
  assign sel_801731 = array_index_801418 == array_index_773104 ? add_801730 : sel_801727;
  assign add_801734 = sel_801731 + 8'h01;
  assign sel_801735 = array_index_801418 == array_index_773110 ? add_801734 : sel_801731;
  assign add_801738 = sel_801735 + 8'h01;
  assign sel_801739 = array_index_801418 == array_index_773116 ? add_801738 : sel_801735;
  assign add_801742 = sel_801739 + 8'h01;
  assign sel_801743 = array_index_801418 == array_index_773122 ? add_801742 : sel_801739;
  assign add_801746 = sel_801743 + 8'h01;
  assign sel_801747 = array_index_801418 == array_index_773128 ? add_801746 : sel_801743;
  assign add_801750 = sel_801747 + 8'h01;
  assign sel_801751 = array_index_801418 == array_index_773134 ? add_801750 : sel_801747;
  assign add_801754 = sel_801751 + 8'h01;
  assign sel_801755 = array_index_801418 == array_index_773140 ? add_801754 : sel_801751;
  assign add_801758 = sel_801755 + 8'h01;
  assign sel_801759 = array_index_801418 == array_index_773146 ? add_801758 : sel_801755;
  assign add_801762 = sel_801759 + 8'h01;
  assign sel_801763 = array_index_801418 == array_index_773152 ? add_801762 : sel_801759;
  assign add_801766 = sel_801763 + 8'h01;
  assign sel_801767 = array_index_801418 == array_index_773158 ? add_801766 : sel_801763;
  assign add_801770 = sel_801767 + 8'h01;
  assign sel_801771 = array_index_801418 == array_index_773164 ? add_801770 : sel_801767;
  assign add_801774 = sel_801771 + 8'h01;
  assign sel_801775 = array_index_801418 == array_index_773170 ? add_801774 : sel_801771;
  assign add_801779 = sel_801775 + 8'h01;
  assign array_index_801780 = set1_unflattened[7'h50];
  assign sel_801781 = array_index_801418 == array_index_773176 ? add_801779 : sel_801775;
  assign add_801784 = sel_801781 + 8'h01;
  assign sel_801785 = array_index_801780 == array_index_772632 ? add_801784 : sel_801781;
  assign add_801788 = sel_801785 + 8'h01;
  assign sel_801789 = array_index_801780 == array_index_772636 ? add_801788 : sel_801785;
  assign add_801792 = sel_801789 + 8'h01;
  assign sel_801793 = array_index_801780 == array_index_772644 ? add_801792 : sel_801789;
  assign add_801796 = sel_801793 + 8'h01;
  assign sel_801797 = array_index_801780 == array_index_772652 ? add_801796 : sel_801793;
  assign add_801800 = sel_801797 + 8'h01;
  assign sel_801801 = array_index_801780 == array_index_772660 ? add_801800 : sel_801797;
  assign add_801804 = sel_801801 + 8'h01;
  assign sel_801805 = array_index_801780 == array_index_772668 ? add_801804 : sel_801801;
  assign add_801808 = sel_801805 + 8'h01;
  assign sel_801809 = array_index_801780 == array_index_772676 ? add_801808 : sel_801805;
  assign add_801812 = sel_801809 + 8'h01;
  assign sel_801813 = array_index_801780 == array_index_772684 ? add_801812 : sel_801809;
  assign add_801816 = sel_801813 + 8'h01;
  assign sel_801817 = array_index_801780 == array_index_772690 ? add_801816 : sel_801813;
  assign add_801820 = sel_801817 + 8'h01;
  assign sel_801821 = array_index_801780 == array_index_772696 ? add_801820 : sel_801817;
  assign add_801824 = sel_801821 + 8'h01;
  assign sel_801825 = array_index_801780 == array_index_772702 ? add_801824 : sel_801821;
  assign add_801828 = sel_801825 + 8'h01;
  assign sel_801829 = array_index_801780 == array_index_772708 ? add_801828 : sel_801825;
  assign add_801832 = sel_801829 + 8'h01;
  assign sel_801833 = array_index_801780 == array_index_772714 ? add_801832 : sel_801829;
  assign add_801836 = sel_801833 + 8'h01;
  assign sel_801837 = array_index_801780 == array_index_772720 ? add_801836 : sel_801833;
  assign add_801840 = sel_801837 + 8'h01;
  assign sel_801841 = array_index_801780 == array_index_772726 ? add_801840 : sel_801837;
  assign add_801844 = sel_801841 + 8'h01;
  assign sel_801845 = array_index_801780 == array_index_772732 ? add_801844 : sel_801841;
  assign add_801848 = sel_801845 + 8'h01;
  assign sel_801849 = array_index_801780 == array_index_772738 ? add_801848 : sel_801845;
  assign add_801852 = sel_801849 + 8'h01;
  assign sel_801853 = array_index_801780 == array_index_772744 ? add_801852 : sel_801849;
  assign add_801856 = sel_801853 + 8'h01;
  assign sel_801857 = array_index_801780 == array_index_772750 ? add_801856 : sel_801853;
  assign add_801860 = sel_801857 + 8'h01;
  assign sel_801861 = array_index_801780 == array_index_772756 ? add_801860 : sel_801857;
  assign add_801864 = sel_801861 + 8'h01;
  assign sel_801865 = array_index_801780 == array_index_772762 ? add_801864 : sel_801861;
  assign add_801868 = sel_801865 + 8'h01;
  assign sel_801869 = array_index_801780 == array_index_772768 ? add_801868 : sel_801865;
  assign add_801872 = sel_801869 + 8'h01;
  assign sel_801873 = array_index_801780 == array_index_772774 ? add_801872 : sel_801869;
  assign add_801876 = sel_801873 + 8'h01;
  assign sel_801877 = array_index_801780 == array_index_772780 ? add_801876 : sel_801873;
  assign add_801880 = sel_801877 + 8'h01;
  assign sel_801881 = array_index_801780 == array_index_772786 ? add_801880 : sel_801877;
  assign add_801884 = sel_801881 + 8'h01;
  assign sel_801885 = array_index_801780 == array_index_772792 ? add_801884 : sel_801881;
  assign add_801888 = sel_801885 + 8'h01;
  assign sel_801889 = array_index_801780 == array_index_772798 ? add_801888 : sel_801885;
  assign add_801892 = sel_801889 + 8'h01;
  assign sel_801893 = array_index_801780 == array_index_772804 ? add_801892 : sel_801889;
  assign add_801896 = sel_801893 + 8'h01;
  assign sel_801897 = array_index_801780 == array_index_772810 ? add_801896 : sel_801893;
  assign add_801900 = sel_801897 + 8'h01;
  assign sel_801901 = array_index_801780 == array_index_772816 ? add_801900 : sel_801897;
  assign add_801904 = sel_801901 + 8'h01;
  assign sel_801905 = array_index_801780 == array_index_772822 ? add_801904 : sel_801901;
  assign add_801908 = sel_801905 + 8'h01;
  assign sel_801909 = array_index_801780 == array_index_772828 ? add_801908 : sel_801905;
  assign add_801912 = sel_801909 + 8'h01;
  assign sel_801913 = array_index_801780 == array_index_772834 ? add_801912 : sel_801909;
  assign add_801916 = sel_801913 + 8'h01;
  assign sel_801917 = array_index_801780 == array_index_772840 ? add_801916 : sel_801913;
  assign add_801920 = sel_801917 + 8'h01;
  assign sel_801921 = array_index_801780 == array_index_772846 ? add_801920 : sel_801917;
  assign add_801924 = sel_801921 + 8'h01;
  assign sel_801925 = array_index_801780 == array_index_772852 ? add_801924 : sel_801921;
  assign add_801928 = sel_801925 + 8'h01;
  assign sel_801929 = array_index_801780 == array_index_772858 ? add_801928 : sel_801925;
  assign add_801932 = sel_801929 + 8'h01;
  assign sel_801933 = array_index_801780 == array_index_772864 ? add_801932 : sel_801929;
  assign add_801936 = sel_801933 + 8'h01;
  assign sel_801937 = array_index_801780 == array_index_772870 ? add_801936 : sel_801933;
  assign add_801940 = sel_801937 + 8'h01;
  assign sel_801941 = array_index_801780 == array_index_772876 ? add_801940 : sel_801937;
  assign add_801944 = sel_801941 + 8'h01;
  assign sel_801945 = array_index_801780 == array_index_772882 ? add_801944 : sel_801941;
  assign add_801948 = sel_801945 + 8'h01;
  assign sel_801949 = array_index_801780 == array_index_772888 ? add_801948 : sel_801945;
  assign add_801952 = sel_801949 + 8'h01;
  assign sel_801953 = array_index_801780 == array_index_772894 ? add_801952 : sel_801949;
  assign add_801956 = sel_801953 + 8'h01;
  assign sel_801957 = array_index_801780 == array_index_772900 ? add_801956 : sel_801953;
  assign add_801960 = sel_801957 + 8'h01;
  assign sel_801961 = array_index_801780 == array_index_772906 ? add_801960 : sel_801957;
  assign add_801964 = sel_801961 + 8'h01;
  assign sel_801965 = array_index_801780 == array_index_772912 ? add_801964 : sel_801961;
  assign add_801968 = sel_801965 + 8'h01;
  assign sel_801969 = array_index_801780 == array_index_772918 ? add_801968 : sel_801965;
  assign add_801972 = sel_801969 + 8'h01;
  assign sel_801973 = array_index_801780 == array_index_772924 ? add_801972 : sel_801969;
  assign add_801976 = sel_801973 + 8'h01;
  assign sel_801977 = array_index_801780 == array_index_772930 ? add_801976 : sel_801973;
  assign add_801980 = sel_801977 + 8'h01;
  assign sel_801981 = array_index_801780 == array_index_772936 ? add_801980 : sel_801977;
  assign add_801984 = sel_801981 + 8'h01;
  assign sel_801985 = array_index_801780 == array_index_772942 ? add_801984 : sel_801981;
  assign add_801988 = sel_801985 + 8'h01;
  assign sel_801989 = array_index_801780 == array_index_772948 ? add_801988 : sel_801985;
  assign add_801992 = sel_801989 + 8'h01;
  assign sel_801993 = array_index_801780 == array_index_772954 ? add_801992 : sel_801989;
  assign add_801996 = sel_801993 + 8'h01;
  assign sel_801997 = array_index_801780 == array_index_772960 ? add_801996 : sel_801993;
  assign add_802000 = sel_801997 + 8'h01;
  assign sel_802001 = array_index_801780 == array_index_772966 ? add_802000 : sel_801997;
  assign add_802004 = sel_802001 + 8'h01;
  assign sel_802005 = array_index_801780 == array_index_772972 ? add_802004 : sel_802001;
  assign add_802008 = sel_802005 + 8'h01;
  assign sel_802009 = array_index_801780 == array_index_772978 ? add_802008 : sel_802005;
  assign add_802012 = sel_802009 + 8'h01;
  assign sel_802013 = array_index_801780 == array_index_772984 ? add_802012 : sel_802009;
  assign add_802016 = sel_802013 + 8'h01;
  assign sel_802017 = array_index_801780 == array_index_772990 ? add_802016 : sel_802013;
  assign add_802020 = sel_802017 + 8'h01;
  assign sel_802021 = array_index_801780 == array_index_772996 ? add_802020 : sel_802017;
  assign add_802024 = sel_802021 + 8'h01;
  assign sel_802025 = array_index_801780 == array_index_773002 ? add_802024 : sel_802021;
  assign add_802028 = sel_802025 + 8'h01;
  assign sel_802029 = array_index_801780 == array_index_773008 ? add_802028 : sel_802025;
  assign add_802032 = sel_802029 + 8'h01;
  assign sel_802033 = array_index_801780 == array_index_773014 ? add_802032 : sel_802029;
  assign add_802036 = sel_802033 + 8'h01;
  assign sel_802037 = array_index_801780 == array_index_773020 ? add_802036 : sel_802033;
  assign add_802040 = sel_802037 + 8'h01;
  assign sel_802041 = array_index_801780 == array_index_773026 ? add_802040 : sel_802037;
  assign add_802044 = sel_802041 + 8'h01;
  assign sel_802045 = array_index_801780 == array_index_773032 ? add_802044 : sel_802041;
  assign add_802048 = sel_802045 + 8'h01;
  assign sel_802049 = array_index_801780 == array_index_773038 ? add_802048 : sel_802045;
  assign add_802052 = sel_802049 + 8'h01;
  assign sel_802053 = array_index_801780 == array_index_773044 ? add_802052 : sel_802049;
  assign add_802056 = sel_802053 + 8'h01;
  assign sel_802057 = array_index_801780 == array_index_773050 ? add_802056 : sel_802053;
  assign add_802060 = sel_802057 + 8'h01;
  assign sel_802061 = array_index_801780 == array_index_773056 ? add_802060 : sel_802057;
  assign add_802064 = sel_802061 + 8'h01;
  assign sel_802065 = array_index_801780 == array_index_773062 ? add_802064 : sel_802061;
  assign add_802068 = sel_802065 + 8'h01;
  assign sel_802069 = array_index_801780 == array_index_773068 ? add_802068 : sel_802065;
  assign add_802072 = sel_802069 + 8'h01;
  assign sel_802073 = array_index_801780 == array_index_773074 ? add_802072 : sel_802069;
  assign add_802076 = sel_802073 + 8'h01;
  assign sel_802077 = array_index_801780 == array_index_773080 ? add_802076 : sel_802073;
  assign add_802080 = sel_802077 + 8'h01;
  assign sel_802081 = array_index_801780 == array_index_773086 ? add_802080 : sel_802077;
  assign add_802084 = sel_802081 + 8'h01;
  assign sel_802085 = array_index_801780 == array_index_773092 ? add_802084 : sel_802081;
  assign add_802088 = sel_802085 + 8'h01;
  assign sel_802089 = array_index_801780 == array_index_773098 ? add_802088 : sel_802085;
  assign add_802092 = sel_802089 + 8'h01;
  assign sel_802093 = array_index_801780 == array_index_773104 ? add_802092 : sel_802089;
  assign add_802096 = sel_802093 + 8'h01;
  assign sel_802097 = array_index_801780 == array_index_773110 ? add_802096 : sel_802093;
  assign add_802100 = sel_802097 + 8'h01;
  assign sel_802101 = array_index_801780 == array_index_773116 ? add_802100 : sel_802097;
  assign add_802104 = sel_802101 + 8'h01;
  assign sel_802105 = array_index_801780 == array_index_773122 ? add_802104 : sel_802101;
  assign add_802108 = sel_802105 + 8'h01;
  assign sel_802109 = array_index_801780 == array_index_773128 ? add_802108 : sel_802105;
  assign add_802112 = sel_802109 + 8'h01;
  assign sel_802113 = array_index_801780 == array_index_773134 ? add_802112 : sel_802109;
  assign add_802116 = sel_802113 + 8'h01;
  assign sel_802117 = array_index_801780 == array_index_773140 ? add_802116 : sel_802113;
  assign add_802120 = sel_802117 + 8'h01;
  assign sel_802121 = array_index_801780 == array_index_773146 ? add_802120 : sel_802117;
  assign add_802124 = sel_802121 + 8'h01;
  assign sel_802125 = array_index_801780 == array_index_773152 ? add_802124 : sel_802121;
  assign add_802128 = sel_802125 + 8'h01;
  assign sel_802129 = array_index_801780 == array_index_773158 ? add_802128 : sel_802125;
  assign add_802132 = sel_802129 + 8'h01;
  assign sel_802133 = array_index_801780 == array_index_773164 ? add_802132 : sel_802129;
  assign add_802136 = sel_802133 + 8'h01;
  assign sel_802137 = array_index_801780 == array_index_773170 ? add_802136 : sel_802133;
  assign add_802141 = sel_802137 + 8'h01;
  assign array_index_802142 = set1_unflattened[7'h51];
  assign sel_802143 = array_index_801780 == array_index_773176 ? add_802141 : sel_802137;
  assign add_802146 = sel_802143 + 8'h01;
  assign sel_802147 = array_index_802142 == array_index_772632 ? add_802146 : sel_802143;
  assign add_802150 = sel_802147 + 8'h01;
  assign sel_802151 = array_index_802142 == array_index_772636 ? add_802150 : sel_802147;
  assign add_802154 = sel_802151 + 8'h01;
  assign sel_802155 = array_index_802142 == array_index_772644 ? add_802154 : sel_802151;
  assign add_802158 = sel_802155 + 8'h01;
  assign sel_802159 = array_index_802142 == array_index_772652 ? add_802158 : sel_802155;
  assign add_802162 = sel_802159 + 8'h01;
  assign sel_802163 = array_index_802142 == array_index_772660 ? add_802162 : sel_802159;
  assign add_802166 = sel_802163 + 8'h01;
  assign sel_802167 = array_index_802142 == array_index_772668 ? add_802166 : sel_802163;
  assign add_802170 = sel_802167 + 8'h01;
  assign sel_802171 = array_index_802142 == array_index_772676 ? add_802170 : sel_802167;
  assign add_802174 = sel_802171 + 8'h01;
  assign sel_802175 = array_index_802142 == array_index_772684 ? add_802174 : sel_802171;
  assign add_802178 = sel_802175 + 8'h01;
  assign sel_802179 = array_index_802142 == array_index_772690 ? add_802178 : sel_802175;
  assign add_802182 = sel_802179 + 8'h01;
  assign sel_802183 = array_index_802142 == array_index_772696 ? add_802182 : sel_802179;
  assign add_802186 = sel_802183 + 8'h01;
  assign sel_802187 = array_index_802142 == array_index_772702 ? add_802186 : sel_802183;
  assign add_802190 = sel_802187 + 8'h01;
  assign sel_802191 = array_index_802142 == array_index_772708 ? add_802190 : sel_802187;
  assign add_802194 = sel_802191 + 8'h01;
  assign sel_802195 = array_index_802142 == array_index_772714 ? add_802194 : sel_802191;
  assign add_802198 = sel_802195 + 8'h01;
  assign sel_802199 = array_index_802142 == array_index_772720 ? add_802198 : sel_802195;
  assign add_802202 = sel_802199 + 8'h01;
  assign sel_802203 = array_index_802142 == array_index_772726 ? add_802202 : sel_802199;
  assign add_802206 = sel_802203 + 8'h01;
  assign sel_802207 = array_index_802142 == array_index_772732 ? add_802206 : sel_802203;
  assign add_802210 = sel_802207 + 8'h01;
  assign sel_802211 = array_index_802142 == array_index_772738 ? add_802210 : sel_802207;
  assign add_802214 = sel_802211 + 8'h01;
  assign sel_802215 = array_index_802142 == array_index_772744 ? add_802214 : sel_802211;
  assign add_802218 = sel_802215 + 8'h01;
  assign sel_802219 = array_index_802142 == array_index_772750 ? add_802218 : sel_802215;
  assign add_802222 = sel_802219 + 8'h01;
  assign sel_802223 = array_index_802142 == array_index_772756 ? add_802222 : sel_802219;
  assign add_802226 = sel_802223 + 8'h01;
  assign sel_802227 = array_index_802142 == array_index_772762 ? add_802226 : sel_802223;
  assign add_802230 = sel_802227 + 8'h01;
  assign sel_802231 = array_index_802142 == array_index_772768 ? add_802230 : sel_802227;
  assign add_802234 = sel_802231 + 8'h01;
  assign sel_802235 = array_index_802142 == array_index_772774 ? add_802234 : sel_802231;
  assign add_802238 = sel_802235 + 8'h01;
  assign sel_802239 = array_index_802142 == array_index_772780 ? add_802238 : sel_802235;
  assign add_802242 = sel_802239 + 8'h01;
  assign sel_802243 = array_index_802142 == array_index_772786 ? add_802242 : sel_802239;
  assign add_802246 = sel_802243 + 8'h01;
  assign sel_802247 = array_index_802142 == array_index_772792 ? add_802246 : sel_802243;
  assign add_802250 = sel_802247 + 8'h01;
  assign sel_802251 = array_index_802142 == array_index_772798 ? add_802250 : sel_802247;
  assign add_802254 = sel_802251 + 8'h01;
  assign sel_802255 = array_index_802142 == array_index_772804 ? add_802254 : sel_802251;
  assign add_802258 = sel_802255 + 8'h01;
  assign sel_802259 = array_index_802142 == array_index_772810 ? add_802258 : sel_802255;
  assign add_802262 = sel_802259 + 8'h01;
  assign sel_802263 = array_index_802142 == array_index_772816 ? add_802262 : sel_802259;
  assign add_802266 = sel_802263 + 8'h01;
  assign sel_802267 = array_index_802142 == array_index_772822 ? add_802266 : sel_802263;
  assign add_802270 = sel_802267 + 8'h01;
  assign sel_802271 = array_index_802142 == array_index_772828 ? add_802270 : sel_802267;
  assign add_802274 = sel_802271 + 8'h01;
  assign sel_802275 = array_index_802142 == array_index_772834 ? add_802274 : sel_802271;
  assign add_802278 = sel_802275 + 8'h01;
  assign sel_802279 = array_index_802142 == array_index_772840 ? add_802278 : sel_802275;
  assign add_802282 = sel_802279 + 8'h01;
  assign sel_802283 = array_index_802142 == array_index_772846 ? add_802282 : sel_802279;
  assign add_802286 = sel_802283 + 8'h01;
  assign sel_802287 = array_index_802142 == array_index_772852 ? add_802286 : sel_802283;
  assign add_802290 = sel_802287 + 8'h01;
  assign sel_802291 = array_index_802142 == array_index_772858 ? add_802290 : sel_802287;
  assign add_802294 = sel_802291 + 8'h01;
  assign sel_802295 = array_index_802142 == array_index_772864 ? add_802294 : sel_802291;
  assign add_802298 = sel_802295 + 8'h01;
  assign sel_802299 = array_index_802142 == array_index_772870 ? add_802298 : sel_802295;
  assign add_802302 = sel_802299 + 8'h01;
  assign sel_802303 = array_index_802142 == array_index_772876 ? add_802302 : sel_802299;
  assign add_802306 = sel_802303 + 8'h01;
  assign sel_802307 = array_index_802142 == array_index_772882 ? add_802306 : sel_802303;
  assign add_802310 = sel_802307 + 8'h01;
  assign sel_802311 = array_index_802142 == array_index_772888 ? add_802310 : sel_802307;
  assign add_802314 = sel_802311 + 8'h01;
  assign sel_802315 = array_index_802142 == array_index_772894 ? add_802314 : sel_802311;
  assign add_802318 = sel_802315 + 8'h01;
  assign sel_802319 = array_index_802142 == array_index_772900 ? add_802318 : sel_802315;
  assign add_802322 = sel_802319 + 8'h01;
  assign sel_802323 = array_index_802142 == array_index_772906 ? add_802322 : sel_802319;
  assign add_802326 = sel_802323 + 8'h01;
  assign sel_802327 = array_index_802142 == array_index_772912 ? add_802326 : sel_802323;
  assign add_802330 = sel_802327 + 8'h01;
  assign sel_802331 = array_index_802142 == array_index_772918 ? add_802330 : sel_802327;
  assign add_802334 = sel_802331 + 8'h01;
  assign sel_802335 = array_index_802142 == array_index_772924 ? add_802334 : sel_802331;
  assign add_802338 = sel_802335 + 8'h01;
  assign sel_802339 = array_index_802142 == array_index_772930 ? add_802338 : sel_802335;
  assign add_802342 = sel_802339 + 8'h01;
  assign sel_802343 = array_index_802142 == array_index_772936 ? add_802342 : sel_802339;
  assign add_802346 = sel_802343 + 8'h01;
  assign sel_802347 = array_index_802142 == array_index_772942 ? add_802346 : sel_802343;
  assign add_802350 = sel_802347 + 8'h01;
  assign sel_802351 = array_index_802142 == array_index_772948 ? add_802350 : sel_802347;
  assign add_802354 = sel_802351 + 8'h01;
  assign sel_802355 = array_index_802142 == array_index_772954 ? add_802354 : sel_802351;
  assign add_802358 = sel_802355 + 8'h01;
  assign sel_802359 = array_index_802142 == array_index_772960 ? add_802358 : sel_802355;
  assign add_802362 = sel_802359 + 8'h01;
  assign sel_802363 = array_index_802142 == array_index_772966 ? add_802362 : sel_802359;
  assign add_802366 = sel_802363 + 8'h01;
  assign sel_802367 = array_index_802142 == array_index_772972 ? add_802366 : sel_802363;
  assign add_802370 = sel_802367 + 8'h01;
  assign sel_802371 = array_index_802142 == array_index_772978 ? add_802370 : sel_802367;
  assign add_802374 = sel_802371 + 8'h01;
  assign sel_802375 = array_index_802142 == array_index_772984 ? add_802374 : sel_802371;
  assign add_802378 = sel_802375 + 8'h01;
  assign sel_802379 = array_index_802142 == array_index_772990 ? add_802378 : sel_802375;
  assign add_802382 = sel_802379 + 8'h01;
  assign sel_802383 = array_index_802142 == array_index_772996 ? add_802382 : sel_802379;
  assign add_802386 = sel_802383 + 8'h01;
  assign sel_802387 = array_index_802142 == array_index_773002 ? add_802386 : sel_802383;
  assign add_802390 = sel_802387 + 8'h01;
  assign sel_802391 = array_index_802142 == array_index_773008 ? add_802390 : sel_802387;
  assign add_802394 = sel_802391 + 8'h01;
  assign sel_802395 = array_index_802142 == array_index_773014 ? add_802394 : sel_802391;
  assign add_802398 = sel_802395 + 8'h01;
  assign sel_802399 = array_index_802142 == array_index_773020 ? add_802398 : sel_802395;
  assign add_802402 = sel_802399 + 8'h01;
  assign sel_802403 = array_index_802142 == array_index_773026 ? add_802402 : sel_802399;
  assign add_802406 = sel_802403 + 8'h01;
  assign sel_802407 = array_index_802142 == array_index_773032 ? add_802406 : sel_802403;
  assign add_802410 = sel_802407 + 8'h01;
  assign sel_802411 = array_index_802142 == array_index_773038 ? add_802410 : sel_802407;
  assign add_802414 = sel_802411 + 8'h01;
  assign sel_802415 = array_index_802142 == array_index_773044 ? add_802414 : sel_802411;
  assign add_802418 = sel_802415 + 8'h01;
  assign sel_802419 = array_index_802142 == array_index_773050 ? add_802418 : sel_802415;
  assign add_802422 = sel_802419 + 8'h01;
  assign sel_802423 = array_index_802142 == array_index_773056 ? add_802422 : sel_802419;
  assign add_802426 = sel_802423 + 8'h01;
  assign sel_802427 = array_index_802142 == array_index_773062 ? add_802426 : sel_802423;
  assign add_802430 = sel_802427 + 8'h01;
  assign sel_802431 = array_index_802142 == array_index_773068 ? add_802430 : sel_802427;
  assign add_802434 = sel_802431 + 8'h01;
  assign sel_802435 = array_index_802142 == array_index_773074 ? add_802434 : sel_802431;
  assign add_802438 = sel_802435 + 8'h01;
  assign sel_802439 = array_index_802142 == array_index_773080 ? add_802438 : sel_802435;
  assign add_802442 = sel_802439 + 8'h01;
  assign sel_802443 = array_index_802142 == array_index_773086 ? add_802442 : sel_802439;
  assign add_802446 = sel_802443 + 8'h01;
  assign sel_802447 = array_index_802142 == array_index_773092 ? add_802446 : sel_802443;
  assign add_802450 = sel_802447 + 8'h01;
  assign sel_802451 = array_index_802142 == array_index_773098 ? add_802450 : sel_802447;
  assign add_802454 = sel_802451 + 8'h01;
  assign sel_802455 = array_index_802142 == array_index_773104 ? add_802454 : sel_802451;
  assign add_802458 = sel_802455 + 8'h01;
  assign sel_802459 = array_index_802142 == array_index_773110 ? add_802458 : sel_802455;
  assign add_802462 = sel_802459 + 8'h01;
  assign sel_802463 = array_index_802142 == array_index_773116 ? add_802462 : sel_802459;
  assign add_802466 = sel_802463 + 8'h01;
  assign sel_802467 = array_index_802142 == array_index_773122 ? add_802466 : sel_802463;
  assign add_802470 = sel_802467 + 8'h01;
  assign sel_802471 = array_index_802142 == array_index_773128 ? add_802470 : sel_802467;
  assign add_802474 = sel_802471 + 8'h01;
  assign sel_802475 = array_index_802142 == array_index_773134 ? add_802474 : sel_802471;
  assign add_802478 = sel_802475 + 8'h01;
  assign sel_802479 = array_index_802142 == array_index_773140 ? add_802478 : sel_802475;
  assign add_802482 = sel_802479 + 8'h01;
  assign sel_802483 = array_index_802142 == array_index_773146 ? add_802482 : sel_802479;
  assign add_802486 = sel_802483 + 8'h01;
  assign sel_802487 = array_index_802142 == array_index_773152 ? add_802486 : sel_802483;
  assign add_802490 = sel_802487 + 8'h01;
  assign sel_802491 = array_index_802142 == array_index_773158 ? add_802490 : sel_802487;
  assign add_802494 = sel_802491 + 8'h01;
  assign sel_802495 = array_index_802142 == array_index_773164 ? add_802494 : sel_802491;
  assign add_802498 = sel_802495 + 8'h01;
  assign sel_802499 = array_index_802142 == array_index_773170 ? add_802498 : sel_802495;
  assign add_802503 = sel_802499 + 8'h01;
  assign array_index_802504 = set1_unflattened[7'h52];
  assign sel_802505 = array_index_802142 == array_index_773176 ? add_802503 : sel_802499;
  assign add_802508 = sel_802505 + 8'h01;
  assign sel_802509 = array_index_802504 == array_index_772632 ? add_802508 : sel_802505;
  assign add_802512 = sel_802509 + 8'h01;
  assign sel_802513 = array_index_802504 == array_index_772636 ? add_802512 : sel_802509;
  assign add_802516 = sel_802513 + 8'h01;
  assign sel_802517 = array_index_802504 == array_index_772644 ? add_802516 : sel_802513;
  assign add_802520 = sel_802517 + 8'h01;
  assign sel_802521 = array_index_802504 == array_index_772652 ? add_802520 : sel_802517;
  assign add_802524 = sel_802521 + 8'h01;
  assign sel_802525 = array_index_802504 == array_index_772660 ? add_802524 : sel_802521;
  assign add_802528 = sel_802525 + 8'h01;
  assign sel_802529 = array_index_802504 == array_index_772668 ? add_802528 : sel_802525;
  assign add_802532 = sel_802529 + 8'h01;
  assign sel_802533 = array_index_802504 == array_index_772676 ? add_802532 : sel_802529;
  assign add_802536 = sel_802533 + 8'h01;
  assign sel_802537 = array_index_802504 == array_index_772684 ? add_802536 : sel_802533;
  assign add_802540 = sel_802537 + 8'h01;
  assign sel_802541 = array_index_802504 == array_index_772690 ? add_802540 : sel_802537;
  assign add_802544 = sel_802541 + 8'h01;
  assign sel_802545 = array_index_802504 == array_index_772696 ? add_802544 : sel_802541;
  assign add_802548 = sel_802545 + 8'h01;
  assign sel_802549 = array_index_802504 == array_index_772702 ? add_802548 : sel_802545;
  assign add_802552 = sel_802549 + 8'h01;
  assign sel_802553 = array_index_802504 == array_index_772708 ? add_802552 : sel_802549;
  assign add_802556 = sel_802553 + 8'h01;
  assign sel_802557 = array_index_802504 == array_index_772714 ? add_802556 : sel_802553;
  assign add_802560 = sel_802557 + 8'h01;
  assign sel_802561 = array_index_802504 == array_index_772720 ? add_802560 : sel_802557;
  assign add_802564 = sel_802561 + 8'h01;
  assign sel_802565 = array_index_802504 == array_index_772726 ? add_802564 : sel_802561;
  assign add_802568 = sel_802565 + 8'h01;
  assign sel_802569 = array_index_802504 == array_index_772732 ? add_802568 : sel_802565;
  assign add_802572 = sel_802569 + 8'h01;
  assign sel_802573 = array_index_802504 == array_index_772738 ? add_802572 : sel_802569;
  assign add_802576 = sel_802573 + 8'h01;
  assign sel_802577 = array_index_802504 == array_index_772744 ? add_802576 : sel_802573;
  assign add_802580 = sel_802577 + 8'h01;
  assign sel_802581 = array_index_802504 == array_index_772750 ? add_802580 : sel_802577;
  assign add_802584 = sel_802581 + 8'h01;
  assign sel_802585 = array_index_802504 == array_index_772756 ? add_802584 : sel_802581;
  assign add_802588 = sel_802585 + 8'h01;
  assign sel_802589 = array_index_802504 == array_index_772762 ? add_802588 : sel_802585;
  assign add_802592 = sel_802589 + 8'h01;
  assign sel_802593 = array_index_802504 == array_index_772768 ? add_802592 : sel_802589;
  assign add_802596 = sel_802593 + 8'h01;
  assign sel_802597 = array_index_802504 == array_index_772774 ? add_802596 : sel_802593;
  assign add_802600 = sel_802597 + 8'h01;
  assign sel_802601 = array_index_802504 == array_index_772780 ? add_802600 : sel_802597;
  assign add_802604 = sel_802601 + 8'h01;
  assign sel_802605 = array_index_802504 == array_index_772786 ? add_802604 : sel_802601;
  assign add_802608 = sel_802605 + 8'h01;
  assign sel_802609 = array_index_802504 == array_index_772792 ? add_802608 : sel_802605;
  assign add_802612 = sel_802609 + 8'h01;
  assign sel_802613 = array_index_802504 == array_index_772798 ? add_802612 : sel_802609;
  assign add_802616 = sel_802613 + 8'h01;
  assign sel_802617 = array_index_802504 == array_index_772804 ? add_802616 : sel_802613;
  assign add_802620 = sel_802617 + 8'h01;
  assign sel_802621 = array_index_802504 == array_index_772810 ? add_802620 : sel_802617;
  assign add_802624 = sel_802621 + 8'h01;
  assign sel_802625 = array_index_802504 == array_index_772816 ? add_802624 : sel_802621;
  assign add_802628 = sel_802625 + 8'h01;
  assign sel_802629 = array_index_802504 == array_index_772822 ? add_802628 : sel_802625;
  assign add_802632 = sel_802629 + 8'h01;
  assign sel_802633 = array_index_802504 == array_index_772828 ? add_802632 : sel_802629;
  assign add_802636 = sel_802633 + 8'h01;
  assign sel_802637 = array_index_802504 == array_index_772834 ? add_802636 : sel_802633;
  assign add_802640 = sel_802637 + 8'h01;
  assign sel_802641 = array_index_802504 == array_index_772840 ? add_802640 : sel_802637;
  assign add_802644 = sel_802641 + 8'h01;
  assign sel_802645 = array_index_802504 == array_index_772846 ? add_802644 : sel_802641;
  assign add_802648 = sel_802645 + 8'h01;
  assign sel_802649 = array_index_802504 == array_index_772852 ? add_802648 : sel_802645;
  assign add_802652 = sel_802649 + 8'h01;
  assign sel_802653 = array_index_802504 == array_index_772858 ? add_802652 : sel_802649;
  assign add_802656 = sel_802653 + 8'h01;
  assign sel_802657 = array_index_802504 == array_index_772864 ? add_802656 : sel_802653;
  assign add_802660 = sel_802657 + 8'h01;
  assign sel_802661 = array_index_802504 == array_index_772870 ? add_802660 : sel_802657;
  assign add_802664 = sel_802661 + 8'h01;
  assign sel_802665 = array_index_802504 == array_index_772876 ? add_802664 : sel_802661;
  assign add_802668 = sel_802665 + 8'h01;
  assign sel_802669 = array_index_802504 == array_index_772882 ? add_802668 : sel_802665;
  assign add_802672 = sel_802669 + 8'h01;
  assign sel_802673 = array_index_802504 == array_index_772888 ? add_802672 : sel_802669;
  assign add_802676 = sel_802673 + 8'h01;
  assign sel_802677 = array_index_802504 == array_index_772894 ? add_802676 : sel_802673;
  assign add_802680 = sel_802677 + 8'h01;
  assign sel_802681 = array_index_802504 == array_index_772900 ? add_802680 : sel_802677;
  assign add_802684 = sel_802681 + 8'h01;
  assign sel_802685 = array_index_802504 == array_index_772906 ? add_802684 : sel_802681;
  assign add_802688 = sel_802685 + 8'h01;
  assign sel_802689 = array_index_802504 == array_index_772912 ? add_802688 : sel_802685;
  assign add_802692 = sel_802689 + 8'h01;
  assign sel_802693 = array_index_802504 == array_index_772918 ? add_802692 : sel_802689;
  assign add_802696 = sel_802693 + 8'h01;
  assign sel_802697 = array_index_802504 == array_index_772924 ? add_802696 : sel_802693;
  assign add_802700 = sel_802697 + 8'h01;
  assign sel_802701 = array_index_802504 == array_index_772930 ? add_802700 : sel_802697;
  assign add_802704 = sel_802701 + 8'h01;
  assign sel_802705 = array_index_802504 == array_index_772936 ? add_802704 : sel_802701;
  assign add_802708 = sel_802705 + 8'h01;
  assign sel_802709 = array_index_802504 == array_index_772942 ? add_802708 : sel_802705;
  assign add_802712 = sel_802709 + 8'h01;
  assign sel_802713 = array_index_802504 == array_index_772948 ? add_802712 : sel_802709;
  assign add_802716 = sel_802713 + 8'h01;
  assign sel_802717 = array_index_802504 == array_index_772954 ? add_802716 : sel_802713;
  assign add_802720 = sel_802717 + 8'h01;
  assign sel_802721 = array_index_802504 == array_index_772960 ? add_802720 : sel_802717;
  assign add_802724 = sel_802721 + 8'h01;
  assign sel_802725 = array_index_802504 == array_index_772966 ? add_802724 : sel_802721;
  assign add_802728 = sel_802725 + 8'h01;
  assign sel_802729 = array_index_802504 == array_index_772972 ? add_802728 : sel_802725;
  assign add_802732 = sel_802729 + 8'h01;
  assign sel_802733 = array_index_802504 == array_index_772978 ? add_802732 : sel_802729;
  assign add_802736 = sel_802733 + 8'h01;
  assign sel_802737 = array_index_802504 == array_index_772984 ? add_802736 : sel_802733;
  assign add_802740 = sel_802737 + 8'h01;
  assign sel_802741 = array_index_802504 == array_index_772990 ? add_802740 : sel_802737;
  assign add_802744 = sel_802741 + 8'h01;
  assign sel_802745 = array_index_802504 == array_index_772996 ? add_802744 : sel_802741;
  assign add_802748 = sel_802745 + 8'h01;
  assign sel_802749 = array_index_802504 == array_index_773002 ? add_802748 : sel_802745;
  assign add_802752 = sel_802749 + 8'h01;
  assign sel_802753 = array_index_802504 == array_index_773008 ? add_802752 : sel_802749;
  assign add_802756 = sel_802753 + 8'h01;
  assign sel_802757 = array_index_802504 == array_index_773014 ? add_802756 : sel_802753;
  assign add_802760 = sel_802757 + 8'h01;
  assign sel_802761 = array_index_802504 == array_index_773020 ? add_802760 : sel_802757;
  assign add_802764 = sel_802761 + 8'h01;
  assign sel_802765 = array_index_802504 == array_index_773026 ? add_802764 : sel_802761;
  assign add_802768 = sel_802765 + 8'h01;
  assign sel_802769 = array_index_802504 == array_index_773032 ? add_802768 : sel_802765;
  assign add_802772 = sel_802769 + 8'h01;
  assign sel_802773 = array_index_802504 == array_index_773038 ? add_802772 : sel_802769;
  assign add_802776 = sel_802773 + 8'h01;
  assign sel_802777 = array_index_802504 == array_index_773044 ? add_802776 : sel_802773;
  assign add_802780 = sel_802777 + 8'h01;
  assign sel_802781 = array_index_802504 == array_index_773050 ? add_802780 : sel_802777;
  assign add_802784 = sel_802781 + 8'h01;
  assign sel_802785 = array_index_802504 == array_index_773056 ? add_802784 : sel_802781;
  assign add_802788 = sel_802785 + 8'h01;
  assign sel_802789 = array_index_802504 == array_index_773062 ? add_802788 : sel_802785;
  assign add_802792 = sel_802789 + 8'h01;
  assign sel_802793 = array_index_802504 == array_index_773068 ? add_802792 : sel_802789;
  assign add_802796 = sel_802793 + 8'h01;
  assign sel_802797 = array_index_802504 == array_index_773074 ? add_802796 : sel_802793;
  assign add_802800 = sel_802797 + 8'h01;
  assign sel_802801 = array_index_802504 == array_index_773080 ? add_802800 : sel_802797;
  assign add_802804 = sel_802801 + 8'h01;
  assign sel_802805 = array_index_802504 == array_index_773086 ? add_802804 : sel_802801;
  assign add_802808 = sel_802805 + 8'h01;
  assign sel_802809 = array_index_802504 == array_index_773092 ? add_802808 : sel_802805;
  assign add_802812 = sel_802809 + 8'h01;
  assign sel_802813 = array_index_802504 == array_index_773098 ? add_802812 : sel_802809;
  assign add_802816 = sel_802813 + 8'h01;
  assign sel_802817 = array_index_802504 == array_index_773104 ? add_802816 : sel_802813;
  assign add_802820 = sel_802817 + 8'h01;
  assign sel_802821 = array_index_802504 == array_index_773110 ? add_802820 : sel_802817;
  assign add_802824 = sel_802821 + 8'h01;
  assign sel_802825 = array_index_802504 == array_index_773116 ? add_802824 : sel_802821;
  assign add_802828 = sel_802825 + 8'h01;
  assign sel_802829 = array_index_802504 == array_index_773122 ? add_802828 : sel_802825;
  assign add_802832 = sel_802829 + 8'h01;
  assign sel_802833 = array_index_802504 == array_index_773128 ? add_802832 : sel_802829;
  assign add_802836 = sel_802833 + 8'h01;
  assign sel_802837 = array_index_802504 == array_index_773134 ? add_802836 : sel_802833;
  assign add_802840 = sel_802837 + 8'h01;
  assign sel_802841 = array_index_802504 == array_index_773140 ? add_802840 : sel_802837;
  assign add_802844 = sel_802841 + 8'h01;
  assign sel_802845 = array_index_802504 == array_index_773146 ? add_802844 : sel_802841;
  assign add_802848 = sel_802845 + 8'h01;
  assign sel_802849 = array_index_802504 == array_index_773152 ? add_802848 : sel_802845;
  assign add_802852 = sel_802849 + 8'h01;
  assign sel_802853 = array_index_802504 == array_index_773158 ? add_802852 : sel_802849;
  assign add_802856 = sel_802853 + 8'h01;
  assign sel_802857 = array_index_802504 == array_index_773164 ? add_802856 : sel_802853;
  assign add_802860 = sel_802857 + 8'h01;
  assign sel_802861 = array_index_802504 == array_index_773170 ? add_802860 : sel_802857;
  assign add_802865 = sel_802861 + 8'h01;
  assign array_index_802866 = set1_unflattened[7'h53];
  assign sel_802867 = array_index_802504 == array_index_773176 ? add_802865 : sel_802861;
  assign add_802870 = sel_802867 + 8'h01;
  assign sel_802871 = array_index_802866 == array_index_772632 ? add_802870 : sel_802867;
  assign add_802874 = sel_802871 + 8'h01;
  assign sel_802875 = array_index_802866 == array_index_772636 ? add_802874 : sel_802871;
  assign add_802878 = sel_802875 + 8'h01;
  assign sel_802879 = array_index_802866 == array_index_772644 ? add_802878 : sel_802875;
  assign add_802882 = sel_802879 + 8'h01;
  assign sel_802883 = array_index_802866 == array_index_772652 ? add_802882 : sel_802879;
  assign add_802886 = sel_802883 + 8'h01;
  assign sel_802887 = array_index_802866 == array_index_772660 ? add_802886 : sel_802883;
  assign add_802890 = sel_802887 + 8'h01;
  assign sel_802891 = array_index_802866 == array_index_772668 ? add_802890 : sel_802887;
  assign add_802894 = sel_802891 + 8'h01;
  assign sel_802895 = array_index_802866 == array_index_772676 ? add_802894 : sel_802891;
  assign add_802898 = sel_802895 + 8'h01;
  assign sel_802899 = array_index_802866 == array_index_772684 ? add_802898 : sel_802895;
  assign add_802902 = sel_802899 + 8'h01;
  assign sel_802903 = array_index_802866 == array_index_772690 ? add_802902 : sel_802899;
  assign add_802906 = sel_802903 + 8'h01;
  assign sel_802907 = array_index_802866 == array_index_772696 ? add_802906 : sel_802903;
  assign add_802910 = sel_802907 + 8'h01;
  assign sel_802911 = array_index_802866 == array_index_772702 ? add_802910 : sel_802907;
  assign add_802914 = sel_802911 + 8'h01;
  assign sel_802915 = array_index_802866 == array_index_772708 ? add_802914 : sel_802911;
  assign add_802918 = sel_802915 + 8'h01;
  assign sel_802919 = array_index_802866 == array_index_772714 ? add_802918 : sel_802915;
  assign add_802922 = sel_802919 + 8'h01;
  assign sel_802923 = array_index_802866 == array_index_772720 ? add_802922 : sel_802919;
  assign add_802926 = sel_802923 + 8'h01;
  assign sel_802927 = array_index_802866 == array_index_772726 ? add_802926 : sel_802923;
  assign add_802930 = sel_802927 + 8'h01;
  assign sel_802931 = array_index_802866 == array_index_772732 ? add_802930 : sel_802927;
  assign add_802934 = sel_802931 + 8'h01;
  assign sel_802935 = array_index_802866 == array_index_772738 ? add_802934 : sel_802931;
  assign add_802938 = sel_802935 + 8'h01;
  assign sel_802939 = array_index_802866 == array_index_772744 ? add_802938 : sel_802935;
  assign add_802942 = sel_802939 + 8'h01;
  assign sel_802943 = array_index_802866 == array_index_772750 ? add_802942 : sel_802939;
  assign add_802946 = sel_802943 + 8'h01;
  assign sel_802947 = array_index_802866 == array_index_772756 ? add_802946 : sel_802943;
  assign add_802950 = sel_802947 + 8'h01;
  assign sel_802951 = array_index_802866 == array_index_772762 ? add_802950 : sel_802947;
  assign add_802954 = sel_802951 + 8'h01;
  assign sel_802955 = array_index_802866 == array_index_772768 ? add_802954 : sel_802951;
  assign add_802958 = sel_802955 + 8'h01;
  assign sel_802959 = array_index_802866 == array_index_772774 ? add_802958 : sel_802955;
  assign add_802962 = sel_802959 + 8'h01;
  assign sel_802963 = array_index_802866 == array_index_772780 ? add_802962 : sel_802959;
  assign add_802966 = sel_802963 + 8'h01;
  assign sel_802967 = array_index_802866 == array_index_772786 ? add_802966 : sel_802963;
  assign add_802970 = sel_802967 + 8'h01;
  assign sel_802971 = array_index_802866 == array_index_772792 ? add_802970 : sel_802967;
  assign add_802974 = sel_802971 + 8'h01;
  assign sel_802975 = array_index_802866 == array_index_772798 ? add_802974 : sel_802971;
  assign add_802978 = sel_802975 + 8'h01;
  assign sel_802979 = array_index_802866 == array_index_772804 ? add_802978 : sel_802975;
  assign add_802982 = sel_802979 + 8'h01;
  assign sel_802983 = array_index_802866 == array_index_772810 ? add_802982 : sel_802979;
  assign add_802986 = sel_802983 + 8'h01;
  assign sel_802987 = array_index_802866 == array_index_772816 ? add_802986 : sel_802983;
  assign add_802990 = sel_802987 + 8'h01;
  assign sel_802991 = array_index_802866 == array_index_772822 ? add_802990 : sel_802987;
  assign add_802994 = sel_802991 + 8'h01;
  assign sel_802995 = array_index_802866 == array_index_772828 ? add_802994 : sel_802991;
  assign add_802998 = sel_802995 + 8'h01;
  assign sel_802999 = array_index_802866 == array_index_772834 ? add_802998 : sel_802995;
  assign add_803002 = sel_802999 + 8'h01;
  assign sel_803003 = array_index_802866 == array_index_772840 ? add_803002 : sel_802999;
  assign add_803006 = sel_803003 + 8'h01;
  assign sel_803007 = array_index_802866 == array_index_772846 ? add_803006 : sel_803003;
  assign add_803010 = sel_803007 + 8'h01;
  assign sel_803011 = array_index_802866 == array_index_772852 ? add_803010 : sel_803007;
  assign add_803014 = sel_803011 + 8'h01;
  assign sel_803015 = array_index_802866 == array_index_772858 ? add_803014 : sel_803011;
  assign add_803018 = sel_803015 + 8'h01;
  assign sel_803019 = array_index_802866 == array_index_772864 ? add_803018 : sel_803015;
  assign add_803022 = sel_803019 + 8'h01;
  assign sel_803023 = array_index_802866 == array_index_772870 ? add_803022 : sel_803019;
  assign add_803026 = sel_803023 + 8'h01;
  assign sel_803027 = array_index_802866 == array_index_772876 ? add_803026 : sel_803023;
  assign add_803030 = sel_803027 + 8'h01;
  assign sel_803031 = array_index_802866 == array_index_772882 ? add_803030 : sel_803027;
  assign add_803034 = sel_803031 + 8'h01;
  assign sel_803035 = array_index_802866 == array_index_772888 ? add_803034 : sel_803031;
  assign add_803038 = sel_803035 + 8'h01;
  assign sel_803039 = array_index_802866 == array_index_772894 ? add_803038 : sel_803035;
  assign add_803042 = sel_803039 + 8'h01;
  assign sel_803043 = array_index_802866 == array_index_772900 ? add_803042 : sel_803039;
  assign add_803046 = sel_803043 + 8'h01;
  assign sel_803047 = array_index_802866 == array_index_772906 ? add_803046 : sel_803043;
  assign add_803050 = sel_803047 + 8'h01;
  assign sel_803051 = array_index_802866 == array_index_772912 ? add_803050 : sel_803047;
  assign add_803054 = sel_803051 + 8'h01;
  assign sel_803055 = array_index_802866 == array_index_772918 ? add_803054 : sel_803051;
  assign add_803058 = sel_803055 + 8'h01;
  assign sel_803059 = array_index_802866 == array_index_772924 ? add_803058 : sel_803055;
  assign add_803062 = sel_803059 + 8'h01;
  assign sel_803063 = array_index_802866 == array_index_772930 ? add_803062 : sel_803059;
  assign add_803066 = sel_803063 + 8'h01;
  assign sel_803067 = array_index_802866 == array_index_772936 ? add_803066 : sel_803063;
  assign add_803070 = sel_803067 + 8'h01;
  assign sel_803071 = array_index_802866 == array_index_772942 ? add_803070 : sel_803067;
  assign add_803074 = sel_803071 + 8'h01;
  assign sel_803075 = array_index_802866 == array_index_772948 ? add_803074 : sel_803071;
  assign add_803078 = sel_803075 + 8'h01;
  assign sel_803079 = array_index_802866 == array_index_772954 ? add_803078 : sel_803075;
  assign add_803082 = sel_803079 + 8'h01;
  assign sel_803083 = array_index_802866 == array_index_772960 ? add_803082 : sel_803079;
  assign add_803086 = sel_803083 + 8'h01;
  assign sel_803087 = array_index_802866 == array_index_772966 ? add_803086 : sel_803083;
  assign add_803090 = sel_803087 + 8'h01;
  assign sel_803091 = array_index_802866 == array_index_772972 ? add_803090 : sel_803087;
  assign add_803094 = sel_803091 + 8'h01;
  assign sel_803095 = array_index_802866 == array_index_772978 ? add_803094 : sel_803091;
  assign add_803098 = sel_803095 + 8'h01;
  assign sel_803099 = array_index_802866 == array_index_772984 ? add_803098 : sel_803095;
  assign add_803102 = sel_803099 + 8'h01;
  assign sel_803103 = array_index_802866 == array_index_772990 ? add_803102 : sel_803099;
  assign add_803106 = sel_803103 + 8'h01;
  assign sel_803107 = array_index_802866 == array_index_772996 ? add_803106 : sel_803103;
  assign add_803110 = sel_803107 + 8'h01;
  assign sel_803111 = array_index_802866 == array_index_773002 ? add_803110 : sel_803107;
  assign add_803114 = sel_803111 + 8'h01;
  assign sel_803115 = array_index_802866 == array_index_773008 ? add_803114 : sel_803111;
  assign add_803118 = sel_803115 + 8'h01;
  assign sel_803119 = array_index_802866 == array_index_773014 ? add_803118 : sel_803115;
  assign add_803122 = sel_803119 + 8'h01;
  assign sel_803123 = array_index_802866 == array_index_773020 ? add_803122 : sel_803119;
  assign add_803126 = sel_803123 + 8'h01;
  assign sel_803127 = array_index_802866 == array_index_773026 ? add_803126 : sel_803123;
  assign add_803130 = sel_803127 + 8'h01;
  assign sel_803131 = array_index_802866 == array_index_773032 ? add_803130 : sel_803127;
  assign add_803134 = sel_803131 + 8'h01;
  assign sel_803135 = array_index_802866 == array_index_773038 ? add_803134 : sel_803131;
  assign add_803138 = sel_803135 + 8'h01;
  assign sel_803139 = array_index_802866 == array_index_773044 ? add_803138 : sel_803135;
  assign add_803142 = sel_803139 + 8'h01;
  assign sel_803143 = array_index_802866 == array_index_773050 ? add_803142 : sel_803139;
  assign add_803146 = sel_803143 + 8'h01;
  assign sel_803147 = array_index_802866 == array_index_773056 ? add_803146 : sel_803143;
  assign add_803150 = sel_803147 + 8'h01;
  assign sel_803151 = array_index_802866 == array_index_773062 ? add_803150 : sel_803147;
  assign add_803154 = sel_803151 + 8'h01;
  assign sel_803155 = array_index_802866 == array_index_773068 ? add_803154 : sel_803151;
  assign add_803158 = sel_803155 + 8'h01;
  assign sel_803159 = array_index_802866 == array_index_773074 ? add_803158 : sel_803155;
  assign add_803162 = sel_803159 + 8'h01;
  assign sel_803163 = array_index_802866 == array_index_773080 ? add_803162 : sel_803159;
  assign add_803166 = sel_803163 + 8'h01;
  assign sel_803167 = array_index_802866 == array_index_773086 ? add_803166 : sel_803163;
  assign add_803170 = sel_803167 + 8'h01;
  assign sel_803171 = array_index_802866 == array_index_773092 ? add_803170 : sel_803167;
  assign add_803174 = sel_803171 + 8'h01;
  assign sel_803175 = array_index_802866 == array_index_773098 ? add_803174 : sel_803171;
  assign add_803178 = sel_803175 + 8'h01;
  assign sel_803179 = array_index_802866 == array_index_773104 ? add_803178 : sel_803175;
  assign add_803182 = sel_803179 + 8'h01;
  assign sel_803183 = array_index_802866 == array_index_773110 ? add_803182 : sel_803179;
  assign add_803186 = sel_803183 + 8'h01;
  assign sel_803187 = array_index_802866 == array_index_773116 ? add_803186 : sel_803183;
  assign add_803190 = sel_803187 + 8'h01;
  assign sel_803191 = array_index_802866 == array_index_773122 ? add_803190 : sel_803187;
  assign add_803194 = sel_803191 + 8'h01;
  assign sel_803195 = array_index_802866 == array_index_773128 ? add_803194 : sel_803191;
  assign add_803198 = sel_803195 + 8'h01;
  assign sel_803199 = array_index_802866 == array_index_773134 ? add_803198 : sel_803195;
  assign add_803202 = sel_803199 + 8'h01;
  assign sel_803203 = array_index_802866 == array_index_773140 ? add_803202 : sel_803199;
  assign add_803206 = sel_803203 + 8'h01;
  assign sel_803207 = array_index_802866 == array_index_773146 ? add_803206 : sel_803203;
  assign add_803210 = sel_803207 + 8'h01;
  assign sel_803211 = array_index_802866 == array_index_773152 ? add_803210 : sel_803207;
  assign add_803214 = sel_803211 + 8'h01;
  assign sel_803215 = array_index_802866 == array_index_773158 ? add_803214 : sel_803211;
  assign add_803218 = sel_803215 + 8'h01;
  assign sel_803219 = array_index_802866 == array_index_773164 ? add_803218 : sel_803215;
  assign add_803222 = sel_803219 + 8'h01;
  assign sel_803223 = array_index_802866 == array_index_773170 ? add_803222 : sel_803219;
  assign add_803227 = sel_803223 + 8'h01;
  assign array_index_803228 = set1_unflattened[7'h54];
  assign sel_803229 = array_index_802866 == array_index_773176 ? add_803227 : sel_803223;
  assign add_803232 = sel_803229 + 8'h01;
  assign sel_803233 = array_index_803228 == array_index_772632 ? add_803232 : sel_803229;
  assign add_803236 = sel_803233 + 8'h01;
  assign sel_803237 = array_index_803228 == array_index_772636 ? add_803236 : sel_803233;
  assign add_803240 = sel_803237 + 8'h01;
  assign sel_803241 = array_index_803228 == array_index_772644 ? add_803240 : sel_803237;
  assign add_803244 = sel_803241 + 8'h01;
  assign sel_803245 = array_index_803228 == array_index_772652 ? add_803244 : sel_803241;
  assign add_803248 = sel_803245 + 8'h01;
  assign sel_803249 = array_index_803228 == array_index_772660 ? add_803248 : sel_803245;
  assign add_803252 = sel_803249 + 8'h01;
  assign sel_803253 = array_index_803228 == array_index_772668 ? add_803252 : sel_803249;
  assign add_803256 = sel_803253 + 8'h01;
  assign sel_803257 = array_index_803228 == array_index_772676 ? add_803256 : sel_803253;
  assign add_803260 = sel_803257 + 8'h01;
  assign sel_803261 = array_index_803228 == array_index_772684 ? add_803260 : sel_803257;
  assign add_803264 = sel_803261 + 8'h01;
  assign sel_803265 = array_index_803228 == array_index_772690 ? add_803264 : sel_803261;
  assign add_803268 = sel_803265 + 8'h01;
  assign sel_803269 = array_index_803228 == array_index_772696 ? add_803268 : sel_803265;
  assign add_803272 = sel_803269 + 8'h01;
  assign sel_803273 = array_index_803228 == array_index_772702 ? add_803272 : sel_803269;
  assign add_803276 = sel_803273 + 8'h01;
  assign sel_803277 = array_index_803228 == array_index_772708 ? add_803276 : sel_803273;
  assign add_803280 = sel_803277 + 8'h01;
  assign sel_803281 = array_index_803228 == array_index_772714 ? add_803280 : sel_803277;
  assign add_803284 = sel_803281 + 8'h01;
  assign sel_803285 = array_index_803228 == array_index_772720 ? add_803284 : sel_803281;
  assign add_803288 = sel_803285 + 8'h01;
  assign sel_803289 = array_index_803228 == array_index_772726 ? add_803288 : sel_803285;
  assign add_803292 = sel_803289 + 8'h01;
  assign sel_803293 = array_index_803228 == array_index_772732 ? add_803292 : sel_803289;
  assign add_803296 = sel_803293 + 8'h01;
  assign sel_803297 = array_index_803228 == array_index_772738 ? add_803296 : sel_803293;
  assign add_803300 = sel_803297 + 8'h01;
  assign sel_803301 = array_index_803228 == array_index_772744 ? add_803300 : sel_803297;
  assign add_803304 = sel_803301 + 8'h01;
  assign sel_803305 = array_index_803228 == array_index_772750 ? add_803304 : sel_803301;
  assign add_803308 = sel_803305 + 8'h01;
  assign sel_803309 = array_index_803228 == array_index_772756 ? add_803308 : sel_803305;
  assign add_803312 = sel_803309 + 8'h01;
  assign sel_803313 = array_index_803228 == array_index_772762 ? add_803312 : sel_803309;
  assign add_803316 = sel_803313 + 8'h01;
  assign sel_803317 = array_index_803228 == array_index_772768 ? add_803316 : sel_803313;
  assign add_803320 = sel_803317 + 8'h01;
  assign sel_803321 = array_index_803228 == array_index_772774 ? add_803320 : sel_803317;
  assign add_803324 = sel_803321 + 8'h01;
  assign sel_803325 = array_index_803228 == array_index_772780 ? add_803324 : sel_803321;
  assign add_803328 = sel_803325 + 8'h01;
  assign sel_803329 = array_index_803228 == array_index_772786 ? add_803328 : sel_803325;
  assign add_803332 = sel_803329 + 8'h01;
  assign sel_803333 = array_index_803228 == array_index_772792 ? add_803332 : sel_803329;
  assign add_803336 = sel_803333 + 8'h01;
  assign sel_803337 = array_index_803228 == array_index_772798 ? add_803336 : sel_803333;
  assign add_803340 = sel_803337 + 8'h01;
  assign sel_803341 = array_index_803228 == array_index_772804 ? add_803340 : sel_803337;
  assign add_803344 = sel_803341 + 8'h01;
  assign sel_803345 = array_index_803228 == array_index_772810 ? add_803344 : sel_803341;
  assign add_803348 = sel_803345 + 8'h01;
  assign sel_803349 = array_index_803228 == array_index_772816 ? add_803348 : sel_803345;
  assign add_803352 = sel_803349 + 8'h01;
  assign sel_803353 = array_index_803228 == array_index_772822 ? add_803352 : sel_803349;
  assign add_803356 = sel_803353 + 8'h01;
  assign sel_803357 = array_index_803228 == array_index_772828 ? add_803356 : sel_803353;
  assign add_803360 = sel_803357 + 8'h01;
  assign sel_803361 = array_index_803228 == array_index_772834 ? add_803360 : sel_803357;
  assign add_803364 = sel_803361 + 8'h01;
  assign sel_803365 = array_index_803228 == array_index_772840 ? add_803364 : sel_803361;
  assign add_803368 = sel_803365 + 8'h01;
  assign sel_803369 = array_index_803228 == array_index_772846 ? add_803368 : sel_803365;
  assign add_803372 = sel_803369 + 8'h01;
  assign sel_803373 = array_index_803228 == array_index_772852 ? add_803372 : sel_803369;
  assign add_803376 = sel_803373 + 8'h01;
  assign sel_803377 = array_index_803228 == array_index_772858 ? add_803376 : sel_803373;
  assign add_803380 = sel_803377 + 8'h01;
  assign sel_803381 = array_index_803228 == array_index_772864 ? add_803380 : sel_803377;
  assign add_803384 = sel_803381 + 8'h01;
  assign sel_803385 = array_index_803228 == array_index_772870 ? add_803384 : sel_803381;
  assign add_803388 = sel_803385 + 8'h01;
  assign sel_803389 = array_index_803228 == array_index_772876 ? add_803388 : sel_803385;
  assign add_803392 = sel_803389 + 8'h01;
  assign sel_803393 = array_index_803228 == array_index_772882 ? add_803392 : sel_803389;
  assign add_803396 = sel_803393 + 8'h01;
  assign sel_803397 = array_index_803228 == array_index_772888 ? add_803396 : sel_803393;
  assign add_803400 = sel_803397 + 8'h01;
  assign sel_803401 = array_index_803228 == array_index_772894 ? add_803400 : sel_803397;
  assign add_803404 = sel_803401 + 8'h01;
  assign sel_803405 = array_index_803228 == array_index_772900 ? add_803404 : sel_803401;
  assign add_803408 = sel_803405 + 8'h01;
  assign sel_803409 = array_index_803228 == array_index_772906 ? add_803408 : sel_803405;
  assign add_803412 = sel_803409 + 8'h01;
  assign sel_803413 = array_index_803228 == array_index_772912 ? add_803412 : sel_803409;
  assign add_803416 = sel_803413 + 8'h01;
  assign sel_803417 = array_index_803228 == array_index_772918 ? add_803416 : sel_803413;
  assign add_803420 = sel_803417 + 8'h01;
  assign sel_803421 = array_index_803228 == array_index_772924 ? add_803420 : sel_803417;
  assign add_803424 = sel_803421 + 8'h01;
  assign sel_803425 = array_index_803228 == array_index_772930 ? add_803424 : sel_803421;
  assign add_803428 = sel_803425 + 8'h01;
  assign sel_803429 = array_index_803228 == array_index_772936 ? add_803428 : sel_803425;
  assign add_803432 = sel_803429 + 8'h01;
  assign sel_803433 = array_index_803228 == array_index_772942 ? add_803432 : sel_803429;
  assign add_803436 = sel_803433 + 8'h01;
  assign sel_803437 = array_index_803228 == array_index_772948 ? add_803436 : sel_803433;
  assign add_803440 = sel_803437 + 8'h01;
  assign sel_803441 = array_index_803228 == array_index_772954 ? add_803440 : sel_803437;
  assign add_803444 = sel_803441 + 8'h01;
  assign sel_803445 = array_index_803228 == array_index_772960 ? add_803444 : sel_803441;
  assign add_803448 = sel_803445 + 8'h01;
  assign sel_803449 = array_index_803228 == array_index_772966 ? add_803448 : sel_803445;
  assign add_803452 = sel_803449 + 8'h01;
  assign sel_803453 = array_index_803228 == array_index_772972 ? add_803452 : sel_803449;
  assign add_803456 = sel_803453 + 8'h01;
  assign sel_803457 = array_index_803228 == array_index_772978 ? add_803456 : sel_803453;
  assign add_803460 = sel_803457 + 8'h01;
  assign sel_803461 = array_index_803228 == array_index_772984 ? add_803460 : sel_803457;
  assign add_803464 = sel_803461 + 8'h01;
  assign sel_803465 = array_index_803228 == array_index_772990 ? add_803464 : sel_803461;
  assign add_803468 = sel_803465 + 8'h01;
  assign sel_803469 = array_index_803228 == array_index_772996 ? add_803468 : sel_803465;
  assign add_803472 = sel_803469 + 8'h01;
  assign sel_803473 = array_index_803228 == array_index_773002 ? add_803472 : sel_803469;
  assign add_803476 = sel_803473 + 8'h01;
  assign sel_803477 = array_index_803228 == array_index_773008 ? add_803476 : sel_803473;
  assign add_803480 = sel_803477 + 8'h01;
  assign sel_803481 = array_index_803228 == array_index_773014 ? add_803480 : sel_803477;
  assign add_803484 = sel_803481 + 8'h01;
  assign sel_803485 = array_index_803228 == array_index_773020 ? add_803484 : sel_803481;
  assign add_803488 = sel_803485 + 8'h01;
  assign sel_803489 = array_index_803228 == array_index_773026 ? add_803488 : sel_803485;
  assign add_803492 = sel_803489 + 8'h01;
  assign sel_803493 = array_index_803228 == array_index_773032 ? add_803492 : sel_803489;
  assign add_803496 = sel_803493 + 8'h01;
  assign sel_803497 = array_index_803228 == array_index_773038 ? add_803496 : sel_803493;
  assign add_803500 = sel_803497 + 8'h01;
  assign sel_803501 = array_index_803228 == array_index_773044 ? add_803500 : sel_803497;
  assign add_803504 = sel_803501 + 8'h01;
  assign sel_803505 = array_index_803228 == array_index_773050 ? add_803504 : sel_803501;
  assign add_803508 = sel_803505 + 8'h01;
  assign sel_803509 = array_index_803228 == array_index_773056 ? add_803508 : sel_803505;
  assign add_803512 = sel_803509 + 8'h01;
  assign sel_803513 = array_index_803228 == array_index_773062 ? add_803512 : sel_803509;
  assign add_803516 = sel_803513 + 8'h01;
  assign sel_803517 = array_index_803228 == array_index_773068 ? add_803516 : sel_803513;
  assign add_803520 = sel_803517 + 8'h01;
  assign sel_803521 = array_index_803228 == array_index_773074 ? add_803520 : sel_803517;
  assign add_803524 = sel_803521 + 8'h01;
  assign sel_803525 = array_index_803228 == array_index_773080 ? add_803524 : sel_803521;
  assign add_803528 = sel_803525 + 8'h01;
  assign sel_803529 = array_index_803228 == array_index_773086 ? add_803528 : sel_803525;
  assign add_803532 = sel_803529 + 8'h01;
  assign sel_803533 = array_index_803228 == array_index_773092 ? add_803532 : sel_803529;
  assign add_803536 = sel_803533 + 8'h01;
  assign sel_803537 = array_index_803228 == array_index_773098 ? add_803536 : sel_803533;
  assign add_803540 = sel_803537 + 8'h01;
  assign sel_803541 = array_index_803228 == array_index_773104 ? add_803540 : sel_803537;
  assign add_803544 = sel_803541 + 8'h01;
  assign sel_803545 = array_index_803228 == array_index_773110 ? add_803544 : sel_803541;
  assign add_803548 = sel_803545 + 8'h01;
  assign sel_803549 = array_index_803228 == array_index_773116 ? add_803548 : sel_803545;
  assign add_803552 = sel_803549 + 8'h01;
  assign sel_803553 = array_index_803228 == array_index_773122 ? add_803552 : sel_803549;
  assign add_803556 = sel_803553 + 8'h01;
  assign sel_803557 = array_index_803228 == array_index_773128 ? add_803556 : sel_803553;
  assign add_803560 = sel_803557 + 8'h01;
  assign sel_803561 = array_index_803228 == array_index_773134 ? add_803560 : sel_803557;
  assign add_803564 = sel_803561 + 8'h01;
  assign sel_803565 = array_index_803228 == array_index_773140 ? add_803564 : sel_803561;
  assign add_803568 = sel_803565 + 8'h01;
  assign sel_803569 = array_index_803228 == array_index_773146 ? add_803568 : sel_803565;
  assign add_803572 = sel_803569 + 8'h01;
  assign sel_803573 = array_index_803228 == array_index_773152 ? add_803572 : sel_803569;
  assign add_803576 = sel_803573 + 8'h01;
  assign sel_803577 = array_index_803228 == array_index_773158 ? add_803576 : sel_803573;
  assign add_803580 = sel_803577 + 8'h01;
  assign sel_803581 = array_index_803228 == array_index_773164 ? add_803580 : sel_803577;
  assign add_803584 = sel_803581 + 8'h01;
  assign sel_803585 = array_index_803228 == array_index_773170 ? add_803584 : sel_803581;
  assign add_803589 = sel_803585 + 8'h01;
  assign array_index_803590 = set1_unflattened[7'h55];
  assign sel_803591 = array_index_803228 == array_index_773176 ? add_803589 : sel_803585;
  assign add_803594 = sel_803591 + 8'h01;
  assign sel_803595 = array_index_803590 == array_index_772632 ? add_803594 : sel_803591;
  assign add_803598 = sel_803595 + 8'h01;
  assign sel_803599 = array_index_803590 == array_index_772636 ? add_803598 : sel_803595;
  assign add_803602 = sel_803599 + 8'h01;
  assign sel_803603 = array_index_803590 == array_index_772644 ? add_803602 : sel_803599;
  assign add_803606 = sel_803603 + 8'h01;
  assign sel_803607 = array_index_803590 == array_index_772652 ? add_803606 : sel_803603;
  assign add_803610 = sel_803607 + 8'h01;
  assign sel_803611 = array_index_803590 == array_index_772660 ? add_803610 : sel_803607;
  assign add_803614 = sel_803611 + 8'h01;
  assign sel_803615 = array_index_803590 == array_index_772668 ? add_803614 : sel_803611;
  assign add_803618 = sel_803615 + 8'h01;
  assign sel_803619 = array_index_803590 == array_index_772676 ? add_803618 : sel_803615;
  assign add_803622 = sel_803619 + 8'h01;
  assign sel_803623 = array_index_803590 == array_index_772684 ? add_803622 : sel_803619;
  assign add_803626 = sel_803623 + 8'h01;
  assign sel_803627 = array_index_803590 == array_index_772690 ? add_803626 : sel_803623;
  assign add_803630 = sel_803627 + 8'h01;
  assign sel_803631 = array_index_803590 == array_index_772696 ? add_803630 : sel_803627;
  assign add_803634 = sel_803631 + 8'h01;
  assign sel_803635 = array_index_803590 == array_index_772702 ? add_803634 : sel_803631;
  assign add_803638 = sel_803635 + 8'h01;
  assign sel_803639 = array_index_803590 == array_index_772708 ? add_803638 : sel_803635;
  assign add_803642 = sel_803639 + 8'h01;
  assign sel_803643 = array_index_803590 == array_index_772714 ? add_803642 : sel_803639;
  assign add_803646 = sel_803643 + 8'h01;
  assign sel_803647 = array_index_803590 == array_index_772720 ? add_803646 : sel_803643;
  assign add_803650 = sel_803647 + 8'h01;
  assign sel_803651 = array_index_803590 == array_index_772726 ? add_803650 : sel_803647;
  assign add_803654 = sel_803651 + 8'h01;
  assign sel_803655 = array_index_803590 == array_index_772732 ? add_803654 : sel_803651;
  assign add_803658 = sel_803655 + 8'h01;
  assign sel_803659 = array_index_803590 == array_index_772738 ? add_803658 : sel_803655;
  assign add_803662 = sel_803659 + 8'h01;
  assign sel_803663 = array_index_803590 == array_index_772744 ? add_803662 : sel_803659;
  assign add_803666 = sel_803663 + 8'h01;
  assign sel_803667 = array_index_803590 == array_index_772750 ? add_803666 : sel_803663;
  assign add_803670 = sel_803667 + 8'h01;
  assign sel_803671 = array_index_803590 == array_index_772756 ? add_803670 : sel_803667;
  assign add_803674 = sel_803671 + 8'h01;
  assign sel_803675 = array_index_803590 == array_index_772762 ? add_803674 : sel_803671;
  assign add_803678 = sel_803675 + 8'h01;
  assign sel_803679 = array_index_803590 == array_index_772768 ? add_803678 : sel_803675;
  assign add_803682 = sel_803679 + 8'h01;
  assign sel_803683 = array_index_803590 == array_index_772774 ? add_803682 : sel_803679;
  assign add_803686 = sel_803683 + 8'h01;
  assign sel_803687 = array_index_803590 == array_index_772780 ? add_803686 : sel_803683;
  assign add_803690 = sel_803687 + 8'h01;
  assign sel_803691 = array_index_803590 == array_index_772786 ? add_803690 : sel_803687;
  assign add_803694 = sel_803691 + 8'h01;
  assign sel_803695 = array_index_803590 == array_index_772792 ? add_803694 : sel_803691;
  assign add_803698 = sel_803695 + 8'h01;
  assign sel_803699 = array_index_803590 == array_index_772798 ? add_803698 : sel_803695;
  assign add_803702 = sel_803699 + 8'h01;
  assign sel_803703 = array_index_803590 == array_index_772804 ? add_803702 : sel_803699;
  assign add_803706 = sel_803703 + 8'h01;
  assign sel_803707 = array_index_803590 == array_index_772810 ? add_803706 : sel_803703;
  assign add_803710 = sel_803707 + 8'h01;
  assign sel_803711 = array_index_803590 == array_index_772816 ? add_803710 : sel_803707;
  assign add_803714 = sel_803711 + 8'h01;
  assign sel_803715 = array_index_803590 == array_index_772822 ? add_803714 : sel_803711;
  assign add_803718 = sel_803715 + 8'h01;
  assign sel_803719 = array_index_803590 == array_index_772828 ? add_803718 : sel_803715;
  assign add_803722 = sel_803719 + 8'h01;
  assign sel_803723 = array_index_803590 == array_index_772834 ? add_803722 : sel_803719;
  assign add_803726 = sel_803723 + 8'h01;
  assign sel_803727 = array_index_803590 == array_index_772840 ? add_803726 : sel_803723;
  assign add_803730 = sel_803727 + 8'h01;
  assign sel_803731 = array_index_803590 == array_index_772846 ? add_803730 : sel_803727;
  assign add_803734 = sel_803731 + 8'h01;
  assign sel_803735 = array_index_803590 == array_index_772852 ? add_803734 : sel_803731;
  assign add_803738 = sel_803735 + 8'h01;
  assign sel_803739 = array_index_803590 == array_index_772858 ? add_803738 : sel_803735;
  assign add_803742 = sel_803739 + 8'h01;
  assign sel_803743 = array_index_803590 == array_index_772864 ? add_803742 : sel_803739;
  assign add_803746 = sel_803743 + 8'h01;
  assign sel_803747 = array_index_803590 == array_index_772870 ? add_803746 : sel_803743;
  assign add_803750 = sel_803747 + 8'h01;
  assign sel_803751 = array_index_803590 == array_index_772876 ? add_803750 : sel_803747;
  assign add_803754 = sel_803751 + 8'h01;
  assign sel_803755 = array_index_803590 == array_index_772882 ? add_803754 : sel_803751;
  assign add_803758 = sel_803755 + 8'h01;
  assign sel_803759 = array_index_803590 == array_index_772888 ? add_803758 : sel_803755;
  assign add_803762 = sel_803759 + 8'h01;
  assign sel_803763 = array_index_803590 == array_index_772894 ? add_803762 : sel_803759;
  assign add_803766 = sel_803763 + 8'h01;
  assign sel_803767 = array_index_803590 == array_index_772900 ? add_803766 : sel_803763;
  assign add_803770 = sel_803767 + 8'h01;
  assign sel_803771 = array_index_803590 == array_index_772906 ? add_803770 : sel_803767;
  assign add_803774 = sel_803771 + 8'h01;
  assign sel_803775 = array_index_803590 == array_index_772912 ? add_803774 : sel_803771;
  assign add_803778 = sel_803775 + 8'h01;
  assign sel_803779 = array_index_803590 == array_index_772918 ? add_803778 : sel_803775;
  assign add_803782 = sel_803779 + 8'h01;
  assign sel_803783 = array_index_803590 == array_index_772924 ? add_803782 : sel_803779;
  assign add_803786 = sel_803783 + 8'h01;
  assign sel_803787 = array_index_803590 == array_index_772930 ? add_803786 : sel_803783;
  assign add_803790 = sel_803787 + 8'h01;
  assign sel_803791 = array_index_803590 == array_index_772936 ? add_803790 : sel_803787;
  assign add_803794 = sel_803791 + 8'h01;
  assign sel_803795 = array_index_803590 == array_index_772942 ? add_803794 : sel_803791;
  assign add_803798 = sel_803795 + 8'h01;
  assign sel_803799 = array_index_803590 == array_index_772948 ? add_803798 : sel_803795;
  assign add_803802 = sel_803799 + 8'h01;
  assign sel_803803 = array_index_803590 == array_index_772954 ? add_803802 : sel_803799;
  assign add_803806 = sel_803803 + 8'h01;
  assign sel_803807 = array_index_803590 == array_index_772960 ? add_803806 : sel_803803;
  assign add_803810 = sel_803807 + 8'h01;
  assign sel_803811 = array_index_803590 == array_index_772966 ? add_803810 : sel_803807;
  assign add_803814 = sel_803811 + 8'h01;
  assign sel_803815 = array_index_803590 == array_index_772972 ? add_803814 : sel_803811;
  assign add_803818 = sel_803815 + 8'h01;
  assign sel_803819 = array_index_803590 == array_index_772978 ? add_803818 : sel_803815;
  assign add_803822 = sel_803819 + 8'h01;
  assign sel_803823 = array_index_803590 == array_index_772984 ? add_803822 : sel_803819;
  assign add_803826 = sel_803823 + 8'h01;
  assign sel_803827 = array_index_803590 == array_index_772990 ? add_803826 : sel_803823;
  assign add_803830 = sel_803827 + 8'h01;
  assign sel_803831 = array_index_803590 == array_index_772996 ? add_803830 : sel_803827;
  assign add_803834 = sel_803831 + 8'h01;
  assign sel_803835 = array_index_803590 == array_index_773002 ? add_803834 : sel_803831;
  assign add_803838 = sel_803835 + 8'h01;
  assign sel_803839 = array_index_803590 == array_index_773008 ? add_803838 : sel_803835;
  assign add_803842 = sel_803839 + 8'h01;
  assign sel_803843 = array_index_803590 == array_index_773014 ? add_803842 : sel_803839;
  assign add_803846 = sel_803843 + 8'h01;
  assign sel_803847 = array_index_803590 == array_index_773020 ? add_803846 : sel_803843;
  assign add_803850 = sel_803847 + 8'h01;
  assign sel_803851 = array_index_803590 == array_index_773026 ? add_803850 : sel_803847;
  assign add_803854 = sel_803851 + 8'h01;
  assign sel_803855 = array_index_803590 == array_index_773032 ? add_803854 : sel_803851;
  assign add_803858 = sel_803855 + 8'h01;
  assign sel_803859 = array_index_803590 == array_index_773038 ? add_803858 : sel_803855;
  assign add_803862 = sel_803859 + 8'h01;
  assign sel_803863 = array_index_803590 == array_index_773044 ? add_803862 : sel_803859;
  assign add_803866 = sel_803863 + 8'h01;
  assign sel_803867 = array_index_803590 == array_index_773050 ? add_803866 : sel_803863;
  assign add_803870 = sel_803867 + 8'h01;
  assign sel_803871 = array_index_803590 == array_index_773056 ? add_803870 : sel_803867;
  assign add_803874 = sel_803871 + 8'h01;
  assign sel_803875 = array_index_803590 == array_index_773062 ? add_803874 : sel_803871;
  assign add_803878 = sel_803875 + 8'h01;
  assign sel_803879 = array_index_803590 == array_index_773068 ? add_803878 : sel_803875;
  assign add_803882 = sel_803879 + 8'h01;
  assign sel_803883 = array_index_803590 == array_index_773074 ? add_803882 : sel_803879;
  assign add_803886 = sel_803883 + 8'h01;
  assign sel_803887 = array_index_803590 == array_index_773080 ? add_803886 : sel_803883;
  assign add_803890 = sel_803887 + 8'h01;
  assign sel_803891 = array_index_803590 == array_index_773086 ? add_803890 : sel_803887;
  assign add_803894 = sel_803891 + 8'h01;
  assign sel_803895 = array_index_803590 == array_index_773092 ? add_803894 : sel_803891;
  assign add_803898 = sel_803895 + 8'h01;
  assign sel_803899 = array_index_803590 == array_index_773098 ? add_803898 : sel_803895;
  assign add_803902 = sel_803899 + 8'h01;
  assign sel_803903 = array_index_803590 == array_index_773104 ? add_803902 : sel_803899;
  assign add_803906 = sel_803903 + 8'h01;
  assign sel_803907 = array_index_803590 == array_index_773110 ? add_803906 : sel_803903;
  assign add_803910 = sel_803907 + 8'h01;
  assign sel_803911 = array_index_803590 == array_index_773116 ? add_803910 : sel_803907;
  assign add_803914 = sel_803911 + 8'h01;
  assign sel_803915 = array_index_803590 == array_index_773122 ? add_803914 : sel_803911;
  assign add_803918 = sel_803915 + 8'h01;
  assign sel_803919 = array_index_803590 == array_index_773128 ? add_803918 : sel_803915;
  assign add_803922 = sel_803919 + 8'h01;
  assign sel_803923 = array_index_803590 == array_index_773134 ? add_803922 : sel_803919;
  assign add_803926 = sel_803923 + 8'h01;
  assign sel_803927 = array_index_803590 == array_index_773140 ? add_803926 : sel_803923;
  assign add_803930 = sel_803927 + 8'h01;
  assign sel_803931 = array_index_803590 == array_index_773146 ? add_803930 : sel_803927;
  assign add_803934 = sel_803931 + 8'h01;
  assign sel_803935 = array_index_803590 == array_index_773152 ? add_803934 : sel_803931;
  assign add_803938 = sel_803935 + 8'h01;
  assign sel_803939 = array_index_803590 == array_index_773158 ? add_803938 : sel_803935;
  assign add_803942 = sel_803939 + 8'h01;
  assign sel_803943 = array_index_803590 == array_index_773164 ? add_803942 : sel_803939;
  assign add_803946 = sel_803943 + 8'h01;
  assign sel_803947 = array_index_803590 == array_index_773170 ? add_803946 : sel_803943;
  assign add_803951 = sel_803947 + 8'h01;
  assign array_index_803952 = set1_unflattened[7'h56];
  assign sel_803953 = array_index_803590 == array_index_773176 ? add_803951 : sel_803947;
  assign add_803956 = sel_803953 + 8'h01;
  assign sel_803957 = array_index_803952 == array_index_772632 ? add_803956 : sel_803953;
  assign add_803960 = sel_803957 + 8'h01;
  assign sel_803961 = array_index_803952 == array_index_772636 ? add_803960 : sel_803957;
  assign add_803964 = sel_803961 + 8'h01;
  assign sel_803965 = array_index_803952 == array_index_772644 ? add_803964 : sel_803961;
  assign add_803968 = sel_803965 + 8'h01;
  assign sel_803969 = array_index_803952 == array_index_772652 ? add_803968 : sel_803965;
  assign add_803972 = sel_803969 + 8'h01;
  assign sel_803973 = array_index_803952 == array_index_772660 ? add_803972 : sel_803969;
  assign add_803976 = sel_803973 + 8'h01;
  assign sel_803977 = array_index_803952 == array_index_772668 ? add_803976 : sel_803973;
  assign add_803980 = sel_803977 + 8'h01;
  assign sel_803981 = array_index_803952 == array_index_772676 ? add_803980 : sel_803977;
  assign add_803984 = sel_803981 + 8'h01;
  assign sel_803985 = array_index_803952 == array_index_772684 ? add_803984 : sel_803981;
  assign add_803988 = sel_803985 + 8'h01;
  assign sel_803989 = array_index_803952 == array_index_772690 ? add_803988 : sel_803985;
  assign add_803992 = sel_803989 + 8'h01;
  assign sel_803993 = array_index_803952 == array_index_772696 ? add_803992 : sel_803989;
  assign add_803996 = sel_803993 + 8'h01;
  assign sel_803997 = array_index_803952 == array_index_772702 ? add_803996 : sel_803993;
  assign add_804000 = sel_803997 + 8'h01;
  assign sel_804001 = array_index_803952 == array_index_772708 ? add_804000 : sel_803997;
  assign add_804004 = sel_804001 + 8'h01;
  assign sel_804005 = array_index_803952 == array_index_772714 ? add_804004 : sel_804001;
  assign add_804008 = sel_804005 + 8'h01;
  assign sel_804009 = array_index_803952 == array_index_772720 ? add_804008 : sel_804005;
  assign add_804012 = sel_804009 + 8'h01;
  assign sel_804013 = array_index_803952 == array_index_772726 ? add_804012 : sel_804009;
  assign add_804016 = sel_804013 + 8'h01;
  assign sel_804017 = array_index_803952 == array_index_772732 ? add_804016 : sel_804013;
  assign add_804020 = sel_804017 + 8'h01;
  assign sel_804021 = array_index_803952 == array_index_772738 ? add_804020 : sel_804017;
  assign add_804024 = sel_804021 + 8'h01;
  assign sel_804025 = array_index_803952 == array_index_772744 ? add_804024 : sel_804021;
  assign add_804028 = sel_804025 + 8'h01;
  assign sel_804029 = array_index_803952 == array_index_772750 ? add_804028 : sel_804025;
  assign add_804032 = sel_804029 + 8'h01;
  assign sel_804033 = array_index_803952 == array_index_772756 ? add_804032 : sel_804029;
  assign add_804036 = sel_804033 + 8'h01;
  assign sel_804037 = array_index_803952 == array_index_772762 ? add_804036 : sel_804033;
  assign add_804040 = sel_804037 + 8'h01;
  assign sel_804041 = array_index_803952 == array_index_772768 ? add_804040 : sel_804037;
  assign add_804044 = sel_804041 + 8'h01;
  assign sel_804045 = array_index_803952 == array_index_772774 ? add_804044 : sel_804041;
  assign add_804048 = sel_804045 + 8'h01;
  assign sel_804049 = array_index_803952 == array_index_772780 ? add_804048 : sel_804045;
  assign add_804052 = sel_804049 + 8'h01;
  assign sel_804053 = array_index_803952 == array_index_772786 ? add_804052 : sel_804049;
  assign add_804056 = sel_804053 + 8'h01;
  assign sel_804057 = array_index_803952 == array_index_772792 ? add_804056 : sel_804053;
  assign add_804060 = sel_804057 + 8'h01;
  assign sel_804061 = array_index_803952 == array_index_772798 ? add_804060 : sel_804057;
  assign add_804064 = sel_804061 + 8'h01;
  assign sel_804065 = array_index_803952 == array_index_772804 ? add_804064 : sel_804061;
  assign add_804068 = sel_804065 + 8'h01;
  assign sel_804069 = array_index_803952 == array_index_772810 ? add_804068 : sel_804065;
  assign add_804072 = sel_804069 + 8'h01;
  assign sel_804073 = array_index_803952 == array_index_772816 ? add_804072 : sel_804069;
  assign add_804076 = sel_804073 + 8'h01;
  assign sel_804077 = array_index_803952 == array_index_772822 ? add_804076 : sel_804073;
  assign add_804080 = sel_804077 + 8'h01;
  assign sel_804081 = array_index_803952 == array_index_772828 ? add_804080 : sel_804077;
  assign add_804084 = sel_804081 + 8'h01;
  assign sel_804085 = array_index_803952 == array_index_772834 ? add_804084 : sel_804081;
  assign add_804088 = sel_804085 + 8'h01;
  assign sel_804089 = array_index_803952 == array_index_772840 ? add_804088 : sel_804085;
  assign add_804092 = sel_804089 + 8'h01;
  assign sel_804093 = array_index_803952 == array_index_772846 ? add_804092 : sel_804089;
  assign add_804096 = sel_804093 + 8'h01;
  assign sel_804097 = array_index_803952 == array_index_772852 ? add_804096 : sel_804093;
  assign add_804100 = sel_804097 + 8'h01;
  assign sel_804101 = array_index_803952 == array_index_772858 ? add_804100 : sel_804097;
  assign add_804104 = sel_804101 + 8'h01;
  assign sel_804105 = array_index_803952 == array_index_772864 ? add_804104 : sel_804101;
  assign add_804108 = sel_804105 + 8'h01;
  assign sel_804109 = array_index_803952 == array_index_772870 ? add_804108 : sel_804105;
  assign add_804112 = sel_804109 + 8'h01;
  assign sel_804113 = array_index_803952 == array_index_772876 ? add_804112 : sel_804109;
  assign add_804116 = sel_804113 + 8'h01;
  assign sel_804117 = array_index_803952 == array_index_772882 ? add_804116 : sel_804113;
  assign add_804120 = sel_804117 + 8'h01;
  assign sel_804121 = array_index_803952 == array_index_772888 ? add_804120 : sel_804117;
  assign add_804124 = sel_804121 + 8'h01;
  assign sel_804125 = array_index_803952 == array_index_772894 ? add_804124 : sel_804121;
  assign add_804128 = sel_804125 + 8'h01;
  assign sel_804129 = array_index_803952 == array_index_772900 ? add_804128 : sel_804125;
  assign add_804132 = sel_804129 + 8'h01;
  assign sel_804133 = array_index_803952 == array_index_772906 ? add_804132 : sel_804129;
  assign add_804136 = sel_804133 + 8'h01;
  assign sel_804137 = array_index_803952 == array_index_772912 ? add_804136 : sel_804133;
  assign add_804140 = sel_804137 + 8'h01;
  assign sel_804141 = array_index_803952 == array_index_772918 ? add_804140 : sel_804137;
  assign add_804144 = sel_804141 + 8'h01;
  assign sel_804145 = array_index_803952 == array_index_772924 ? add_804144 : sel_804141;
  assign add_804148 = sel_804145 + 8'h01;
  assign sel_804149 = array_index_803952 == array_index_772930 ? add_804148 : sel_804145;
  assign add_804152 = sel_804149 + 8'h01;
  assign sel_804153 = array_index_803952 == array_index_772936 ? add_804152 : sel_804149;
  assign add_804156 = sel_804153 + 8'h01;
  assign sel_804157 = array_index_803952 == array_index_772942 ? add_804156 : sel_804153;
  assign add_804160 = sel_804157 + 8'h01;
  assign sel_804161 = array_index_803952 == array_index_772948 ? add_804160 : sel_804157;
  assign add_804164 = sel_804161 + 8'h01;
  assign sel_804165 = array_index_803952 == array_index_772954 ? add_804164 : sel_804161;
  assign add_804168 = sel_804165 + 8'h01;
  assign sel_804169 = array_index_803952 == array_index_772960 ? add_804168 : sel_804165;
  assign add_804172 = sel_804169 + 8'h01;
  assign sel_804173 = array_index_803952 == array_index_772966 ? add_804172 : sel_804169;
  assign add_804176 = sel_804173 + 8'h01;
  assign sel_804177 = array_index_803952 == array_index_772972 ? add_804176 : sel_804173;
  assign add_804180 = sel_804177 + 8'h01;
  assign sel_804181 = array_index_803952 == array_index_772978 ? add_804180 : sel_804177;
  assign add_804184 = sel_804181 + 8'h01;
  assign sel_804185 = array_index_803952 == array_index_772984 ? add_804184 : sel_804181;
  assign add_804188 = sel_804185 + 8'h01;
  assign sel_804189 = array_index_803952 == array_index_772990 ? add_804188 : sel_804185;
  assign add_804192 = sel_804189 + 8'h01;
  assign sel_804193 = array_index_803952 == array_index_772996 ? add_804192 : sel_804189;
  assign add_804196 = sel_804193 + 8'h01;
  assign sel_804197 = array_index_803952 == array_index_773002 ? add_804196 : sel_804193;
  assign add_804200 = sel_804197 + 8'h01;
  assign sel_804201 = array_index_803952 == array_index_773008 ? add_804200 : sel_804197;
  assign add_804204 = sel_804201 + 8'h01;
  assign sel_804205 = array_index_803952 == array_index_773014 ? add_804204 : sel_804201;
  assign add_804208 = sel_804205 + 8'h01;
  assign sel_804209 = array_index_803952 == array_index_773020 ? add_804208 : sel_804205;
  assign add_804212 = sel_804209 + 8'h01;
  assign sel_804213 = array_index_803952 == array_index_773026 ? add_804212 : sel_804209;
  assign add_804216 = sel_804213 + 8'h01;
  assign sel_804217 = array_index_803952 == array_index_773032 ? add_804216 : sel_804213;
  assign add_804220 = sel_804217 + 8'h01;
  assign sel_804221 = array_index_803952 == array_index_773038 ? add_804220 : sel_804217;
  assign add_804224 = sel_804221 + 8'h01;
  assign sel_804225 = array_index_803952 == array_index_773044 ? add_804224 : sel_804221;
  assign add_804228 = sel_804225 + 8'h01;
  assign sel_804229 = array_index_803952 == array_index_773050 ? add_804228 : sel_804225;
  assign add_804232 = sel_804229 + 8'h01;
  assign sel_804233 = array_index_803952 == array_index_773056 ? add_804232 : sel_804229;
  assign add_804236 = sel_804233 + 8'h01;
  assign sel_804237 = array_index_803952 == array_index_773062 ? add_804236 : sel_804233;
  assign add_804240 = sel_804237 + 8'h01;
  assign sel_804241 = array_index_803952 == array_index_773068 ? add_804240 : sel_804237;
  assign add_804244 = sel_804241 + 8'h01;
  assign sel_804245 = array_index_803952 == array_index_773074 ? add_804244 : sel_804241;
  assign add_804248 = sel_804245 + 8'h01;
  assign sel_804249 = array_index_803952 == array_index_773080 ? add_804248 : sel_804245;
  assign add_804252 = sel_804249 + 8'h01;
  assign sel_804253 = array_index_803952 == array_index_773086 ? add_804252 : sel_804249;
  assign add_804256 = sel_804253 + 8'h01;
  assign sel_804257 = array_index_803952 == array_index_773092 ? add_804256 : sel_804253;
  assign add_804260 = sel_804257 + 8'h01;
  assign sel_804261 = array_index_803952 == array_index_773098 ? add_804260 : sel_804257;
  assign add_804264 = sel_804261 + 8'h01;
  assign sel_804265 = array_index_803952 == array_index_773104 ? add_804264 : sel_804261;
  assign add_804268 = sel_804265 + 8'h01;
  assign sel_804269 = array_index_803952 == array_index_773110 ? add_804268 : sel_804265;
  assign add_804272 = sel_804269 + 8'h01;
  assign sel_804273 = array_index_803952 == array_index_773116 ? add_804272 : sel_804269;
  assign add_804276 = sel_804273 + 8'h01;
  assign sel_804277 = array_index_803952 == array_index_773122 ? add_804276 : sel_804273;
  assign add_804280 = sel_804277 + 8'h01;
  assign sel_804281 = array_index_803952 == array_index_773128 ? add_804280 : sel_804277;
  assign add_804284 = sel_804281 + 8'h01;
  assign sel_804285 = array_index_803952 == array_index_773134 ? add_804284 : sel_804281;
  assign add_804288 = sel_804285 + 8'h01;
  assign sel_804289 = array_index_803952 == array_index_773140 ? add_804288 : sel_804285;
  assign add_804292 = sel_804289 + 8'h01;
  assign sel_804293 = array_index_803952 == array_index_773146 ? add_804292 : sel_804289;
  assign add_804296 = sel_804293 + 8'h01;
  assign sel_804297 = array_index_803952 == array_index_773152 ? add_804296 : sel_804293;
  assign add_804300 = sel_804297 + 8'h01;
  assign sel_804301 = array_index_803952 == array_index_773158 ? add_804300 : sel_804297;
  assign add_804304 = sel_804301 + 8'h01;
  assign sel_804305 = array_index_803952 == array_index_773164 ? add_804304 : sel_804301;
  assign add_804308 = sel_804305 + 8'h01;
  assign sel_804309 = array_index_803952 == array_index_773170 ? add_804308 : sel_804305;
  assign add_804313 = sel_804309 + 8'h01;
  assign array_index_804314 = set1_unflattened[7'h57];
  assign sel_804315 = array_index_803952 == array_index_773176 ? add_804313 : sel_804309;
  assign add_804318 = sel_804315 + 8'h01;
  assign sel_804319 = array_index_804314 == array_index_772632 ? add_804318 : sel_804315;
  assign add_804322 = sel_804319 + 8'h01;
  assign sel_804323 = array_index_804314 == array_index_772636 ? add_804322 : sel_804319;
  assign add_804326 = sel_804323 + 8'h01;
  assign sel_804327 = array_index_804314 == array_index_772644 ? add_804326 : sel_804323;
  assign add_804330 = sel_804327 + 8'h01;
  assign sel_804331 = array_index_804314 == array_index_772652 ? add_804330 : sel_804327;
  assign add_804334 = sel_804331 + 8'h01;
  assign sel_804335 = array_index_804314 == array_index_772660 ? add_804334 : sel_804331;
  assign add_804338 = sel_804335 + 8'h01;
  assign sel_804339 = array_index_804314 == array_index_772668 ? add_804338 : sel_804335;
  assign add_804342 = sel_804339 + 8'h01;
  assign sel_804343 = array_index_804314 == array_index_772676 ? add_804342 : sel_804339;
  assign add_804346 = sel_804343 + 8'h01;
  assign sel_804347 = array_index_804314 == array_index_772684 ? add_804346 : sel_804343;
  assign add_804350 = sel_804347 + 8'h01;
  assign sel_804351 = array_index_804314 == array_index_772690 ? add_804350 : sel_804347;
  assign add_804354 = sel_804351 + 8'h01;
  assign sel_804355 = array_index_804314 == array_index_772696 ? add_804354 : sel_804351;
  assign add_804358 = sel_804355 + 8'h01;
  assign sel_804359 = array_index_804314 == array_index_772702 ? add_804358 : sel_804355;
  assign add_804362 = sel_804359 + 8'h01;
  assign sel_804363 = array_index_804314 == array_index_772708 ? add_804362 : sel_804359;
  assign add_804366 = sel_804363 + 8'h01;
  assign sel_804367 = array_index_804314 == array_index_772714 ? add_804366 : sel_804363;
  assign add_804370 = sel_804367 + 8'h01;
  assign sel_804371 = array_index_804314 == array_index_772720 ? add_804370 : sel_804367;
  assign add_804374 = sel_804371 + 8'h01;
  assign sel_804375 = array_index_804314 == array_index_772726 ? add_804374 : sel_804371;
  assign add_804378 = sel_804375 + 8'h01;
  assign sel_804379 = array_index_804314 == array_index_772732 ? add_804378 : sel_804375;
  assign add_804382 = sel_804379 + 8'h01;
  assign sel_804383 = array_index_804314 == array_index_772738 ? add_804382 : sel_804379;
  assign add_804386 = sel_804383 + 8'h01;
  assign sel_804387 = array_index_804314 == array_index_772744 ? add_804386 : sel_804383;
  assign add_804390 = sel_804387 + 8'h01;
  assign sel_804391 = array_index_804314 == array_index_772750 ? add_804390 : sel_804387;
  assign add_804394 = sel_804391 + 8'h01;
  assign sel_804395 = array_index_804314 == array_index_772756 ? add_804394 : sel_804391;
  assign add_804398 = sel_804395 + 8'h01;
  assign sel_804399 = array_index_804314 == array_index_772762 ? add_804398 : sel_804395;
  assign add_804402 = sel_804399 + 8'h01;
  assign sel_804403 = array_index_804314 == array_index_772768 ? add_804402 : sel_804399;
  assign add_804406 = sel_804403 + 8'h01;
  assign sel_804407 = array_index_804314 == array_index_772774 ? add_804406 : sel_804403;
  assign add_804410 = sel_804407 + 8'h01;
  assign sel_804411 = array_index_804314 == array_index_772780 ? add_804410 : sel_804407;
  assign add_804414 = sel_804411 + 8'h01;
  assign sel_804415 = array_index_804314 == array_index_772786 ? add_804414 : sel_804411;
  assign add_804418 = sel_804415 + 8'h01;
  assign sel_804419 = array_index_804314 == array_index_772792 ? add_804418 : sel_804415;
  assign add_804422 = sel_804419 + 8'h01;
  assign sel_804423 = array_index_804314 == array_index_772798 ? add_804422 : sel_804419;
  assign add_804426 = sel_804423 + 8'h01;
  assign sel_804427 = array_index_804314 == array_index_772804 ? add_804426 : sel_804423;
  assign add_804430 = sel_804427 + 8'h01;
  assign sel_804431 = array_index_804314 == array_index_772810 ? add_804430 : sel_804427;
  assign add_804434 = sel_804431 + 8'h01;
  assign sel_804435 = array_index_804314 == array_index_772816 ? add_804434 : sel_804431;
  assign add_804438 = sel_804435 + 8'h01;
  assign sel_804439 = array_index_804314 == array_index_772822 ? add_804438 : sel_804435;
  assign add_804442 = sel_804439 + 8'h01;
  assign sel_804443 = array_index_804314 == array_index_772828 ? add_804442 : sel_804439;
  assign add_804446 = sel_804443 + 8'h01;
  assign sel_804447 = array_index_804314 == array_index_772834 ? add_804446 : sel_804443;
  assign add_804450 = sel_804447 + 8'h01;
  assign sel_804451 = array_index_804314 == array_index_772840 ? add_804450 : sel_804447;
  assign add_804454 = sel_804451 + 8'h01;
  assign sel_804455 = array_index_804314 == array_index_772846 ? add_804454 : sel_804451;
  assign add_804458 = sel_804455 + 8'h01;
  assign sel_804459 = array_index_804314 == array_index_772852 ? add_804458 : sel_804455;
  assign add_804462 = sel_804459 + 8'h01;
  assign sel_804463 = array_index_804314 == array_index_772858 ? add_804462 : sel_804459;
  assign add_804466 = sel_804463 + 8'h01;
  assign sel_804467 = array_index_804314 == array_index_772864 ? add_804466 : sel_804463;
  assign add_804470 = sel_804467 + 8'h01;
  assign sel_804471 = array_index_804314 == array_index_772870 ? add_804470 : sel_804467;
  assign add_804474 = sel_804471 + 8'h01;
  assign sel_804475 = array_index_804314 == array_index_772876 ? add_804474 : sel_804471;
  assign add_804478 = sel_804475 + 8'h01;
  assign sel_804479 = array_index_804314 == array_index_772882 ? add_804478 : sel_804475;
  assign add_804482 = sel_804479 + 8'h01;
  assign sel_804483 = array_index_804314 == array_index_772888 ? add_804482 : sel_804479;
  assign add_804486 = sel_804483 + 8'h01;
  assign sel_804487 = array_index_804314 == array_index_772894 ? add_804486 : sel_804483;
  assign add_804490 = sel_804487 + 8'h01;
  assign sel_804491 = array_index_804314 == array_index_772900 ? add_804490 : sel_804487;
  assign add_804494 = sel_804491 + 8'h01;
  assign sel_804495 = array_index_804314 == array_index_772906 ? add_804494 : sel_804491;
  assign add_804498 = sel_804495 + 8'h01;
  assign sel_804499 = array_index_804314 == array_index_772912 ? add_804498 : sel_804495;
  assign add_804502 = sel_804499 + 8'h01;
  assign sel_804503 = array_index_804314 == array_index_772918 ? add_804502 : sel_804499;
  assign add_804506 = sel_804503 + 8'h01;
  assign sel_804507 = array_index_804314 == array_index_772924 ? add_804506 : sel_804503;
  assign add_804510 = sel_804507 + 8'h01;
  assign sel_804511 = array_index_804314 == array_index_772930 ? add_804510 : sel_804507;
  assign add_804514 = sel_804511 + 8'h01;
  assign sel_804515 = array_index_804314 == array_index_772936 ? add_804514 : sel_804511;
  assign add_804518 = sel_804515 + 8'h01;
  assign sel_804519 = array_index_804314 == array_index_772942 ? add_804518 : sel_804515;
  assign add_804522 = sel_804519 + 8'h01;
  assign sel_804523 = array_index_804314 == array_index_772948 ? add_804522 : sel_804519;
  assign add_804526 = sel_804523 + 8'h01;
  assign sel_804527 = array_index_804314 == array_index_772954 ? add_804526 : sel_804523;
  assign add_804530 = sel_804527 + 8'h01;
  assign sel_804531 = array_index_804314 == array_index_772960 ? add_804530 : sel_804527;
  assign add_804534 = sel_804531 + 8'h01;
  assign sel_804535 = array_index_804314 == array_index_772966 ? add_804534 : sel_804531;
  assign add_804538 = sel_804535 + 8'h01;
  assign sel_804539 = array_index_804314 == array_index_772972 ? add_804538 : sel_804535;
  assign add_804542 = sel_804539 + 8'h01;
  assign sel_804543 = array_index_804314 == array_index_772978 ? add_804542 : sel_804539;
  assign add_804546 = sel_804543 + 8'h01;
  assign sel_804547 = array_index_804314 == array_index_772984 ? add_804546 : sel_804543;
  assign add_804550 = sel_804547 + 8'h01;
  assign sel_804551 = array_index_804314 == array_index_772990 ? add_804550 : sel_804547;
  assign add_804554 = sel_804551 + 8'h01;
  assign sel_804555 = array_index_804314 == array_index_772996 ? add_804554 : sel_804551;
  assign add_804558 = sel_804555 + 8'h01;
  assign sel_804559 = array_index_804314 == array_index_773002 ? add_804558 : sel_804555;
  assign add_804562 = sel_804559 + 8'h01;
  assign sel_804563 = array_index_804314 == array_index_773008 ? add_804562 : sel_804559;
  assign add_804566 = sel_804563 + 8'h01;
  assign sel_804567 = array_index_804314 == array_index_773014 ? add_804566 : sel_804563;
  assign add_804570 = sel_804567 + 8'h01;
  assign sel_804571 = array_index_804314 == array_index_773020 ? add_804570 : sel_804567;
  assign add_804574 = sel_804571 + 8'h01;
  assign sel_804575 = array_index_804314 == array_index_773026 ? add_804574 : sel_804571;
  assign add_804578 = sel_804575 + 8'h01;
  assign sel_804579 = array_index_804314 == array_index_773032 ? add_804578 : sel_804575;
  assign add_804582 = sel_804579 + 8'h01;
  assign sel_804583 = array_index_804314 == array_index_773038 ? add_804582 : sel_804579;
  assign add_804586 = sel_804583 + 8'h01;
  assign sel_804587 = array_index_804314 == array_index_773044 ? add_804586 : sel_804583;
  assign add_804590 = sel_804587 + 8'h01;
  assign sel_804591 = array_index_804314 == array_index_773050 ? add_804590 : sel_804587;
  assign add_804594 = sel_804591 + 8'h01;
  assign sel_804595 = array_index_804314 == array_index_773056 ? add_804594 : sel_804591;
  assign add_804598 = sel_804595 + 8'h01;
  assign sel_804599 = array_index_804314 == array_index_773062 ? add_804598 : sel_804595;
  assign add_804602 = sel_804599 + 8'h01;
  assign sel_804603 = array_index_804314 == array_index_773068 ? add_804602 : sel_804599;
  assign add_804606 = sel_804603 + 8'h01;
  assign sel_804607 = array_index_804314 == array_index_773074 ? add_804606 : sel_804603;
  assign add_804610 = sel_804607 + 8'h01;
  assign sel_804611 = array_index_804314 == array_index_773080 ? add_804610 : sel_804607;
  assign add_804614 = sel_804611 + 8'h01;
  assign sel_804615 = array_index_804314 == array_index_773086 ? add_804614 : sel_804611;
  assign add_804618 = sel_804615 + 8'h01;
  assign sel_804619 = array_index_804314 == array_index_773092 ? add_804618 : sel_804615;
  assign add_804622 = sel_804619 + 8'h01;
  assign sel_804623 = array_index_804314 == array_index_773098 ? add_804622 : sel_804619;
  assign add_804626 = sel_804623 + 8'h01;
  assign sel_804627 = array_index_804314 == array_index_773104 ? add_804626 : sel_804623;
  assign add_804630 = sel_804627 + 8'h01;
  assign sel_804631 = array_index_804314 == array_index_773110 ? add_804630 : sel_804627;
  assign add_804634 = sel_804631 + 8'h01;
  assign sel_804635 = array_index_804314 == array_index_773116 ? add_804634 : sel_804631;
  assign add_804638 = sel_804635 + 8'h01;
  assign sel_804639 = array_index_804314 == array_index_773122 ? add_804638 : sel_804635;
  assign add_804642 = sel_804639 + 8'h01;
  assign sel_804643 = array_index_804314 == array_index_773128 ? add_804642 : sel_804639;
  assign add_804646 = sel_804643 + 8'h01;
  assign sel_804647 = array_index_804314 == array_index_773134 ? add_804646 : sel_804643;
  assign add_804650 = sel_804647 + 8'h01;
  assign sel_804651 = array_index_804314 == array_index_773140 ? add_804650 : sel_804647;
  assign add_804654 = sel_804651 + 8'h01;
  assign sel_804655 = array_index_804314 == array_index_773146 ? add_804654 : sel_804651;
  assign add_804658 = sel_804655 + 8'h01;
  assign sel_804659 = array_index_804314 == array_index_773152 ? add_804658 : sel_804655;
  assign add_804662 = sel_804659 + 8'h01;
  assign sel_804663 = array_index_804314 == array_index_773158 ? add_804662 : sel_804659;
  assign add_804666 = sel_804663 + 8'h01;
  assign sel_804667 = array_index_804314 == array_index_773164 ? add_804666 : sel_804663;
  assign add_804670 = sel_804667 + 8'h01;
  assign sel_804671 = array_index_804314 == array_index_773170 ? add_804670 : sel_804667;
  assign add_804675 = sel_804671 + 8'h01;
  assign array_index_804676 = set1_unflattened[7'h58];
  assign sel_804677 = array_index_804314 == array_index_773176 ? add_804675 : sel_804671;
  assign add_804680 = sel_804677 + 8'h01;
  assign sel_804681 = array_index_804676 == array_index_772632 ? add_804680 : sel_804677;
  assign add_804684 = sel_804681 + 8'h01;
  assign sel_804685 = array_index_804676 == array_index_772636 ? add_804684 : sel_804681;
  assign add_804688 = sel_804685 + 8'h01;
  assign sel_804689 = array_index_804676 == array_index_772644 ? add_804688 : sel_804685;
  assign add_804692 = sel_804689 + 8'h01;
  assign sel_804693 = array_index_804676 == array_index_772652 ? add_804692 : sel_804689;
  assign add_804696 = sel_804693 + 8'h01;
  assign sel_804697 = array_index_804676 == array_index_772660 ? add_804696 : sel_804693;
  assign add_804700 = sel_804697 + 8'h01;
  assign sel_804701 = array_index_804676 == array_index_772668 ? add_804700 : sel_804697;
  assign add_804704 = sel_804701 + 8'h01;
  assign sel_804705 = array_index_804676 == array_index_772676 ? add_804704 : sel_804701;
  assign add_804708 = sel_804705 + 8'h01;
  assign sel_804709 = array_index_804676 == array_index_772684 ? add_804708 : sel_804705;
  assign add_804712 = sel_804709 + 8'h01;
  assign sel_804713 = array_index_804676 == array_index_772690 ? add_804712 : sel_804709;
  assign add_804716 = sel_804713 + 8'h01;
  assign sel_804717 = array_index_804676 == array_index_772696 ? add_804716 : sel_804713;
  assign add_804720 = sel_804717 + 8'h01;
  assign sel_804721 = array_index_804676 == array_index_772702 ? add_804720 : sel_804717;
  assign add_804724 = sel_804721 + 8'h01;
  assign sel_804725 = array_index_804676 == array_index_772708 ? add_804724 : sel_804721;
  assign add_804728 = sel_804725 + 8'h01;
  assign sel_804729 = array_index_804676 == array_index_772714 ? add_804728 : sel_804725;
  assign add_804732 = sel_804729 + 8'h01;
  assign sel_804733 = array_index_804676 == array_index_772720 ? add_804732 : sel_804729;
  assign add_804736 = sel_804733 + 8'h01;
  assign sel_804737 = array_index_804676 == array_index_772726 ? add_804736 : sel_804733;
  assign add_804740 = sel_804737 + 8'h01;
  assign sel_804741 = array_index_804676 == array_index_772732 ? add_804740 : sel_804737;
  assign add_804744 = sel_804741 + 8'h01;
  assign sel_804745 = array_index_804676 == array_index_772738 ? add_804744 : sel_804741;
  assign add_804748 = sel_804745 + 8'h01;
  assign sel_804749 = array_index_804676 == array_index_772744 ? add_804748 : sel_804745;
  assign add_804752 = sel_804749 + 8'h01;
  assign sel_804753 = array_index_804676 == array_index_772750 ? add_804752 : sel_804749;
  assign add_804756 = sel_804753 + 8'h01;
  assign sel_804757 = array_index_804676 == array_index_772756 ? add_804756 : sel_804753;
  assign add_804760 = sel_804757 + 8'h01;
  assign sel_804761 = array_index_804676 == array_index_772762 ? add_804760 : sel_804757;
  assign add_804764 = sel_804761 + 8'h01;
  assign sel_804765 = array_index_804676 == array_index_772768 ? add_804764 : sel_804761;
  assign add_804768 = sel_804765 + 8'h01;
  assign sel_804769 = array_index_804676 == array_index_772774 ? add_804768 : sel_804765;
  assign add_804772 = sel_804769 + 8'h01;
  assign sel_804773 = array_index_804676 == array_index_772780 ? add_804772 : sel_804769;
  assign add_804776 = sel_804773 + 8'h01;
  assign sel_804777 = array_index_804676 == array_index_772786 ? add_804776 : sel_804773;
  assign add_804780 = sel_804777 + 8'h01;
  assign sel_804781 = array_index_804676 == array_index_772792 ? add_804780 : sel_804777;
  assign add_804784 = sel_804781 + 8'h01;
  assign sel_804785 = array_index_804676 == array_index_772798 ? add_804784 : sel_804781;
  assign add_804788 = sel_804785 + 8'h01;
  assign sel_804789 = array_index_804676 == array_index_772804 ? add_804788 : sel_804785;
  assign add_804792 = sel_804789 + 8'h01;
  assign sel_804793 = array_index_804676 == array_index_772810 ? add_804792 : sel_804789;
  assign add_804796 = sel_804793 + 8'h01;
  assign sel_804797 = array_index_804676 == array_index_772816 ? add_804796 : sel_804793;
  assign add_804800 = sel_804797 + 8'h01;
  assign sel_804801 = array_index_804676 == array_index_772822 ? add_804800 : sel_804797;
  assign add_804804 = sel_804801 + 8'h01;
  assign sel_804805 = array_index_804676 == array_index_772828 ? add_804804 : sel_804801;
  assign add_804808 = sel_804805 + 8'h01;
  assign sel_804809 = array_index_804676 == array_index_772834 ? add_804808 : sel_804805;
  assign add_804812 = sel_804809 + 8'h01;
  assign sel_804813 = array_index_804676 == array_index_772840 ? add_804812 : sel_804809;
  assign add_804816 = sel_804813 + 8'h01;
  assign sel_804817 = array_index_804676 == array_index_772846 ? add_804816 : sel_804813;
  assign add_804820 = sel_804817 + 8'h01;
  assign sel_804821 = array_index_804676 == array_index_772852 ? add_804820 : sel_804817;
  assign add_804824 = sel_804821 + 8'h01;
  assign sel_804825 = array_index_804676 == array_index_772858 ? add_804824 : sel_804821;
  assign add_804828 = sel_804825 + 8'h01;
  assign sel_804829 = array_index_804676 == array_index_772864 ? add_804828 : sel_804825;
  assign add_804832 = sel_804829 + 8'h01;
  assign sel_804833 = array_index_804676 == array_index_772870 ? add_804832 : sel_804829;
  assign add_804836 = sel_804833 + 8'h01;
  assign sel_804837 = array_index_804676 == array_index_772876 ? add_804836 : sel_804833;
  assign add_804840 = sel_804837 + 8'h01;
  assign sel_804841 = array_index_804676 == array_index_772882 ? add_804840 : sel_804837;
  assign add_804844 = sel_804841 + 8'h01;
  assign sel_804845 = array_index_804676 == array_index_772888 ? add_804844 : sel_804841;
  assign add_804848 = sel_804845 + 8'h01;
  assign sel_804849 = array_index_804676 == array_index_772894 ? add_804848 : sel_804845;
  assign add_804852 = sel_804849 + 8'h01;
  assign sel_804853 = array_index_804676 == array_index_772900 ? add_804852 : sel_804849;
  assign add_804856 = sel_804853 + 8'h01;
  assign sel_804857 = array_index_804676 == array_index_772906 ? add_804856 : sel_804853;
  assign add_804860 = sel_804857 + 8'h01;
  assign sel_804861 = array_index_804676 == array_index_772912 ? add_804860 : sel_804857;
  assign add_804864 = sel_804861 + 8'h01;
  assign sel_804865 = array_index_804676 == array_index_772918 ? add_804864 : sel_804861;
  assign add_804868 = sel_804865 + 8'h01;
  assign sel_804869 = array_index_804676 == array_index_772924 ? add_804868 : sel_804865;
  assign add_804872 = sel_804869 + 8'h01;
  assign sel_804873 = array_index_804676 == array_index_772930 ? add_804872 : sel_804869;
  assign add_804876 = sel_804873 + 8'h01;
  assign sel_804877 = array_index_804676 == array_index_772936 ? add_804876 : sel_804873;
  assign add_804880 = sel_804877 + 8'h01;
  assign sel_804881 = array_index_804676 == array_index_772942 ? add_804880 : sel_804877;
  assign add_804884 = sel_804881 + 8'h01;
  assign sel_804885 = array_index_804676 == array_index_772948 ? add_804884 : sel_804881;
  assign add_804888 = sel_804885 + 8'h01;
  assign sel_804889 = array_index_804676 == array_index_772954 ? add_804888 : sel_804885;
  assign add_804892 = sel_804889 + 8'h01;
  assign sel_804893 = array_index_804676 == array_index_772960 ? add_804892 : sel_804889;
  assign add_804896 = sel_804893 + 8'h01;
  assign sel_804897 = array_index_804676 == array_index_772966 ? add_804896 : sel_804893;
  assign add_804900 = sel_804897 + 8'h01;
  assign sel_804901 = array_index_804676 == array_index_772972 ? add_804900 : sel_804897;
  assign add_804904 = sel_804901 + 8'h01;
  assign sel_804905 = array_index_804676 == array_index_772978 ? add_804904 : sel_804901;
  assign add_804908 = sel_804905 + 8'h01;
  assign sel_804909 = array_index_804676 == array_index_772984 ? add_804908 : sel_804905;
  assign add_804912 = sel_804909 + 8'h01;
  assign sel_804913 = array_index_804676 == array_index_772990 ? add_804912 : sel_804909;
  assign add_804916 = sel_804913 + 8'h01;
  assign sel_804917 = array_index_804676 == array_index_772996 ? add_804916 : sel_804913;
  assign add_804920 = sel_804917 + 8'h01;
  assign sel_804921 = array_index_804676 == array_index_773002 ? add_804920 : sel_804917;
  assign add_804924 = sel_804921 + 8'h01;
  assign sel_804925 = array_index_804676 == array_index_773008 ? add_804924 : sel_804921;
  assign add_804928 = sel_804925 + 8'h01;
  assign sel_804929 = array_index_804676 == array_index_773014 ? add_804928 : sel_804925;
  assign add_804932 = sel_804929 + 8'h01;
  assign sel_804933 = array_index_804676 == array_index_773020 ? add_804932 : sel_804929;
  assign add_804936 = sel_804933 + 8'h01;
  assign sel_804937 = array_index_804676 == array_index_773026 ? add_804936 : sel_804933;
  assign add_804940 = sel_804937 + 8'h01;
  assign sel_804941 = array_index_804676 == array_index_773032 ? add_804940 : sel_804937;
  assign add_804944 = sel_804941 + 8'h01;
  assign sel_804945 = array_index_804676 == array_index_773038 ? add_804944 : sel_804941;
  assign add_804948 = sel_804945 + 8'h01;
  assign sel_804949 = array_index_804676 == array_index_773044 ? add_804948 : sel_804945;
  assign add_804952 = sel_804949 + 8'h01;
  assign sel_804953 = array_index_804676 == array_index_773050 ? add_804952 : sel_804949;
  assign add_804956 = sel_804953 + 8'h01;
  assign sel_804957 = array_index_804676 == array_index_773056 ? add_804956 : sel_804953;
  assign add_804960 = sel_804957 + 8'h01;
  assign sel_804961 = array_index_804676 == array_index_773062 ? add_804960 : sel_804957;
  assign add_804964 = sel_804961 + 8'h01;
  assign sel_804965 = array_index_804676 == array_index_773068 ? add_804964 : sel_804961;
  assign add_804968 = sel_804965 + 8'h01;
  assign sel_804969 = array_index_804676 == array_index_773074 ? add_804968 : sel_804965;
  assign add_804972 = sel_804969 + 8'h01;
  assign sel_804973 = array_index_804676 == array_index_773080 ? add_804972 : sel_804969;
  assign add_804976 = sel_804973 + 8'h01;
  assign sel_804977 = array_index_804676 == array_index_773086 ? add_804976 : sel_804973;
  assign add_804980 = sel_804977 + 8'h01;
  assign sel_804981 = array_index_804676 == array_index_773092 ? add_804980 : sel_804977;
  assign add_804984 = sel_804981 + 8'h01;
  assign sel_804985 = array_index_804676 == array_index_773098 ? add_804984 : sel_804981;
  assign add_804988 = sel_804985 + 8'h01;
  assign sel_804989 = array_index_804676 == array_index_773104 ? add_804988 : sel_804985;
  assign add_804992 = sel_804989 + 8'h01;
  assign sel_804993 = array_index_804676 == array_index_773110 ? add_804992 : sel_804989;
  assign add_804996 = sel_804993 + 8'h01;
  assign sel_804997 = array_index_804676 == array_index_773116 ? add_804996 : sel_804993;
  assign add_805000 = sel_804997 + 8'h01;
  assign sel_805001 = array_index_804676 == array_index_773122 ? add_805000 : sel_804997;
  assign add_805004 = sel_805001 + 8'h01;
  assign sel_805005 = array_index_804676 == array_index_773128 ? add_805004 : sel_805001;
  assign add_805008 = sel_805005 + 8'h01;
  assign sel_805009 = array_index_804676 == array_index_773134 ? add_805008 : sel_805005;
  assign add_805012 = sel_805009 + 8'h01;
  assign sel_805013 = array_index_804676 == array_index_773140 ? add_805012 : sel_805009;
  assign add_805016 = sel_805013 + 8'h01;
  assign sel_805017 = array_index_804676 == array_index_773146 ? add_805016 : sel_805013;
  assign add_805020 = sel_805017 + 8'h01;
  assign sel_805021 = array_index_804676 == array_index_773152 ? add_805020 : sel_805017;
  assign add_805024 = sel_805021 + 8'h01;
  assign sel_805025 = array_index_804676 == array_index_773158 ? add_805024 : sel_805021;
  assign add_805028 = sel_805025 + 8'h01;
  assign sel_805029 = array_index_804676 == array_index_773164 ? add_805028 : sel_805025;
  assign add_805032 = sel_805029 + 8'h01;
  assign sel_805033 = array_index_804676 == array_index_773170 ? add_805032 : sel_805029;
  assign add_805037 = sel_805033 + 8'h01;
  assign array_index_805038 = set1_unflattened[7'h59];
  assign sel_805039 = array_index_804676 == array_index_773176 ? add_805037 : sel_805033;
  assign add_805042 = sel_805039 + 8'h01;
  assign sel_805043 = array_index_805038 == array_index_772632 ? add_805042 : sel_805039;
  assign add_805046 = sel_805043 + 8'h01;
  assign sel_805047 = array_index_805038 == array_index_772636 ? add_805046 : sel_805043;
  assign add_805050 = sel_805047 + 8'h01;
  assign sel_805051 = array_index_805038 == array_index_772644 ? add_805050 : sel_805047;
  assign add_805054 = sel_805051 + 8'h01;
  assign sel_805055 = array_index_805038 == array_index_772652 ? add_805054 : sel_805051;
  assign add_805058 = sel_805055 + 8'h01;
  assign sel_805059 = array_index_805038 == array_index_772660 ? add_805058 : sel_805055;
  assign add_805062 = sel_805059 + 8'h01;
  assign sel_805063 = array_index_805038 == array_index_772668 ? add_805062 : sel_805059;
  assign add_805066 = sel_805063 + 8'h01;
  assign sel_805067 = array_index_805038 == array_index_772676 ? add_805066 : sel_805063;
  assign add_805070 = sel_805067 + 8'h01;
  assign sel_805071 = array_index_805038 == array_index_772684 ? add_805070 : sel_805067;
  assign add_805074 = sel_805071 + 8'h01;
  assign sel_805075 = array_index_805038 == array_index_772690 ? add_805074 : sel_805071;
  assign add_805078 = sel_805075 + 8'h01;
  assign sel_805079 = array_index_805038 == array_index_772696 ? add_805078 : sel_805075;
  assign add_805082 = sel_805079 + 8'h01;
  assign sel_805083 = array_index_805038 == array_index_772702 ? add_805082 : sel_805079;
  assign add_805086 = sel_805083 + 8'h01;
  assign sel_805087 = array_index_805038 == array_index_772708 ? add_805086 : sel_805083;
  assign add_805090 = sel_805087 + 8'h01;
  assign sel_805091 = array_index_805038 == array_index_772714 ? add_805090 : sel_805087;
  assign add_805094 = sel_805091 + 8'h01;
  assign sel_805095 = array_index_805038 == array_index_772720 ? add_805094 : sel_805091;
  assign add_805098 = sel_805095 + 8'h01;
  assign sel_805099 = array_index_805038 == array_index_772726 ? add_805098 : sel_805095;
  assign add_805102 = sel_805099 + 8'h01;
  assign sel_805103 = array_index_805038 == array_index_772732 ? add_805102 : sel_805099;
  assign add_805106 = sel_805103 + 8'h01;
  assign sel_805107 = array_index_805038 == array_index_772738 ? add_805106 : sel_805103;
  assign add_805110 = sel_805107 + 8'h01;
  assign sel_805111 = array_index_805038 == array_index_772744 ? add_805110 : sel_805107;
  assign add_805114 = sel_805111 + 8'h01;
  assign sel_805115 = array_index_805038 == array_index_772750 ? add_805114 : sel_805111;
  assign add_805118 = sel_805115 + 8'h01;
  assign sel_805119 = array_index_805038 == array_index_772756 ? add_805118 : sel_805115;
  assign add_805122 = sel_805119 + 8'h01;
  assign sel_805123 = array_index_805038 == array_index_772762 ? add_805122 : sel_805119;
  assign add_805126 = sel_805123 + 8'h01;
  assign sel_805127 = array_index_805038 == array_index_772768 ? add_805126 : sel_805123;
  assign add_805130 = sel_805127 + 8'h01;
  assign sel_805131 = array_index_805038 == array_index_772774 ? add_805130 : sel_805127;
  assign add_805134 = sel_805131 + 8'h01;
  assign sel_805135 = array_index_805038 == array_index_772780 ? add_805134 : sel_805131;
  assign add_805138 = sel_805135 + 8'h01;
  assign sel_805139 = array_index_805038 == array_index_772786 ? add_805138 : sel_805135;
  assign add_805142 = sel_805139 + 8'h01;
  assign sel_805143 = array_index_805038 == array_index_772792 ? add_805142 : sel_805139;
  assign add_805146 = sel_805143 + 8'h01;
  assign sel_805147 = array_index_805038 == array_index_772798 ? add_805146 : sel_805143;
  assign add_805150 = sel_805147 + 8'h01;
  assign sel_805151 = array_index_805038 == array_index_772804 ? add_805150 : sel_805147;
  assign add_805154 = sel_805151 + 8'h01;
  assign sel_805155 = array_index_805038 == array_index_772810 ? add_805154 : sel_805151;
  assign add_805158 = sel_805155 + 8'h01;
  assign sel_805159 = array_index_805038 == array_index_772816 ? add_805158 : sel_805155;
  assign add_805162 = sel_805159 + 8'h01;
  assign sel_805163 = array_index_805038 == array_index_772822 ? add_805162 : sel_805159;
  assign add_805166 = sel_805163 + 8'h01;
  assign sel_805167 = array_index_805038 == array_index_772828 ? add_805166 : sel_805163;
  assign add_805170 = sel_805167 + 8'h01;
  assign sel_805171 = array_index_805038 == array_index_772834 ? add_805170 : sel_805167;
  assign add_805174 = sel_805171 + 8'h01;
  assign sel_805175 = array_index_805038 == array_index_772840 ? add_805174 : sel_805171;
  assign add_805178 = sel_805175 + 8'h01;
  assign sel_805179 = array_index_805038 == array_index_772846 ? add_805178 : sel_805175;
  assign add_805182 = sel_805179 + 8'h01;
  assign sel_805183 = array_index_805038 == array_index_772852 ? add_805182 : sel_805179;
  assign add_805186 = sel_805183 + 8'h01;
  assign sel_805187 = array_index_805038 == array_index_772858 ? add_805186 : sel_805183;
  assign add_805190 = sel_805187 + 8'h01;
  assign sel_805191 = array_index_805038 == array_index_772864 ? add_805190 : sel_805187;
  assign add_805194 = sel_805191 + 8'h01;
  assign sel_805195 = array_index_805038 == array_index_772870 ? add_805194 : sel_805191;
  assign add_805198 = sel_805195 + 8'h01;
  assign sel_805199 = array_index_805038 == array_index_772876 ? add_805198 : sel_805195;
  assign add_805202 = sel_805199 + 8'h01;
  assign sel_805203 = array_index_805038 == array_index_772882 ? add_805202 : sel_805199;
  assign add_805206 = sel_805203 + 8'h01;
  assign sel_805207 = array_index_805038 == array_index_772888 ? add_805206 : sel_805203;
  assign add_805210 = sel_805207 + 8'h01;
  assign sel_805211 = array_index_805038 == array_index_772894 ? add_805210 : sel_805207;
  assign add_805214 = sel_805211 + 8'h01;
  assign sel_805215 = array_index_805038 == array_index_772900 ? add_805214 : sel_805211;
  assign add_805218 = sel_805215 + 8'h01;
  assign sel_805219 = array_index_805038 == array_index_772906 ? add_805218 : sel_805215;
  assign add_805222 = sel_805219 + 8'h01;
  assign sel_805223 = array_index_805038 == array_index_772912 ? add_805222 : sel_805219;
  assign add_805226 = sel_805223 + 8'h01;
  assign sel_805227 = array_index_805038 == array_index_772918 ? add_805226 : sel_805223;
  assign add_805230 = sel_805227 + 8'h01;
  assign sel_805231 = array_index_805038 == array_index_772924 ? add_805230 : sel_805227;
  assign add_805234 = sel_805231 + 8'h01;
  assign sel_805235 = array_index_805038 == array_index_772930 ? add_805234 : sel_805231;
  assign add_805238 = sel_805235 + 8'h01;
  assign sel_805239 = array_index_805038 == array_index_772936 ? add_805238 : sel_805235;
  assign add_805242 = sel_805239 + 8'h01;
  assign sel_805243 = array_index_805038 == array_index_772942 ? add_805242 : sel_805239;
  assign add_805246 = sel_805243 + 8'h01;
  assign sel_805247 = array_index_805038 == array_index_772948 ? add_805246 : sel_805243;
  assign add_805250 = sel_805247 + 8'h01;
  assign sel_805251 = array_index_805038 == array_index_772954 ? add_805250 : sel_805247;
  assign add_805254 = sel_805251 + 8'h01;
  assign sel_805255 = array_index_805038 == array_index_772960 ? add_805254 : sel_805251;
  assign add_805258 = sel_805255 + 8'h01;
  assign sel_805259 = array_index_805038 == array_index_772966 ? add_805258 : sel_805255;
  assign add_805262 = sel_805259 + 8'h01;
  assign sel_805263 = array_index_805038 == array_index_772972 ? add_805262 : sel_805259;
  assign add_805266 = sel_805263 + 8'h01;
  assign sel_805267 = array_index_805038 == array_index_772978 ? add_805266 : sel_805263;
  assign add_805270 = sel_805267 + 8'h01;
  assign sel_805271 = array_index_805038 == array_index_772984 ? add_805270 : sel_805267;
  assign add_805274 = sel_805271 + 8'h01;
  assign sel_805275 = array_index_805038 == array_index_772990 ? add_805274 : sel_805271;
  assign add_805278 = sel_805275 + 8'h01;
  assign sel_805279 = array_index_805038 == array_index_772996 ? add_805278 : sel_805275;
  assign add_805282 = sel_805279 + 8'h01;
  assign sel_805283 = array_index_805038 == array_index_773002 ? add_805282 : sel_805279;
  assign add_805286 = sel_805283 + 8'h01;
  assign sel_805287 = array_index_805038 == array_index_773008 ? add_805286 : sel_805283;
  assign add_805290 = sel_805287 + 8'h01;
  assign sel_805291 = array_index_805038 == array_index_773014 ? add_805290 : sel_805287;
  assign add_805294 = sel_805291 + 8'h01;
  assign sel_805295 = array_index_805038 == array_index_773020 ? add_805294 : sel_805291;
  assign add_805298 = sel_805295 + 8'h01;
  assign sel_805299 = array_index_805038 == array_index_773026 ? add_805298 : sel_805295;
  assign add_805302 = sel_805299 + 8'h01;
  assign sel_805303 = array_index_805038 == array_index_773032 ? add_805302 : sel_805299;
  assign add_805306 = sel_805303 + 8'h01;
  assign sel_805307 = array_index_805038 == array_index_773038 ? add_805306 : sel_805303;
  assign add_805310 = sel_805307 + 8'h01;
  assign sel_805311 = array_index_805038 == array_index_773044 ? add_805310 : sel_805307;
  assign add_805314 = sel_805311 + 8'h01;
  assign sel_805315 = array_index_805038 == array_index_773050 ? add_805314 : sel_805311;
  assign add_805318 = sel_805315 + 8'h01;
  assign sel_805319 = array_index_805038 == array_index_773056 ? add_805318 : sel_805315;
  assign add_805322 = sel_805319 + 8'h01;
  assign sel_805323 = array_index_805038 == array_index_773062 ? add_805322 : sel_805319;
  assign add_805326 = sel_805323 + 8'h01;
  assign sel_805327 = array_index_805038 == array_index_773068 ? add_805326 : sel_805323;
  assign add_805330 = sel_805327 + 8'h01;
  assign sel_805331 = array_index_805038 == array_index_773074 ? add_805330 : sel_805327;
  assign add_805334 = sel_805331 + 8'h01;
  assign sel_805335 = array_index_805038 == array_index_773080 ? add_805334 : sel_805331;
  assign add_805338 = sel_805335 + 8'h01;
  assign sel_805339 = array_index_805038 == array_index_773086 ? add_805338 : sel_805335;
  assign add_805342 = sel_805339 + 8'h01;
  assign sel_805343 = array_index_805038 == array_index_773092 ? add_805342 : sel_805339;
  assign add_805346 = sel_805343 + 8'h01;
  assign sel_805347 = array_index_805038 == array_index_773098 ? add_805346 : sel_805343;
  assign add_805350 = sel_805347 + 8'h01;
  assign sel_805351 = array_index_805038 == array_index_773104 ? add_805350 : sel_805347;
  assign add_805354 = sel_805351 + 8'h01;
  assign sel_805355 = array_index_805038 == array_index_773110 ? add_805354 : sel_805351;
  assign add_805358 = sel_805355 + 8'h01;
  assign sel_805359 = array_index_805038 == array_index_773116 ? add_805358 : sel_805355;
  assign add_805362 = sel_805359 + 8'h01;
  assign sel_805363 = array_index_805038 == array_index_773122 ? add_805362 : sel_805359;
  assign add_805366 = sel_805363 + 8'h01;
  assign sel_805367 = array_index_805038 == array_index_773128 ? add_805366 : sel_805363;
  assign add_805370 = sel_805367 + 8'h01;
  assign sel_805371 = array_index_805038 == array_index_773134 ? add_805370 : sel_805367;
  assign add_805374 = sel_805371 + 8'h01;
  assign sel_805375 = array_index_805038 == array_index_773140 ? add_805374 : sel_805371;
  assign add_805378 = sel_805375 + 8'h01;
  assign sel_805379 = array_index_805038 == array_index_773146 ? add_805378 : sel_805375;
  assign add_805382 = sel_805379 + 8'h01;
  assign sel_805383 = array_index_805038 == array_index_773152 ? add_805382 : sel_805379;
  assign add_805386 = sel_805383 + 8'h01;
  assign sel_805387 = array_index_805038 == array_index_773158 ? add_805386 : sel_805383;
  assign add_805390 = sel_805387 + 8'h01;
  assign sel_805391 = array_index_805038 == array_index_773164 ? add_805390 : sel_805387;
  assign add_805394 = sel_805391 + 8'h01;
  assign sel_805395 = array_index_805038 == array_index_773170 ? add_805394 : sel_805391;
  assign add_805398 = sel_805395 + 8'h01;
  assign out = {array_index_805038 == array_index_773176 ? add_805398 : sel_805395, {set1_unflattened[89], set1_unflattened[88], set1_unflattened[87], set1_unflattened[86], set1_unflattened[85], set1_unflattened[84], set1_unflattened[83], set1_unflattened[82], set1_unflattened[81], set1_unflattened[80], set1_unflattened[79], set1_unflattened[78], set1_unflattened[77], set1_unflattened[76], set1_unflattened[75], set1_unflattened[74], set1_unflattened[73], set1_unflattened[72], set1_unflattened[71], set1_unflattened[70], set1_unflattened[69], set1_unflattened[68], set1_unflattened[67], set1_unflattened[66], set1_unflattened[65], set1_unflattened[64], set1_unflattened[63], set1_unflattened[62], set1_unflattened[61], set1_unflattened[60], set1_unflattened[59], set1_unflattened[58], set1_unflattened[57], set1_unflattened[56], set1_unflattened[55], set1_unflattened[54], set1_unflattened[53], set1_unflattened[52], set1_unflattened[51], set1_unflattened[50], set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[89], set2_unflattened[88], set2_unflattened[87], set2_unflattened[86], set2_unflattened[85], set2_unflattened[84], set2_unflattened[83], set2_unflattened[82], set2_unflattened[81], set2_unflattened[80], set2_unflattened[79], set2_unflattened[78], set2_unflattened[77], set2_unflattened[76], set2_unflattened[75], set2_unflattened[74], set2_unflattened[73], set2_unflattened[72], set2_unflattened[71], set2_unflattened[70], set2_unflattened[69], set2_unflattened[68], set2_unflattened[67], set2_unflattened[66], set2_unflattened[65], set2_unflattened[64], set2_unflattened[63], set2_unflattened[62], set2_unflattened[61], set2_unflattened[60], set2_unflattened[59], set2_unflattened[58], set2_unflattened[57], set2_unflattened[56], set2_unflattened[55], set2_unflattened[54], set2_unflattened[53], set2_unflattened[52], set2_unflattened[51], set2_unflattened[50], set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
