module min_hash(set1, set2, out);
  wire _00000_, _00001_, _00002_, _00003_, _00004_, _00005_, _00006_, _00007_, _00008_, _00009_, _00010_, _00011_, _00012_, _00013_, _00014_, _00015_, _00016_, _00017_, _00018_, _00019_, _00020_, _00021_, _00022_, _00023_, _00024_, _00025_, _00026_, _00027_, _00028_, _00029_, _00030_, _00031_, _00032_, _00033_, _00034_, _00035_, _00036_, _00037_, _00038_, _00039_, _00040_, _00041_, _00042_, _00043_, _00044_, _00045_, _00046_, _00047_, _00048_, _00049_, _00050_, _00051_, _00052_, _00053_, _00054_, _00055_, _00056_, _00057_, _00058_, _00059_, _00060_, _00061_, _00062_, _00063_, _00064_, _00065_, _00066_, _00067_, _00068_, _00069_, _00070_, _00071_, _00072_, _00073_, _00074_, _00075_, _00076_, _00077_, _00078_, _00079_, _00080_, _00081_, _00082_, _00083_, _00084_, _00085_, _00086_, _00087_, _00088_, _00089_, _00090_, _00091_, _00092_, _00093_, _00094_, _00095_, _00096_, _00097_, _00098_, _00099_, _00100_, _00101_, _00102_, _00103_, _00104_, _00105_, _00106_, _00107_, _00108_, _00109_, _00110_, _00111_, _00112_, _00113_, _00114_, _00115_, _00116_, _00117_, _00118_, _00119_, _00120_, _00121_, _00122_, _00123_, _00124_, _00125_, _00126_, _00127_, _00128_, _00129_, _00130_, _00131_, _00132_, _00133_, _00134_, _00135_, _00136_, _00137_, _00138_, _00139_, _00140_, _00141_, _00142_, _00143_, _00144_, _00145_, _00146_, _00147_, _00148_, _00149_, _00150_, _00151_, _00152_, _00153_, _00154_, _00155_, _00156_, _00157_, _00158_, _00159_, _00160_, _00161_, _00162_, _00163_, _00164_, _00165_, _00166_, _00167_, _00168_, _00169_, _00170_, _00171_, _00172_, _00173_, _00174_, _00175_, _00176_, _00177_, _00178_, _00179_, _00180_, _00181_, _00182_, _00183_, _00184_, _00185_, _00186_, _00187_, _00188_, _00189_, _00190_, _00191_, _00192_, _00193_, _00194_, _00195_, _00196_, _00197_, _00198_, _00199_, _00200_, _00201_, _00202_, _00203_, _00204_, _00205_, _00206_, _00207_, _00208_, _00209_, _00210_, _00211_, _00212_, _00213_, _00214_, _00215_, _00216_, _00217_, _00218_, _00219_, _00220_, _00221_, _00222_, _00223_, _00224_, _00225_, _00226_, _00227_, _00228_, _00229_, _00230_, _00231_, _00232_, _00233_, _00234_, _00235_, _00236_, _00237_, _00238_, _00239_, _00240_, _00241_, _00242_, _00243_, _00244_, _00245_, _00246_, _00247_, _00248_, _00249_, _00250_, _00251_, _00252_, _00253_, _00254_, _00255_, _00256_, _00257_, _00258_, _00259_, _00260_, _00261_, _00262_, _00263_, _00264_, _00265_, _00266_, _00267_, _00268_, _00269_, _00270_, _00271_, _00272_, _00273_, _00274_, _00275_, _00276_, _00277_, _00278_, _00279_, _00280_, _00281_, _00282_, _00283_, _00284_, _00285_, _00286_, _00287_, _00288_, _00289_, _00290_, _00291_, _00292_, _00293_, _00294_, _00295_, _00296_, _00297_, _00298_, _00299_, _00300_, _00301_, _00302_, _00303_, _00304_, _00305_, _00306_, _00307_, _00308_, _00309_, _00310_, _00311_, _00312_, _00313_, _00314_, _00315_, _00316_, _00317_, _00318_, _00319_, _00320_, _00321_, _00322_, _00323_, _00324_, _00325_, _00326_, _00327_, _00328_, _00329_, _00330_, _00331_, _00332_, _00333_, _00334_, _00335_, _00336_, _00337_, _00338_, _00339_, _00340_, _00341_, _00342_, _00343_, _00344_, _00345_, _00346_, _00347_, _00348_, _00349_, _00350_, _00351_, _00352_, _00353_, _00354_, _00355_, _00356_, _00357_, _00358_, _00359_, _00360_, _00361_, _00362_, _00363_, _00364_, _00365_, _00366_, _00367_, _00368_, _00369_, _00370_, _00371_, _00372_, _00373_, _00374_, _00375_, _00376_, _00377_, _00378_, _00379_, _00380_, _00381_, _00382_, _00383_, _00384_, _00385_, _00386_, _00387_, _00388_, _00389_, _00390_, _00391_, _00392_, _00393_, _00394_, _00395_, _00396_, _00397_, _00398_, _00399_, _00400_, _00401_, _00402_, _00403_, _00404_, _00405_, _00406_, _00407_, _00408_, _00409_, _00410_, _00411_, _00412_, _00413_, _00414_, _00415_, _00416_, _00417_, _00418_, _00419_, _00420_, _00421_, _00422_, _00423_, _00424_, _00425_, _00426_, _00427_, _00428_, _00429_, _00430_, _00431_, _00432_, _00433_, _00434_, _00435_, _00436_, _00437_, _00438_, _00439_, _00440_, _00441_, _00442_, _00443_, _00444_, _00445_, _00446_, _00447_, _00448_, _00449_, _00450_, _00451_, _00452_, _00453_, _00454_, _00455_, _00456_, _00457_, _00458_, _00459_, _00460_, _00461_, _00462_, _00463_, _00464_, _00465_, _00466_, _00467_, _00468_, _00469_, _00470_, _00471_, _00472_, _00473_, _00474_, _00475_, _00476_, _00477_, _00478_, _00479_, _00480_, _00481_, _00482_, _00483_, _00484_, _00485_, _00486_, _00487_, _00488_, _00489_, _00490_, _00491_, _00492_, _00493_, _00494_, _00495_, _00496_, _00497_, _00498_, _00499_, _00500_, _00501_, _00502_, _00503_, _00504_, _00505_, _00506_, _00507_, _00508_, _00509_, _00510_, _00511_, _00512_, _00513_, _00514_, _00515_, _00516_, _00517_, _00518_, _00519_, _00520_, _00521_, _00522_, _00523_, _00524_, _00525_, _00526_, _00527_, _00528_, _00529_, _00530_, _00531_, _00532_, _00533_, _00534_, _00535_, _00536_, _00537_, _00538_, _00539_, _00540_, _00541_, _00542_, _00543_, _00544_, _00545_, _00546_, _00547_, _00548_, _00549_, _00550_, _00551_, _00552_, _00553_, _00554_, _00555_, _00556_, _00557_, _00558_, _00559_, _00560_, _00561_, _00562_, _00563_, _00564_, _00565_, _00566_, _00567_, _00568_, _00569_, _00570_, _00571_, _00572_, _00573_, _00574_, _00575_, _00576_, _00577_, _00578_, _00579_, _00580_, _00581_, _00582_, _00583_, _00584_, _00585_, _00586_, _00587_, _00588_, _00589_, _00590_, _00591_, _00592_, _00593_, _00594_, _00595_, _00596_, _00597_, _00598_, _00599_, _00600_, _00601_, _00602_, _00603_, _00604_, _00605_, _00606_, _00607_, _00608_, _00609_, _00610_, _00611_, _00612_, _00613_, _00614_, _00615_, _00616_, _00617_, _00618_, _00619_, _00620_, _00621_, _00622_, _00623_, _00624_, _00625_, _00626_, _00627_, _00628_, _00629_, _00630_, _00631_, _00632_, _00633_, _00634_, _00635_, _00636_, _00637_, _00638_, _00639_, _00640_, _00641_, _00642_, _00643_, _00644_, _00645_, _00646_, _00647_, _00648_, _00649_, _00650_, _00651_, _00652_, _00653_, _00654_, _00655_, _00656_, _00657_, _00658_, _00659_, _00660_, _00661_, _00662_, _00663_, _00664_, _00665_, _00666_, _00667_, _00668_, _00669_, _00670_, _00671_, _00672_, _00673_, _00674_, _00675_, _00676_, _00677_, _00678_, _00679_, _00680_, _00681_, _00682_, _00683_, _00684_, _00685_, _00686_, _00687_, _00688_, _00689_, _00690_, _00691_, _00692_, _00693_, _00694_, _00695_, _00696_, _00697_, _00698_, _00699_, _00700_, _00701_, _00702_, _00703_, _00704_, _00705_, _00706_, _00707_, _00708_, _00709_, _00710_, _00711_, _00712_, _00713_, _00714_, _00715_, _00716_, _00717_, _00718_, _00719_, _00720_, _00721_, _00722_, _00723_, _00724_, _00725_, _00726_, _00727_, _00728_, _00729_, _00730_, _00731_, _00732_, _00733_, _00734_, _00735_, _00736_, _00737_, _00738_, _00739_, _00740_, _00741_, _00742_, _00743_, _00744_, _00745_, _00746_, _00747_, _00748_, _00749_, _00750_, _00751_, _00752_, _00753_, _00754_, _00755_, _00756_, _00757_, _00758_, _00759_, _00760_, _00761_, _00762_, _00763_, _00764_, _00765_, _00766_, _00767_, _00768_, _00769_, _00770_, _00771_, _00772_, _00773_, _00774_, _00775_, _00776_, _00777_, _00778_, _00779_, _00780_, _00781_, _00782_, _00783_, _00784_, _00785_, _00786_, _00787_, _00788_, _00789_, _00790_, _00791_, _00792_, _00793_, _00794_, _00795_, _00796_, _00797_, _00798_, _00799_, _00800_, _00801_, _00802_, _00803_, _00804_, _00805_, _00806_, _00807_, _00808_, _00809_, _00810_, _00811_, _00812_, _00813_, _00814_, _00815_, _00816_, _00817_, _00818_, _00819_, _00820_, _00821_, _00822_, _00823_, _00824_, _00825_, _00826_, _00827_, _00828_, _00829_, _00830_, _00831_, _00832_, _00833_, _00834_, _00835_, _00836_, _00837_, _00838_, _00839_, _00840_, _00841_, _00842_, _00843_, _00844_, _00845_, _00846_, _00847_, _00848_, _00849_, _00850_, _00851_, _00852_, _00853_, _00854_, _00855_, _00856_, _00857_, _00858_, _00859_, _00860_, _00861_, _00862_, _00863_, _00864_, _00865_, _00866_, _00867_, _00868_, _00869_, _00870_, _00871_, _00872_, _00873_, _00874_, _00875_, _00876_, _00877_, _00878_, _00879_, _00880_, _00881_, _00882_, _00883_, _00884_, _00885_, _00886_, _00887_, _00888_, _00889_, _00890_, _00891_, _00892_, _00893_, _00894_, _00895_, _00896_, _00897_, _00898_, _00899_, _00900_, _00901_, _00902_, _00903_, _00904_, _00905_, _00906_, _00907_, _00908_, _00909_, _00910_, _00911_, _00912_, _00913_, _00914_, _00915_, _00916_, _00917_, _00918_, _00919_, _00920_, _00921_, _00922_, _00923_, _00924_, _00925_, _00926_, _00927_, _00928_, _00929_, _00930_, _00931_, _00932_, _00933_, _00934_, _00935_, _00936_, _00937_, _00938_, _00939_, _00940_, _00941_, _00942_, _00943_, _00944_, _00945_, _00946_, _00947_, _00948_, _00949_, _00950_, _00951_, _00952_, _00953_, _00954_, _00955_, _00956_, _00957_, _00958_, _00959_, _00960_, _00961_, _00962_, _00963_, _00964_, _00965_, _00966_, _00967_, _00968_, _00969_, _00970_, _00971_, _00972_, _00973_, _00974_, _00975_, _00976_, _00977_, _00978_, _00979_, _00980_, _00981_, _00982_, _00983_, _00984_, _00985_, _00986_, _00987_, _00988_, _00989_, _00990_, _00991_, _00992_, _00993_, _00994_, _00995_, _00996_, _00997_, _00998_, _00999_, _01000_, _01001_, _01002_, _01003_, _01004_, _01005_, _01006_, _01007_, _01008_, _01009_, _01010_, _01011_, _01012_, _01013_, _01014_, _01015_, _01016_, _01017_, _01018_, _01019_, _01020_, _01021_, _01022_, _01023_, _01024_, _01025_, _01026_, _01027_, _01028_, _01029_, _01030_, _01031_, _01032_, _01033_, _01034_, _01035_, _01036_, _01037_, _01038_, _01039_, _01040_, _01041_, _01042_, _01043_, _01044_, _01045_, _01046_, _01047_, _01048_, _01049_, _01050_, _01051_, _01052_, _01053_, _01054_, _01055_, _01056_, _01057_, _01058_, _01059_, _01060_, _01061_, _01062_, _01063_, _01064_, _01065_, _01066_, _01067_, _01068_, _01069_, _01070_, _01071_, _01072_, _01073_, _01074_, _01075_, _01076_, _01077_, _01078_, _01079_, _01080_, _01081_, _01082_, _01083_, _01084_, _01085_, _01086_, _01087_, _01088_, _01089_, _01090_, _01091_, _01092_, _01093_, _01094_, _01095_, _01096_, _01097_, _01098_, _01099_, _01100_, _01101_, _01102_, _01103_, _01104_, _01105_, _01106_, _01107_, _01108_, _01109_, _01110_, _01111_, _01112_, _01113_, _01114_, _01115_, _01116_, _01117_, _01118_, _01119_, _01120_, _01121_, _01122_, _01123_, _01124_, _01125_, _01126_, _01127_, _01128_, _01129_, _01130_, _01131_, _01132_, _01133_, _01134_, _01135_, _01136_, _01137_, _01138_, _01139_, _01140_, _01141_, _01142_, _01143_, _01144_, _01145_, _01146_, _01147_, _01148_, _01149_, _01150_, _01151_, _01152_, _01153_, _01154_, _01155_, _01156_, _01157_, _01158_, _01159_, _01160_, _01161_, _01162_, _01163_, _01164_, _01165_, _01166_, _01167_, _01168_, _01169_, _01170_, _01171_, _01172_, _01173_, _01174_, _01175_, _01176_, _01177_, _01178_, _01179_, _01180_, _01181_, _01182_, _01183_, _01184_, _01185_, _01186_, _01187_, _01188_, _01189_, _01190_, _01191_, _01192_, _01193_, _01194_, _01195_, _01196_, _01197_, _01198_, _01199_, _01200_, _01201_, _01202_, _01203_, _01204_, _01205_, _01206_, _01207_, _01208_, _01209_, _01210_, _01211_, _01212_, _01213_, _01214_, _01215_, _01216_, _01217_, _01218_, _01219_, _01220_, _01221_, _01222_, _01223_, _01224_, _01225_, _01226_, _01227_, _01228_, _01229_, _01230_, _01231_, _01232_, _01233_, _01234_, _01235_, _01236_, _01237_, _01238_, _01239_, _01240_, _01241_, _01242_, _01243_, _01244_, _01245_, _01246_, _01247_, _01248_, _01249_, _01250_, _01251_, _01252_, _01253_, _01254_, _01255_, _01256_, _01257_, _01258_, _01259_, _01260_, _01261_, _01262_, _01263_, _01264_, _01265_, _01266_, _01267_, _01268_, _01269_, _01270_, _01271_, _01272_, _01273_, _01274_, _01275_, _01276_, _01277_, _01278_, _01279_, _01280_, _01281_, _01282_, _01283_, _01284_, _01285_, _01286_, _01287_, _01288_, _01289_, _01290_, _01291_, _01292_, _01293_, _01294_, _01295_, _01296_, _01297_, _01298_, _01299_, _01300_, _01301_, _01302_, _01303_, _01304_, _01305_, _01306_, _01307_, _01308_, _01309_, _01310_, _01311_, _01312_, _01313_, _01314_, _01315_, _01316_, _01317_, _01318_, _01319_, _01320_, _01321_, _01322_, _01323_, _01324_, _01325_, _01326_, _01327_, _01328_, _01329_, _01330_, _01331_, _01332_, _01333_, _01334_, _01335_, _01336_, _01337_, _01338_, _01339_, _01340_, _01341_, _01342_, _01343_, _01344_, _01345_, _01346_, _01347_, _01348_, _01349_, _01350_, _01351_, _01352_, _01353_, _01354_, _01355_, _01356_, _01357_, _01358_, _01359_, _01360_, _01361_, _01362_, _01363_, _01364_, _01365_, _01366_, _01367_, _01368_, _01369_, _01370_, _01371_, _01372_, _01373_, _01374_, _01375_, _01376_, _01377_, _01378_, _01379_, _01380_, _01381_, _01382_, _01383_, _01384_, _01385_, _01386_, _01387_, _01388_, _01389_, _01390_, _01391_, _01392_, _01393_, _01394_, _01395_, _01396_, _01397_, _01398_, _01399_, _01400_, _01401_, _01402_, _01403_, _01404_, _01405_, _01406_, _01407_, _01408_, _01409_, _01410_, _01411_, _01412_, _01413_, _01414_, _01415_, _01416_, _01417_, _01418_, _01419_, _01420_, _01421_, _01422_, _01423_, _01424_, _01425_, _01426_, _01427_, _01428_, _01429_, _01430_, _01431_, _01432_, _01433_, _01434_, _01435_, _01436_, _01437_, _01438_, _01439_, _01440_, _01441_, _01442_, _01443_, _01444_, _01445_, _01446_, _01447_, _01448_, _01449_, _01450_, _01451_, _01452_, _01453_, _01454_, _01455_, _01456_, _01457_, _01458_, _01459_, _01460_, _01461_, _01462_, _01463_, _01464_, _01465_, _01466_, _01467_, _01468_, _01469_, _01470_, _01471_, _01472_, _01473_, _01474_, _01475_, _01476_, _01477_, _01478_, _01479_, _01480_, _01481_, _01482_, _01483_, _01484_, _01485_, _01486_, _01487_, _01488_, _01489_, _01490_, _01491_, _01492_, _01493_, _01494_, _01495_, _01496_, _01497_, _01498_, _01499_, _01500_, _01501_, _01502_, _01503_, _01504_, _01505_, _01506_, _01507_, _01508_, _01509_, _01510_, _01511_, _01512_, _01513_, _01514_, _01515_, _01516_, _01517_, _01518_, _01519_, _01520_, _01521_, _01522_, _01523_, _01524_, _01525_, _01526_, _01527_, _01528_, _01529_, _01530_, _01531_, _01532_, _01533_, _01534_, _01535_, _01536_, _01537_, _01538_, _01539_, _01540_, _01541_, _01542_, _01543_, _01544_, _01545_, _01546_, _01547_, _01548_, _01549_, _01550_, _01551_, _01552_, _01553_, _01554_, _01555_, _01556_, _01557_, _01558_, _01559_, _01560_, _01561_, _01562_, _01563_, _01564_, _01565_, _01566_, _01567_, _01568_, _01569_, _01570_, _01571_, _01572_, _01573_, _01574_, _01575_, _01576_, _01577_, _01578_, _01579_, _01580_, _01581_, _01582_, _01583_, _01584_, _01585_, _01586_, _01587_, _01588_, _01589_, _01590_, _01591_, _01592_, _01593_, _01594_, _01595_, _01596_, _01597_, _01598_, _01599_, _01600_, _01601_, _01602_, _01603_, _01604_, _01605_, _01606_, _01607_, _01608_, _01609_, _01610_, _01611_, _01612_, _01613_, _01614_, _01615_, _01616_, _01617_, _01618_, _01619_, _01620_, _01621_, _01622_, _01623_, _01624_, _01625_, _01626_, _01627_, _01628_, _01629_, _01630_, _01631_, _01632_, _01633_, _01634_, _01635_, _01636_, _01637_, _01638_, _01639_, _01640_, _01641_, _01642_, _01643_, _01644_, _01645_, _01646_, _01647_, _01648_, _01649_, _01650_, _01651_, _01652_, _01653_, _01654_, _01655_, _01656_, _01657_, _01658_, _01659_, _01660_, _01661_, _01662_, _01663_, _01664_, _01665_, _01666_, _01667_, _01668_, _01669_, _01670_, _01671_, _01672_, _01673_, _01674_, _01675_, _01676_, _01677_, _01678_, _01679_, _01680_, _01681_, _01682_, _01683_, _01684_, _01685_, _01686_, _01687_, _01688_, _01689_, _01690_, _01691_, _01692_, _01693_, _01694_, _01695_, _01696_, _01697_, _01698_, _01699_, _01700_, _01701_, _01702_, _01703_, _01704_, _01705_, _01706_, _01707_, _01708_, _01709_, _01710_, _01711_, _01712_, _01713_, _01714_, _01715_, _01716_, _01717_, _01718_, _01719_, _01720_, _01721_, _01722_, _01723_, _01724_, _01725_, _01726_, _01727_, _01728_, _01729_, _01730_, _01731_, _01732_, _01733_, _01734_, _01735_, _01736_, _01737_, _01738_, _01739_, _01740_, _01741_, _01742_, _01743_, _01744_, _01745_, _01746_, _01747_, _01748_, _01749_, _01750_, _01751_, _01752_, _01753_, _01754_, _01755_, _01756_, _01757_, _01758_, _01759_, _01760_, _01761_, _01762_, _01763_, _01764_, _01765_, _01766_, _01767_, _01768_, _01769_, _01770_, _01771_, _01772_, _01773_, _01774_, _01775_, _01776_, _01777_, _01778_, _01779_, _01780_, _01781_, _01782_, _01783_, _01784_, _01785_, _01786_, _01787_, _01788_, _01789_, _01790_, _01791_, _01792_, _01793_, _01794_, _01795_, _01796_, _01797_, _01798_, _01799_, _01800_, _01801_, _01802_, _01803_, _01804_, _01805_, _01806_, _01807_, _01808_, _01809_, _01810_, _01811_, _01812_, _01813_, _01814_, _01815_, _01816_, _01817_, _01818_, _01819_, _01820_, _01821_, _01822_, _01823_, _01824_, _01825_, _01826_, _01827_, _01828_, _01829_, _01830_, _01831_, _01832_, _01833_, _01834_, _01835_, _01836_, _01837_, _01838_, _01839_, _01840_, _01841_, _01842_, _01843_, _01844_, _01845_, _01846_, _01847_, _01848_, _01849_, _01850_, _01851_, _01852_, _01853_, _01854_, _01855_, _01856_, _01857_, _01858_, _01859_, _01860_, _01861_, _01862_, _01863_, _01864_, _01865_, _01866_, _01867_, _01868_, _01869_, _01870_, _01871_, _01872_, _01873_, _01874_, _01875_, _01876_, _01877_, _01878_, _01879_, _01880_, _01881_, _01882_, _01883_, _01884_, _01885_, _01886_, _01887_, _01888_, _01889_, _01890_, _01891_, _01892_, _01893_, _01894_, _01895_, _01896_, _01897_, _01898_, _01899_, _01900_, _01901_, _01902_, _01903_, _01904_, _01905_, _01906_, _01907_, _01908_, _01909_, _01910_, _01911_, _01912_, _01913_, _01914_, _01915_, _01916_, _01917_, _01918_, _01919_, _01920_, _01921_, _01922_, _01923_, _01924_, _01925_, _01926_, _01927_, _01928_, _01929_, _01930_, _01931_, _01932_, _01933_, _01934_, _01935_, _01936_, _01937_, _01938_, _01939_, _01940_, _01941_, _01942_, _01943_, _01944_, _01945_, _01946_, _01947_, _01948_, _01949_, _01950_, _01951_, _01952_, _01953_, _01954_, _01955_, _01956_, _01957_, _01958_, _01959_, _01960_, _01961_, _01962_, _01963_, _01964_, _01965_, _01966_, _01967_, _01968_, _01969_, _01970_, _01971_, _01972_, _01973_, _01974_, _01975_, _01976_, _01977_, _01978_, _01979_, _01980_, _01981_, _01982_, _01983_, _01984_, _01985_, _01986_, _01987_, _01988_, _01989_, _01990_, _01991_, _01992_, _01993_, _01994_, _01995_, _01996_, _01997_, _01998_, _01999_, _02000_, _02001_, _02002_, _02003_, _02004_, _02005_, _02006_, _02007_, _02008_, _02009_, _02010_, _02011_, _02012_, _02013_, _02014_, _02015_, _02016_, _02017_, _02018_, _02019_, _02020_, _02021_, _02022_, _02023_, _02024_, _02025_, _02026_, _02027_, _02028_, _02029_, _02030_, _02031_, _02032_, _02033_, _02034_, _02035_, _02036_, _02037_, _02038_, _02039_, _02040_, _02041_, _02042_, _02043_, _02044_, _02045_, _02046_, _02047_, _02048_, _02049_, _02050_, _02051_, _02052_, _02053_, _02054_, _02055_, _02056_, _02057_, _02058_, _02059_, _02060_, _02061_, _02062_, _02063_, _02064_, _02065_, _02066_, _02067_, _02068_, _02069_, _02070_, _02071_, _02072_, _02073_, _02074_, _02075_, _02076_, _02077_, _02078_, _02079_, _02080_, _02081_, _02082_, _02083_, _02084_, _02085_, _02086_, _02087_, _02088_, _02089_, _02090_, _02091_, _02092_, _02093_, _02094_, _02095_, _02096_, _02097_, _02098_, _02099_, _02100_, _02101_, _02102_, _02103_, _02104_, _02105_, _02106_, _02107_, _02108_, _02109_, _02110_, _02111_, _02112_, _02113_, _02114_, _02115_, _02116_, _02117_, _02118_, _02119_, _02120_, _02121_, _02122_, _02123_, _02124_, _02125_, _02126_, _02127_, _02128_, _02129_, _02130_, _02131_, _02132_, _02133_, _02134_, _02135_, _02136_, _02137_, _02138_, _02139_, _02140_, _02141_, _02142_, _02143_, _02144_, _02145_, _02146_, _02147_, _02148_, _02149_, _02150_, _02151_, _02152_, _02153_, _02154_, _02155_, _02156_, _02157_, _02158_, _02159_, _02160_, _02161_, _02162_, _02163_, _02164_, _02165_, _02166_, _02167_, _02168_, _02169_, _02170_, _02171_, _02172_, _02173_, _02174_, _02175_, _02176_, _02177_, _02178_, _02179_, _02180_, _02181_, _02182_, _02183_, _02184_, _02185_, _02186_, _02187_, _02188_, _02189_, _02190_, _02191_, _02192_, _02193_, _02194_, _02195_, _02196_, _02197_, _02198_, _02199_, _02200_, _02201_, _02202_, _02203_, _02204_, _02205_, _02206_, _02207_, _02208_, _02209_, _02210_, _02211_, _02212_, _02213_, _02214_, _02215_, _02216_, _02217_, _02218_, _02219_, _02220_, _02221_, _02222_, _02223_, _02224_, _02225_, _02226_, _02227_, _02228_, _02229_, _02230_, _02231_, _02232_, _02233_, _02234_, _02235_, _02236_, _02237_, _02238_, _02239_, _02240_, _02241_, _02242_, _02243_, _02244_, _02245_, _02246_, _02247_, _02248_, _02249_, _02250_, _02251_, _02252_, _02253_, _02254_, _02255_, _02256_, _02257_, _02258_, _02259_, _02260_, _02261_, _02262_, _02263_, _02264_, _02265_, _02266_, _02267_, _02268_, _02269_, _02270_, _02271_, _02272_, _02273_, _02274_, _02275_, _02276_, _02277_, _02278_, _02279_, _02280_, _02281_, _02282_, _02283_, _02284_, _02285_, _02286_, _02287_, _02288_, _02289_, _02290_, _02291_, _02292_, _02293_, _02294_, _02295_, _02296_, _02297_, _02298_, _02299_, _02300_, _02301_, _02302_, _02303_, _02304_, _02305_, _02306_, _02307_, _02308_, _02309_, _02310_, _02311_, _02312_, _02313_, _02314_, _02315_, _02316_, _02317_, _02318_, _02319_, _02320_, _02321_, _02322_, _02323_, _02324_, _02325_, _02326_, _02327_, _02328_, _02329_, _02330_, _02331_, _02332_, _02333_, _02334_, _02335_, _02336_, _02337_, _02338_, _02339_, _02340_, _02341_, _02342_, _02343_, _02344_, _02345_, _02346_, _02347_, _02348_, _02349_, _02350_, _02351_, _02352_, _02353_, _02354_, _02355_, _02356_, _02357_, _02358_, _02359_, _02360_, _02361_, _02362_, _02363_, _02364_, _02365_, _02366_, _02367_, _02368_, _02369_, _02370_, _02371_, _02372_, _02373_, _02374_, _02375_, _02376_, _02377_, _02378_, _02379_, _02380_, _02381_, _02382_, _02383_, _02384_, _02385_, _02386_, _02387_, _02388_, _02389_, _02390_, _02391_, _02392_, _02393_, _02394_, _02395_, _02396_, _02397_, _02398_, _02399_, _02400_, _02401_, _02402_, _02403_, _02404_, _02405_, _02406_, _02407_, _02408_, _02409_, _02410_, _02411_, _02412_, _02413_, _02414_, _02415_, _02416_, _02417_, _02418_, _02419_, _02420_, _02421_, _02422_, _02423_, _02424_, _02425_, _02426_, _02427_, _02428_, _02429_, _02430_, _02431_, _02432_, _02433_, _02434_, _02435_, _02436_, _02437_, _02438_, _02439_, _02440_, _02441_, _02442_, _02443_, _02444_, _02445_, _02446_, _02447_, _02448_, _02449_, _02450_, _02451_, _02452_, _02453_, _02454_, _02455_, _02456_, _02457_, _02458_, _02459_, _02460_, _02461_, _02462_, _02463_, _02464_, _02465_, _02466_, _02467_, _02468_, _02469_, _02470_, _02471_, _02472_, _02473_, _02474_, _02475_, _02476_, _02477_, _02478_, _02479_, _02480_, _02481_, _02482_, _02483_, _02484_, _02485_, _02486_, _02487_, _02488_, _02489_, _02490_, _02491_, _02492_, _02493_, _02494_, _02495_, _02496_, _02497_, _02498_, _02499_, _02500_, _02501_, _02502_, _02503_, _02504_, _02505_, _02506_, _02507_, _02508_, _02509_, _02510_, _02511_, _02512_, _02513_, _02514_, _02515_, _02516_, _02517_, _02518_, _02519_, _02520_, _02521_, _02522_, _02523_, _02524_, _02525_, _02526_, _02527_, _02528_, _02529_, _02530_, _02531_, _02532_, _02533_, _02534_, _02535_, _02536_, _02537_, _02538_, _02539_, _02540_, _02541_, _02542_, _02543_, _02544_, _02545_, _02546_, _02547_, _02548_, _02549_, _02550_, _02551_, _02552_, _02553_, _02554_, _02555_, _02556_, _02557_, _02558_, _02559_, _02560_, _02561_, _02562_, _02563_, _02564_, _02565_, _02566_, _02567_, _02568_, _02569_, _02570_, _02571_, _02572_, _02573_, _02574_, _02575_, _02576_, _02577_, _02578_, _02579_, _02580_, _02581_, _02582_, _02583_, _02584_, _02585_, _02586_, _02587_, _02588_, _02589_, _02590_, _02591_, _02592_, _02593_, _02594_, _02595_, _02596_, _02597_, _02598_, _02599_, _02600_, _02601_, _02602_, _02603_, _02604_, _02605_, _02606_, _02607_, _02608_, _02609_, _02610_, _02611_, _02612_, _02613_, _02614_, _02615_, _02616_, _02617_, _02618_, _02619_, _02620_, _02621_, _02622_, _02623_, _02624_, _02625_, _02626_, _02627_, _02628_, _02629_, _02630_, _02631_, _02632_, _02633_, _02634_, _02635_, _02636_, _02637_, _02638_, _02639_, _02640_, _02641_, _02642_, _02643_, _02644_, _02645_, _02646_, _02647_, _02648_, _02649_, _02650_, _02651_, _02652_, _02653_, _02654_, _02655_, _02656_, _02657_, _02658_, _02659_, _02660_, _02661_, _02662_, _02663_, _02664_, _02665_, _02666_, _02667_, _02668_, _02669_, _02670_, _02671_, _02672_, _02673_, _02674_, _02675_, _02676_, _02677_, _02678_, _02679_, _02680_, _02681_, _02682_, _02683_, _02684_, _02685_, _02686_, _02687_, _02688_, _02689_, _02690_, _02691_, _02692_, _02693_, _02694_, _02695_, _02696_, _02697_, _02698_, _02699_, _02700_, _02701_, _02702_, _02703_, _02704_, _02705_, _02706_, _02707_, _02708_, _02709_, _02710_, _02711_, _02712_, _02713_, _02714_, _02715_, _02716_, _02717_, _02718_, _02719_, _02720_, _02721_, _02722_, _02723_, _02724_, _02725_, _02726_, _02727_, _02728_, _02729_, _02730_, _02731_, _02732_, _02733_, _02734_, _02735_, _02736_, _02737_, _02738_, _02739_, _02740_, _02741_, _02742_, _02743_, _02744_, _02745_, _02746_, _02747_, _02748_, _02749_, _02750_, _02751_, _02752_, _02753_, _02754_, _02755_, _02756_, _02757_, _02758_, _02759_, _02760_, _02761_, _02762_, _02763_, _02764_, _02765_, _02766_, _02767_, _02768_, _02769_, _02770_, _02771_, _02772_, _02773_, _02774_, _02775_, _02776_, _02777_, _02778_, _02779_, _02780_, _02781_, _02782_, _02783_, _02784_, _02785_, _02786_, _02787_, _02788_, _02789_, _02790_, _02791_, _02792_, _02793_, _02794_, _02795_, _02796_, _02797_, _02798_, _02799_, _02800_, _02801_, _02802_, _02803_, _02804_, _02805_, _02806_, _02807_, _02808_, _02809_, _02810_, _02811_, _02812_, _02813_, _02814_, _02815_, _02816_, _02817_, _02818_, _02819_, _02820_, _02821_, _02822_, _02823_, _02824_, _02825_, _02826_, _02827_, _02828_, _02829_, _02830_, _02831_, _02832_, _02833_, _02834_, _02835_, _02836_, _02837_, _02838_, _02839_, _02840_, _02841_, _02842_, _02843_, _02844_, _02845_, _02846_, _02847_, _02848_, _02849_, _02850_, _02851_, _02852_, _02853_, _02854_, _02855_, _02856_, _02857_, _02858_, _02859_, _02860_, _02861_, _02862_, _02863_, _02864_, _02865_, _02866_, _02867_, _02868_, _02869_, _02870_, _02871_, _02872_, _02873_, _02874_, _02875_, _02876_, _02877_, _02878_, _02879_, _02880_, _02881_, _02882_, _02883_, _02884_, _02885_, _02886_, _02887_, _02888_, _02889_, _02890_, _02891_, _02892_, _02893_, _02894_, _02895_, _02896_, _02897_, _02898_, _02899_, _02900_, _02901_, _02902_, _02903_, _02904_, _02905_, _02906_, _02907_, _02908_, _02909_, _02910_, _02911_, _02912_, _02913_, _02914_, _02915_, _02916_, _02917_, _02918_, _02919_, _02920_, _02921_, _02922_, _02923_, _02924_, _02925_, _02926_, _02927_, _02928_, _02929_, _02930_, _02931_, _02932_, _02933_, _02934_, _02935_, _02936_, _02937_, _02938_, _02939_, _02940_, _02941_, _02942_, _02943_, _02944_, _02945_, _02946_, _02947_, _02948_, _02949_, _02950_, _02951_, _02952_, _02953_, _02954_, _02955_, _02956_, _02957_, _02958_, _02959_, _02960_, _02961_, _02962_, _02963_, _02964_, _02965_, _02966_, _02967_, _02968_, _02969_, _02970_, _02971_, _02972_, _02973_, _02974_, _02975_, _02976_, _02977_, _02978_, _02979_, _02980_, _02981_, _02982_, _02983_, _02984_, _02985_, _02986_, _02987_, _02988_, _02989_, _02990_, _02991_, _02992_, _02993_, _02994_, _02995_, _02996_, _02997_, _02998_, _02999_, _03000_, _03001_, _03002_, _03003_, _03004_, _03005_, _03006_, _03007_, _03008_, _03009_, _03010_, _03011_, _03012_, _03013_, _03014_, _03015_, _03016_, _03017_, _03018_, _03019_, _03020_, _03021_, _03022_, _03023_, _03024_, _03025_, _03026_, _03027_, _03028_, _03029_, _03030_, _03031_, _03032_, _03033_, _03034_, _03035_, _03036_, _03037_, _03038_, _03039_, _03040_, _03041_, _03042_, _03043_, _03044_, _03045_, _03046_, _03047_, _03048_, _03049_, _03050_, _03051_, _03052_, _03053_, _03054_, _03055_, _03056_, _03057_, _03058_, _03059_, _03060_, _03061_, _03062_, _03063_, _03064_, _03065_, _03066_, _03067_, _03068_, _03069_, _03070_, _03071_, _03072_, _03073_, _03074_, _03075_, _03076_, _03077_, _03078_, _03079_, _03080_, _03081_, _03082_, _03083_, _03084_, _03085_, _03086_, _03087_, _03088_, _03089_, _03090_, _03091_, _03092_, _03093_, _03094_, _03095_, _03096_, _03097_, _03098_, _03099_, _03100_, _03101_, _03102_, _03103_, _03104_, _03105_, _03106_, _03107_, _03108_, _03109_, _03110_, _03111_, _03112_, _03113_, _03114_, _03115_, _03116_, _03117_, _03118_, _03119_, _03120_, _03121_, _03122_, _03123_, _03124_, _03125_, _03126_, _03127_, _03128_, _03129_, _03130_, _03131_, _03132_, _03133_, _03134_, _03135_, _03136_, _03137_, _03138_, _03139_, _03140_, _03141_, _03142_, _03143_, _03144_, _03145_, _03146_, _03147_, _03148_, _03149_, _03150_, _03151_, _03152_, _03153_, _03154_, _03155_, _03156_, _03157_, _03158_, _03159_, _03160_, _03161_, _03162_, _03163_, _03164_, _03165_, _03166_, _03167_, _03168_, _03169_, _03170_, _03171_, _03172_, _03173_, _03174_, _03175_, _03176_, _03177_, _03178_, _03179_, _03180_, _03181_, _03182_, _03183_, _03184_, _03185_, _03186_, _03187_, _03188_, _03189_, _03190_, _03191_, _03192_, _03193_, _03194_, _03195_, _03196_, _03197_, _03198_, _03199_, _03200_, _03201_, _03202_, _03203_, _03204_, _03205_, _03206_, _03207_, _03208_, _03209_, _03210_, _03211_, _03212_, _03213_, _03214_, _03215_, _03216_, _03217_, _03218_, _03219_, _03220_, _03221_, _03222_, _03223_, _03224_, _03225_, _03226_, _03227_, _03228_, _03229_, _03230_, _03231_, _03232_, _03233_, _03234_, _03235_, _03236_, _03237_, _03238_, _03239_, _03240_, _03241_, _03242_, _03243_, _03244_, _03245_, _03246_, _03247_, _03248_, _03249_, _03250_, _03251_, _03252_, _03253_, _03254_, _03255_, _03256_, _03257_, _03258_, _03259_, _03260_, _03261_, _03262_, _03263_, _03264_, _03265_, _03266_, _03267_, _03268_, _03269_, _03270_, _03271_, _03272_, _03273_, _03274_, _03275_, _03276_, _03277_, _03278_, _03279_, _03280_, _03281_, _03282_, _03283_, _03284_, _03285_, _03286_, _03287_, _03288_, _03289_, _03290_, _03291_, _03292_, _03293_, _03294_, _03295_, _03296_, _03297_, _03298_, _03299_, _03300_, _03301_, _03302_, _03303_, _03304_, _03305_, _03306_, _03307_, _03308_, _03309_, _03310_, _03311_, _03312_, _03313_, _03314_, _03315_, _03316_, _03317_, _03318_, _03319_, _03320_, _03321_, _03322_, _03323_, _03324_, _03325_, _03326_, _03327_, _03328_, _03329_, _03330_, _03331_, _03332_, _03333_, _03334_, _03335_, _03336_, _03337_, _03338_, _03339_, _03340_, _03341_, _03342_, _03343_, _03344_, _03345_, _03346_, _03347_, _03348_, _03349_, _03350_, _03351_, _03352_, _03353_, _03354_, _03355_, _03356_, _03357_, _03358_, _03359_, _03360_, _03361_, _03362_, _03363_, _03364_, _03365_, _03366_, _03367_, _03368_, _03369_, _03370_, _03371_, _03372_, _03373_, _03374_, _03375_, _03376_, _03377_, _03378_, _03379_, _03380_, _03381_, _03382_, _03383_, _03384_, _03385_, _03386_, _03387_, _03388_, _03389_, _03390_, _03391_, _03392_, _03393_, _03394_, _03395_, _03396_, _03397_, _03398_, _03399_, _03400_, _03401_, _03402_, _03403_, _03404_, _03405_, _03406_, _03407_, _03408_, _03409_, _03410_, _03411_, _03412_, _03413_, _03414_, _03415_, _03416_, _03417_, _03418_, _03419_, _03420_, _03421_, _03422_, _03423_, _03424_, _03425_, _03426_, _03427_, _03428_, _03429_, _03430_, _03431_, _03432_, _03433_, _03434_, _03435_, _03436_, _03437_, _03438_, _03439_, _03440_, _03441_, _03442_, _03443_, _03444_, _03445_, _03446_, _03447_, _03448_, _03449_, _03450_, _03451_, _03452_, _03453_, _03454_, _03455_, _03456_, _03457_, _03458_, _03459_, _03460_, _03461_, _03462_, _03463_, _03464_, _03465_, _03466_, _03467_, _03468_, _03469_, _03470_, _03471_, _03472_, _03473_, _03474_, _03475_, _03476_, _03477_, _03478_, _03479_, _03480_, _03481_, _03482_, _03483_, _03484_, _03485_, _03486_, _03487_, _03488_, _03489_, _03490_, _03491_, _03492_, _03493_, _03494_, _03495_, _03496_, _03497_, _03498_, _03499_, _03500_, _03501_, _03502_, _03503_, _03504_, _03505_, _03506_, _03507_, _03508_, _03509_, _03510_, _03511_, _03512_, _03513_, _03514_, _03515_, _03516_, _03517_, _03518_, _03519_, _03520_, _03521_, _03522_, _03523_, _03524_, _03525_, _03526_, _03527_, _03528_, _03529_, _03530_, _03531_, _03532_, _03533_, _03534_, _03535_, _03536_, _03537_, _03538_, _03539_, _03540_, _03541_, _03542_, _03543_, _03544_, _03545_, _03546_, _03547_, _03548_, _03549_, _03550_, _03551_, _03552_, _03553_, _03554_, _03555_, _03556_, _03557_, _03558_, _03559_, _03560_, _03561_, _03562_, _03563_, _03564_, _03565_, _03566_, _03567_, _03568_, _03569_, _03570_, _03571_, _03572_, _03573_, _03574_, _03575_, _03576_, _03577_, _03578_, _03579_, _03580_, _03581_, _03582_, _03583_, _03584_, _03585_, _03586_, _03587_, _03588_, _03589_, _03590_, _03591_, _03592_, _03593_, _03594_, _03595_, _03596_, _03597_, _03598_, _03599_, _03600_, _03601_, _03602_, _03603_, _03604_, _03605_, _03606_, _03607_, _03608_, _03609_, _03610_, _03611_, _03612_, _03613_, _03614_, _03615_, _03616_, _03617_, _03618_, _03619_, _03620_, _03621_, _03622_, _03623_, _03624_, _03625_, _03626_, _03627_, _03628_, _03629_, _03630_, _03631_, _03632_, _03633_, _03634_, _03635_, _03636_, _03637_, _03638_, _03639_, _03640_, _03641_, _03642_, _03643_, _03644_, _03645_, _03646_, _03647_, _03648_, _03649_, _03650_, _03651_, _03652_, _03653_, _03654_, _03655_, _03656_, _03657_, _03658_, _03659_, _03660_, _03661_, _03662_, _03663_, _03664_, _03665_, _03666_, _03667_, _03668_, _03669_, _03670_, _03671_, _03672_, _03673_, _03674_, _03675_, _03676_, _03677_, _03678_, _03679_, _03680_, _03681_, _03682_, _03683_, _03684_, _03685_, _03686_, _03687_, _03688_, _03689_, _03690_, _03691_, _03692_, _03693_, _03694_, _03695_, _03696_, _03697_, _03698_, _03699_, _03700_, _03701_, _03702_, _03703_, _03704_, _03705_, _03706_, _03707_, _03708_, _03709_, _03710_, _03711_, _03712_, _03713_, _03714_, _03715_, _03716_, _03717_, _03718_, _03719_, _03720_, _03721_, _03722_, _03723_, _03724_, _03725_, _03726_, _03727_, _03728_, _03729_, _03730_, _03731_, _03732_, _03733_, _03734_, _03735_, _03736_, _03737_, _03738_, _03739_, _03740_, _03741_, _03742_, _03743_, _03744_, _03745_, _03746_, _03747_, _03748_, _03749_, _03750_, _03751_, _03752_, _03753_, _03754_, _03755_, _03756_, _03757_, _03758_, _03759_, _03760_, _03761_, _03762_, _03763_, _03764_, _03765_, _03766_, _03767_, _03768_, _03769_, _03770_, _03771_, _03772_, _03773_, _03774_, _03775_, _03776_, _03777_, _03778_, _03779_, _03780_, _03781_, _03782_, _03783_, _03784_, _03785_, _03786_, _03787_, _03788_, _03789_, _03790_, _03791_, _03792_, _03793_, _03794_, _03795_, _03796_, _03797_, _03798_, _03799_, _03800_, _03801_, _03802_, _03803_, _03804_, _03805_, _03806_, _03807_, _03808_, _03809_, _03810_, _03811_, _03812_, _03813_, _03814_, _03815_, _03816_, _03817_, _03818_, _03819_, _03820_, _03821_, _03822_, _03823_, _03824_, _03825_, _03826_, _03827_, _03828_, _03829_, _03830_, _03831_, _03832_, _03833_, _03834_, _03835_, _03836_, _03837_, _03838_, _03839_, _03840_, _03841_, _03842_, _03843_, _03844_, _03845_, _03846_, _03847_, _03848_, _03849_, _03850_, _03851_, _03852_, _03853_, _03854_, _03855_, _03856_, _03857_, _03858_, _03859_, _03860_, _03861_, _03862_, _03863_, _03864_, _03865_, _03866_, _03867_, _03868_, _03869_, _03870_, _03871_, _03872_, _03873_, _03874_, _03875_, _03876_, _03877_, _03878_, _03879_, _03880_, _03881_, _03882_, _03883_, _03884_, _03885_, _03886_, _03887_, _03888_, _03889_, _03890_, _03891_, _03892_, _03893_, _03894_, _03895_, _03896_, _03897_, _03898_, _03899_, _03900_, _03901_, _03902_, _03903_, _03904_, _03905_, _03906_, _03907_, _03908_, _03909_, _03910_, _03911_, _03912_, _03913_, _03914_, _03915_, _03916_, _03917_, _03918_, _03919_, _03920_, _03921_, _03922_, _03923_, _03924_, _03925_, _03926_, _03927_, _03928_, _03929_, _03930_, _03931_, _03932_, _03933_, _03934_, _03935_, _03936_, _03937_, _03938_, _03939_, _03940_, _03941_, _03942_, _03943_, _03944_, _03945_, _03946_, _03947_, _03948_, _03949_, _03950_, _03951_, _03952_, _03953_, _03954_, _03955_, _03956_, _03957_, _03958_, _03959_, _03960_, _03961_, _03962_, _03963_, _03964_, _03965_, _03966_, _03967_, _03968_, _03969_, _03970_, _03971_, _03972_, _03973_, _03974_, _03975_, _03976_, _03977_, _03978_, _03979_, _03980_, _03981_, _03982_, _03983_, _03984_, _03985_, _03986_, _03987_, _03988_, _03989_, _03990_, _03991_, _03992_, _03993_, _03994_, _03995_, _03996_, _03997_, _03998_, _03999_, _04000_, _04001_, _04002_, _04003_, _04004_, _04005_, _04006_, _04007_, _04008_, _04009_, _04010_, _04011_, _04012_, _04013_, _04014_, _04015_, _04016_, _04017_, _04018_, _04019_, _04020_, _04021_, _04022_, _04023_, _04024_, _04025_, _04026_, _04027_, _04028_, _04029_, _04030_, _04031_, _04032_, _04033_, _04034_, _04035_, _04036_, _04037_, _04038_, _04039_, _04040_, _04041_, _04042_, _04043_, _04044_, _04045_, _04046_, _04047_, _04048_, _04049_, _04050_, _04051_, _04052_, _04053_, _04054_, _04055_, _04056_, _04057_, _04058_, _04059_, _04060_, _04061_, _04062_, _04063_, _04064_, _04065_, _04066_, _04067_, _04068_, _04069_, _04070_, _04071_, _04072_, _04073_, _04074_, _04075_, _04076_, _04077_, _04078_, _04079_, _04080_, _04081_, _04082_, _04083_, _04084_, _04085_, _04086_, _04087_, _04088_, _04089_, _04090_, _04091_, _04092_, _04093_, _04094_, _04095_, _04096_, _04097_, _04098_, _04099_, _04100_, _04101_, _04102_, _04103_, _04104_, _04105_, _04106_, _04107_, _04108_, _04109_, _04110_, _04111_, _04112_, _04113_, _04114_, _04115_, _04116_, _04117_, _04118_, _04119_, _04120_, _04121_, _04122_, _04123_, _04124_, _04125_, _04126_, _04127_, _04128_, _04129_, _04130_, _04131_, _04132_, _04133_, _04134_, _04135_, _04136_, _04137_, _04138_, _04139_, _04140_, _04141_, _04142_, _04143_, _04144_, _04145_, _04146_, _04147_, _04148_, _04149_, _04150_, _04151_, _04152_, _04153_, _04154_, _04155_, _04156_, _04157_, _04158_, _04159_, _04160_, _04161_, _04162_, _04163_, _04164_, _04165_, _04166_, _04167_, _04168_, _04169_, _04170_, _04171_, _04172_, _04173_, _04174_, _04175_, _04176_, _04177_, _04178_, _04179_, _04180_, _04181_, _04182_, _04183_, _04184_, _04185_, _04186_, _04187_, _04188_, _04189_, _04190_, _04191_, _04192_, _04193_, _04194_, _04195_, _04196_, _04197_, _04198_, _04199_, _04200_, _04201_, _04202_, _04203_, _04204_, _04205_, _04206_, _04207_, _04208_, _04209_, _04210_, _04211_, _04212_, _04213_, _04214_, _04215_, _04216_, _04217_, _04218_, _04219_, _04220_, _04221_, _04222_, _04223_, _04224_, _04225_, _04226_, _04227_, _04228_, _04229_, _04230_, _04231_, _04232_, _04233_, _04234_, _04235_, _04236_, _04237_, _04238_, _04239_, _04240_, _04241_, _04242_, _04243_, _04244_, _04245_, _04246_, _04247_, _04248_, _04249_, _04250_, _04251_, _04252_, _04253_, _04254_, _04255_, _04256_, _04257_, _04258_, _04259_, _04260_, _04261_, _04262_, _04263_, _04264_, _04265_, _04266_, _04267_, _04268_, _04269_, _04270_, _04271_, _04272_, _04273_, _04274_, _04275_, _04276_, _04277_, _04278_, _04279_, _04280_, _04281_, _04282_, _04283_, _04284_, _04285_, _04286_, _04287_, _04288_, _04289_, _04290_, _04291_, _04292_, _04293_, _04294_, _04295_, _04296_, _04297_, _04298_, _04299_, _04300_, _04301_, _04302_, _04303_, _04304_, _04305_, _04306_, _04307_, _04308_, _04309_, _04310_, _04311_, _04312_, _04313_, _04314_, _04315_, _04316_, _04317_, _04318_, _04319_, _04320_, _04321_, _04322_, _04323_, _04324_, _04325_, _04326_, _04327_, _04328_, _04329_, _04330_, _04331_, _04332_, _04333_, _04334_, _04335_, _04336_, _04337_, _04338_, _04339_, _04340_, _04341_, _04342_, _04343_, _04344_, _04345_, _04346_, _04347_, _04348_, _04349_, _04350_, _04351_, _04352_, _04353_, _04354_, _04355_, _04356_, _04357_, _04358_, _04359_, _04360_, _04361_, _04362_, _04363_, _04364_, _04365_, _04366_, _04367_, _04368_, _04369_, _04370_, _04371_, _04372_, _04373_, _04374_, _04375_, _04376_, _04377_, _04378_, _04379_, _04380_, _04381_, _04382_, _04383_, _04384_, _04385_, _04386_, _04387_, _04388_, _04389_, _04390_, _04391_, _04392_, _04393_, _04394_, _04395_, _04396_, _04397_, _04398_, _04399_, _04400_, _04401_, _04402_, _04403_, _04404_, _04405_, _04406_, _04407_, _04408_, _04409_, _04410_, _04411_, _04412_, _04413_, _04414_, _04415_, _04416_, _04417_, _04418_, _04419_, _04420_, _04421_, _04422_, _04423_, _04424_, _04425_, _04426_, _04427_, _04428_, _04429_, _04430_, _04431_, _04432_, _04433_, _04434_, _04435_, _04436_, _04437_, _04438_, _04439_, _04440_, _04441_, _04442_, _04443_, _04444_, _04445_, _04446_, _04447_, _04448_, _04449_, _04450_, _04451_, _04452_, _04453_, _04454_, _04455_, _04456_, _04457_, _04458_, _04459_, _04460_, _04461_, _04462_, _04463_, _04464_, _04465_, _04466_, _04467_, _04468_, _04469_, _04470_, _04471_, _04472_, _04473_, _04474_, _04475_, _04476_, _04477_, _04478_, _04479_, _04480_, _04481_, _04482_, _04483_, _04484_, _04485_, _04486_, _04487_, _04488_, _04489_, _04490_, _04491_, _04492_, _04493_, _04494_, _04495_, _04496_, _04497_, _04498_, _04499_, _04500_, _04501_, _04502_, _04503_, _04504_, _04505_, _04506_, _04507_, _04508_, _04509_, _04510_, _04511_, _04512_, _04513_, _04514_, _04515_, _04516_, _04517_, _04518_, _04519_, _04520_, _04521_, _04522_, _04523_, _04524_, _04525_, _04526_, _04527_, _04528_, _04529_, _04530_, _04531_, _04532_, _04533_, _04534_, _04535_, _04536_, _04537_, _04538_, _04539_, _04540_, _04541_, _04542_, _04543_, _04544_, _04545_, _04546_, _04547_, _04548_, _04549_, _04550_, _04551_, _04552_, _04553_, _04554_, _04555_, _04556_, _04557_, _04558_, _04559_, _04560_, _04561_, _04562_, _04563_, _04564_, _04565_, _04566_, _04567_, _04568_, _04569_, _04570_, _04571_, _04572_, _04573_, _04574_, _04575_, _04576_, _04577_, _04578_, _04579_, _04580_, _04581_, _04582_, _04583_, _04584_, _04585_, _04586_, _04587_, _04588_, _04589_, _04590_, _04591_, _04592_, _04593_, _04594_, _04595_, _04596_, _04597_, _04598_, _04599_, _04600_, _04601_, _04602_, _04603_, _04604_, _04605_, _04606_, _04607_, _04608_, _04609_, _04610_, _04611_, _04612_, _04613_, _04614_, _04615_, _04616_, _04617_, _04618_, _04619_, _04620_, _04621_, _04622_, _04623_, _04624_, _04625_, _04626_, _04627_, _04628_, _04629_, _04630_, _04631_, _04632_, _04633_, _04634_, _04635_, _04636_, _04637_, _04638_, _04639_, _04640_, _04641_, _04642_, _04643_, _04644_, _04645_, _04646_, _04647_, _04648_, _04649_, _04650_, _04651_, _04652_, _04653_, _04654_, _04655_, _04656_, _04657_, _04658_, _04659_, _04660_, _04661_, _04662_, _04663_, _04664_, _04665_, _04666_, _04667_, _04668_, _04669_, _04670_, _04671_, _04672_, _04673_, _04674_, _04675_, _04676_, _04677_, _04678_, _04679_, _04680_, _04681_, _04682_, _04683_, _04684_, _04685_, _04686_, _04687_, _04688_, _04689_, _04690_, _04691_, _04692_, _04693_, _04694_, _04695_, _04696_, _04697_, _04698_, _04699_, _04700_, _04701_, _04702_, _04703_, _04704_, _04705_, _04706_, _04707_, _04708_, _04709_, _04710_, _04711_, _04712_, _04713_, _04714_, _04715_, _04716_, _04717_, _04718_, _04719_, _04720_, _04721_, _04722_, _04723_, _04724_, _04725_, _04726_, _04727_, _04728_, _04729_, _04730_, _04731_, _04732_, _04733_, _04734_, _04735_, _04736_, _04737_, _04738_, _04739_, _04740_, _04741_, _04742_, _04743_, _04744_, _04745_, _04746_, _04747_, _04748_, _04749_, _04750_, _04751_, _04752_, _04753_, _04754_, _04755_, _04756_, _04757_, _04758_, _04759_, _04760_, _04761_, _04762_, _04763_, _04764_, _04765_, _04766_, _04767_, _04768_, _04769_, _04770_, _04771_, _04772_, _04773_, _04774_, _04775_, _04776_, _04777_, _04778_, _04779_, _04780_, _04781_, _04782_, _04783_, _04784_, _04785_, _04786_, _04787_, _04788_, _04789_, _04790_, _04791_, _04792_, _04793_, _04794_, _04795_, _04796_, _04797_, _04798_, _04799_, _04800_, _04801_, _04802_, _04803_, _04804_, _04805_, _04806_, _04807_, _04808_, _04809_, _04810_, _04811_, _04812_, _04813_, _04814_, _04815_, _04816_, _04817_, _04818_, _04819_, _04820_, _04821_, _04822_, _04823_, _04824_, _04825_, _04826_, _04827_, _04828_, _04829_, _04830_, _04831_, _04832_, _04833_, _04834_, _04835_, _04836_, _04837_, _04838_, _04839_, _04840_, _04841_, _04842_, _04843_, _04844_, _04845_, _04846_, _04847_, _04848_, _04849_, _04850_, _04851_, _04852_, _04853_, _04854_, _04855_, _04856_, _04857_, _04858_, _04859_, _04860_, _04861_, _04862_, _04863_, _04864_, _04865_, _04866_, _04867_, _04868_, _04869_, _04870_, _04871_, _04872_, _04873_, _04874_, _04875_, _04876_, _04877_, _04878_, _04879_, _04880_, _04881_, _04882_, _04883_, _04884_, _04885_, _04886_, _04887_, _04888_, _04889_, _04890_, _04891_, _04892_, _04893_, _04894_, _04895_, _04896_, _04897_, _04898_, _04899_, _04900_, _04901_, _04902_, _04903_, _04904_, _04905_, _04906_, _04907_, _04908_, _04909_, _04910_, _04911_, _04912_, _04913_, _04914_, _04915_, _04916_, _04917_, _04918_, _04919_, _04920_, _04921_, _04922_, _04923_, _04924_, _04925_, _04926_, _04927_, _04928_, _04929_, _04930_, _04931_, _04932_, _04933_, _04934_, _04935_, _04936_, _04937_, _04938_, _04939_, _04940_, _04941_, _04942_, _04943_, _04944_, _04945_, _04946_, _04947_, _04948_, _04949_, _04950_, _04951_, _04952_, _04953_, _04954_, _04955_, _04956_, _04957_, _04958_, _04959_, _04960_, _04961_, _04962_, _04963_, _04964_, _04965_, _04966_, _04967_, _04968_, _04969_, _04970_, _04971_, _04972_, _04973_, _04974_, _04975_, _04976_, _04977_, _04978_, _04979_, _04980_, _04981_, _04982_, _04983_, _04984_, _04985_, _04986_, _04987_, _04988_, _04989_, _04990_, _04991_, _04992_, _04993_, _04994_, _04995_, _04996_, _04997_, _04998_, _04999_, _05000_, _05001_, _05002_, _05003_, _05004_, _05005_, _05006_, _05007_, _05008_, _05009_, _05010_, _05011_, _05012_, _05013_, _05014_, _05015_, _05016_, _05017_, _05018_, _05019_, _05020_, _05021_, _05022_, _05023_, _05024_, _05025_, _05026_, _05027_, _05028_, _05029_, _05030_, _05031_, _05032_, _05033_, _05034_, _05035_, _05036_, _05037_, _05038_, _05039_, _05040_, _05041_, _05042_, _05043_, _05044_, _05045_, _05046_, _05047_, _05048_, _05049_, _05050_, _05051_, _05052_, _05053_, _05054_, _05055_, _05056_, _05057_, _05058_, _05059_, _05060_, _05061_, _05062_, _05063_, _05064_, _05065_, _05066_, _05067_, _05068_, _05069_, _05070_, _05071_, _05072_, _05073_, _05074_, _05075_, _05076_, _05077_, _05078_, _05079_, _05080_, _05081_, _05082_, _05083_, _05084_, _05085_, _05086_, _05087_, _05088_, _05089_, _05090_, _05091_, _05092_, _05093_, _05094_, _05095_, _05096_, _05097_, _05098_, _05099_, _05100_, _05101_, _05102_, _05103_, _05104_, _05105_, _05106_, _05107_, _05108_, _05109_, _05110_, _05111_, _05112_, _05113_, _05114_, _05115_, _05116_, _05117_, _05118_, _05119_, _05120_, _05121_, _05122_, _05123_, _05124_, _05125_, _05126_, _05127_, _05128_, _05129_, _05130_, _05131_, _05132_, _05133_, _05134_, _05135_, _05136_, _05137_, _05138_, _05139_, _05140_, _05141_, _05142_, _05143_, _05144_, _05145_, _05146_, _05147_, _05148_, _05149_, _05150_, _05151_, _05152_, _05153_, _05154_, _05155_, _05156_, _05157_, _05158_, _05159_, _05160_, _05161_, _05162_, _05163_, _05164_, _05165_, _05166_, _05167_, _05168_, _05169_, _05170_, _05171_, _05172_, _05173_, _05174_, _05175_, _05176_, _05177_, _05178_, _05179_, _05180_, _05181_, _05182_, _05183_, _05184_, _05185_, _05186_, _05187_, _05188_, _05189_, _05190_, _05191_, _05192_, _05193_, _05194_, _05195_, _05196_, _05197_, _05198_, _05199_, _05200_, _05201_, _05202_, _05203_, _05204_, _05205_, _05206_, _05207_, _05208_, _05209_, _05210_, _05211_, _05212_, _05213_, _05214_, _05215_, _05216_, _05217_, _05218_, _05219_, _05220_, _05221_, _05222_, _05223_, _05224_, _05225_, _05226_, _05227_, _05228_, _05229_, _05230_, _05231_, _05232_, _05233_, _05234_, _05235_, _05236_, _05237_, _05238_, _05239_, _05240_, _05241_, _05242_, _05243_, _05244_, _05245_, _05246_, _05247_, _05248_, _05249_, _05250_, _05251_, _05252_, _05253_, _05254_, _05255_, _05256_, _05257_, _05258_, _05259_, _05260_, _05261_, _05262_, _05263_, _05264_, _05265_, _05266_, _05267_, _05268_, _05269_, _05270_, _05271_, _05272_, _05273_, _05274_, _05275_, _05276_, _05277_, _05278_, _05279_, _05280_, _05281_, _05282_, _05283_, _05284_, _05285_, _05286_, _05287_, _05288_, _05289_, _05290_, _05291_, _05292_, _05293_, _05294_, _05295_, _05296_, _05297_, _05298_, _05299_, _05300_, _05301_, _05302_, _05303_, _05304_, _05305_, _05306_, _05307_, _05308_, _05309_, _05310_, _05311_, _05312_, _05313_, _05314_, _05315_, _05316_, _05317_, _05318_, _05319_, _05320_, _05321_, _05322_, _05323_, _05324_, _05325_, _05326_, _05327_, _05328_, _05329_, _05330_, _05331_, _05332_, _05333_, _05334_, _05335_, _05336_, _05337_, _05338_, _05339_, _05340_, _05341_, _05342_, _05343_, _05344_, _05345_, _05346_, _05347_, _05348_, _05349_, _05350_, _05351_, _05352_, _05353_, _05354_, _05355_, _05356_, _05357_, _05358_, _05359_, _05360_, _05361_, _05362_, _05363_, _05364_, _05365_, _05366_, _05367_, _05368_, _05369_, _05370_, _05371_, _05372_, _05373_, _05374_, _05375_, _05376_, _05377_, _05378_, _05379_, _05380_, _05381_, _05382_, _05383_, _05384_, _05385_, _05386_, _05387_, _05388_, _05389_, _05390_, _05391_, _05392_, _05393_, _05394_, _05395_, _05396_, _05397_, _05398_, _05399_, _05400_, _05401_, _05402_, _05403_, _05404_, _05405_, _05406_, _05407_, _05408_, _05409_, _05410_, _05411_, _05412_, _05413_, _05414_, _05415_, _05416_, _05417_, _05418_, _05419_, _05420_, _05421_, _05422_, _05423_, _05424_, _05425_, _05426_, _05427_, _05428_, _05429_, _05430_, _05431_, _05432_, _05433_, _05434_, _05435_, _05436_, _05437_, _05438_, _05439_, _05440_, _05441_, _05442_, _05443_, _05444_, _05445_, _05446_, _05447_, _05448_, _05449_, _05450_, _05451_, _05452_, _05453_, _05454_, _05455_, _05456_, _05457_, _05458_, _05459_, _05460_, _05461_, _05462_, _05463_, _05464_, _05465_, _05466_, _05467_, _05468_, _05469_, _05470_, _05471_, _05472_, _05473_, _05474_, _05475_, _05476_, _05477_, _05478_, _05479_, _05480_, _05481_, _05482_, _05483_, _05484_, _05485_, _05486_, _05487_, _05488_, _05489_, _05490_, _05491_, _05492_, _05493_, _05494_, _05495_, _05496_, _05497_, _05498_, _05499_, _05500_, _05501_, _05502_, _05503_, _05504_, _05505_, _05506_, _05507_, _05508_, _05509_, _05510_, _05511_, _05512_, _05513_, _05514_, _05515_, _05516_, _05517_, _05518_, _05519_, _05520_, _05521_, _05522_, _05523_, _05524_, _05525_, _05526_, _05527_, _05528_, _05529_, _05530_, _05531_, _05532_, _05533_, _05534_, _05535_, _05536_, _05537_, _05538_, _05539_, _05540_, _05541_, _05542_, _05543_, _05544_, _05545_, _05546_, _05547_, _05548_, _05549_, _05550_, _05551_, _05552_, _05553_, _05554_, _05555_, _05556_, _05557_, _05558_, _05559_, _05560_, _05561_, _05562_, _05563_, _05564_, _05565_, _05566_, _05567_, _05568_, _05569_, _05570_, _05571_, _05572_, _05573_, _05574_, _05575_, _05576_, _05577_, _05578_, _05579_, _05580_, _05581_, _05582_, _05583_, _05584_, _05585_, _05586_, _05587_, _05588_, _05589_, _05590_, _05591_, _05592_, _05593_, _05594_, _05595_, _05596_, _05597_, _05598_, _05599_, _05600_, _05601_, _05602_, _05603_, _05604_, _05605_, _05606_, _05607_, _05608_, _05609_, _05610_, _05611_, _05612_, _05613_, _05614_, _05615_, _05616_, _05617_, _05618_, _05619_, _05620_, _05621_, _05622_, _05623_, _05624_, _05625_, _05626_, _05627_, _05628_, _05629_, _05630_, _05631_, _05632_, _05633_, _05634_, _05635_, _05636_, _05637_, _05638_, _05639_, _05640_, _05641_, _05642_, _05643_, _05644_, _05645_, _05646_, _05647_, _05648_, _05649_, _05650_, _05651_, _05652_, _05653_, _05654_, _05655_, _05656_, _05657_, _05658_, _05659_, _05660_, _05661_, _05662_, _05663_, _05664_, _05665_, _05666_, _05667_, _05668_, _05669_, _05670_, _05671_, _05672_, _05673_, _05674_, _05675_, _05676_, _05677_, _05678_, _05679_, _05680_, _05681_, _05682_, _05683_, _05684_, _05685_, _05686_, _05687_, _05688_, _05689_, _05690_, _05691_, _05692_, _05693_, _05694_, _05695_, _05696_, _05697_, _05698_, _05699_, _05700_, _05701_, _05702_, _05703_, _05704_, _05705_, _05706_, _05707_, _05708_, _05709_, _05710_, _05711_, _05712_, _05713_, _05714_, _05715_, _05716_, _05717_, _05718_, _05719_, _05720_, _05721_, _05722_, _05723_, _05724_, _05725_, _05726_, _05727_, _05728_, _05729_, _05730_, _05731_, _05732_, _05733_, _05734_, _05735_, _05736_, _05737_, _05738_, _05739_, _05740_, _05741_, _05742_, _05743_, _05744_, _05745_, _05746_, _05747_, _05748_, _05749_, _05750_, _05751_, _05752_, _05753_, _05754_, _05755_, _05756_, _05757_, _05758_, _05759_, _05760_, _05761_, _05762_, _05763_, _05764_, _05765_, _05766_, _05767_, _05768_, _05769_, _05770_, _05771_, _05772_, _05773_, _05774_, _05775_, _05776_, _05777_, _05778_, _05779_, _05780_, _05781_, _05782_, _05783_, _05784_, _05785_, _05786_, _05787_, _05788_, _05789_, _05790_, _05791_, _05792_, _05793_, _05794_, _05795_, _05796_, _05797_, _05798_, _05799_, _05800_, _05801_, _05802_, _05803_, _05804_, _05805_, _05806_, _05807_, _05808_, _05809_, _05810_, _05811_, _05812_, _05813_, _05814_, _05815_, _05816_, _05817_, _05818_, _05819_, _05820_, _05821_, _05822_, _05823_, _05824_, _05825_, _05826_, _05827_, _05828_, _05829_, _05830_, _05831_, _05832_, _05833_, _05834_, _05835_, _05836_, _05837_, _05838_, _05839_, _05840_, _05841_, _05842_, _05843_, _05844_, _05845_, _05846_, _05847_, _05848_, _05849_, _05850_, _05851_, _05852_, _05853_, _05854_, _05855_, _05856_, _05857_, _05858_, _05859_, _05860_, _05861_, _05862_, _05863_, _05864_, _05865_, _05866_, _05867_, _05868_, _05869_, _05870_, _05871_, _05872_, _05873_, _05874_, _05875_, _05876_, _05877_, _05878_, _05879_, _05880_, _05881_, _05882_, _05883_, _05884_, _05885_, _05886_, _05887_, _05888_, _05889_, _05890_, _05891_, _05892_, _05893_, _05894_, _05895_, _05896_, _05897_, _05898_, _05899_, _05900_, _05901_, _05902_, _05903_, _05904_, _05905_, _05906_, _05907_, _05908_, _05909_, _05910_, _05911_, _05912_, _05913_, _05914_, _05915_, _05916_, _05917_, _05918_, _05919_, _05920_, _05921_, _05922_, _05923_, _05924_, _05925_, _05926_, _05927_, _05928_, _05929_, _05930_, _05931_, _05932_, _05933_, _05934_, _05935_, _05936_, _05937_, _05938_, _05939_, _05940_, _05941_, _05942_, _05943_, _05944_, _05945_, _05946_, _05947_, _05948_, _05949_, _05950_, _05951_, _05952_, _05953_, _05954_, _05955_, _05956_, _05957_, _05958_, _05959_, _05960_, _05961_, _05962_, _05963_, _05964_, _05965_, _05966_, _05967_, _05968_, _05969_, _05970_, _05971_, _05972_, _05973_, _05974_, _05975_, _05976_, _05977_, _05978_, _05979_, _05980_, _05981_, _05982_, _05983_, _05984_, _05985_, _05986_, _05987_, _05988_, _05989_, _05990_, _05991_, _05992_, _05993_, _05994_, _05995_, _05996_, _05997_, _05998_, _05999_, _06000_, _06001_, _06002_, _06003_, _06004_, _06005_, _06006_, _06007_, _06008_, _06009_, _06010_, _06011_, _06012_, _06013_, _06014_, _06015_, _06016_, _06017_, _06018_, _06019_, _06020_, _06021_, _06022_, _06023_, _06024_, _06025_, _06026_, _06027_, _06028_, _06029_, _06030_, _06031_, _06032_, _06033_, _06034_, _06035_, _06036_, _06037_, _06038_, _06039_, _06040_, _06041_, _06042_, _06043_, _06044_, _06045_, _06046_, _06047_, _06048_, _06049_, _06050_, _06051_, _06052_, _06053_, _06054_, _06055_, _06056_, _06057_, _06058_, _06059_, _06060_, _06061_, _06062_, _06063_, _06064_, _06065_, _06066_, _06067_, _06068_, _06069_, _06070_, _06071_, _06072_, _06073_, _06074_, _06075_, _06076_, _06077_, _06078_, _06079_, _06080_, _06081_, _06082_, _06083_, _06084_, _06085_, _06086_, _06087_, _06088_, _06089_, _06090_, _06091_, _06092_, _06093_, _06094_, _06095_, _06096_, _06097_, _06098_, _06099_, _06100_, _06101_, _06102_, _06103_, _06104_, _06105_, _06106_, _06107_, _06108_, _06109_, _06110_, _06111_, _06112_, _06113_, _06114_, _06115_, _06116_, _06117_, _06118_, _06119_, _06120_, _06121_, _06122_, _06123_, _06124_, _06125_, _06126_, _06127_, _06128_, _06129_, _06130_, _06131_, _06132_, _06133_, _06134_, _06135_, _06136_, _06137_, _06138_, _06139_, _06140_, _06141_, _06142_, _06143_, _06144_, _06145_, _06146_, _06147_, _06148_, _06149_, _06150_, _06151_, _06152_, _06153_, _06154_, _06155_, _06156_, _06157_, _06158_, _06159_, _06160_, _06161_, _06162_, _06163_, _06164_, _06165_, _06166_, _06167_, _06168_, _06169_, _06170_, _06171_, _06172_, _06173_, _06174_, _06175_, _06176_, _06177_, _06178_, _06179_, _06180_, _06181_, _06182_, _06183_, _06184_, _06185_, _06186_, _06187_, _06188_, _06189_, _06190_, _06191_, _06192_, _06193_, _06194_, _06195_, _06196_, _06197_, _06198_, _06199_, _06200_, _06201_, _06202_, _06203_, _06204_, _06205_, _06206_, _06207_, _06208_, _06209_, _06210_, _06211_, _06212_, _06213_, _06214_, _06215_, _06216_, _06217_, _06218_, _06219_, _06220_, _06221_, _06222_, _06223_, _06224_, _06225_, _06226_, _06227_, _06228_, _06229_, _06230_, _06231_, _06232_, _06233_, _06234_, _06235_, _06236_, _06237_, _06238_, _06239_, _06240_, _06241_, _06242_, _06243_, _06244_, _06245_, _06246_, _06247_, _06248_, _06249_, _06250_, _06251_, _06252_, _06253_, _06254_, _06255_, _06256_, _06257_, _06258_, _06259_, _06260_, _06261_, _06262_, _06263_, _06264_, _06265_, _06266_, _06267_, _06268_, _06269_, _06270_, _06271_, _06272_, _06273_, _06274_, _06275_, _06276_, _06277_, _06278_, _06279_, _06280_, _06281_, _06282_, _06283_, _06284_, _06285_, _06286_, _06287_, _06288_, _06289_, _06290_, _06291_, _06292_, _06293_, _06294_, _06295_, _06296_, _06297_, _06298_, _06299_, _06300_, _06301_, _06302_, _06303_, _06304_, _06305_, _06306_, _06307_, _06308_, _06309_, _06310_, _06311_, _06312_, _06313_, _06314_, _06315_, _06316_, _06317_, _06318_, _06319_, _06320_, _06321_, _06322_, _06323_, _06324_, _06325_, _06326_, _06327_, _06328_, _06329_, _06330_, _06331_, _06332_, _06333_, _06334_, _06335_, _06336_, _06337_, _06338_, _06339_, _06340_, _06341_, _06342_, _06343_, _06344_, _06345_, _06346_, _06347_, _06348_, _06349_, _06350_, _06351_, _06352_, _06353_, _06354_, _06355_, _06356_, _06357_, _06358_, _06359_, _06360_, _06361_, _06362_, _06363_, _06364_, _06365_, _06366_, _06367_, _06368_, _06369_, _06370_, _06371_, _06372_, _06373_, _06374_, _06375_, _06376_, _06377_, _06378_, _06379_, _06380_, _06381_, _06382_, _06383_, _06384_, _06385_, _06386_, _06387_, _06388_, _06389_, _06390_, _06391_, _06392_, _06393_, _06394_, _06395_, _06396_, _06397_, _06398_, _06399_, _06400_, _06401_, _06402_, _06403_, _06404_, _06405_, _06406_, _06407_, _06408_, _06409_, _06410_, _06411_, _06412_, _06413_, _06414_, _06415_, _06416_, _06417_, _06418_, _06419_, _06420_, _06421_, _06422_, _06423_, _06424_, _06425_, _06426_, _06427_, _06428_, _06429_, _06430_, _06431_, _06432_, _06433_, _06434_, _06435_, _06436_, _06437_, _06438_, _06439_, _06440_, _06441_, _06442_, _06443_, _06444_, _06445_, _06446_, _06447_, _06448_, _06449_, _06450_, _06451_, _06452_, _06453_, _06454_, _06455_, _06456_, _06457_, _06458_, _06459_, _06460_, _06461_, _06462_, _06463_, _06464_, _06465_, _06466_, _06467_, _06468_, _06469_, _06470_, _06471_, _06472_, _06473_, _06474_, _06475_, _06476_, _06477_, _06478_, _06479_, _06480_, _06481_, _06482_, _06483_, _06484_, _06485_, _06486_, _06487_, _06488_, _06489_, _06490_, _06491_, _06492_, _06493_, _06494_, _06495_, _06496_, _06497_, _06498_, _06499_, _06500_, _06501_, _06502_, _06503_, _06504_, _06505_, _06506_, _06507_, _06508_, _06509_, _06510_, _06511_, _06512_, _06513_, _06514_, _06515_, _06516_, _06517_, _06518_, _06519_, _06520_, _06521_, _06522_, _06523_, _06524_, _06525_, _06526_, _06527_, _06528_, _06529_, _06530_, _06531_, _06532_, _06533_, _06534_, _06535_, _06536_, _06537_, _06538_, _06539_, _06540_, _06541_, _06542_, _06543_, _06544_, _06545_, _06546_, _06547_, _06548_, _06549_, _06550_, _06551_, _06552_, _06553_, _06554_, _06555_, _06556_, _06557_, _06558_, _06559_, _06560_, _06561_, _06562_, _06563_, _06564_, _06565_, _06566_, _06567_, _06568_, _06569_, _06570_, _06571_, _06572_, _06573_, _06574_, _06575_, _06576_, _06577_, _06578_, _06579_, _06580_, _06581_, _06582_, _06583_, _06584_, _06585_, _06586_, _06587_, _06588_, _06589_, _06590_, _06591_, _06592_, _06593_, _06594_, _06595_, _06596_, _06597_, _06598_, _06599_, _06600_, _06601_, _06602_, _06603_, _06604_, _06605_, _06606_, _06607_, _06608_, _06609_, _06610_, _06611_, _06612_, _06613_, _06614_, _06615_, _06616_, _06617_, _06618_, _06619_, _06620_, _06621_, _06622_, _06623_, _06624_, _06625_, _06626_, _06627_, _06628_, _06629_, _06630_, _06631_, _06632_, _06633_, _06634_, _06635_, _06636_, _06637_, _06638_, _06639_, _06640_, _06641_, _06642_, _06643_, _06644_, _06645_, _06646_, _06647_, _06648_, _06649_, _06650_, _06651_, _06652_, _06653_, _06654_, _06655_, _06656_, _06657_, _06658_, _06659_, _06660_, _06661_, _06662_, _06663_, _06664_, _06665_, _06666_, _06667_, _06668_, _06669_, _06670_, _06671_, _06672_, _06673_, _06674_, _06675_, _06676_, _06677_, _06678_, _06679_, _06680_, _06681_, _06682_, _06683_, _06684_, _06685_, _06686_, _06687_, _06688_, _06689_, _06690_, _06691_, _06692_, _06693_, _06694_, _06695_, _06696_, _06697_, _06698_, _06699_, _06700_, _06701_, _06702_, _06703_, _06704_, _06705_, _06706_, _06707_, _06708_, _06709_, _06710_, _06711_, _06712_, _06713_, _06714_, _06715_, _06716_, _06717_, _06718_, _06719_, _06720_, _06721_, _06722_, _06723_, _06724_, _06725_, _06726_, _06727_, _06728_, _06729_, _06730_, _06731_, _06732_, _06733_, _06734_, _06735_, _06736_, _06737_, _06738_, _06739_, _06740_, _06741_, _06742_, _06743_, _06744_, _06745_, _06746_, _06747_, _06748_, _06749_, _06750_, _06751_, _06752_, _06753_, _06754_, _06755_, _06756_, _06757_, _06758_, _06759_, _06760_, _06761_, _06762_, _06763_, _06764_, _06765_, _06766_, _06767_, _06768_, _06769_, _06770_, _06771_, _06772_, _06773_, _06774_, _06775_, _06776_, _06777_, _06778_, _06779_, _06780_, _06781_, _06782_, _06783_, _06784_, _06785_, _06786_, _06787_, _06788_, _06789_, _06790_, _06791_, _06792_, _06793_, _06794_, _06795_, _06796_, _06797_, _06798_, _06799_, _06800_, _06801_, _06802_, _06803_, _06804_, _06805_, _06806_, _06807_, _06808_, _06809_, _06810_, _06811_, _06812_, _06813_, _06814_, _06815_, _06816_, _06817_, _06818_, _06819_, _06820_, _06821_, _06822_, _06823_, _06824_, _06825_, _06826_, _06827_, _06828_, _06829_, _06830_, _06831_, _06832_, _06833_, _06834_, _06835_, _06836_, _06837_, _06838_, _06839_, _06840_, _06841_, _06842_, _06843_, _06844_, _06845_, _06846_, _06847_, _06848_, _06849_, _06850_, _06851_, _06852_, _06853_, _06854_, _06855_, _06856_, _06857_, _06858_, _06859_, _06860_, _06861_, _06862_, _06863_, _06864_, _06865_, _06866_, _06867_, _06868_, _06869_, _06870_, _06871_, _06872_, _06873_, _06874_, _06875_, _06876_, _06877_, _06878_, _06879_, _06880_, _06881_, _06882_, _06883_, _06884_, _06885_, _06886_, _06887_, _06888_, _06889_, _06890_, _06891_, _06892_, _06893_, _06894_, _06895_, _06896_, _06897_, _06898_, _06899_, _06900_, _06901_, _06902_, _06903_, _06904_, _06905_, _06906_, _06907_, _06908_, _06909_, _06910_, _06911_, _06912_, _06913_, _06914_, _06915_, _06916_, _06917_, _06918_, _06919_, _06920_, _06921_, _06922_, _06923_, _06924_, _06925_, _06926_, _06927_, _06928_, _06929_, _06930_, _06931_, _06932_, _06933_, _06934_, _06935_, _06936_, _06937_, _06938_, _06939_, _06940_, _06941_, _06942_, _06943_, _06944_, _06945_, _06946_, _06947_, _06948_, _06949_, _06950_, _06951_, _06952_, _06953_, _06954_, _06955_, _06956_, _06957_, _06958_, _06959_, _06960_, _06961_, _06962_, _06963_, _06964_, _06965_, _06966_, _06967_, _06968_, _06969_, _06970_, _06971_, _06972_, _06973_, _06974_, _06975_, _06976_, _06977_, _06978_, _06979_, _06980_, _06981_, _06982_, _06983_, _06984_, _06985_, _06986_, _06987_, _06988_, _06989_, _06990_, _06991_, _06992_, _06993_, _06994_, _06995_, _06996_, _06997_, _06998_, _06999_, _07000_, _07001_, _07002_, _07003_, _07004_, _07005_, _07006_, _07007_, _07008_, _07009_, _07010_, _07011_, _07012_, _07013_, _07014_, _07015_, _07016_, _07017_, _07018_, _07019_, _07020_, _07021_, _07022_, _07023_, _07024_, _07025_, _07026_, _07027_, _07028_, _07029_, _07030_, _07031_, _07032_, _07033_, _07034_, _07035_, _07036_, _07037_, _07038_, _07039_, _07040_, _07041_, _07042_, _07043_, _07044_, _07045_, _07046_, _07047_, _07048_, _07049_, _07050_, _07051_, _07052_, _07053_, _07054_, _07055_, _07056_, _07057_, _07058_, _07059_, _07060_, _07061_, _07062_, _07063_, _07064_, _07065_, _07066_, _07067_, _07068_, _07069_, _07070_, _07071_, _07072_, _07073_, _07074_, _07075_, _07076_, _07077_, _07078_, _07079_, _07080_, _07081_, _07082_, _07083_, _07084_, _07085_, _07086_, _07087_, _07088_, _07089_, _07090_, _07091_, _07092_, _07093_, _07094_, _07095_, _07096_, _07097_, _07098_, _07099_, _07100_, _07101_, _07102_, _07103_, _07104_, _07105_, _07106_, _07107_, _07108_, _07109_, _07110_, _07111_, _07112_, _07113_, _07114_, _07115_, _07116_, _07117_, _07118_, _07119_, _07120_, _07121_, _07122_, _07123_, _07124_, _07125_, _07126_, _07127_, _07128_, _07129_, _07130_, _07131_, _07132_, _07133_, _07134_, _07135_, _07136_, _07137_, _07138_, _07139_, _07140_, _07141_, _07142_, _07143_, _07144_, _07145_, _07146_, _07147_, _07148_, _07149_, _07150_, _07151_, _07152_, _07153_, _07154_, _07155_, _07156_, _07157_, _07158_, _07159_, _07160_, _07161_, _07162_, _07163_, _07164_, _07165_, _07166_, _07167_, _07168_, _07169_, _07170_, _07171_, _07172_, _07173_, _07174_, _07175_, _07176_, _07177_, _07178_, _07179_, _07180_, _07181_, _07182_, _07183_, _07184_, _07185_, _07186_, _07187_, _07188_, _07189_, _07190_, _07191_, _07192_, _07193_, _07194_, _07195_, _07196_, _07197_, _07198_, _07199_, _07200_, _07201_, _07202_, _07203_, _07204_, _07205_, _07206_, _07207_, _07208_, _07209_, _07210_, _07211_, _07212_, _07213_, _07214_, _07215_, _07216_, _07217_, _07218_, _07219_, _07220_, _07221_, _07222_, _07223_, _07224_, _07225_, _07226_, _07227_, _07228_, _07229_, _07230_, _07231_, _07232_, _07233_, _07234_, _07235_, _07236_, _07237_, _07238_, _07239_, _07240_, _07241_, _07242_, _07243_, _07244_, _07245_, _07246_, _07247_, _07248_, _07249_, _07250_, _07251_, _07252_, _07253_, _07254_, _07255_, _07256_, _07257_, _07258_, _07259_, _07260_, _07261_, _07262_, _07263_, _07264_, _07265_, _07266_, _07267_, _07268_, _07269_, _07270_, _07271_, _07272_, _07273_, _07274_, _07275_, _07276_, _07277_, _07278_, _07279_, _07280_, _07281_, _07282_, _07283_, _07284_, _07285_, _07286_, _07287_, _07288_, _07289_, _07290_, _07291_, _07292_, _07293_, _07294_, _07295_, _07296_, _07297_, _07298_, _07299_, _07300_, _07301_, _07302_, _07303_, _07304_, _07305_, _07306_, _07307_, _07308_, _07309_, _07310_, _07311_, _07312_, _07313_, _07314_, _07315_, _07316_, _07317_, _07318_, _07319_, _07320_, _07321_, _07322_, _07323_, _07324_, _07325_, _07326_, _07327_, _07328_, _07329_, _07330_, _07331_, _07332_, _07333_, _07334_, _07335_, _07336_, _07337_, _07338_, _07339_, _07340_, _07341_, _07342_, _07343_, _07344_, _07345_, _07346_, _07347_, _07348_, _07349_, _07350_, _07351_, _07352_, _07353_, _07354_, _07355_, _07356_, _07357_, _07358_, _07359_, _07360_, _07361_, _07362_, _07363_, _07364_, _07365_, _07366_, _07367_, _07368_, _07369_, _07370_, _07371_, _07372_, _07373_, _07374_, _07375_, _07376_, _07377_, _07378_, _07379_, _07380_, _07381_, _07382_, _07383_, _07384_, _07385_, _07386_, _07387_, _07388_, _07389_, _07390_, _07391_, _07392_, _07393_, _07394_, _07395_, _07396_, _07397_, _07398_, _07399_, _07400_, _07401_, _07402_, _07403_, _07404_, _07405_, _07406_, _07407_, _07408_, _07409_, _07410_, _07411_, _07412_, _07413_, _07414_, _07415_, _07416_, _07417_, _07418_, _07419_, _07420_, _07421_, _07422_, _07423_, _07424_, _07425_, _07426_, _07427_, _07428_, _07429_, _07430_, _07431_, _07432_, _07433_, _07434_, _07435_, _07436_, _07437_, _07438_, _07439_, _07440_, _07441_, _07442_, _07443_, _07444_, _07445_, _07446_, _07447_, _07448_, _07449_, _07450_, _07451_, _07452_, _07453_, _07454_, _07455_, _07456_, _07457_, _07458_, _07459_, _07460_, _07461_, _07462_, _07463_, _07464_, _07465_, _07466_, _07467_, _07468_, _07469_, _07470_, _07471_, _07472_, _07473_, _07474_, _07475_, _07476_, _07477_, _07478_, _07479_, _07480_, _07481_, _07482_, _07483_, _07484_, _07485_, _07486_, _07487_, _07488_, _07489_, _07490_, _07491_, _07492_, _07493_, _07494_, _07495_, _07496_, _07497_, _07498_, _07499_, _07500_, _07501_, _07502_, _07503_, _07504_, _07505_, _07506_, _07507_, _07508_, _07509_, _07510_, _07511_, _07512_, _07513_, _07514_, _07515_, _07516_, _07517_, _07518_, _07519_, _07520_, _07521_, _07522_, _07523_, _07524_, _07525_, _07526_, _07527_, _07528_, _07529_, _07530_, _07531_, _07532_, _07533_, _07534_, _07535_, _07536_, _07537_, _07538_, _07539_, _07540_, _07541_, _07542_, _07543_, _07544_, _07545_, _07546_, _07547_, _07548_, _07549_, _07550_, _07551_, _07552_, _07553_, _07554_, _07555_, _07556_, _07557_, _07558_, _07559_, _07560_, _07561_, _07562_, _07563_, _07564_, _07565_, _07566_, _07567_, _07568_, _07569_, _07570_, _07571_, _07572_, _07573_, _07574_, _07575_, _07576_, _07577_, _07578_, _07579_, _07580_, _07581_, _07582_, _07583_, _07584_, _07585_, _07586_, _07587_, _07588_, _07589_, _07590_, _07591_, _07592_, _07593_, _07594_, _07595_, _07596_, _07597_, _07598_, _07599_, _07600_, _07601_, _07602_, _07603_, _07604_, _07605_, _07606_, _07607_, _07608_, _07609_, _07610_, _07611_, _07612_, _07613_, _07614_, _07615_, _07616_, _07617_, _07618_, _07619_, _07620_, _07621_, _07622_, _07623_, _07624_, _07625_, _07626_, _07627_, _07628_, _07629_, _07630_, _07631_, _07632_, _07633_, _07634_, _07635_, _07636_, _07637_, _07638_, _07639_, _07640_, _07641_, _07642_, _07643_, _07644_, _07645_, _07646_, _07647_, _07648_, _07649_, _07650_, _07651_, _07652_, _07653_, _07654_, _07655_, _07656_, _07657_, _07658_, _07659_, _07660_, _07661_, _07662_, _07663_, _07664_, _07665_, _07666_, _07667_, _07668_, _07669_, _07670_, _07671_, _07672_, _07673_, _07674_, _07675_, _07676_, _07677_, _07678_, _07679_, _07680_, _07681_, _07682_, _07683_, _07684_, _07685_, _07686_, _07687_, _07688_, _07689_, _07690_, _07691_, _07692_, _07693_, _07694_, _07695_, _07696_, _07697_, _07698_, _07699_, _07700_, _07701_, _07702_, _07703_, _07704_, _07705_, _07706_, _07707_, _07708_, _07709_, _07710_, _07711_, _07712_, _07713_, _07714_, _07715_, _07716_, _07717_, _07718_, _07719_, _07720_, _07721_, _07722_, _07723_, _07724_, _07725_, _07726_, _07727_, _07728_, _07729_, _07730_, _07731_, _07732_, _07733_, _07734_, _07735_, _07736_, _07737_, _07738_, _07739_, _07740_, _07741_, _07742_, _07743_, _07744_, _07745_, _07746_, _07747_, _07748_, _07749_, _07750_, _07751_, _07752_, _07753_, _07754_, _07755_, _07756_, _07757_, _07758_, _07759_, _07760_, _07761_, _07762_, _07763_, _07764_, _07765_, _07766_, _07767_, _07768_, _07769_, _07770_, _07771_, _07772_, _07773_, _07774_, _07775_, _07776_, _07777_, _07778_, _07779_, _07780_, _07781_, _07782_, _07783_, _07784_, _07785_, _07786_, _07787_, _07788_, _07789_, _07790_, _07791_, _07792_, _07793_, _07794_, _07795_, _07796_, _07797_, _07798_, _07799_, _07800_, _07801_, _07802_, _07803_, _07804_, _07805_, _07806_, _07807_, _07808_, _07809_, _07810_, _07811_, _07812_, _07813_, _07814_, _07815_, _07816_, _07817_, _07818_, _07819_, _07820_, _07821_, _07822_, _07823_, _07824_, _07825_, _07826_, _07827_, _07828_, _07829_, _07830_, _07831_, _07832_, _07833_, _07834_, _07835_, _07836_, _07837_, _07838_, _07839_, _07840_, _07841_, _07842_, _07843_, _07844_, _07845_, _07846_, _07847_, _07848_, _07849_, _07850_, _07851_, _07852_, _07853_, _07854_, _07855_, _07856_, _07857_, _07858_, _07859_, _07860_, _07861_, _07862_, _07863_, _07864_, _07865_, _07866_, _07867_, _07868_, _07869_, _07870_, _07871_, _07872_, _07873_, _07874_, _07875_, _07876_, _07877_, _07878_, _07879_, _07880_, _07881_, _07882_, _07883_, _07884_, _07885_, _07886_, _07887_, _07888_, _07889_, _07890_, _07891_, _07892_, _07893_, _07894_, _07895_, _07896_, _07897_, _07898_, _07899_, _07900_, _07901_, _07902_, _07903_, _07904_, _07905_, _07906_, _07907_, _07908_, _07909_, _07910_, _07911_, _07912_, _07913_, _07914_, _07915_, _07916_, _07917_, _07918_, _07919_, _07920_, _07921_, _07922_, _07923_, _07924_, _07925_, _07926_, _07927_, _07928_, _07929_, _07930_, _07931_, _07932_, _07933_, _07934_, _07935_, _07936_, _07937_, _07938_, _07939_, _07940_, _07941_, _07942_, _07943_, _07944_, _07945_, _07946_, _07947_, _07948_, _07949_, _07950_, _07951_, _07952_, _07953_, _07954_, _07955_, _07956_, _07957_, _07958_, _07959_, _07960_, _07961_, _07962_, _07963_, _07964_, _07965_, _07966_, _07967_, _07968_, _07969_, _07970_, _07971_, _07972_, _07973_, _07974_, _07975_, _07976_, _07977_, _07978_, _07979_, _07980_, _07981_, _07982_, _07983_, _07984_, _07985_, _07986_, _07987_, _07988_, _07989_, _07990_, _07991_, _07992_, _07993_, _07994_, _07995_, _07996_, _07997_, _07998_, _07999_, _08000_, _08001_, _08002_, _08003_, _08004_, _08005_, _08006_, _08007_, _08008_, _08009_, _08010_, _08011_, _08012_, _08013_, _08014_, _08015_, _08016_, _08017_, _08018_, _08019_, _08020_, _08021_, _08022_, _08023_, _08024_, _08025_, _08026_, _08027_, _08028_, _08029_, _08030_, _08031_, _08032_, _08033_, _08034_, _08035_, _08036_, _08037_, _08038_, _08039_, _08040_, _08041_, _08042_, _08043_, _08044_, _08045_, _08046_, _08047_, _08048_, _08049_, _08050_, _08051_, _08052_, _08053_, _08054_, _08055_, _08056_, _08057_, _08058_, _08059_, _08060_, _08061_, _08062_, _08063_, _08064_, _08065_, _08066_, _08067_, _08068_, _08069_, _08070_, _08071_, _08072_, _08073_, _08074_, _08075_, _08076_, _08077_, _08078_, _08079_, _08080_, _08081_, _08082_, _08083_, _08084_, _08085_, _08086_, _08087_, _08088_, _08089_, _08090_, _08091_, _08092_, _08093_, _08094_, _08095_, _08096_, _08097_, _08098_, _08099_, _08100_, _08101_, _08102_, _08103_, _08104_, _08105_, _08106_, _08107_, _08108_, _08109_, _08110_, _08111_, _08112_, _08113_, _08114_, _08115_, _08116_, _08117_, _08118_, _08119_, _08120_, _08121_, _08122_, _08123_, _08124_, _08125_, _08126_, _08127_, _08128_, _08129_, _08130_, _08131_, _08132_, _08133_, _08134_, _08135_, _08136_, _08137_, _08138_, _08139_, _08140_, _08141_, _08142_, _08143_, _08144_, _08145_, _08146_, _08147_, _08148_, _08149_, _08150_, _08151_, _08152_, _08153_, _08154_, _08155_, _08156_, _08157_, _08158_, _08159_, _08160_, _08161_, _08162_, _08163_, _08164_, _08165_, _08166_, _08167_, _08168_, _08169_, _08170_, _08171_, _08172_, _08173_, _08174_, _08175_, _08176_, _08177_, _08178_, _08179_, _08180_, _08181_, _08182_, _08183_, _08184_, _08185_, _08186_, _08187_, _08188_, _08189_, _08190_, _08191_, _08192_, _08193_, _08194_, _08195_, _08196_, _08197_, _08198_, _08199_, _08200_, _08201_, _08202_, _08203_, _08204_, _08205_, _08206_, _08207_, _08208_, _08209_, _08210_, _08211_, _08212_, _08213_, _08214_, _08215_, _08216_, _08217_, _08218_, _08219_, _08220_, _08221_, _08222_, _08223_, _08224_, _08225_, _08226_, _08227_, _08228_, _08229_, _08230_, _08231_, _08232_, _08233_, _08234_, _08235_, _08236_, _08237_, _08238_, _08239_, _08240_, _08241_, _08242_, _08243_, _08244_, _08245_, _08246_, _08247_, _08248_, _08249_, _08250_, _08251_, _08252_, _08253_, _08254_, _08255_, _08256_, _08257_, _08258_, _08259_, _08260_, _08261_, _08262_, _08263_, _08264_, _08265_, _08266_, _08267_, _08268_, _08269_, _08270_, _08271_, _08272_, _08273_, _08274_, _08275_, _08276_, _08277_, _08278_, _08279_, _08280_, _08281_, _08282_, _08283_, _08284_, _08285_, _08286_, _08287_, _08288_, _08289_, _08290_, _08291_, _08292_, _08293_, _08294_, _08295_, _08296_, _08297_, _08298_, _08299_, _08300_, _08301_, _08302_, _08303_, _08304_, _08305_, _08306_, _08307_, _08308_, _08309_, _08310_, _08311_, _08312_, _08313_, _08314_, _08315_, _08316_, _08317_, _08318_, _08319_, _08320_, _08321_, _08322_, _08323_, _08324_, _08325_, _08326_, _08327_, _08328_, _08329_, _08330_, _08331_, _08332_, _08333_, _08334_, _08335_, _08336_, _08337_, _08338_, _08339_, _08340_, _08341_, _08342_, _08343_, _08344_, _08345_, _08346_, _08347_, _08348_, _08349_, _08350_, _08351_, _08352_, _08353_, _08354_, _08355_, _08356_, _08357_, _08358_, _08359_, _08360_, _08361_, _08362_, _08363_, _08364_, _08365_, _08366_, _08367_, _08368_, _08369_, _08370_, _08371_, _08372_, _08373_, _08374_, _08375_, _08376_, _08377_, _08378_, _08379_, _08380_, _08381_, _08382_, _08383_, _08384_, _08385_, _08386_, _08387_, _08388_, _08389_, _08390_, _08391_, _08392_, _08393_, _08394_, _08395_, _08396_, _08397_, _08398_, _08399_, _08400_, _08401_, _08402_, _08403_, _08404_, _08405_, _08406_, _08407_, _08408_, _08409_, _08410_, _08411_, _08412_, _08413_, _08414_, _08415_, _08416_, _08417_, _08418_, _08419_, _08420_, _08421_, _08422_, _08423_, _08424_, _08425_, _08426_, _08427_, _08428_, _08429_, _08430_, _08431_, _08432_, _08433_, _08434_, _08435_, _08436_, _08437_, _08438_, _08439_, _08440_, _08441_, _08442_, _08443_, _08444_, _08445_, _08446_, _08447_, _08448_, _08449_, _08450_, _08451_, _08452_, _08453_, _08454_, _08455_, _08456_, _08457_, _08458_, _08459_, _08460_, _08461_, _08462_, _08463_, _08464_, _08465_, _08466_, _08467_, _08468_, _08469_, _08470_, _08471_, _08472_, _08473_, _08474_, _08475_, _08476_, _08477_, _08478_, _08479_, _08480_, _08481_, _08482_, _08483_, _08484_, _08485_, _08486_, _08487_, _08488_, _08489_, _08490_, _08491_, _08492_, _08493_, _08494_, _08495_, _08496_, _08497_, _08498_, _08499_, _08500_, _08501_, _08502_, _08503_, _08504_, _08505_, _08506_, _08507_, _08508_, _08509_, _08510_, _08511_, _08512_, _08513_, _08514_, _08515_, _08516_, _08517_, _08518_, _08519_, _08520_, _08521_, _08522_, _08523_, _08524_, _08525_, _08526_, _08527_, _08528_, _08529_, _08530_, _08531_, _08532_, _08533_, _08534_, _08535_, _08536_, _08537_, _08538_, _08539_, _08540_, _08541_, _08542_, _08543_, _08544_, _08545_, _08546_, _08547_, _08548_, _08549_, _08550_, _08551_, _08552_, _08553_, _08554_, _08555_, _08556_, _08557_, _08558_, _08559_, _08560_, _08561_, _08562_, _08563_, _08564_, _08565_, _08566_, _08567_, _08568_, _08569_, _08570_, _08571_, _08572_, _08573_, _08574_, _08575_, _08576_, _08577_, _08578_, _08579_, _08580_, _08581_, _08582_, _08583_, _08584_, _08585_, _08586_, _08587_, _08588_, _08589_, _08590_, _08591_, _08592_, _08593_, _08594_, _08595_, _08596_, _08597_, _08598_, _08599_, _08600_, _08601_, _08602_, _08603_, _08604_, _08605_, _08606_, _08607_, _08608_, _08609_, _08610_, _08611_, _08612_, _08613_, _08614_, _08615_, _08616_, _08617_, _08618_, _08619_, _08620_, _08621_, _08622_, _08623_, _08624_, _08625_, _08626_, _08627_, _08628_, _08629_, _08630_, _08631_, _08632_, _08633_, _08634_, _08635_, _08636_, _08637_, _08638_, _08639_, _08640_, _08641_, _08642_, _08643_, _08644_, _08645_, _08646_, _08647_, _08648_, _08649_, _08650_, _08651_, _08652_, _08653_, _08654_, _08655_, _08656_, _08657_, _08658_, _08659_, _08660_, _08661_, _08662_, _08663_, _08664_, _08665_, _08666_, _08667_, _08668_, _08669_, _08670_, _08671_, _08672_, _08673_, _08674_, _08675_, _08676_, _08677_, _08678_, _08679_, _08680_, _08681_, _08682_, _08683_, _08684_, _08685_, _08686_, _08687_, _08688_, _08689_, _08690_, _08691_, _08692_, _08693_, _08694_, _08695_, _08696_, _08697_, _08698_, _08699_, _08700_, _08701_, _08702_, _08703_, _08704_, _08705_, _08706_, _08707_, _08708_, _08709_, _08710_, _08711_, _08712_, _08713_, _08714_, _08715_, _08716_, _08717_, _08718_, _08719_, _08720_, _08721_, _08722_, _08723_, _08724_, _08725_, _08726_, _08727_, _08728_, _08729_, _08730_, _08731_, _08732_, _08733_, _08734_, _08735_, _08736_, _08737_, _08738_, _08739_, _08740_, _08741_, _08742_, _08743_, _08744_, _08745_, _08746_, _08747_, _08748_, _08749_, _08750_, _08751_, _08752_, _08753_, _08754_, _08755_, _08756_, _08757_, _08758_, _08759_, _08760_, _08761_, _08762_, _08763_, _08764_, _08765_, _08766_, _08767_, _08768_, _08769_, _08770_, _08771_, _08772_, _08773_, _08774_, _08775_, _08776_, _08777_, _08778_, _08779_, _08780_, _08781_, _08782_, _08783_, _08784_, _08785_, _08786_, _08787_, _08788_, _08789_, _08790_, _08791_, _08792_, _08793_, _08794_, _08795_, _08796_, _08797_, _08798_, _08799_, _08800_, _08801_, _08802_, _08803_, _08804_, _08805_, _08806_, _08807_, _08808_, _08809_, _08810_, _08811_, _08812_, _08813_, _08814_, _08815_, _08816_, _08817_, _08818_, _08819_, _08820_, _08821_, _08822_, _08823_, _08824_, _08825_, _08826_, _08827_, _08828_, _08829_, _08830_, _08831_, _08832_, _08833_, _08834_, _08835_, _08836_, _08837_, _08838_, _08839_, _08840_, _08841_, _08842_, _08843_, _08844_, _08845_, _08846_, _08847_, _08848_, _08849_, _08850_, _08851_, _08852_, _08853_, _08854_, _08855_, _08856_, _08857_, _08858_, _08859_, _08860_, _08861_, _08862_, _08863_, _08864_, _08865_, _08866_, _08867_, _08868_, _08869_, _08870_, _08871_, _08872_, _08873_, _08874_, _08875_, _08876_, _08877_, _08878_, _08879_, _08880_, _08881_, _08882_, _08883_, _08884_, _08885_, _08886_, _08887_, _08888_, _08889_, _08890_, _08891_, _08892_, _08893_, _08894_, _08895_, _08896_, _08897_, _08898_, _08899_, _08900_, _08901_, _08902_, _08903_, _08904_, _08905_, _08906_, _08907_, _08908_, _08909_, _08910_, _08911_, _08912_, _08913_, _08914_, _08915_, _08916_, _08917_, _08918_, _08919_, _08920_, _08921_, _08922_, _08923_, _08924_, _08925_, _08926_, _08927_, _08928_, _08929_, _08930_, _08931_, _08932_, _08933_, _08934_, _08935_, _08936_, _08937_, _08938_, _08939_, _08940_, _08941_, _08942_, _08943_, _08944_, _08945_, _08946_, _08947_, _08948_, _08949_, _08950_, _08951_, _08952_, _08953_, _08954_, _08955_, _08956_, _08957_, _08958_, _08959_, _08960_, _08961_, _08962_, _08963_, _08964_, _08965_, _08966_, _08967_, _08968_, _08969_, _08970_, _08971_, _08972_, _08973_, _08974_, _08975_, _08976_, _08977_, _08978_, _08979_, _08980_, _08981_, _08982_, _08983_, _08984_, _08985_, _08986_, _08987_, _08988_, _08989_, _08990_, _08991_, _08992_, _08993_, _08994_, _08995_, _08996_, _08997_, _08998_, _08999_, _09000_, _09001_, _09002_, _09003_, _09004_, _09005_, _09006_, _09007_, _09008_, _09009_, _09010_, _09011_, _09012_, _09013_, _09014_, _09015_, _09016_, _09017_, _09018_, _09019_, _09020_, _09021_, _09022_, _09023_, _09024_, _09025_, _09026_, _09027_, _09028_, _09029_, _09030_, _09031_, _09032_, _09033_, _09034_, _09035_, _09036_, _09037_, _09038_, _09039_, _09040_, _09041_, _09042_, _09043_, _09044_, _09045_, _09046_, _09047_, _09048_, _09049_, _09050_, _09051_, _09052_, _09053_, _09054_, _09055_, _09056_, _09057_, _09058_, _09059_, _09060_, _09061_, _09062_, _09063_, _09064_, _09065_, _09066_, _09067_, _09068_, _09069_, _09070_, _09071_, _09072_, _09073_, _09074_, _09075_, _09076_, _09077_, _09078_, _09079_, _09080_, _09081_, _09082_, _09083_, _09084_, _09085_, _09086_, _09087_, _09088_, _09089_, _09090_, _09091_, _09092_, _09093_, _09094_, _09095_, _09096_, _09097_, _09098_, _09099_, _09100_, _09101_, _09102_, _09103_, _09104_, _09105_, _09106_, _09107_, _09108_, _09109_, _09110_, _09111_, _09112_, _09113_, _09114_, _09115_, _09116_, _09117_, _09118_, _09119_, _09120_, _09121_, _09122_, _09123_, _09124_, _09125_, _09126_, _09127_, _09128_, _09129_, _09130_, _09131_, _09132_, _09133_, _09134_, _09135_, _09136_, _09137_, _09138_, _09139_, _09140_, _09141_, _09142_, _09143_, _09144_, _09145_, _09146_, _09147_, _09148_, _09149_, _09150_, _09151_, _09152_, _09153_, _09154_, _09155_, _09156_, _09157_, _09158_, _09159_, _09160_, _09161_, _09162_, _09163_, _09164_, _09165_, _09166_, _09167_, _09168_, _09169_, _09170_, _09171_, _09172_, _09173_, _09174_, _09175_, _09176_, _09177_, _09178_, _09179_, _09180_, _09181_, _09182_, _09183_, _09184_, _09185_, _09186_, _09187_, _09188_, _09189_, _09190_, _09191_, _09192_, _09193_, _09194_, _09195_, _09196_, _09197_, _09198_, _09199_, _09200_, _09201_, _09202_, _09203_, _09204_, _09205_, _09206_, _09207_, _09208_, _09209_, _09210_, _09211_, _09212_, _09213_, _09214_, _09215_, _09216_, _09217_, _09218_, _09219_, _09220_, _09221_, _09222_, _09223_, _09224_, _09225_, _09226_, _09227_, _09228_, _09229_, _09230_, _09231_, _09232_, _09233_, _09234_, _09235_, _09236_, _09237_, _09238_, _09239_, _09240_, _09241_, _09242_, _09243_, _09244_, _09245_, _09246_, _09247_, _09248_, _09249_, _09250_, _09251_, _09252_, _09253_, _09254_, _09255_, _09256_, _09257_, _09258_, _09259_, _09260_, _09261_, _09262_, _09263_, _09264_, _09265_, _09266_, _09267_, _09268_, _09269_, _09270_, _09271_, _09272_, _09273_, _09274_, _09275_, _09276_, _09277_, _09278_, _09279_, _09280_, _09281_, _09282_, _09283_, _09284_, _09285_, _09286_, _09287_, _09288_, _09289_, _09290_, _09291_, _09292_, _09293_, _09294_, _09295_, _09296_, _09297_, _09298_, _09299_, _09300_, _09301_, _09302_, _09303_, _09304_, _09305_, _09306_, _09307_, _09308_, _09309_, _09310_, _09311_, _09312_, _09313_, _09314_, _09315_, _09316_, _09317_, _09318_, _09319_, _09320_, _09321_, _09322_, _09323_, _09324_, _09325_, _09326_, _09327_, _09328_, _09329_, _09330_, _09331_, _09332_, _09333_, _09334_, _09335_, _09336_, _09337_, _09338_, _09339_, _09340_, _09341_, _09342_, _09343_, _09344_, _09345_, _09346_, _09347_, _09348_, _09349_, _09350_, _09351_, _09352_, _09353_, _09354_, _09355_, _09356_, _09357_, _09358_, _09359_, _09360_, _09361_, _09362_, _09363_, _09364_, _09365_, _09366_, _09367_, _09368_, _09369_, _09370_, _09371_, _09372_, _09373_, _09374_, _09375_, _09376_, _09377_, _09378_, _09379_, _09380_, _09381_, _09382_, _09383_, _09384_, _09385_, _09386_, _09387_, _09388_, _09389_, _09390_, _09391_, _09392_, _09393_, _09394_, _09395_, _09396_, _09397_, _09398_, _09399_, _09400_, _09401_, _09402_, _09403_, _09404_, _09405_, _09406_, _09407_, _09408_, _09409_, _09410_, _09411_, _09412_, _09413_, _09414_, _09415_, _09416_, _09417_, _09418_, _09419_, _09420_, _09421_, _09422_, _09423_, _09424_, _09425_, _09426_, _09427_, _09428_, _09429_, _09430_, _09431_, _09432_, _09433_, _09434_, _09435_, _09436_, _09437_, _09438_, _09439_, _09440_, _09441_, _09442_, _09443_, _09444_, _09445_, _09446_, _09447_, _09448_, _09449_, _09450_, _09451_, _09452_, _09453_, _09454_, _09455_, _09456_, _09457_, _09458_, _09459_, _09460_, _09461_, _09462_, _09463_, _09464_, _09465_, _09466_, _09467_, _09468_, _09469_, _09470_, _09471_, _09472_, _09473_, _09474_, _09475_, _09476_, _09477_, _09478_, _09479_, _09480_, _09481_, _09482_, _09483_, _09484_, _09485_, _09486_, _09487_, _09488_, _09489_, _09490_, _09491_, _09492_, _09493_, _09494_, _09495_, _09496_, _09497_, _09498_, _09499_, _09500_, _09501_, _09502_, _09503_, _09504_, _09505_, _09506_, _09507_, _09508_, _09509_, _09510_, _09511_, _09512_, _09513_, _09514_, _09515_, _09516_, _09517_, _09518_, _09519_, _09520_, _09521_, _09522_, _09523_, _09524_, _09525_, _09526_, _09527_, _09528_, _09529_, _09530_, _09531_, _09532_, _09533_, _09534_, _09535_, _09536_, _09537_, _09538_, _09539_, _09540_, _09541_, _09542_, _09543_, _09544_, _09545_, _09546_, _09547_, _09548_, _09549_, _09550_, _09551_, _09552_, _09553_, _09554_, _09555_, _09556_, _09557_, _09558_, _09559_, _09560_, _09561_, _09562_, _09563_, _09564_, _09565_, _09566_, _09567_, _09568_, _09569_, _09570_, _09571_, _09572_, _09573_, _09574_, _09575_, _09576_, _09577_, _09578_, _09579_, _09580_, _09581_, _09582_, _09583_, _09584_, _09585_, _09586_, _09587_, _09588_, _09589_, _09590_, _09591_, _09592_, _09593_, _09594_, _09595_, _09596_, _09597_, _09598_, _09599_, _09600_, _09601_, _09602_, _09603_, _09604_, _09605_, _09606_, _09607_, _09608_, _09609_, _09610_, _09611_, _09612_, _09613_, _09614_, _09615_, _09616_, _09617_, _09618_, _09619_, _09620_, _09621_, _09622_, _09623_, _09624_, _09625_, _09626_, _09627_, _09628_, _09629_, _09630_, _09631_, _09632_, _09633_, _09634_, _09635_, _09636_, _09637_, _09638_, _09639_, _09640_, _09641_, _09642_, _09643_, _09644_, _09645_, _09646_, _09647_, _09648_, _09649_, _09650_, _09651_, _09652_, _09653_, _09654_, _09655_, _09656_, _09657_, _09658_, _09659_, _09660_, _09661_, _09662_, _09663_, _09664_, _09665_, _09666_, _09667_, _09668_, _09669_, _09670_, _09671_, _09672_, _09673_, _09674_, _09675_, _09676_, _09677_, _09678_, _09679_, _09680_, _09681_, _09682_, _09683_, _09684_, _09685_, _09686_, _09687_, _09688_, _09689_, _09690_, _09691_, _09692_, _09693_, _09694_, _09695_, _09696_, _09697_, _09698_, _09699_, _09700_, _09701_, _09702_, _09703_, _09704_, _09705_, _09706_, _09707_, _09708_, _09709_, _09710_, _09711_, _09712_, _09713_, _09714_, _09715_, _09716_, _09717_, _09718_, _09719_, _09720_, _09721_, _09722_, _09723_, _09724_, _09725_, _09726_, _09727_, _09728_, _09729_, _09730_, _09731_, _09732_, _09733_, _09734_, _09735_, _09736_, _09737_, _09738_, _09739_, _09740_, _09741_, _09742_, _09743_, _09744_, _09745_, _09746_, _09747_, _09748_, _09749_, _09750_, _09751_, _09752_, _09753_, _09754_, _09755_, _09756_, _09757_, _09758_, _09759_, _09760_, _09761_, _09762_, _09763_, _09764_, _09765_, _09766_, _09767_, _09768_, _09769_, _09770_, _09771_, _09772_, _09773_, _09774_, _09775_, _09776_, _09777_, _09778_, _09779_, _09780_, _09781_, _09782_, _09783_, _09784_, _09785_, _09786_, _09787_, _09788_, _09789_, _09790_, _09791_, _09792_, _09793_, _09794_, _09795_, _09796_, _09797_, _09798_, _09799_, _09800_, _09801_, _09802_, _09803_, _09804_, _09805_, _09806_, _09807_, _09808_, _09809_, _09810_, _09811_, _09812_, _09813_, _09814_, _09815_, _09816_, _09817_, _09818_, _09819_, _09820_, _09821_, _09822_, _09823_, _09824_, _09825_, _09826_, _09827_, _09828_, _09829_, _09830_, _09831_, _09832_, _09833_, _09834_, _09835_, _09836_, _09837_, _09838_, _09839_, _09840_, _09841_, _09842_, _09843_, _09844_, _09845_, _09846_, _09847_, _09848_, _09849_, _09850_, _09851_, _09852_, _09853_, _09854_, _09855_, _09856_, _09857_, _09858_, _09859_, _09860_, _09861_, _09862_, _09863_, _09864_, _09865_, _09866_, _09867_, _09868_, _09869_, _09870_, _09871_, _09872_, _09873_, _09874_, _09875_, _09876_, _09877_, _09878_, _09879_, _09880_, _09881_, _09882_, _09883_, _09884_, _09885_, _09886_, _09887_, _09888_, _09889_, _09890_, _09891_, _09892_, _09893_, _09894_, _09895_, _09896_, _09897_, _09898_, _09899_, _09900_, _09901_, _09902_, _09903_, _09904_, _09905_, _09906_, _09907_, _09908_, _09909_, _09910_, _09911_, _09912_, _09913_, _09914_, _09915_, _09916_, _09917_, _09918_, _09919_, _09920_, _09921_, _09922_, _09923_, _09924_, _09925_, _09926_, _09927_, _09928_, _09929_, _09930_, _09931_, _09932_, _09933_, _09934_, _09935_, _09936_, _09937_, _09938_, _09939_, _09940_, _09941_, _09942_, _09943_, _09944_, _09945_, _09946_, _09947_, _09948_, _09949_, _09950_, _09951_, _09952_, _09953_, _09954_, _09955_, _09956_, _09957_, _09958_, _09959_, _09960_, _09961_, _09962_, _09963_, _09964_, _09965_, _09966_, _09967_, _09968_, _09969_, _09970_, _09971_, _09972_, _09973_, _09974_, _09975_, _09976_, _09977_, _09978_, _09979_, _09980_, _09981_, _09982_, _09983_, _09984_, _09985_, _09986_, _09987_, _09988_, _09989_, _09990_, _09991_, _09992_, _09993_, _09994_, _09995_, _09996_, _09997_, _09998_, _09999_, _10000_, _10001_, _10002_, _10003_, _10004_, _10005_, _10006_, _10007_, _10008_, _10009_, _10010_, _10011_, _10012_, _10013_, _10014_, _10015_, _10016_, _10017_, _10018_, _10019_, _10020_, _10021_, _10022_, _10023_, _10024_, _10025_, _10026_, _10027_, _10028_, _10029_, _10030_, _10031_, _10032_, _10033_, _10034_, _10035_, _10036_, _10037_, _10038_, _10039_, _10040_, _10041_, _10042_, _10043_, _10044_, _10045_, _10046_, _10047_, _10048_, _10049_, _10050_, _10051_, _10052_, _10053_, _10054_, _10055_, _10056_, _10057_, _10058_, _10059_, _10060_, _10061_, _10062_, _10063_, _10064_, _10065_, _10066_, _10067_, _10068_, _10069_, _10070_, _10071_, _10072_, _10073_, _10074_, _10075_, _10076_, _10077_, _10078_, _10079_, _10080_, _10081_, _10082_, _10083_, _10084_, _10085_, _10086_, _10087_, _10088_, _10089_, _10090_, _10091_, _10092_, _10093_, _10094_, _10095_, _10096_, _10097_, _10098_, _10099_, _10100_, _10101_, _10102_, _10103_, _10104_, _10105_, _10106_, _10107_, _10108_, _10109_, _10110_, _10111_, _10112_, _10113_, _10114_, _10115_, _10116_, _10117_, _10118_, _10119_, _10120_, _10121_, _10122_, _10123_, _10124_, _10125_, _10126_, _10127_, _10128_, _10129_, _10130_, _10131_, _10132_, _10133_, _10134_, _10135_, _10136_, _10137_, _10138_, _10139_, _10140_, _10141_, _10142_, _10143_, _10144_, _10145_, _10146_, _10147_, _10148_, _10149_, _10150_, _10151_, _10152_, _10153_, _10154_, _10155_, _10156_, _10157_, _10158_, _10159_, _10160_, _10161_, _10162_, _10163_, _10164_, _10165_, _10166_, _10167_, _10168_, _10169_, _10170_, _10171_, _10172_, _10173_, _10174_, _10175_, _10176_, _10177_, _10178_, _10179_, _10180_, _10181_, _10182_, _10183_, _10184_, _10185_, _10186_, _10187_, _10188_, _10189_, _10190_, _10191_, _10192_, _10193_, _10194_, _10195_, _10196_, _10197_, _10198_, _10199_, _10200_, _10201_, _10202_, _10203_, _10204_, _10205_, _10206_, _10207_, _10208_, _10209_, _10210_, _10211_, _10212_, _10213_, _10214_, _10215_, _10216_, _10217_, _10218_, _10219_, _10220_, _10221_, _10222_, _10223_, _10224_, _10225_, _10226_, _10227_, _10228_, _10229_, _10230_, _10231_, _10232_, _10233_, _10234_, _10235_, _10236_, _10237_, _10238_, _10239_, _10240_, _10241_, _10242_, _10243_, _10244_, _10245_, _10246_, _10247_, _10248_, _10249_, _10250_, _10251_, _10252_, _10253_, _10254_, _10255_, _10256_, _10257_, _10258_, _10259_, _10260_, _10261_, _10262_, _10263_, _10264_, _10265_, _10266_, _10267_, _10268_, _10269_, _10270_, _10271_, _10272_, _10273_, _10274_, _10275_, _10276_, _10277_, _10278_, _10279_, _10280_, _10281_, _10282_, _10283_, _10284_, _10285_, _10286_, _10287_, _10288_, _10289_, _10290_, _10291_, _10292_, _10293_, _10294_, _10295_, _10296_, _10297_, _10298_, _10299_, _10300_, _10301_, _10302_, _10303_, _10304_, _10305_, _10306_, _10307_, _10308_, _10309_, _10310_, _10311_, _10312_, _10313_, _10314_, _10315_, _10316_, _10317_, _10318_, _10319_, _10320_, _10321_, _10322_, _10323_, _10324_, _10325_, _10326_, _10327_, _10328_, _10329_, _10330_, _10331_, _10332_, _10333_, _10334_, _10335_, _10336_, _10337_, _10338_, _10339_, _10340_, _10341_, _10342_, _10343_, _10344_, _10345_, _10346_, _10347_, _10348_, _10349_, _10350_, _10351_, _10352_, _10353_, _10354_, _10355_, _10356_, _10357_, _10358_, _10359_, _10360_, _10361_, _10362_, _10363_, _10364_, _10365_, _10366_, _10367_, _10368_, _10369_, _10370_, _10371_, _10372_, _10373_, _10374_, _10375_, _10376_, _10377_, _10378_, _10379_, _10380_, _10381_, _10382_, _10383_, _10384_, _10385_, _10386_, _10387_, _10388_, _10389_, _10390_, _10391_, _10392_, _10393_, _10394_, _10395_, _10396_, _10397_, _10398_, _10399_, _10400_, _10401_, _10402_, _10403_, _10404_, _10405_, _10406_, _10407_, _10408_, _10409_, _10410_, _10411_, _10412_, _10413_, _10414_, _10415_, _10416_, _10417_, _10418_, _10419_, _10420_, _10421_, _10422_, _10423_, _10424_, _10425_, _10426_, _10427_, _10428_, _10429_, _10430_, _10431_, _10432_, _10433_, _10434_, _10435_, _10436_, _10437_, _10438_, _10439_, _10440_, _10441_, _10442_, _10443_, _10444_, _10445_, _10446_, _10447_, _10448_, _10449_, _10450_, _10451_, _10452_, _10453_, _10454_, _10455_, _10456_, _10457_, _10458_, _10459_, _10460_, _10461_, _10462_, _10463_, _10464_, _10465_, _10466_, _10467_, _10468_, _10469_, _10470_, _10471_, _10472_, _10473_, _10474_, _10475_, _10476_, _10477_, _10478_, _10479_, _10480_, _10481_, _10482_, _10483_, _10484_, _10485_, _10486_, _10487_, _10488_, _10489_, _10490_, _10491_, _10492_, _10493_, _10494_, _10495_, _10496_, _10497_, _10498_, _10499_, _10500_, _10501_, _10502_, _10503_, _10504_, _10505_, _10506_, _10507_, _10508_, _10509_, _10510_, _10511_, _10512_, _10513_, _10514_, _10515_, _10516_, _10517_, _10518_, _10519_, _10520_, _10521_, _10522_, _10523_, _10524_, _10525_, _10526_, _10527_, _10528_, _10529_, _10530_, _10531_, _10532_, _10533_, _10534_, _10535_, _10536_, _10537_, _10538_, _10539_, _10540_, _10541_, _10542_, _10543_, _10544_, _10545_, _10546_, _10547_, _10548_, _10549_, _10550_, _10551_, _10552_, _10553_, _10554_, _10555_, _10556_, _10557_, _10558_, _10559_, _10560_, _10561_, _10562_, _10563_, _10564_, _10565_, _10566_, _10567_, _10568_, _10569_, _10570_, _10571_, _10572_, _10573_, _10574_, _10575_, _10576_, _10577_, _10578_, _10579_, _10580_, _10581_, _10582_, _10583_, _10584_, _10585_, _10586_, _10587_, _10588_, _10589_, _10590_, _10591_, _10592_, _10593_, _10594_, _10595_, _10596_, , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , ;
  input [159:0] set1;
  input [159:0] set2;
  input set1[0], set1[1], set1[2], set1[3], set1[4], set1[5], set1[6], set1[7], set1[8], set1[9], set1[10], set1[11], set1[12], set1[13], set1[14], set1[15], set1[16], set1[17], set1[18], set1[19], set1[20], set1[21], set1[22], set1[23], set1[24], set1[25], set1[26], set1[27], set1[28], set1[29], set1[30], set1[31], set1[32], set1[33], set1[34], set1[35], set1[36], set1[37], set1[38], set1[39], set1[40], set1[41], set1[42], set1[43], set1[44], set1[45], set1[46], set1[47], set1[48], set1[49], set1[50], set1[51], set1[52], set1[53], set1[54], set1[55], set1[56], set1[57], set1[58], set1[59], set1[60], set1[61], set1[62], set1[63], set1[64], set1[65], set1[66], set1[67], set1[68], set1[69], set1[70], set1[71], set1[72], set1[73], set1[74], set1[75], set1[76], set1[77], set1[78], set1[79], set1[80], set1[81], set1[82], set1[83], set1[84], set1[85], set1[86], set1[87], set1[88], set1[89], set1[90], set1[91], set1[92], set1[93], set1[94], set1[95], set1[96], set1[97], set1[98], set1[99], set1[100], set1[101], set1[102], set1[103], set1[104], set1[105], set1[106], set1[107], set1[108], set1[109], set1[110], set1[111], set1[112], set1[113], set1[114], set1[115], set1[116], set1[117], set1[118], set1[119], set1[120], set1[121], set1[122], set1[123], set1[124], set1[125], set1[126], set1[127], set1[128], set1[129], set1[130], set1[131], set1[132], set1[133], set1[134], set1[135], set1[136], set1[137], set1[138], set1[139], set1[140], set1[141], set1[142], set1[143], set1[144], set1[145], set1[146], set1[147], set1[148], set1[149], set1[150], set1[151], set1[152], set1[153], set1[154], set1[155], set1[156], set1[157], set1[158], set1[159], set2[0], set2[1], set2[2], set2[3], set2[4], set2[5], set2[6], set2[7], set2[8], set2[9], set2[10], set2[11], set2[12], set2[13], set2[14], set2[15], set2[16], set2[17], set2[18], set2[19], set2[20], set2[21], set2[22], set2[23], set2[24], set2[25], set2[26], set2[27], set2[28], set2[29], set2[30], set2[31], set2[32], set2[33], set2[34], set2[35], set2[36], set2[37], set2[38], set2[39], set2[40], set2[41], set2[42], set2[43], set2[44], set2[45], set2[46], set2[47], set2[48], set2[49], set2[50], set2[51], set2[52], set2[53], set2[54], set2[55], set2[56], set2[57], set2[58], set2[59], set2[60], set2[61], set2[62], set2[63], set2[64], set2[65], set2[66], set2[67], set2[68], set2[69], set2[70], set2[71], set2[72], set2[73], set2[74], set2[75], set2[76], set2[77], set2[78], set2[79], set2[80], set2[81], set2[82], set2[83], set2[84], set2[85], set2[86], set2[87], set2[88], set2[89], set2[90], set2[91], set2[92], set2[93], set2[94], set2[95], set2[96], set2[97], set2[98], set2[99], set2[100], set2[101], set2[102], set2[103], set2[104], set2[105], set2[106], set2[107], set2[108], set2[109], set2[110], set2[111], set2[112], set2[113], set2[114], set2[115], set2[116], set2[117], set2[118], set2[119], set2[120], set2[121], set2[122], set2[123], set2[124], set2[125], set2[126], set2[127], set2[128], set2[129], set2[130], set2[131], set2[132], set2[133], set2[134], set2[135], set2[136], set2[137], set2[138], set2[139], set2[140], set2[141], set2[142], set2[143], set2[144], set2[145], set2[146], set2[147], set2[148], set2[149], set2[150], set2[151], set2[152], set2[153], set2[154], set2[155], set2[156], set2[157], set2[158], set2[159];
  output out[0], out[1], out[2], out[3], out[4], out[5], out[6], out[7], out[8], out[9], out[10], out[11], out[12], out[13], out[14], out[15], out[16], out[17], out[18], out[19], out[20], out[21], out[22], out[23], out[24], out[25], out[26], out[27], out[28], out[29], out[30], out[31], out[32], out[33], out[34], out[35], out[36], out[37], out[38], out[39], out[40], out[41], out[42], out[43], out[44], out[45], out[46], out[47], out[48], out[49], out[50], out[51], out[52], out[53], out[54], out[55], out[56], out[57], out[58], out[59], out[60], out[61], out[62], out[63], out[64], out[65], out[66], out[67], out[68], out[69], out[70], out[71], out[72], out[73], out[74], out[75], out[76], out[77], out[78], out[79], out[80], out[81], out[82], out[83], out[84], out[85], out[86], out[87], out[88], out[89], out[90], out[91], out[92], out[93], out[94], out[95], out[96], out[97], out[98], out[99], out[100], out[101], out[102], out[103], out[104], out[105], out[106], out[107], out[108], out[109], out[110], out[111], out[112], out[113], out[114], out[115], out[116], out[117], out[118], out[119], out[120], out[121], out[122], out[123], out[124], out[125], out[126], out[127], out[128], out[129], out[130], out[131], out[132], out[133], out[134], out[135], out[136], out[137], out[138], out[139], out[140], out[141], out[142], out[143], out[144], out[145], out[146], out[147], out[148], out[149], out[150], out[151], out[152], out[153], out[154], out[155], out[156], out[157], out[158], out[159], out[160], out[161], out[162], out[163], out[164], out[165], out[166], out[167], out[168], out[169], out[170], out[171], out[172], out[173], out[174], out[175], out[176], out[177], out[178], out[179], out[180], out[181], out[182], out[183], out[184], out[185], out[186], out[187], out[188], out[189], out[190], out[191], out[192], out[193], out[194], out[195], out[196], out[197], out[198], out[199], out[200], out[201], out[202], out[203], out[204], out[205], out[206], out[207], out[208], out[209], out[210], out[211], out[212], out[213], out[214], out[215], out[216], out[217], out[218], out[219], out[220], out[221], out[222], out[223], out[224], out[225], out[226], out[227], out[228], out[229], out[230], out[231], out[232], out[233], out[234], out[235], out[236], out[237], out[238], out[239], out[240], out[241], out[242], out[243], out[244], out[245], out[246], out[247], out[248], out[249], out[250], out[251], out[252], out[253], out[254], out[255], out[256], out[257], out[258], out[259], out[260], out[261], out[262], out[263], out[264], out[265], out[266], out[267], out[268], out[269], out[270], out[271], out[272], out[273], out[274], out[275], out[276], out[277], out[278], out[279], out[280], out[281], out[282], out[283], out[284], out[285], out[286], out[287], out[288], out[289], out[290], out[291], out[292], out[293], out[294], out[295], out[296], out[297], out[298], out[299], out[300], out[301], out[302], out[303], out[304], out[305], out[306], out[307], out[308], out[309], out[310], out[311], out[312], out[313], out[314], out[315], out[316], out[317], out[318], out[319], out[320], out[321], out[322], out[323], out[324], out[325], out[326], out[327];
  not g_10597_(out[7], _07700_);
  not g_10598_(out[167], _07711_);
  not g_10599_(out[11], _07722_);
  not g_10600_(out[171], _07733_);
  not g_10601_(out[172], _07744_);
  not g_10602_(out[27], _07755_);
  not g_10603_(out[28], _07766_);
  not g_10604_(out[39], _07777_);
  not g_10605_(out[43], _07788_);
  not g_10606_(out[59], _07799_);
  not g_10607_(out[75], _07810_);
  not g_10608_(out[91], _07821_);
  not g_10609_(out[107], _07832_);
  not g_10610_(out[123], _07843_);
  not g_10611_(out[139], _07854_);
  not g_10612_(out[151], _07865_);
  not g_10613_(out[155], _07876_);
  not g_10614_(out[187], _07887_);
  not g_10615_(out[203], _07898_);
  not g_10616_(out[219], _07909_);
  not g_10617_(out[235], _07920_);
  not g_10618_(out[251], _07931_);
  not g_10619_(out[267], _07942_);
  not g_10620_(out[283], _07953_);
  not g_10621_(out[299], _07964_);
  not g_10622_(out[311], _07975_);
  not g_10623_(out[315], _07986_);
  xor g_10624_(out[146], out[306], _07997_);
  and g_10625_(_07865_, out[311], _08008_);
  xor g_10626_(out[149], out[309], _08019_);
  xor g_10627_(out[155], out[315], _08030_);
  or g_10628_(_08019_, _08030_, _08041_);
  xor g_10629_(out[147], out[307], _08052_);
  xor g_10630_(out[157], out[317], _08063_);
  xor g_10631_(out[148], out[308], _08074_);
  xor g_10632_(out[154], out[314], _08085_);
  xor g_10633_(out[150], out[310], _08096_);
  xor g_10634_(out[153], out[313], _08107_);
  and g_10635_(out[151], _07975_, _08118_);
  or g_10636_(_08052_, _08074_, _08129_);
  xor g_10637_(out[156], out[316], _08140_);
  xor g_10638_(out[145], out[305], _08151_);
  xor g_10639_(out[144], out[304], _08162_);
  xor g_10640_(out[158], out[318], _08173_);
  xor g_10641_(out[152], out[312], _08184_);
  or g_10642_(_08085_, _08096_, _08195_);
  or g_10643_(_08129_, _08195_, _08206_);
  or g_10644_(_08041_, _08063_, _08217_);
  or g_10645_(_08206_, _08217_, _08228_);
  or g_10646_(_08140_, _08162_, _08239_);
  or g_10647_(_08228_, _08239_, _08250_);
  or g_10648_(_07997_, _08008_, _08261_);
  xor g_10649_(out[159], out[319], _08272_);
  or g_10650_(_08173_, _08272_, _08283_);
  or g_10651_(_08261_, _08283_, _08294_);
  or g_10652_(_08107_, _08118_, _08305_);
  or g_10653_(_08151_, _08305_, _08316_);
  or g_10654_(_08294_, _08316_, _08327_);
  or g_10655_(_08184_, _08327_, _08338_);
  or g_10656_(_08250_, _08338_, _08349_);
  xor g_10657_(out[135], out[311], _08360_);
  and g_10658_(_07854_, out[315], _08371_);
  xor g_10659_(out[142], out[318], _08382_);
  xor g_10660_(out[136], out[312], _08393_);
  xor g_10661_(out[129], out[305], _08404_);
  xor g_10662_(out[141], out[317], _08415_);
  xor g_10663_(out[137], out[313], _08425_);
  xor g_10664_(out[132], out[308], _08436_);
  xor g_10665_(out[130], out[306], _08447_);
  and g_10666_(out[139], _07986_, _08458_);
  xor g_10667_(out[131], out[307], _08469_);
  xor g_10668_(out[134], out[310], _08480_);
  xor g_10669_(out[143], out[319], _08491_);
  xor g_10670_(out[138], out[314], _08502_);
  xor g_10671_(out[133], out[309], _08513_);
  xor g_10672_(out[128], out[304], _08524_);
  or g_10673_(_08382_, _08436_, _08535_);
  or g_10674_(_08393_, _08415_, _08546_);
  or g_10675_(_08447_, _08502_, _08557_);
  or g_10676_(_08546_, _08557_, _08568_);
  or g_10677_(_08425_, _08469_, _08579_);
  or g_10678_(_08513_, _08524_, _08590_);
  or g_10679_(_08579_, _08590_, _08601_);
  or g_10680_(_08568_, _08601_, _08612_);
  xor g_10681_(out[140], out[316], _08623_);
  or g_10682_(_08371_, _08623_, _08634_);
  or g_10683_(_08360_, _08480_, _08645_);
  or g_10684_(_08634_, _08645_, _08656_);
  or g_10685_(_08404_, _08458_, _08667_);
  or g_10686_(_08491_, _08667_, _08678_);
  or g_10687_(_08656_, _08678_, _08689_);
  or g_10688_(_08612_, _08689_, _08700_);
  or g_10689_(_08535_, _08700_, _08711_);
  xor g_10690_(out[122], out[314], _08722_);
  xor g_10691_(out[120], out[312], _08732_);
  xor g_10692_(out[113], out[305], _08743_);
  and g_10693_(_07843_, out[315], _08754_);
  and g_10694_(out[123], _07986_, _08765_);
  xor g_10695_(out[114], out[306], _08776_);
  xor g_10696_(out[117], out[309], _08787_);
  xor g_10697_(out[121], out[313], _08798_);
  xor g_10698_(out[124], out[316], _08809_);
  xor g_10699_(out[125], out[317], _08820_);
  xor g_10700_(out[127], out[319], _08831_);
  xor g_10701_(out[116], out[308], _08842_);
  xor g_10702_(out[118], out[310], _08853_);
  xor g_10703_(out[115], out[307], _08864_);
  xor g_10704_(out[112], out[304], _08875_);
  xor g_10705_(out[126], out[318], _08886_);
  or g_10706_(_08842_, _08886_, _08897_);
  or g_10707_(_08732_, _08820_, _08908_);
  or g_10708_(_08722_, _08776_, _08919_);
  or g_10709_(_08908_, _08919_, _08930_);
  or g_10710_(_08798_, _08864_, _08941_);
  or g_10711_(_08787_, _08875_, _08952_);
  or g_10712_(_08941_, _08952_, _08963_);
  or g_10713_(_08930_, _08963_, _08974_);
  or g_10714_(_08754_, _08809_, _08985_);
  xor g_10715_(out[119], out[311], _08996_);
  or g_10716_(_08853_, _08996_, _09007_);
  or g_10717_(_08985_, _09007_, _09018_);
  or g_10718_(_08743_, _08765_, _09029_);
  or g_10719_(_08831_, _09029_, _09040_);
  or g_10720_(_09018_, _09040_, _09050_);
  or g_10721_(_08974_, _09050_, _09061_);
  or g_10722_(_08897_, _09061_, _09072_);
  xor g_10723_(out[103], out[311], _09083_);
  and g_10724_(_07832_, out[315], _09094_);
  xor g_10725_(out[110], out[318], _09105_);
  xor g_10726_(out[104], out[312], _09116_);
  xor g_10727_(out[97], out[305], _09127_);
  xor g_10728_(out[109], out[317], _09138_);
  xor g_10729_(out[105], out[313], _09149_);
  xor g_10730_(out[100], out[308], _09160_);
  xor g_10731_(out[98], out[306], _09171_);
  and g_10732_(out[107], _07986_, _09182_);
  xor g_10733_(out[99], out[307], _09193_);
  xor g_10734_(out[102], out[310], _09204_);
  xor g_10735_(out[111], out[319], _09215_);
  xor g_10736_(out[106], out[314], _09226_);
  xor g_10737_(out[101], out[309], _09237_);
  xor g_10738_(out[96], out[304], _09248_);
  or g_10739_(_09105_, _09160_, _09259_);
  or g_10740_(_09116_, _09138_, _09270_);
  or g_10741_(_09171_, _09226_, _09281_);
  or g_10742_(_09270_, _09281_, _09292_);
  or g_10743_(_09149_, _09193_, _09303_);
  or g_10744_(_09237_, _09248_, _09314_);
  or g_10745_(_09303_, _09314_, _09325_);
  or g_10746_(_09292_, _09325_, _09335_);
  xor g_10747_(out[108], out[316], _09346_);
  or g_10748_(_09094_, _09346_, _09357_);
  or g_10749_(_09083_, _09204_, _09368_);
  or g_10750_(_09357_, _09368_, _09379_);
  or g_10751_(_09127_, _09182_, _09390_);
  or g_10752_(_09215_, _09390_, _09401_);
  or g_10753_(_09379_, _09401_, _09412_);
  or g_10754_(_09335_, _09412_, _09423_);
  or g_10755_(_09259_, _09423_, _09434_);
  xor g_10756_(out[81], out[305], _09445_);
  and g_10757_(out[91], _07986_, _09456_);
  xor g_10758_(out[89], out[313], _09467_);
  xor g_10759_(out[80], out[304], _09478_);
  xor g_10760_(out[94], out[318], _09489_);
  xor g_10761_(out[84], out[308], _09500_);
  or g_10762_(_09489_, _09500_, _09511_);
  xor g_10763_(out[93], out[317], _09522_);
  xor g_10764_(out[83], out[307], _09533_);
  and g_10765_(_07821_, out[315], _09544_);
  xor g_10766_(out[86], out[310], _09555_);
  xor g_10767_(out[90], out[314], _09566_);
  xor g_10768_(out[85], out[309], _09576_);
  xor g_10769_(out[95], out[319], _09587_);
  xor g_10770_(out[88], out[312], _09598_);
  or g_10771_(_09522_, _09598_, _09609_);
  xor g_10772_(out[82], out[306], _09620_);
  or g_10773_(_09566_, _09620_, _09631_);
  or g_10774_(_09609_, _09631_, _09642_);
  or g_10775_(_09467_, _09533_, _09653_);
  or g_10776_(_09576_, _09653_, _09664_);
  or g_10777_(_09642_, _09664_, _09675_);
  or g_10778_(_09511_, _09675_, _09686_);
  xor g_10779_(out[92], out[316], _09697_);
  or g_10780_(_09544_, _09697_, _09708_);
  xor g_10781_(out[87], out[311], _09719_);
  or g_10782_(_09555_, _09719_, _09730_);
  or g_10783_(_09708_, _09730_, _09740_);
  or g_10784_(_09445_, _09456_, _09751_);
  or g_10785_(_09587_, _09751_, _09762_);
  or g_10786_(_09740_, _09762_, _09773_);
  or g_10787_(_09478_, _09773_, _09784_);
  or g_10788_(_09686_, _09784_, _09790_);
  xor g_10789_(out[71], out[311], _09791_);
  and g_10790_(_07810_, out[315], _09792_);
  xor g_10791_(out[78], out[318], _09793_);
  xor g_10792_(out[72], out[312], _09794_);
  xor g_10793_(out[65], out[305], _09795_);
  xor g_10794_(out[77], out[317], _09796_);
  xor g_10795_(out[73], out[313], _09797_);
  xor g_10796_(out[68], out[308], _09798_);
  xor g_10797_(out[66], out[306], _09799_);
  and g_10798_(out[75], _07986_, _09800_);
  xor g_10799_(out[67], out[307], _09801_);
  xor g_10800_(out[70], out[310], _09802_);
  xor g_10801_(out[79], out[319], _09803_);
  xor g_10802_(out[74], out[314], _09804_);
  xor g_10803_(out[69], out[309], _09805_);
  xor g_10804_(out[64], out[304], _09806_);
  or g_10805_(_09793_, _09798_, _09807_);
  or g_10806_(_09794_, _09796_, _09808_);
  or g_10807_(_09799_, _09804_, _09809_);
  or g_10808_(_09808_, _09809_, _09810_);
  or g_10809_(_09797_, _09801_, _09811_);
  or g_10810_(_09805_, _09806_, _09812_);
  or g_10811_(_09811_, _09812_, _09813_);
  or g_10812_(_09810_, _09813_, _09814_);
  xor g_10813_(out[76], out[316], _09815_);
  or g_10814_(_09792_, _09815_, _09816_);
  or g_10815_(_09791_, _09802_, _09817_);
  or g_10816_(_09816_, _09817_, _09818_);
  or g_10817_(_09795_, _09800_, _09819_);
  or g_10818_(_09803_, _09819_, _09820_);
  or g_10819_(_09818_, _09820_, _09821_);
  or g_10820_(_09814_, _09821_, _09822_);
  or g_10821_(_09807_, _09822_, _09823_);
  not g_10822_(_09823_, _09824_);
  xor g_10823_(out[60], out[316], _09825_);
  and g_10824_(_07799_, out[315], _09826_);
  xor g_10825_(out[56], out[312], _09827_);
  xor g_10826_(out[54], out[310], _09828_);
  xor g_10827_(out[61], out[317], _09829_);
  xor g_10828_(out[62], out[318], _09830_);
  xor g_10829_(out[50], out[306], _09831_);
  xor g_10830_(out[57], out[313], _09832_);
  xor g_10831_(out[53], out[309], _09833_);
  xor g_10832_(out[49], out[305], _09834_);
  and g_10833_(out[59], _07986_, _09835_);
  or g_10834_(_09827_, _09829_, _09836_);
  xor g_10835_(out[63], out[319], _09837_);
  xor g_10836_(out[58], out[314], _09838_);
  xor g_10837_(out[52], out[308], _09839_);
  xor g_10838_(out[51], out[307], _09840_);
  xor g_10839_(out[48], out[304], _09841_);
  or g_10840_(_09831_, _09838_, _09842_);
  or g_10841_(_09836_, _09842_, _09843_);
  or g_10842_(_09832_, _09840_, _09844_);
  or g_10843_(_09833_, _09844_, _09845_);
  or g_10844_(_09843_, _09845_, _09846_);
  or g_10845_(_09830_, _09839_, _09847_);
  or g_10846_(_09846_, _09847_, _09848_);
  or g_10847_(_09825_, _09826_, _09849_);
  xor g_10848_(out[55], out[311], _09850_);
  or g_10849_(_09828_, _09850_, _09851_);
  or g_10850_(_09849_, _09851_, _09852_);
  or g_10851_(_09834_, _09835_, _09853_);
  or g_10852_(_09837_, _09853_, _09854_);
  or g_10853_(_09852_, _09854_, _09855_);
  or g_10854_(_09841_, _09855_, _09856_);
  or g_10855_(_09848_, _09856_, _09857_);
  not g_10856_(_09857_, _09858_);
  xor g_10857_(out[39], out[311], _09859_);
  and g_10858_(_07788_, out[315], _09860_);
  xor g_10859_(out[46], out[318], _09861_);
  xor g_10860_(out[40], out[312], _09862_);
  xor g_10861_(out[33], out[305], _09863_);
  xor g_10862_(out[45], out[317], _09864_);
  xor g_10863_(out[41], out[313], _09865_);
  xor g_10864_(out[36], out[308], _09866_);
  xor g_10865_(out[34], out[306], _09867_);
  and g_10866_(out[43], _07986_, _09868_);
  xor g_10867_(out[35], out[307], _09869_);
  xor g_10868_(out[38], out[310], _09870_);
  xor g_10869_(out[47], out[319], _09871_);
  xor g_10870_(out[42], out[314], _09872_);
  xor g_10871_(out[37], out[309], _09873_);
  xor g_10872_(out[32], out[304], _09874_);
  or g_10873_(_09861_, _09866_, _09875_);
  or g_10874_(_09862_, _09864_, _09876_);
  or g_10875_(_09867_, _09872_, _09877_);
  or g_10876_(_09876_, _09877_, _09878_);
  or g_10877_(_09865_, _09869_, _09879_);
  or g_10878_(_09873_, _09874_, _09880_);
  or g_10879_(_09879_, _09880_, _09881_);
  or g_10880_(_09878_, _09881_, _09882_);
  xor g_10881_(out[44], out[316], _09883_);
  or g_10882_(_09860_, _09883_, _09884_);
  or g_10883_(_09859_, _09870_, _09885_);
  or g_10884_(_09884_, _09885_, _09886_);
  or g_10885_(_09863_, _09868_, _09887_);
  or g_10886_(_09871_, _09887_, _09888_);
  or g_10887_(_09886_, _09888_, _09889_);
  or g_10888_(_09882_, _09889_, _09890_);
  or g_10889_(_09875_, _09890_, _09891_);
  xor g_10890_(out[17], out[305], _09892_);
  and g_10891_(out[27], _07986_, _09893_);
  xor g_10892_(out[25], out[313], _09894_);
  xor g_10893_(out[16], out[304], _09895_);
  xor g_10894_(out[30], out[318], _09896_);
  xor g_10895_(out[20], out[308], _09897_);
  or g_10896_(_09896_, _09897_, _09898_);
  xor g_10897_(out[29], out[317], _09899_);
  xor g_10898_(out[19], out[307], _09900_);
  and g_10899_(_07755_, out[315], _09901_);
  xor g_10900_(out[22], out[310], _09902_);
  xor g_10901_(out[26], out[314], _09903_);
  xor g_10902_(out[21], out[309], _09904_);
  xor g_10903_(out[31], out[319], _09905_);
  xor g_10904_(out[24], out[312], _09906_);
  or g_10905_(_09899_, _09906_, _09907_);
  xor g_10906_(out[18], out[306], _09908_);
  or g_10907_(_09903_, _09908_, _09909_);
  or g_10908_(_09907_, _09909_, _09910_);
  or g_10909_(_09894_, _09900_, _09911_);
  or g_10910_(_09904_, _09911_, _09912_);
  or g_10911_(_09910_, _09912_, _09913_);
  or g_10912_(_09898_, _09913_, _09914_);
  xor g_10913_(out[28], out[316], _09915_);
  or g_10914_(_09901_, _09915_, _09916_);
  xor g_10915_(out[23], out[311], _09917_);
  or g_10916_(_09902_, _09917_, _09918_);
  or g_10917_(_09916_, _09918_, _09919_);
  or g_10918_(_09892_, _09893_, _09920_);
  or g_10919_(_09905_, _09920_, _09921_);
  or g_10920_(_09919_, _09921_, _09922_);
  or g_10921_(_09895_, _09922_, _09923_);
  or g_10922_(_09914_, _09923_, _09924_);
  xor g_10923_(out[2], out[306], _09925_);
  xor g_10924_(out[0], out[304], _09926_);
  xor g_10925_(out[9], out[313], _09927_);
  xor g_10926_(out[8], out[312], _09928_);
  xor g_10927_(out[5], out[309], _09929_);
  xor g_10928_(out[14], out[318], _09930_);
  xor g_10929_(out[13], out[317], _09931_);
  xor g_10930_(out[15], out[319], _09932_);
  xor g_10931_(out[10], out[314], _09933_);
  xor g_10932_(out[6], out[310], _09934_);
  xor g_10933_(out[3], out[307], _09935_);
  and g_10934_(_07722_, out[315], _09936_);
  and g_10935_(out[11], _07986_, _09937_);
  xor g_10936_(out[4], out[308], _09938_);
  xor g_10937_(out[1], out[305], _09939_);
  or g_10938_(_09930_, _09938_, _09940_);
  or g_10939_(_09928_, _09931_, _09941_);
  or g_10940_(_09925_, _09933_, _09942_);
  or g_10941_(_09941_, _09942_, _09943_);
  or g_10942_(_09927_, _09935_, _09944_);
  or g_10943_(_09926_, _09929_, _09945_);
  or g_10944_(_09944_, _09945_, _09946_);
  or g_10945_(_09943_, _09946_, _09947_);
  xor g_10946_(out[12], out[316], _09948_);
  or g_10947_(_09936_, _09948_, _09949_);
  xor g_10948_(out[7], out[311], _09950_);
  or g_10949_(_09934_, _09950_, _09951_);
  or g_10950_(_09949_, _09951_, _09952_);
  or g_10951_(_09937_, _09939_, _09953_);
  or g_10952_(_09932_, _09953_, _09954_);
  or g_10953_(_09952_, _09954_, _09955_);
  or g_10954_(_09947_, _09955_, _09956_);
  or g_10955_(_09940_, _09956_, _09957_);
  xor g_10956_(out[151], out[295], _09958_);
  and g_10957_(_07876_, out[299], _09959_);
  xor g_10958_(out[158], out[302], _09960_);
  xor g_10959_(out[152], out[296], _09961_);
  xor g_10960_(out[145], out[289], _09962_);
  xor g_10961_(out[157], out[301], _09963_);
  xor g_10962_(out[153], out[297], _09964_);
  xor g_10963_(out[148], out[292], _09965_);
  xor g_10964_(out[146], out[290], _09966_);
  and g_10965_(out[155], _07964_, _09967_);
  xor g_10966_(out[147], out[291], _09968_);
  xor g_10967_(out[150], out[294], _09969_);
  xor g_10968_(out[159], out[303], _09970_);
  xor g_10969_(out[154], out[298], _09971_);
  xor g_10970_(out[149], out[293], _09972_);
  xor g_10971_(out[144], out[288], _09973_);
  or g_10972_(_09960_, _09965_, _09974_);
  or g_10973_(_09961_, _09963_, _09975_);
  or g_10974_(_09966_, _09971_, _09976_);
  or g_10975_(_09975_, _09976_, _09977_);
  or g_10976_(_09964_, _09968_, _09978_);
  or g_10977_(_09972_, _09973_, _09979_);
  or g_10978_(_09978_, _09979_, _09980_);
  or g_10979_(_09977_, _09980_, _09981_);
  xor g_10980_(out[156], out[300], _09982_);
  or g_10981_(_09959_, _09982_, _09983_);
  or g_10982_(_09958_, _09969_, _09984_);
  or g_10983_(_09983_, _09984_, _09985_);
  or g_10984_(_09962_, _09967_, _09986_);
  or g_10985_(_09970_, _09986_, _09987_);
  or g_10986_(_09985_, _09987_, _09988_);
  or g_10987_(_09981_, _09988_, _09989_);
  or g_10988_(_09974_, _09989_, _09990_);
  xor g_10989_(out[129], out[289], _09991_);
  and g_10990_(_07854_, out[299], _09992_);
  and g_10991_(out[139], _07964_, _09993_);
  xor g_10992_(out[137], out[297], _09994_);
  xor g_10993_(out[128], out[288], _09995_);
  xor g_10994_(out[142], out[302], _09996_);
  xor g_10995_(out[132], out[292], _09997_);
  or g_10996_(_09996_, _09997_, _09998_);
  xor g_10997_(out[141], out[301], _09999_);
  xor g_10998_(out[131], out[291], _10000_);
  xor g_10999_(out[140], out[300], _10001_);
  xor g_11000_(out[134], out[294], _10002_);
  xor g_11001_(out[138], out[298], _10003_);
  xor g_11002_(out[133], out[293], _10004_);
  xor g_11003_(out[143], out[303], _10005_);
  xor g_11004_(out[136], out[296], _10006_);
  or g_11005_(_09999_, _10006_, _10007_);
  xor g_11006_(out[130], out[290], _10008_);
  or g_11007_(_10003_, _10008_, _10009_);
  or g_11008_(_10007_, _10009_, _10010_);
  or g_11009_(_09994_, _10000_, _10011_);
  or g_11010_(_10004_, _10011_, _10012_);
  or g_11011_(_10010_, _10012_, _10013_);
  or g_11012_(_09998_, _10013_, _10014_);
  or g_11013_(_09992_, _10001_, _10015_);
  xor g_11014_(out[135], out[295], _10016_);
  or g_11015_(_10002_, _10016_, _10017_);
  or g_11016_(_10015_, _10017_, _10018_);
  or g_11017_(_09991_, _09993_, _10019_);
  or g_11018_(_10005_, _10019_, _10020_);
  or g_11019_(_10018_, _10020_, _10021_);
  or g_11020_(_09995_, _10021_, _10022_);
  or g_11021_(_10014_, _10022_, _10023_);
  xor g_11022_(out[119], out[295], _10024_);
  and g_11023_(_07843_, out[299], _10025_);
  xor g_11024_(out[126], out[302], _10026_);
  xor g_11025_(out[120], out[296], _10027_);
  xor g_11026_(out[113], out[289], _10028_);
  xor g_11027_(out[125], out[301], _10029_);
  xor g_11028_(out[121], out[297], _10030_);
  xor g_11029_(out[116], out[292], _10031_);
  xor g_11030_(out[114], out[290], _10032_);
  and g_11031_(out[123], _07964_, _10033_);
  xor g_11032_(out[115], out[291], _10034_);
  xor g_11033_(out[118], out[294], _10035_);
  xor g_11034_(out[127], out[303], _10036_);
  xor g_11035_(out[122], out[298], _10037_);
  xor g_11036_(out[117], out[293], _10038_);
  xor g_11037_(out[112], out[288], _10039_);
  or g_11038_(_10026_, _10031_, _10040_);
  or g_11039_(_10027_, _10029_, _10041_);
  or g_11040_(_10032_, _10037_, _10042_);
  or g_11041_(_10041_, _10042_, _10043_);
  or g_11042_(_10030_, _10034_, _10044_);
  or g_11043_(_10038_, _10039_, _10045_);
  or g_11044_(_10044_, _10045_, _10046_);
  or g_11045_(_10043_, _10046_, _10047_);
  xor g_11046_(out[124], out[300], _10048_);
  or g_11047_(_10025_, _10048_, _10049_);
  or g_11048_(_10024_, _10035_, _10050_);
  or g_11049_(_10049_, _10050_, _10051_);
  or g_11050_(_10028_, _10033_, _10052_);
  or g_11051_(_10036_, _10052_, _10053_);
  or g_11052_(_10051_, _10053_, _10054_);
  or g_11053_(_10047_, _10054_, _10055_);
  or g_11054_(_10040_, _10055_, _10056_);
  xor g_11055_(out[97], out[289], _10057_);
  and g_11056_(out[107], _07964_, _10058_);
  xor g_11057_(out[105], out[297], _10059_);
  xor g_11058_(out[96], out[288], _10060_);
  xor g_11059_(out[110], out[302], _10061_);
  xor g_11060_(out[100], out[292], _10062_);
  or g_11061_(_10061_, _10062_, _10063_);
  xor g_11062_(out[109], out[301], _10064_);
  xor g_11063_(out[99], out[291], _10065_);
  and g_11064_(_07832_, out[299], _10066_);
  xor g_11065_(out[102], out[294], _10067_);
  xor g_11066_(out[106], out[298], _10068_);
  xor g_11067_(out[101], out[293], _10069_);
  xor g_11068_(out[111], out[303], _10070_);
  xor g_11069_(out[104], out[296], _10071_);
  or g_11070_(_10064_, _10071_, _10072_);
  xor g_11071_(out[98], out[290], _10073_);
  or g_11072_(_10068_, _10073_, _10074_);
  or g_11073_(_10072_, _10074_, _10075_);
  or g_11074_(_10059_, _10065_, _10076_);
  or g_11075_(_10069_, _10076_, _10077_);
  or g_11076_(_10075_, _10077_, _10078_);
  or g_11077_(_10063_, _10078_, _10079_);
  xor g_11078_(out[108], out[300], _10080_);
  or g_11079_(_10066_, _10080_, _10081_);
  xor g_11080_(out[103], out[295], _10082_);
  or g_11081_(_10067_, _10082_, _10083_);
  or g_11082_(_10081_, _10083_, _10084_);
  or g_11083_(_10057_, _10058_, _10085_);
  or g_11084_(_10070_, _10085_, _10086_);
  or g_11085_(_10084_, _10086_, _10087_);
  or g_11086_(_10060_, _10087_, _10088_);
  or g_11087_(_10079_, _10088_, _10089_);
  xor g_11088_(out[87], out[295], _10090_);
  and g_11089_(_07821_, out[299], _10091_);
  xor g_11090_(out[94], out[302], _10092_);
  xor g_11091_(out[88], out[296], _10093_);
  xor g_11092_(out[81], out[289], _10094_);
  xor g_11093_(out[93], out[301], _10095_);
  xor g_11094_(out[89], out[297], _10096_);
  xor g_11095_(out[84], out[292], _10097_);
  xor g_11096_(out[82], out[290], _10098_);
  and g_11097_(out[91], _07964_, _10099_);
  xor g_11098_(out[83], out[291], _10100_);
  xor g_11099_(out[86], out[294], _10101_);
  xor g_11100_(out[95], out[303], _10102_);
  xor g_11101_(out[90], out[298], _10103_);
  xor g_11102_(out[85], out[293], _10104_);
  xor g_11103_(out[80], out[288], _10105_);
  or g_11104_(_10092_, _10097_, _10106_);
  or g_11105_(_10093_, _10095_, _10107_);
  or g_11106_(_10098_, _10103_, _10108_);
  or g_11107_(_10107_, _10108_, _10109_);
  or g_11108_(_10096_, _10100_, _10110_);
  or g_11109_(_10104_, _10105_, _10111_);
  or g_11110_(_10110_, _10111_, _10112_);
  or g_11111_(_10109_, _10112_, _10113_);
  xor g_11112_(out[92], out[300], _10114_);
  or g_11113_(_10091_, _10114_, _10115_);
  or g_11114_(_10090_, _10101_, _10116_);
  or g_11115_(_10115_, _10116_, _10117_);
  or g_11116_(_10094_, _10099_, _10118_);
  or g_11117_(_10102_, _10118_, _10119_);
  or g_11118_(_10117_, _10119_, _10120_);
  or g_11119_(_10113_, _10120_, _10121_);
  or g_11120_(_10106_, _10121_, _10122_);
  xor g_11121_(out[65], out[289], _10123_);
  and g_11122_(out[75], _07964_, _10124_);
  xor g_11123_(out[73], out[297], _10125_);
  xor g_11124_(out[64], out[288], _10126_);
  xor g_11125_(out[78], out[302], _10127_);
  xor g_11126_(out[68], out[292], _10128_);
  or g_11127_(_10127_, _10128_, _10129_);
  xor g_11128_(out[77], out[301], _10130_);
  xor g_11129_(out[67], out[291], _10131_);
  and g_11130_(_07810_, out[299], _10132_);
  xor g_11131_(out[70], out[294], _10133_);
  xor g_11132_(out[74], out[298], _10134_);
  xor g_11133_(out[69], out[293], _10135_);
  xor g_11134_(out[79], out[303], _10136_);
  xor g_11135_(out[72], out[296], _10137_);
  or g_11136_(_10130_, _10137_, _10138_);
  xor g_11137_(out[66], out[290], _10139_);
  or g_11138_(_10134_, _10139_, _10140_);
  or g_11139_(_10138_, _10140_, _10141_);
  or g_11140_(_10125_, _10131_, _10142_);
  or g_11141_(_10135_, _10142_, _10143_);
  or g_11142_(_10141_, _10143_, _10144_);
  or g_11143_(_10129_, _10144_, _10145_);
  xor g_11144_(out[76], out[300], _10146_);
  or g_11145_(_10132_, _10146_, _10147_);
  xor g_11146_(out[71], out[295], _10148_);
  or g_11147_(_10133_, _10148_, _10149_);
  or g_11148_(_10147_, _10149_, _10150_);
  or g_11149_(_10123_, _10124_, _10151_);
  or g_11150_(_10136_, _10151_, _10152_);
  or g_11151_(_10150_, _10152_, _10153_);
  or g_11152_(_10126_, _10153_, _10154_);
  or g_11153_(_10145_, _10154_, _10155_);
  xor g_11154_(out[55], out[295], _10156_);
  and g_11155_(_07799_, out[299], _10157_);
  xor g_11156_(out[62], out[302], _10158_);
  xor g_11157_(out[56], out[296], _10159_);
  xor g_11158_(out[49], out[289], _10160_);
  xor g_11159_(out[61], out[301], _10161_);
  xor g_11160_(out[57], out[297], _10162_);
  xor g_11161_(out[52], out[292], _10163_);
  xor g_11162_(out[50], out[290], _10164_);
  and g_11163_(out[59], _07964_, _10165_);
  xor g_11164_(out[51], out[291], _10166_);
  xor g_11165_(out[54], out[294], _10167_);
  xor g_11166_(out[63], out[303], _10168_);
  xor g_11167_(out[58], out[298], _10169_);
  xor g_11168_(out[53], out[293], _10170_);
  xor g_11169_(out[48], out[288], _10171_);
  or g_11170_(_10158_, _10163_, _10172_);
  or g_11171_(_10159_, _10161_, _10173_);
  or g_11172_(_10164_, _10169_, _10174_);
  or g_11173_(_10173_, _10174_, _10175_);
  or g_11174_(_10162_, _10166_, _10176_);
  or g_11175_(_10170_, _10171_, _10177_);
  or g_11176_(_10176_, _10177_, _10178_);
  or g_11177_(_10175_, _10178_, _10179_);
  xor g_11178_(out[60], out[300], _10180_);
  or g_11179_(_10157_, _10180_, _10181_);
  or g_11180_(_10156_, _10167_, _10182_);
  or g_11181_(_10181_, _10182_, _10183_);
  or g_11182_(_10160_, _10165_, _10184_);
  or g_11183_(_10168_, _10184_, _10185_);
  or g_11184_(_10183_, _10185_, _10186_);
  or g_11185_(_10179_, _10186_, _10187_);
  or g_11186_(_10172_, _10187_, _10188_);
  xor g_11187_(out[33], out[289], _10189_);
  and g_11188_(out[43], _07964_, _10190_);
  xor g_11189_(out[41], out[297], _10191_);
  xor g_11190_(out[32], out[288], _10192_);
  xor g_11191_(out[46], out[302], _10193_);
  xor g_11192_(out[36], out[292], _10194_);
  or g_11193_(_10193_, _10194_, _10195_);
  xor g_11194_(out[45], out[301], _10196_);
  xor g_11195_(out[35], out[291], _10197_);
  and g_11196_(_07788_, out[299], _10198_);
  xor g_11197_(out[38], out[294], _10199_);
  xor g_11198_(out[42], out[298], _10200_);
  xor g_11199_(out[37], out[293], _10201_);
  xor g_11200_(out[47], out[303], _10202_);
  xor g_11201_(out[40], out[296], _10203_);
  or g_11202_(_10196_, _10203_, _10204_);
  xor g_11203_(out[34], out[290], _10205_);
  or g_11204_(_10200_, _10205_, _10206_);
  or g_11205_(_10204_, _10206_, _10207_);
  or g_11206_(_10191_, _10197_, _10208_);
  or g_11207_(_10201_, _10208_, _10209_);
  or g_11208_(_10207_, _10209_, _10210_);
  or g_11209_(_10195_, _10210_, _10211_);
  xor g_11210_(out[44], out[300], _10212_);
  or g_11211_(_10198_, _10212_, _10213_);
  xor g_11212_(out[39], out[295], _10214_);
  or g_11213_(_10199_, _10214_, _10215_);
  or g_11214_(_10213_, _10215_, _10216_);
  or g_11215_(_10189_, _10190_, _10217_);
  or g_11216_(_10202_, _10217_, _10218_);
  or g_11217_(_10216_, _10218_, _10219_);
  or g_11218_(_10192_, _10219_, _10220_);
  or g_11219_(_10211_, _10220_, _10221_);
  xor g_11220_(out[23], out[295], _10222_);
  and g_11221_(_07755_, out[299], _10223_);
  xor g_11222_(out[30], out[302], _10224_);
  xor g_11223_(out[24], out[296], _10225_);
  xor g_11224_(out[17], out[289], _10226_);
  xor g_11225_(out[29], out[301], _10227_);
  xor g_11226_(out[25], out[297], _10228_);
  xor g_11227_(out[20], out[292], _10229_);
  xor g_11228_(out[18], out[290], _10230_);
  and g_11229_(out[27], _07964_, _10231_);
  xor g_11230_(out[19], out[291], _10232_);
  xor g_11231_(out[22], out[294], _10233_);
  xor g_11232_(out[31], out[303], _10234_);
  xor g_11233_(out[26], out[298], _10235_);
  xor g_11234_(out[21], out[293], _10236_);
  xor g_11235_(out[16], out[288], _10237_);
  or g_11236_(_10224_, _10229_, _10238_);
  or g_11237_(_10225_, _10227_, _10239_);
  or g_11238_(_10230_, _10235_, _10240_);
  or g_11239_(_10239_, _10240_, _10241_);
  or g_11240_(_10228_, _10232_, _10242_);
  or g_11241_(_10236_, _10237_, _10243_);
  or g_11242_(_10242_, _10243_, _10244_);
  or g_11243_(_10241_, _10244_, _10245_);
  xor g_11244_(out[28], out[300], _10246_);
  or g_11245_(_10223_, _10246_, _10247_);
  or g_11246_(_10222_, _10233_, _10248_);
  or g_11247_(_10247_, _10248_, _10249_);
  or g_11248_(_10226_, _10231_, _10250_);
  or g_11249_(_10234_, _10250_, _10251_);
  or g_11250_(_10249_, _10251_, _10252_);
  or g_11251_(_10245_, _10252_, _10253_);
  or g_11252_(_10238_, _10253_, _10254_);
  xor g_11253_(out[1], out[289], _10255_);
  and g_11254_(out[11], _07964_, _10256_);
  xor g_11255_(out[14], out[302], _10257_);
  xor g_11256_(out[3], out[291], _10258_);
  xor g_11257_(out[4], out[292], _10259_);
  xor g_11258_(out[2], out[290], _10260_);
  xor g_11259_(out[9], out[297], _10261_);
  xor g_11260_(out[0], out[288], _10262_);
  and g_11261_(_07722_, out[299], _10263_);
  xor g_11262_(out[6], out[294], _10264_);
  xor g_11263_(out[10], out[298], _10265_);
  xor g_11264_(out[5], out[293], _10266_);
  xor g_11265_(out[15], out[303], _10267_);
  xor g_11266_(out[13], out[301], _10268_);
  xor g_11267_(out[8], out[296], _05390_);
  or g_11268_(_10257_, _10259_, _05391_);
  or g_11269_(_10268_, _05390_, _05392_);
  or g_11270_(_10260_, _10265_, _05393_);
  or g_11271_(_05392_, _05393_, _05394_);
  or g_11272_(_10258_, _10261_, _05395_);
  or g_11273_(_10262_, _10266_, _05396_);
  or g_11274_(_05395_, _05396_, _05397_);
  or g_11275_(_05394_, _05397_, _05398_);
  xor g_11276_(out[12], out[300], _05399_);
  or g_11277_(_10263_, _05399_, _05400_);
  xor g_11278_(out[7], out[295], _05401_);
  or g_11279_(_10264_, _05401_, _05402_);
  or g_11280_(_05400_, _05402_, _05403_);
  or g_11281_(_10255_, _10256_, _05404_);
  or g_11282_(_10267_, _05404_, _05405_);
  or g_11283_(_05403_, _05405_, _05406_);
  or g_11284_(_05398_, _05406_, _05407_);
  or g_11285_(_05391_, _05407_, _05408_);
  not g_11286_(_05408_, _05409_);
  and g_11287_(out[155], _07953_, _05410_);
  xor g_11288_(out[148], out[276], _05411_);
  xor g_11289_(out[146], out[274], _05412_);
  xor g_11290_(out[153], out[281], _05413_);
  xor g_11291_(out[144], out[272], _05414_);
  xor g_11292_(out[147], out[275], _05415_);
  and g_11293_(_07876_, out[283], _05416_);
  xor g_11294_(out[154], out[282], _05417_);
  xor g_11295_(out[159], out[287], _05418_);
  xor g_11296_(out[150], out[278], _05419_);
  xor g_11297_(out[149], out[277], _05420_);
  xor g_11298_(out[157], out[285], _05421_);
  xor g_11299_(out[158], out[286], _05422_);
  xor g_11300_(out[152], out[280], _05423_);
  xor g_11301_(out[145], out[273], _05424_);
  or g_11302_(_05411_, _05422_, _05425_);
  or g_11303_(_05421_, _05423_, _05426_);
  or g_11304_(_05412_, _05417_, _05427_);
  or g_11305_(_05426_, _05427_, _05428_);
  or g_11306_(_05413_, _05415_, _05429_);
  or g_11307_(_05414_, _05420_, _05430_);
  or g_11308_(_05429_, _05430_, _05431_);
  or g_11309_(_05428_, _05431_, _05432_);
  xor g_11310_(out[156], out[284], _05433_);
  or g_11311_(_05416_, _05433_, _05434_);
  xor g_11312_(out[151], out[279], _05435_);
  or g_11313_(_05419_, _05435_, _05436_);
  or g_11314_(_05434_, _05436_, _05437_);
  or g_11315_(_05410_, _05424_, _05438_);
  or g_11316_(_05418_, _05438_, _05439_);
  or g_11317_(_05437_, _05439_, _05440_);
  or g_11318_(_05432_, _05440_, _05441_);
  or g_11319_(_05425_, _05441_, _05442_);
  xor g_11320_(out[135], out[279], _05443_);
  and g_11321_(_07854_, out[283], _05444_);
  xor g_11322_(out[142], out[286], _05445_);
  xor g_11323_(out[136], out[280], _05446_);
  xor g_11324_(out[129], out[273], _05447_);
  xor g_11325_(out[141], out[285], _05448_);
  xor g_11326_(out[137], out[281], _05449_);
  xor g_11327_(out[132], out[276], _05450_);
  xor g_11328_(out[130], out[274], _05451_);
  and g_11329_(out[139], _07953_, _05452_);
  xor g_11330_(out[131], out[275], _05453_);
  xor g_11331_(out[134], out[278], _05454_);
  xor g_11332_(out[143], out[287], _05455_);
  xor g_11333_(out[138], out[282], _05456_);
  xor g_11334_(out[133], out[277], _05457_);
  xor g_11335_(out[128], out[272], _05458_);
  or g_11336_(_05445_, _05450_, _05459_);
  or g_11337_(_05446_, _05448_, _05460_);
  or g_11338_(_05451_, _05456_, _05461_);
  or g_11339_(_05460_, _05461_, _05462_);
  or g_11340_(_05449_, _05453_, _05463_);
  or g_11341_(_05457_, _05458_, _05464_);
  or g_11342_(_05463_, _05464_, _05465_);
  or g_11343_(_05462_, _05465_, _05466_);
  xor g_11344_(out[140], out[284], _05467_);
  or g_11345_(_05444_, _05467_, _05468_);
  or g_11346_(_05443_, _05454_, _05469_);
  or g_11347_(_05468_, _05469_, _05470_);
  or g_11348_(_05447_, _05452_, _05471_);
  or g_11349_(_05455_, _05471_, _05472_);
  or g_11350_(_05470_, _05472_, _05473_);
  or g_11351_(_05466_, _05473_, _05474_);
  or g_11352_(_05459_, _05474_, _05475_);
  not g_11353_(_05475_, _05476_);
  xor g_11354_(out[113], out[273], _05477_);
  and g_11355_(out[123], _07953_, _05478_);
  xor g_11356_(out[121], out[281], _05479_);
  xor g_11357_(out[112], out[272], _05480_);
  xor g_11358_(out[126], out[286], _05481_);
  xor g_11359_(out[116], out[276], _05482_);
  or g_11360_(_05481_, _05482_, _05483_);
  xor g_11361_(out[125], out[285], _05484_);
  xor g_11362_(out[115], out[275], _05485_);
  and g_11363_(_07843_, out[283], _05486_);
  xor g_11364_(out[118], out[278], _05487_);
  xor g_11365_(out[122], out[282], _05488_);
  xor g_11366_(out[117], out[277], _05489_);
  xor g_11367_(out[127], out[287], _05490_);
  xor g_11368_(out[120], out[280], _05491_);
  or g_11369_(_05484_, _05491_, _05492_);
  xor g_11370_(out[114], out[274], _05493_);
  or g_11371_(_05488_, _05493_, _05494_);
  or g_11372_(_05492_, _05494_, _05495_);
  or g_11373_(_05479_, _05485_, _05496_);
  or g_11374_(_05489_, _05496_, _05497_);
  or g_11375_(_05495_, _05497_, _05498_);
  or g_11376_(_05483_, _05498_, _05499_);
  xor g_11377_(out[124], out[284], _05500_);
  or g_11378_(_05486_, _05500_, _05501_);
  xor g_11379_(out[119], out[279], _05502_);
  or g_11380_(_05487_, _05502_, _05503_);
  or g_11381_(_05501_, _05503_, _05504_);
  or g_11382_(_05477_, _05478_, _05505_);
  or g_11383_(_05490_, _05505_, _05506_);
  or g_11384_(_05504_, _05506_, _05507_);
  or g_11385_(_05480_, _05507_, _05508_);
  or g_11386_(_05499_, _05508_, _05509_);
  xor g_11387_(out[103], out[279], _05510_);
  and g_11388_(_07832_, out[283], _05511_);
  xor g_11389_(out[110], out[286], _05512_);
  xor g_11390_(out[104], out[280], _05513_);
  xor g_11391_(out[97], out[273], _05514_);
  xor g_11392_(out[109], out[285], _05515_);
  xor g_11393_(out[105], out[281], _05516_);
  xor g_11394_(out[100], out[276], _05517_);
  xor g_11395_(out[98], out[274], _05518_);
  and g_11396_(out[107], _07953_, _05519_);
  xor g_11397_(out[99], out[275], _05520_);
  xor g_11398_(out[102], out[278], _05521_);
  xor g_11399_(out[111], out[287], _05522_);
  xor g_11400_(out[106], out[282], _05523_);
  xor g_11401_(out[101], out[277], _05524_);
  xor g_11402_(out[96], out[272], _05525_);
  or g_11403_(_05512_, _05517_, _05526_);
  or g_11404_(_05513_, _05515_, _05527_);
  or g_11405_(_05518_, _05523_, _05528_);
  or g_11406_(_05527_, _05528_, _05529_);
  or g_11407_(_05516_, _05520_, _05530_);
  or g_11408_(_05524_, _05525_, _05531_);
  or g_11409_(_05530_, _05531_, _05532_);
  or g_11410_(_05529_, _05532_, _05533_);
  xor g_11411_(out[108], out[284], _05534_);
  or g_11412_(_05511_, _05534_, _05535_);
  or g_11413_(_05510_, _05521_, _05536_);
  or g_11414_(_05535_, _05536_, _05537_);
  or g_11415_(_05514_, _05519_, _05538_);
  or g_11416_(_05522_, _05538_, _05539_);
  or g_11417_(_05537_, _05539_, _05540_);
  or g_11418_(_05533_, _05540_, _05541_);
  or g_11419_(_05526_, _05541_, _05542_);
  xor g_11420_(out[90], out[282], _05543_);
  xor g_11421_(out[82], out[274], _05544_);
  xor g_11422_(out[81], out[273], _05545_);
  and g_11423_(_07821_, out[283], _05546_);
  and g_11424_(out[91], _07953_, _05547_);
  xor g_11425_(out[93], out[285], _05548_);
  xor g_11426_(out[83], out[275], _05549_);
  xor g_11427_(out[94], out[286], _05550_);
  xor g_11428_(out[92], out[284], _05551_);
  xor g_11429_(out[88], out[280], _05552_);
  xor g_11430_(out[95], out[287], _05553_);
  xor g_11431_(out[85], out[277], _05554_);
  xor g_11432_(out[86], out[278], _05555_);
  xor g_11433_(out[80], out[272], _05556_);
  xor g_11434_(out[84], out[276], _05557_);
  or g_11435_(_05548_, _05552_, _05558_);
  xor g_11436_(out[89], out[281], _05559_);
  or g_11437_(_05543_, _05544_, _05560_);
  or g_11438_(_05558_, _05560_, _05561_);
  or g_11439_(_05549_, _05559_, _05562_);
  or g_11440_(_05554_, _05562_, _05563_);
  or g_11441_(_05561_, _05563_, _05564_);
  or g_11442_(_05550_, _05557_, _05565_);
  or g_11443_(_05564_, _05565_, _05566_);
  or g_11444_(_05546_, _05551_, _05567_);
  xor g_11445_(out[87], out[279], _05568_);
  or g_11446_(_05555_, _05568_, _05569_);
  or g_11447_(_05567_, _05569_, _05570_);
  or g_11448_(_05545_, _05547_, _05571_);
  or g_11449_(_05553_, _05571_, _05572_);
  or g_11450_(_05570_, _05572_, _05573_);
  or g_11451_(_05556_, _05573_, _05574_);
  or g_11452_(_05566_, _05574_, _05575_);
  not g_11453_(_05575_, _05576_);
  xor g_11454_(out[71], out[279], _05577_);
  and g_11455_(_07810_, out[283], _05578_);
  xor g_11456_(out[78], out[286], _05579_);
  xor g_11457_(out[72], out[280], _05580_);
  xor g_11458_(out[65], out[273], _05581_);
  xor g_11459_(out[77], out[285], _05582_);
  xor g_11460_(out[73], out[281], _05583_);
  xor g_11461_(out[68], out[276], _05584_);
  xor g_11462_(out[66], out[274], _05585_);
  and g_11463_(out[75], _07953_, _05586_);
  xor g_11464_(out[67], out[275], _05587_);
  xor g_11465_(out[70], out[278], _05588_);
  xor g_11466_(out[79], out[287], _05589_);
  xor g_11467_(out[74], out[282], _05590_);
  xor g_11468_(out[69], out[277], _05591_);
  xor g_11469_(out[64], out[272], _05592_);
  or g_11470_(_05579_, _05584_, _05593_);
  or g_11471_(_05580_, _05582_, _05594_);
  or g_11472_(_05585_, _05590_, _05595_);
  or g_11473_(_05594_, _05595_, _05596_);
  or g_11474_(_05583_, _05587_, _05597_);
  or g_11475_(_05591_, _05592_, _05598_);
  or g_11476_(_05597_, _05598_, _05599_);
  or g_11477_(_05596_, _05599_, _05600_);
  xor g_11478_(out[76], out[284], _05601_);
  or g_11479_(_05578_, _05601_, _05602_);
  or g_11480_(_05577_, _05588_, _05603_);
  or g_11481_(_05602_, _05603_, _05604_);
  or g_11482_(_05581_, _05586_, _05605_);
  or g_11483_(_05589_, _05605_, _05606_);
  or g_11484_(_05604_, _05606_, _05607_);
  or g_11485_(_05600_, _05607_, _05608_);
  or g_11486_(_05593_, _05608_, _05609_);
  xor g_11487_(out[50], out[274], _05610_);
  xor g_11488_(out[48], out[272], _05611_);
  xor g_11489_(out[57], out[281], _05612_);
  xor g_11490_(out[56], out[280], _05613_);
  xor g_11491_(out[53], out[277], _05614_);
  xor g_11492_(out[62], out[286], _05615_);
  xor g_11493_(out[61], out[285], _05616_);
  xor g_11494_(out[63], out[287], _05617_);
  xor g_11495_(out[58], out[282], _05618_);
  xor g_11496_(out[54], out[278], _05619_);
  xor g_11497_(out[51], out[275], _05620_);
  and g_11498_(_07799_, out[283], _05621_);
  and g_11499_(out[59], _07953_, _05622_);
  xor g_11500_(out[52], out[276], _05623_);
  xor g_11501_(out[49], out[273], _05624_);
  or g_11502_(_05615_, _05623_, _05625_);
  or g_11503_(_05613_, _05616_, _05626_);
  or g_11504_(_05610_, _05618_, _05627_);
  or g_11505_(_05626_, _05627_, _05628_);
  or g_11506_(_05612_, _05620_, _05629_);
  or g_11507_(_05611_, _05614_, _05630_);
  or g_11508_(_05629_, _05630_, _05631_);
  or g_11509_(_05628_, _05631_, _05632_);
  xor g_11510_(out[60], out[284], _05633_);
  or g_11511_(_05621_, _05633_, _05634_);
  xor g_11512_(out[55], out[279], _05635_);
  or g_11513_(_05619_, _05635_, _05636_);
  or g_11514_(_05634_, _05636_, _05637_);
  or g_11515_(_05622_, _05624_, _05638_);
  or g_11516_(_05617_, _05638_, _05639_);
  or g_11517_(_05637_, _05639_, _05640_);
  or g_11518_(_05632_, _05640_, _05641_);
  or g_11519_(_05625_, _05641_, _05642_);
  xor g_11520_(out[39], out[279], _05643_);
  and g_11521_(_07788_, out[283], _05644_);
  xor g_11522_(out[46], out[286], _05645_);
  xor g_11523_(out[40], out[280], _05646_);
  xor g_11524_(out[33], out[273], _05647_);
  xor g_11525_(out[45], out[285], _05648_);
  xor g_11526_(out[41], out[281], _05649_);
  xor g_11527_(out[36], out[276], _05650_);
  xor g_11528_(out[34], out[274], _05651_);
  and g_11529_(out[43], _07953_, _05652_);
  xor g_11530_(out[35], out[275], _05653_);
  xor g_11531_(out[38], out[278], _05654_);
  xor g_11532_(out[47], out[287], _05655_);
  xor g_11533_(out[42], out[282], _05656_);
  xor g_11534_(out[37], out[277], _05657_);
  xor g_11535_(out[32], out[272], _05658_);
  or g_11536_(_05645_, _05650_, _05659_);
  or g_11537_(_05646_, _05648_, _05660_);
  or g_11538_(_05651_, _05656_, _05661_);
  or g_11539_(_05660_, _05661_, _05662_);
  or g_11540_(_05649_, _05653_, _05663_);
  or g_11541_(_05657_, _05658_, _05664_);
  or g_11542_(_05663_, _05664_, _05665_);
  or g_11543_(_05662_, _05665_, _05666_);
  xor g_11544_(out[44], out[284], _05667_);
  or g_11545_(_05644_, _05667_, _05668_);
  or g_11546_(_05643_, _05654_, _05669_);
  or g_11547_(_05668_, _05669_, _05670_);
  or g_11548_(_05647_, _05652_, _05671_);
  or g_11549_(_05655_, _05671_, _05672_);
  or g_11550_(_05670_, _05672_, _05673_);
  or g_11551_(_05666_, _05673_, _05674_);
  or g_11552_(_05659_, _05674_, _05675_);
  not g_11553_(_05675_, _05676_);
  xor g_11554_(out[17], out[273], _05677_);
  and g_11555_(out[27], _07953_, _05678_);
  xor g_11556_(out[30], out[286], _05679_);
  xor g_11557_(out[19], out[275], _05680_);
  xor g_11558_(out[20], out[276], _05681_);
  xor g_11559_(out[18], out[274], _05682_);
  xor g_11560_(out[25], out[281], _05683_);
  xor g_11561_(out[16], out[272], _05684_);
  and g_11562_(_07755_, out[283], _05685_);
  xor g_11563_(out[22], out[278], _05686_);
  xor g_11564_(out[26], out[282], _05687_);
  xor g_11565_(out[21], out[277], _05688_);
  xor g_11566_(out[31], out[287], _05689_);
  xor g_11567_(out[29], out[285], _05690_);
  xor g_11568_(out[24], out[280], _05691_);
  or g_11569_(_05679_, _05681_, _05692_);
  or g_11570_(_05690_, _05691_, _05693_);
  or g_11571_(_05682_, _05687_, _05694_);
  or g_11572_(_05693_, _05694_, _05695_);
  or g_11573_(_05680_, _05683_, _05696_);
  or g_11574_(_05684_, _05688_, _05697_);
  or g_11575_(_05696_, _05697_, _05698_);
  or g_11576_(_05695_, _05698_, _05699_);
  xor g_11577_(out[28], out[284], _05700_);
  or g_11578_(_05685_, _05700_, _05701_);
  xor g_11579_(out[23], out[279], _05702_);
  or g_11580_(_05686_, _05702_, _05703_);
  or g_11581_(_05701_, _05703_, _05704_);
  or g_11582_(_05677_, _05678_, _05705_);
  or g_11583_(_05689_, _05705_, _05706_);
  or g_11584_(_05704_, _05706_, _05707_);
  or g_11585_(_05699_, _05707_, _05708_);
  or g_11586_(_05692_, _05708_, _05709_);
  and g_11587_(out[11], _07953_, _05710_);
  and g_11588_(_07722_, out[283], _05711_);
  xor g_11589_(out[8], out[280], _05712_);
  xor g_11590_(out[15], out[287], _05713_);
  xor g_11591_(out[1], out[273], _05714_);
  xor g_11592_(out[2], out[274], _05715_);
  xor g_11593_(out[4], out[276], _05716_);
  xor g_11594_(out[5], out[277], _05717_);
  xor g_11595_(out[9], out[281], _05718_);
  xor g_11596_(out[3], out[275], _05719_);
  xor g_11597_(out[14], out[286], _05720_);
  xor g_11598_(out[0], out[272], _05721_);
  xor g_11599_(out[10], out[282], _05722_);
  xor g_11600_(out[13], out[285], _05723_);
  or g_11601_(_05712_, _05723_, _05724_);
  xor g_11602_(out[6], out[278], _05725_);
  or g_11603_(_05715_, _05722_, _05726_);
  or g_11604_(_05724_, _05726_, _05727_);
  or g_11605_(_05718_, _05719_, _05728_);
  or g_11606_(_05717_, _05728_, _05729_);
  or g_11607_(_05727_, _05729_, _05730_);
  or g_11608_(_05716_, _05720_, _05731_);
  or g_11609_(_05730_, _05731_, _05732_);
  xor g_11610_(out[12], out[284], _05733_);
  or g_11611_(_05711_, _05733_, _05734_);
  xor g_11612_(out[7], out[279], _05735_);
  or g_11613_(_05725_, _05735_, _05736_);
  or g_11614_(_05734_, _05736_, _05737_);
  or g_11615_(_05710_, _05714_, _05738_);
  or g_11616_(_05713_, _05738_, _05739_);
  or g_11617_(_05737_, _05739_, _05740_);
  or g_11618_(_05721_, _05740_, _05741_);
  or g_11619_(_05732_, _05741_, _05742_);
  xor g_11620_(out[151], out[263], _05743_);
  and g_11621_(_07876_, out[267], _05744_);
  xor g_11622_(out[158], out[270], _05745_);
  xor g_11623_(out[152], out[264], _05746_);
  xor g_11624_(out[145], out[257], _05747_);
  xor g_11625_(out[157], out[269], _05748_);
  xor g_11626_(out[153], out[265], _05749_);
  xor g_11627_(out[148], out[260], _05750_);
  xor g_11628_(out[146], out[258], _05751_);
  and g_11629_(out[155], _07942_, _05752_);
  xor g_11630_(out[147], out[259], _05753_);
  xor g_11631_(out[150], out[262], _05754_);
  xor g_11632_(out[159], out[271], _05755_);
  xor g_11633_(out[154], out[266], _05756_);
  xor g_11634_(out[149], out[261], _05757_);
  xor g_11635_(out[144], out[256], _05758_);
  or g_11636_(_05745_, _05750_, _05759_);
  or g_11637_(_05746_, _05748_, _05760_);
  or g_11638_(_05751_, _05756_, _05761_);
  or g_11639_(_05760_, _05761_, _05762_);
  or g_11640_(_05749_, _05753_, _05763_);
  or g_11641_(_05757_, _05758_, _05764_);
  or g_11642_(_05763_, _05764_, _05765_);
  or g_11643_(_05762_, _05765_, _05766_);
  xor g_11644_(out[156], out[268], _05767_);
  or g_11645_(_05744_, _05767_, _05768_);
  or g_11646_(_05743_, _05754_, _05769_);
  or g_11647_(_05768_, _05769_, _05770_);
  or g_11648_(_05747_, _05752_, _05771_);
  or g_11649_(_05755_, _05771_, _05772_);
  or g_11650_(_05770_, _05772_, _05773_);
  or g_11651_(_05766_, _05773_, _05774_);
  or g_11652_(_05759_, _05774_, _05775_);
  xor g_11653_(out[129], out[257], _05776_);
  and g_11654_(out[139], _07942_, _05777_);
  xor g_11655_(out[137], out[265], _05778_);
  xor g_11656_(out[128], out[256], _05779_);
  xor g_11657_(out[142], out[270], _05780_);
  xor g_11658_(out[132], out[260], _05781_);
  or g_11659_(_05780_, _05781_, _05782_);
  xor g_11660_(out[141], out[269], _05783_);
  xor g_11661_(out[131], out[259], _05784_);
  and g_11662_(_07854_, out[267], _05785_);
  xor g_11663_(out[134], out[262], _05786_);
  xor g_11664_(out[138], out[266], _05787_);
  xor g_11665_(out[133], out[261], _05788_);
  xor g_11666_(out[143], out[271], _05789_);
  xor g_11667_(out[136], out[264], _05790_);
  or g_11668_(_05783_, _05790_, _05791_);
  xor g_11669_(out[130], out[258], _05792_);
  or g_11670_(_05787_, _05792_, _05793_);
  or g_11671_(_05791_, _05793_, _05794_);
  or g_11672_(_05778_, _05784_, _05795_);
  or g_11673_(_05788_, _05795_, _05796_);
  or g_11674_(_05794_, _05796_, _05797_);
  or g_11675_(_05782_, _05797_, _05798_);
  xor g_11676_(out[140], out[268], _05799_);
  or g_11677_(_05785_, _05799_, _05800_);
  xor g_11678_(out[135], out[263], _05801_);
  or g_11679_(_05786_, _05801_, _05802_);
  or g_11680_(_05800_, _05802_, _05803_);
  or g_11681_(_05776_, _05777_, _05804_);
  or g_11682_(_05789_, _05804_, _05805_);
  or g_11683_(_05803_, _05805_, _05806_);
  or g_11684_(_05779_, _05806_, _05807_);
  or g_11685_(_05798_, _05807_, _05808_);
  xor g_11686_(out[119], out[263], _05809_);
  and g_11687_(_07843_, out[267], _05810_);
  xor g_11688_(out[126], out[270], _05811_);
  xor g_11689_(out[120], out[264], _05812_);
  xor g_11690_(out[113], out[257], _05813_);
  xor g_11691_(out[125], out[269], _05814_);
  xor g_11692_(out[121], out[265], _05815_);
  xor g_11693_(out[116], out[260], _05816_);
  xor g_11694_(out[114], out[258], _05817_);
  and g_11695_(out[123], _07942_, _05818_);
  xor g_11696_(out[115], out[259], _05819_);
  xor g_11697_(out[118], out[262], _05820_);
  xor g_11698_(out[127], out[271], _05821_);
  xor g_11699_(out[122], out[266], _05822_);
  xor g_11700_(out[117], out[261], _05823_);
  xor g_11701_(out[112], out[256], _05824_);
  or g_11702_(_05811_, _05816_, _05825_);
  or g_11703_(_05812_, _05814_, _05826_);
  or g_11704_(_05817_, _05822_, _05827_);
  or g_11705_(_05826_, _05827_, _05828_);
  or g_11706_(_05815_, _05819_, _05829_);
  or g_11707_(_05823_, _05824_, _05830_);
  or g_11708_(_05829_, _05830_, _05831_);
  or g_11709_(_05828_, _05831_, _05832_);
  xor g_11710_(out[124], out[268], _05833_);
  or g_11711_(_05810_, _05833_, _05834_);
  or g_11712_(_05809_, _05820_, _05835_);
  or g_11713_(_05834_, _05835_, _05836_);
  or g_11714_(_05813_, _05818_, _05837_);
  or g_11715_(_05821_, _05837_, _05838_);
  or g_11716_(_05836_, _05838_, _05839_);
  or g_11717_(_05832_, _05839_, _05840_);
  or g_11718_(_05825_, _05840_, _05841_);
  xor g_11719_(out[100], out[260], _05842_);
  xor g_11720_(out[108], out[268], _05843_);
  and g_11721_(_07832_, out[267], _05844_);
  xor g_11722_(out[106], out[266], _05845_);
  xor g_11723_(out[102], out[262], _05846_);
  xor g_11724_(out[101], out[261], _05847_);
  xor g_11725_(out[99], out[259], _05848_);
  xor g_11726_(out[109], out[269], _05849_);
  xor g_11727_(out[110], out[270], _05850_);
  xor g_11728_(out[97], out[257], _05851_);
  xor g_11729_(out[98], out[258], _05852_);
  and g_11730_(out[107], _07942_, _05853_);
  xor g_11731_(out[96], out[256], _05854_);
  xor g_11732_(out[111], out[271], _05855_);
  xor g_11733_(out[104], out[264], _05856_);
  or g_11734_(_05849_, _05856_, _05857_);
  xor g_11735_(out[105], out[265], _05858_);
  or g_11736_(_05845_, _05852_, _05859_);
  or g_11737_(_05857_, _05859_, _05860_);
  or g_11738_(_05848_, _05858_, _05861_);
  or g_11739_(_05847_, _05861_, _05862_);
  or g_11740_(_05860_, _05862_, _05863_);
  or g_11741_(_05842_, _05850_, _05864_);
  or g_11742_(_05863_, _05864_, _05865_);
  or g_11743_(_05843_, _05844_, _05866_);
  xor g_11744_(out[103], out[263], _05867_);
  or g_11745_(_05846_, _05867_, _05868_);
  or g_11746_(_05866_, _05868_, _05869_);
  or g_11747_(_05851_, _05853_, _05870_);
  or g_11748_(_05855_, _05870_, _05871_);
  or g_11749_(_05869_, _05871_, _05872_);
  or g_11750_(_05854_, _05872_, _05873_);
  or g_11751_(_05865_, _05873_, _05874_);
  xor g_11752_(out[87], out[263], _05875_);
  and g_11753_(_07821_, out[267], _05876_);
  xor g_11754_(out[94], out[270], _05877_);
  xor g_11755_(out[88], out[264], _05878_);
  xor g_11756_(out[81], out[257], _05879_);
  xor g_11757_(out[93], out[269], _05880_);
  xor g_11758_(out[89], out[265], _05881_);
  xor g_11759_(out[84], out[260], _05882_);
  xor g_11760_(out[82], out[258], _05883_);
  and g_11761_(out[91], _07942_, _05884_);
  xor g_11762_(out[83], out[259], _05885_);
  xor g_11763_(out[86], out[262], _05886_);
  xor g_11764_(out[95], out[271], _05887_);
  xor g_11765_(out[90], out[266], _05888_);
  xor g_11766_(out[85], out[261], _05889_);
  xor g_11767_(out[80], out[256], _05890_);
  or g_11768_(_05877_, _05882_, _05891_);
  or g_11769_(_05878_, _05880_, _05892_);
  or g_11770_(_05883_, _05888_, _05893_);
  or g_11771_(_05892_, _05893_, _05894_);
  or g_11772_(_05881_, _05885_, _05895_);
  or g_11773_(_05889_, _05890_, _05896_);
  or g_11774_(_05895_, _05896_, _05897_);
  or g_11775_(_05894_, _05897_, _05898_);
  xor g_11776_(out[92], out[268], _05899_);
  or g_11777_(_05876_, _05899_, _05900_);
  or g_11778_(_05875_, _05886_, _05901_);
  or g_11779_(_05900_, _05901_, _05902_);
  or g_11780_(_05879_, _05884_, _05903_);
  or g_11781_(_05887_, _05903_, _05904_);
  or g_11782_(_05902_, _05904_, _05905_);
  or g_11783_(_05898_, _05905_, _05906_);
  or g_11784_(_05891_, _05906_, _05907_);
  xor g_11785_(out[74], out[266], _05908_);
  xor g_11786_(out[66], out[258], _05909_);
  xor g_11787_(out[65], out[257], _05910_);
  and g_11788_(_07810_, out[267], _05911_);
  and g_11789_(out[75], _07942_, _05912_);
  xor g_11790_(out[77], out[269], _05913_);
  xor g_11791_(out[67], out[259], _05914_);
  xor g_11792_(out[78], out[270], _05915_);
  xor g_11793_(out[76], out[268], _05916_);
  xor g_11794_(out[72], out[264], _05917_);
  xor g_11795_(out[79], out[271], _05918_);
  xor g_11796_(out[69], out[261], _05919_);
  xor g_11797_(out[70], out[262], _05920_);
  xor g_11798_(out[64], out[256], _05921_);
  xor g_11799_(out[68], out[260], _05922_);
  or g_11800_(_05913_, _05917_, _05923_);
  xor g_11801_(out[73], out[265], _05924_);
  or g_11802_(_05908_, _05909_, _05925_);
  or g_11803_(_05923_, _05925_, _05926_);
  or g_11804_(_05914_, _05924_, _05927_);
  or g_11805_(_05919_, _05927_, _05928_);
  or g_11806_(_05926_, _05928_, _05929_);
  or g_11807_(_05915_, _05922_, _05930_);
  or g_11808_(_05929_, _05930_, _05931_);
  or g_11809_(_05911_, _05916_, _05932_);
  xor g_11810_(out[71], out[263], _05933_);
  or g_11811_(_05920_, _05933_, _05934_);
  or g_11812_(_05932_, _05934_, _05935_);
  or g_11813_(_05910_, _05912_, _05936_);
  or g_11814_(_05918_, _05936_, _05937_);
  or g_11815_(_05935_, _05937_, _05938_);
  or g_11816_(_05921_, _05938_, _05939_);
  or g_11817_(_05931_, _05939_, _05940_);
  not g_11818_(_05940_, _05941_);
  xor g_11819_(out[55], out[263], _05942_);
  and g_11820_(_07799_, out[267], _05943_);
  xor g_11821_(out[62], out[270], _05944_);
  xor g_11822_(out[56], out[264], _05945_);
  xor g_11823_(out[49], out[257], _05946_);
  xor g_11824_(out[61], out[269], _05947_);
  xor g_11825_(out[57], out[265], _05948_);
  xor g_11826_(out[52], out[260], _05949_);
  xor g_11827_(out[50], out[258], _05950_);
  and g_11828_(out[59], _07942_, _05951_);
  xor g_11829_(out[51], out[259], _05952_);
  xor g_11830_(out[54], out[262], _05953_);
  xor g_11831_(out[63], out[271], _05954_);
  xor g_11832_(out[58], out[266], _05955_);
  xor g_11833_(out[53], out[261], _05956_);
  xor g_11834_(out[48], out[256], _05957_);
  or g_11835_(_05944_, _05949_, _05958_);
  or g_11836_(_05945_, _05947_, _05959_);
  or g_11837_(_05950_, _05955_, _05960_);
  or g_11838_(_05959_, _05960_, _05961_);
  or g_11839_(_05948_, _05952_, _05962_);
  or g_11840_(_05956_, _05957_, _05963_);
  or g_11841_(_05962_, _05963_, _05964_);
  or g_11842_(_05961_, _05964_, _05965_);
  xor g_11843_(out[60], out[268], _05966_);
  or g_11844_(_05943_, _05966_, _05967_);
  or g_11845_(_05942_, _05953_, _05968_);
  or g_11846_(_05967_, _05968_, _05969_);
  or g_11847_(_05946_, _05951_, _05970_);
  or g_11848_(_05954_, _05970_, _05971_);
  or g_11849_(_05969_, _05971_, _05972_);
  or g_11850_(_05965_, _05972_, _05973_);
  or g_11851_(_05958_, _05973_, _05974_);
  not g_11852_(_05974_, _05975_);
  xor g_11853_(out[33], out[257], _05976_);
  and g_11854_(_07788_, out[267], _05977_);
  and g_11855_(out[43], _07942_, _05978_);
  xor g_11856_(out[40], out[264], _05979_);
  xor g_11857_(out[42], out[266], _05980_);
  xor g_11858_(out[34], out[258], _05981_);
  xor g_11859_(out[36], out[260], _05982_);
  xor g_11860_(out[45], out[269], _05983_);
  xor g_11861_(out[41], out[265], _05984_);
  xor g_11862_(out[35], out[259], _05985_);
  xor g_11863_(out[37], out[261], _05986_);
  xor g_11864_(out[46], out[270], _05987_);
  xor g_11865_(out[32], out[256], _05988_);
  xor g_11866_(out[47], out[271], _05989_);
  or g_11867_(_05979_, _05983_, _05990_);
  xor g_11868_(out[38], out[262], _05991_);
  or g_11869_(_05980_, _05981_, _05992_);
  or g_11870_(_05990_, _05992_, _05993_);
  or g_11871_(_05984_, _05985_, _05994_);
  or g_11872_(_05986_, _05994_, _05995_);
  or g_11873_(_05993_, _05995_, _05996_);
  or g_11874_(_05982_, _05987_, _05997_);
  or g_11875_(_05996_, _05997_, _05998_);
  xor g_11876_(out[44], out[268], _05999_);
  or g_11877_(_05977_, _05999_, _06000_);
  xor g_11878_(out[39], out[263], _06001_);
  or g_11879_(_05991_, _06001_, _06002_);
  or g_11880_(_06000_, _06002_, _06003_);
  or g_11881_(_05976_, _05978_, _06004_);
  or g_11882_(_05989_, _06004_, _06005_);
  or g_11883_(_06003_, _06005_, _06006_);
  or g_11884_(_05988_, _06006_, _06007_);
  or g_11885_(_05998_, _06007_, _06008_);
  xor g_11886_(out[23], out[263], _06009_);
  and g_11887_(_07755_, out[267], _06010_);
  xor g_11888_(out[30], out[270], _06011_);
  xor g_11889_(out[24], out[264], _06012_);
  xor g_11890_(out[17], out[257], _06013_);
  xor g_11891_(out[29], out[269], _06014_);
  xor g_11892_(out[25], out[265], _06015_);
  xor g_11893_(out[20], out[260], _06016_);
  xor g_11894_(out[18], out[258], _06017_);
  and g_11895_(out[27], _07942_, _06018_);
  xor g_11896_(out[19], out[259], _06019_);
  xor g_11897_(out[22], out[262], _06020_);
  xor g_11898_(out[31], out[271], _06021_);
  xor g_11899_(out[26], out[266], _06022_);
  xor g_11900_(out[21], out[261], _06023_);
  xor g_11901_(out[16], out[256], _06024_);
  or g_11902_(_06011_, _06016_, _06025_);
  or g_11903_(_06012_, _06014_, _06026_);
  or g_11904_(_06017_, _06022_, _06027_);
  or g_11905_(_06026_, _06027_, _06028_);
  or g_11906_(_06015_, _06019_, _06029_);
  or g_11907_(_06023_, _06024_, _06030_);
  or g_11908_(_06029_, _06030_, _06031_);
  or g_11909_(_06028_, _06031_, _06032_);
  xor g_11910_(out[28], out[268], _06033_);
  or g_11911_(_06010_, _06033_, _06034_);
  or g_11912_(_06009_, _06020_, _06035_);
  or g_11913_(_06034_, _06035_, _06036_);
  or g_11914_(_06013_, _06018_, _06037_);
  or g_11915_(_06021_, _06037_, _06038_);
  or g_11916_(_06036_, _06038_, _06039_);
  or g_11917_(_06032_, _06039_, _06040_);
  or g_11918_(_06025_, _06040_, _06041_);
  and g_11919_(out[11], _07942_, _06042_);
  and g_11920_(_07722_, out[267], _06043_);
  xor g_11921_(out[8], out[264], _06044_);
  xor g_11922_(out[15], out[271], _06045_);
  xor g_11923_(out[1], out[257], _06046_);
  xor g_11924_(out[2], out[258], _06047_);
  xor g_11925_(out[4], out[260], _06048_);
  xor g_11926_(out[5], out[261], _06049_);
  xor g_11927_(out[9], out[265], _06050_);
  xor g_11928_(out[3], out[259], _06051_);
  xor g_11929_(out[14], out[270], _06052_);
  xor g_11930_(out[0], out[256], _06053_);
  xor g_11931_(out[10], out[266], _06054_);
  xor g_11932_(out[13], out[269], _06055_);
  or g_11933_(_06044_, _06055_, _06056_);
  xor g_11934_(out[6], out[262], _06057_);
  or g_11935_(_06047_, _06054_, _06058_);
  or g_11936_(_06056_, _06058_, _06059_);
  or g_11937_(_06050_, _06051_, _06060_);
  or g_11938_(_06049_, _06060_, _06061_);
  or g_11939_(_06059_, _06061_, _06062_);
  or g_11940_(_06048_, _06052_, _06063_);
  or g_11941_(_06062_, _06063_, _06064_);
  xor g_11942_(out[12], out[268], _06065_);
  or g_11943_(_06043_, _06065_, _06066_);
  xor g_11944_(out[7], out[263], _06067_);
  or g_11945_(_06057_, _06067_, _06068_);
  or g_11946_(_06066_, _06068_, _06069_);
  or g_11947_(_06042_, _06046_, _06070_);
  or g_11948_(_06045_, _06070_, _06071_);
  or g_11949_(_06069_, _06071_, _06072_);
  or g_11950_(_06053_, _06072_, _06073_);
  or g_11951_(_06064_, _06073_, _06074_);
  xor g_11952_(out[146], out[242], _06075_);
  xor g_11953_(out[144], out[240], _06076_);
  xor g_11954_(out[153], out[249], _06077_);
  xor g_11955_(out[152], out[248], _06078_);
  xor g_11956_(out[149], out[245], _06079_);
  xor g_11957_(out[158], out[254], _06080_);
  xor g_11958_(out[157], out[253], _06081_);
  xor g_11959_(out[159], out[255], _06082_);
  xor g_11960_(out[154], out[250], _06083_);
  xor g_11961_(out[150], out[246], _06084_);
  xor g_11962_(out[147], out[243], _06085_);
  and g_11963_(_07876_, out[251], _06086_);
  and g_11964_(out[155], _07931_, _06087_);
  xor g_11965_(out[148], out[244], _06088_);
  xor g_11966_(out[145], out[241], _06089_);
  or g_11967_(_06080_, _06088_, _06090_);
  or g_11968_(_06078_, _06081_, _06091_);
  or g_11969_(_06075_, _06083_, _06092_);
  or g_11970_(_06091_, _06092_, _06093_);
  or g_11971_(_06077_, _06085_, _06094_);
  or g_11972_(_06076_, _06079_, _06095_);
  or g_11973_(_06094_, _06095_, _06096_);
  or g_11974_(_06093_, _06096_, _06097_);
  xor g_11975_(out[156], out[252], _06098_);
  or g_11976_(_06086_, _06098_, _06099_);
  xor g_11977_(out[151], out[247], _06100_);
  or g_11978_(_06084_, _06100_, _06101_);
  or g_11979_(_06099_, _06101_, _06102_);
  or g_11980_(_06087_, _06089_, _06103_);
  or g_11981_(_06082_, _06103_, _06104_);
  or g_11982_(_06102_, _06104_, _06105_);
  or g_11983_(_06097_, _06105_, _06106_);
  or g_11984_(_06090_, _06106_, _06107_);
  xor g_11985_(out[135], out[247], _06108_);
  and g_11986_(_07854_, out[251], _06109_);
  xor g_11987_(out[142], out[254], _06110_);
  xor g_11988_(out[136], out[248], _06111_);
  xor g_11989_(out[129], out[241], _06112_);
  xor g_11990_(out[141], out[253], _06113_);
  xor g_11991_(out[137], out[249], _06114_);
  xor g_11992_(out[132], out[244], _06115_);
  xor g_11993_(out[130], out[242], _06116_);
  and g_11994_(out[139], _07931_, _06117_);
  xor g_11995_(out[131], out[243], _06118_);
  xor g_11996_(out[134], out[246], _06119_);
  xor g_11997_(out[143], out[255], _06120_);
  xor g_11998_(out[138], out[250], _06121_);
  xor g_11999_(out[133], out[245], _06122_);
  xor g_12000_(out[128], out[240], _06123_);
  or g_12001_(_06110_, _06115_, _06124_);
  or g_12002_(_06111_, _06113_, _06125_);
  or g_12003_(_06116_, _06121_, _06126_);
  or g_12004_(_06125_, _06126_, _06127_);
  or g_12005_(_06114_, _06118_, _06128_);
  or g_12006_(_06122_, _06123_, _06129_);
  or g_12007_(_06128_, _06129_, _06130_);
  or g_12008_(_06127_, _06130_, _06131_);
  xor g_12009_(out[140], out[252], _06132_);
  or g_12010_(_06109_, _06132_, _06133_);
  or g_12011_(_06108_, _06119_, _06134_);
  or g_12012_(_06133_, _06134_, _06135_);
  or g_12013_(_06112_, _06117_, _06136_);
  or g_12014_(_06120_, _06136_, _06137_);
  or g_12015_(_06135_, _06137_, _06138_);
  or g_12016_(_06131_, _06138_, _06139_);
  or g_12017_(_06124_, _06139_, _06140_);
  not g_12018_(_06140_, _06141_);
  xor g_12019_(out[124], out[252], _06142_);
  and g_12020_(_07843_, out[251], _06143_);
  xor g_12021_(out[120], out[248], _06144_);
  xor g_12022_(out[118], out[246], _06145_);
  xor g_12023_(out[125], out[253], _06146_);
  xor g_12024_(out[126], out[254], _06147_);
  xor g_12025_(out[114], out[242], _06148_);
  xor g_12026_(out[121], out[249], _06149_);
  xor g_12027_(out[117], out[245], _06150_);
  xor g_12028_(out[113], out[241], _06151_);
  and g_12029_(out[123], _07931_, _06152_);
  or g_12030_(_06144_, _06146_, _06153_);
  xor g_12031_(out[127], out[255], _06154_);
  xor g_12032_(out[122], out[250], _06155_);
  xor g_12033_(out[116], out[244], _06156_);
  xor g_12034_(out[115], out[243], _06157_);
  xor g_12035_(out[112], out[240], _06158_);
  or g_12036_(_06148_, _06155_, _06159_);
  or g_12037_(_06153_, _06159_, _06160_);
  or g_12038_(_06149_, _06157_, _06161_);
  or g_12039_(_06150_, _06161_, _06162_);
  or g_12040_(_06160_, _06162_, _06163_);
  or g_12041_(_06147_, _06156_, _06164_);
  or g_12042_(_06163_, _06164_, _06165_);
  or g_12043_(_06142_, _06143_, _06166_);
  xor g_12044_(out[119], out[247], _06167_);
  or g_12045_(_06145_, _06167_, _06168_);
  or g_12046_(_06166_, _06168_, _06169_);
  or g_12047_(_06151_, _06152_, _06170_);
  or g_12048_(_06154_, _06170_, _06171_);
  or g_12049_(_06169_, _06171_, _06172_);
  or g_12050_(_06158_, _06172_, _06173_);
  or g_12051_(_06165_, _06173_, _06174_);
  not g_12052_(_06174_, _06175_);
  xor g_12053_(out[103], out[247], _06176_);
  and g_12054_(_07832_, out[251], _06177_);
  xor g_12055_(out[110], out[254], _06178_);
  xor g_12056_(out[104], out[248], _06179_);
  xor g_12057_(out[97], out[241], _06180_);
  xor g_12058_(out[109], out[253], _06181_);
  xor g_12059_(out[105], out[249], _06182_);
  xor g_12060_(out[100], out[244], _06183_);
  xor g_12061_(out[98], out[242], _06184_);
  and g_12062_(out[107], _07931_, _06185_);
  xor g_12063_(out[99], out[243], _06186_);
  xor g_12064_(out[102], out[246], _06187_);
  xor g_12065_(out[111], out[255], _06188_);
  xor g_12066_(out[106], out[250], _06189_);
  xor g_12067_(out[101], out[245], _06190_);
  xor g_12068_(out[96], out[240], _06191_);
  or g_12069_(_06178_, _06183_, _06192_);
  or g_12070_(_06179_, _06181_, _06193_);
  or g_12071_(_06184_, _06189_, _06194_);
  or g_12072_(_06193_, _06194_, _06195_);
  or g_12073_(_06182_, _06186_, _06196_);
  or g_12074_(_06190_, _06191_, _06197_);
  or g_12075_(_06196_, _06197_, _06198_);
  or g_12076_(_06195_, _06198_, _06199_);
  xor g_12077_(out[108], out[252], _06200_);
  or g_12078_(_06177_, _06200_, _06201_);
  or g_12079_(_06176_, _06187_, _06202_);
  or g_12080_(_06201_, _06202_, _06203_);
  or g_12081_(_06180_, _06185_, _06204_);
  or g_12082_(_06188_, _06204_, _06205_);
  or g_12083_(_06203_, _06205_, _06206_);
  or g_12084_(_06199_, _06206_, _06207_);
  or g_12085_(_06192_, _06207_, _06208_);
  not g_12086_(_06208_, _06209_);
  xor g_12087_(out[83], out[243], _06210_);
  xor g_12088_(out[84], out[244], _06211_);
  xor g_12089_(out[94], out[254], _06212_);
  xor g_12090_(out[82], out[242], _06213_);
  xor g_12091_(out[85], out[245], _06214_);
  xor g_12092_(out[89], out[249], _06215_);
  xor g_12093_(out[88], out[248], _06216_);
  xor g_12094_(out[95], out[255], _06217_);
  xor g_12095_(out[90], out[250], _06218_);
  xor g_12096_(out[86], out[246], _06219_);
  xor g_12097_(out[80], out[240], _06220_);
  and g_12098_(_07821_, out[251], _06221_);
  and g_12099_(out[91], _07931_, _06222_);
  xor g_12100_(out[93], out[253], _06223_);
  or g_12101_(_06216_, _06223_, _06224_);
  xor g_12102_(out[81], out[241], _06225_);
  or g_12103_(_06213_, _06218_, _06226_);
  or g_12104_(_06224_, _06226_, _06227_);
  or g_12105_(_06210_, _06215_, _06228_);
  or g_12106_(_06214_, _06228_, _06229_);
  or g_12107_(_06227_, _06229_, _06230_);
  or g_12108_(_06211_, _06212_, _06231_);
  or g_12109_(_06230_, _06231_, _06232_);
  xor g_12110_(out[92], out[252], _06233_);
  or g_12111_(_06221_, _06233_, _06234_);
  xor g_12112_(out[87], out[247], _06235_);
  or g_12113_(_06219_, _06235_, _06236_);
  or g_12114_(_06234_, _06236_, _06237_);
  or g_12115_(_06222_, _06225_, _06238_);
  or g_12116_(_06217_, _06238_, _06239_);
  or g_12117_(_06237_, _06239_, _06240_);
  or g_12118_(_06220_, _06240_, _06241_);
  or g_12119_(_06232_, _06241_, _06242_);
  not g_12120_(_06242_, _06243_);
  xor g_12121_(out[71], out[247], _06244_);
  and g_12122_(_07810_, out[251], _06245_);
  xor g_12123_(out[78], out[254], _06246_);
  xor g_12124_(out[72], out[248], _06247_);
  xor g_12125_(out[65], out[241], _06248_);
  xor g_12126_(out[77], out[253], _06249_);
  xor g_12127_(out[73], out[249], _06250_);
  xor g_12128_(out[68], out[244], _06251_);
  xor g_12129_(out[66], out[242], _06252_);
  and g_12130_(out[75], _07931_, _06253_);
  xor g_12131_(out[67], out[243], _06254_);
  xor g_12132_(out[70], out[246], _06255_);
  xor g_12133_(out[79], out[255], _06256_);
  xor g_12134_(out[74], out[250], _06257_);
  xor g_12135_(out[69], out[245], _06258_);
  xor g_12136_(out[64], out[240], _06259_);
  or g_12137_(_06246_, _06251_, _06260_);
  or g_12138_(_06247_, _06249_, _06261_);
  or g_12139_(_06252_, _06257_, _06262_);
  or g_12140_(_06261_, _06262_, _06263_);
  or g_12141_(_06250_, _06254_, _06264_);
  or g_12142_(_06258_, _06259_, _06265_);
  or g_12143_(_06264_, _06265_, _06266_);
  or g_12144_(_06263_, _06266_, _06267_);
  xor g_12145_(out[76], out[252], _06268_);
  or g_12146_(_06245_, _06268_, _06269_);
  or g_12147_(_06244_, _06255_, _06270_);
  or g_12148_(_06269_, _06270_, _06271_);
  or g_12149_(_06248_, _06253_, _06272_);
  or g_12150_(_06256_, _06272_, _06273_);
  or g_12151_(_06271_, _06273_, _06274_);
  or g_12152_(_06267_, _06274_, _06275_);
  or g_12153_(_06260_, _06275_, _06276_);
  xor g_12154_(out[60], out[252], _06277_);
  and g_12155_(_07799_, out[251], _06278_);
  xor g_12156_(out[61], out[253], _06279_);
  xor g_12157_(out[54], out[246], _06280_);
  xor g_12158_(out[56], out[248], _06281_);
  xor g_12159_(out[57], out[249], _06282_);
  xor g_12160_(out[62], out[254], _06283_);
  xor g_12161_(out[52], out[244], _06284_);
  or g_12162_(_06283_, _06284_, _06285_);
  xor g_12163_(out[53], out[245], _06286_);
  xor g_12164_(out[49], out[241], _06287_);
  and g_12165_(out[59], _07931_, _06288_);
  xor g_12166_(out[63], out[255], _06289_);
  xor g_12167_(out[58], out[250], _06290_);
  xor g_12168_(out[48], out[240], _06291_);
  xor g_12169_(out[50], out[242], _06292_);
  xor g_12170_(out[51], out[243], _06293_);
  or g_12171_(_06279_, _06281_, _06294_);
  or g_12172_(_06290_, _06292_, _06295_);
  or g_12173_(_06294_, _06295_, _06296_);
  or g_12174_(_06282_, _06293_, _06297_);
  or g_12175_(_06286_, _06291_, _06298_);
  or g_12176_(_06297_, _06298_, _06299_);
  or g_12177_(_06296_, _06299_, _06300_);
  or g_12178_(_06277_, _06278_, _06301_);
  xor g_12179_(out[55], out[247], _06302_);
  or g_12180_(_06280_, _06302_, _06303_);
  or g_12181_(_06301_, _06303_, _06304_);
  or g_12182_(_06287_, _06288_, _06305_);
  or g_12183_(_06289_, _06305_, _06306_);
  or g_12184_(_06304_, _06306_, _06307_);
  or g_12185_(_06300_, _06307_, _06308_);
  or g_12186_(_06285_, _06308_, _06309_);
  xor g_12187_(out[39], out[247], _06310_);
  and g_12188_(_07788_, out[251], _06311_);
  xor g_12189_(out[46], out[254], _06312_);
  xor g_12190_(out[40], out[248], _06313_);
  xor g_12191_(out[33], out[241], _06314_);
  xor g_12192_(out[45], out[253], _06315_);
  xor g_12193_(out[41], out[249], _06316_);
  xor g_12194_(out[36], out[244], _06317_);
  xor g_12195_(out[34], out[242], _06318_);
  and g_12196_(out[43], _07931_, _06319_);
  xor g_12197_(out[35], out[243], _06320_);
  xor g_12198_(out[38], out[246], _06321_);
  xor g_12199_(out[47], out[255], _06322_);
  xor g_12200_(out[42], out[250], _06323_);
  xor g_12201_(out[37], out[245], _06324_);
  xor g_12202_(out[32], out[240], _06325_);
  or g_12203_(_06312_, _06317_, _06326_);
  or g_12204_(_06313_, _06315_, _06327_);
  or g_12205_(_06318_, _06323_, _06328_);
  or g_12206_(_06327_, _06328_, _06329_);
  or g_12207_(_06316_, _06320_, _06330_);
  or g_12208_(_06324_, _06325_, _06331_);
  or g_12209_(_06330_, _06331_, _06332_);
  or g_12210_(_06329_, _06332_, _06333_);
  xor g_12211_(out[44], out[252], _06334_);
  or g_12212_(_06311_, _06334_, _06335_);
  or g_12213_(_06310_, _06321_, _06336_);
  or g_12214_(_06335_, _06336_, _06337_);
  or g_12215_(_06314_, _06319_, _06338_);
  or g_12216_(_06322_, _06338_, _06339_);
  or g_12217_(_06337_, _06339_, _06340_);
  or g_12218_(_06333_, _06340_, _06341_);
  or g_12219_(_06326_, _06341_, _06342_);
  not g_12220_(_06342_, _06343_);
  xor g_12221_(out[17], out[241], _06344_);
  and g_12222_(out[27], _07931_, _06345_);
  xor g_12223_(out[25], out[249], _06346_);
  xor g_12224_(out[16], out[240], _06347_);
  xor g_12225_(out[30], out[254], _06348_);
  xor g_12226_(out[20], out[244], _06349_);
  or g_12227_(_06348_, _06349_, _06350_);
  xor g_12228_(out[29], out[253], _06351_);
  xor g_12229_(out[19], out[243], _06352_);
  and g_12230_(_07755_, out[251], _06353_);
  xor g_12231_(out[22], out[246], _06354_);
  xor g_12232_(out[26], out[250], _06355_);
  xor g_12233_(out[21], out[245], _06356_);
  xor g_12234_(out[31], out[255], _06357_);
  xor g_12235_(out[24], out[248], _06358_);
  or g_12236_(_06351_, _06358_, _06359_);
  xor g_12237_(out[18], out[242], _06360_);
  or g_12238_(_06355_, _06360_, _06361_);
  or g_12239_(_06359_, _06361_, _06362_);
  or g_12240_(_06346_, _06352_, _06363_);
  or g_12241_(_06356_, _06363_, _06364_);
  or g_12242_(_06362_, _06364_, _06365_);
  or g_12243_(_06350_, _06365_, _06366_);
  xor g_12244_(out[28], out[252], _06367_);
  or g_12245_(_06353_, _06367_, _06368_);
  xor g_12246_(out[23], out[247], _06369_);
  or g_12247_(_06354_, _06369_, _06370_);
  or g_12248_(_06368_, _06370_, _06371_);
  or g_12249_(_06344_, _06345_, _06372_);
  or g_12250_(_06357_, _06372_, _06373_);
  or g_12251_(_06371_, _06373_, _06374_);
  or g_12252_(_06347_, _06374_, _06375_);
  or g_12253_(_06366_, _06375_, _06376_);
  xor g_12254_(out[8], out[248], _06377_);
  xor g_12255_(out[5], out[245], _06378_);
  xor g_12256_(out[3], out[243], _06379_);
  xor g_12257_(out[14], out[254], _06380_);
  xor g_12258_(out[13], out[253], _06381_);
  xor g_12259_(out[2], out[242], _06382_);
  xor g_12260_(out[9], out[249], _06383_);
  xor g_12261_(out[6], out[246], _06384_);
  xor g_12262_(out[15], out[255], _06385_);
  xor g_12263_(out[10], out[250], _06386_);
  xor g_12264_(out[4], out[244], _06387_);
  xor g_12265_(out[0], out[240], _06388_);
  and g_12266_(_07722_, out[251], _06389_);
  and g_12267_(out[11], _07931_, _06390_);
  or g_12268_(_06377_, _06381_, _06391_);
  xor g_12269_(out[1], out[241], _06392_);
  or g_12270_(_06382_, _06386_, _06393_);
  or g_12271_(_06391_, _06393_, _06394_);
  or g_12272_(_06379_, _06383_, _06395_);
  or g_12273_(_06378_, _06395_, _06396_);
  or g_12274_(_06394_, _06396_, _06397_);
  or g_12275_(_06380_, _06387_, _06398_);
  or g_12276_(_06397_, _06398_, _06399_);
  xor g_12277_(out[12], out[252], _06400_);
  or g_12278_(_06389_, _06400_, _06401_);
  xor g_12279_(out[7], out[247], _06402_);
  or g_12280_(_06384_, _06402_, _06403_);
  or g_12281_(_06401_, _06403_, _06404_);
  or g_12282_(_06390_, _06392_, _06405_);
  or g_12283_(_06385_, _06405_, _06406_);
  or g_12284_(_06404_, _06406_, _06407_);
  or g_12285_(_06388_, _06407_, _06408_);
  or g_12286_(_06399_, _06408_, _06409_);
  not g_12287_(_06409_, _06410_);
  xor g_12288_(out[151], out[231], _06411_);
  and g_12289_(_07876_, out[235], _06412_);
  xor g_12290_(out[158], out[238], _06413_);
  xor g_12291_(out[152], out[232], _06414_);
  xor g_12292_(out[145], out[225], _06415_);
  xor g_12293_(out[157], out[237], _06416_);
  xor g_12294_(out[153], out[233], _06417_);
  xor g_12295_(out[148], out[228], _06418_);
  xor g_12296_(out[146], out[226], _06419_);
  and g_12297_(out[155], _07920_, _06420_);
  xor g_12298_(out[147], out[227], _06421_);
  xor g_12299_(out[150], out[230], _06422_);
  xor g_12300_(out[159], out[239], _06423_);
  xor g_12301_(out[154], out[234], _06424_);
  xor g_12302_(out[149], out[229], _06425_);
  xor g_12303_(out[144], out[224], _06426_);
  or g_12304_(_06413_, _06418_, _06427_);
  or g_12305_(_06414_, _06416_, _06428_);
  or g_12306_(_06419_, _06424_, _06429_);
  or g_12307_(_06428_, _06429_, _06430_);
  or g_12308_(_06417_, _06421_, _06431_);
  or g_12309_(_06425_, _06426_, _06432_);
  or g_12310_(_06431_, _06432_, _06433_);
  or g_12311_(_06430_, _06433_, _06434_);
  xor g_12312_(out[156], out[236], _06435_);
  or g_12313_(_06412_, _06435_, _06436_);
  or g_12314_(_06411_, _06422_, _06437_);
  or g_12315_(_06436_, _06437_, _06438_);
  or g_12316_(_06415_, _06420_, _06439_);
  or g_12317_(_06423_, _06439_, _06440_);
  or g_12318_(_06438_, _06440_, _06441_);
  or g_12319_(_06434_, _06441_, _06442_);
  or g_12320_(_06427_, _06442_, _06443_);
  not g_12321_(_06443_, _06444_);
  xor g_12322_(out[131], out[227], _06445_);
  xor g_12323_(out[132], out[228], _06446_);
  xor g_12324_(out[142], out[238], _06447_);
  xor g_12325_(out[130], out[226], _06448_);
  xor g_12326_(out[133], out[229], _06449_);
  xor g_12327_(out[137], out[233], _06450_);
  xor g_12328_(out[136], out[232], _06451_);
  xor g_12329_(out[143], out[239], _06452_);
  xor g_12330_(out[138], out[234], _06453_);
  xor g_12331_(out[134], out[230], _06454_);
  xor g_12332_(out[128], out[224], _06455_);
  and g_12333_(_07854_, out[235], _06456_);
  and g_12334_(out[139], _07920_, _06457_);
  xor g_12335_(out[141], out[237], _06458_);
  or g_12336_(_06451_, _06458_, _06459_);
  xor g_12337_(out[129], out[225], _06460_);
  or g_12338_(_06448_, _06453_, _06461_);
  or g_12339_(_06459_, _06461_, _06462_);
  or g_12340_(_06445_, _06450_, _06463_);
  or g_12341_(_06449_, _06463_, _06464_);
  or g_12342_(_06462_, _06464_, _06465_);
  or g_12343_(_06446_, _06447_, _06466_);
  or g_12344_(_06465_, _06466_, _06467_);
  xor g_12345_(out[140], out[236], _06468_);
  or g_12346_(_06456_, _06468_, _06469_);
  xor g_12347_(out[135], out[231], _06470_);
  or g_12348_(_06454_, _06470_, _06471_);
  or g_12349_(_06469_, _06471_, _06472_);
  or g_12350_(_06457_, _06460_, _06473_);
  or g_12351_(_06452_, _06473_, _06474_);
  or g_12352_(_06472_, _06474_, _06475_);
  or g_12353_(_06455_, _06475_, _06476_);
  or g_12354_(_06467_, _06476_, _06477_);
  not g_12355_(_06477_, _06478_);
  xor g_12356_(out[119], out[231], _06479_);
  and g_12357_(_07843_, out[235], _06480_);
  xor g_12358_(out[126], out[238], _06481_);
  xor g_12359_(out[120], out[232], _06482_);
  xor g_12360_(out[113], out[225], _06483_);
  xor g_12361_(out[125], out[237], _06484_);
  xor g_12362_(out[121], out[233], _06485_);
  xor g_12363_(out[116], out[228], _06486_);
  xor g_12364_(out[114], out[226], _06487_);
  and g_12365_(out[123], _07920_, _06488_);
  xor g_12366_(out[115], out[227], _06489_);
  xor g_12367_(out[118], out[230], _06490_);
  xor g_12368_(out[127], out[239], _06491_);
  xor g_12369_(out[122], out[234], _06492_);
  xor g_12370_(out[117], out[229], _06493_);
  xor g_12371_(out[112], out[224], _06494_);
  or g_12372_(_06481_, _06486_, _06495_);
  or g_12373_(_06482_, _06484_, _06496_);
  or g_12374_(_06487_, _06492_, _06497_);
  or g_12375_(_06496_, _06497_, _06498_);
  or g_12376_(_06485_, _06489_, _06499_);
  or g_12377_(_06493_, _06494_, _06500_);
  or g_12378_(_06499_, _06500_, _06501_);
  or g_12379_(_06498_, _06501_, _06502_);
  xor g_12380_(out[124], out[236], _06503_);
  or g_12381_(_06480_, _06503_, _06504_);
  or g_12382_(_06479_, _06490_, _06505_);
  or g_12383_(_06504_, _06505_, _06506_);
  or g_12384_(_06483_, _06488_, _06507_);
  or g_12385_(_06491_, _06507_, _06508_);
  or g_12386_(_06506_, _06508_, _06509_);
  or g_12387_(_06502_, _06509_, _06510_);
  or g_12388_(_06495_, _06510_, _06511_);
  not g_12389_(_06511_, _06512_);
  xor g_12390_(out[97], out[225], _06513_);
  and g_12391_(out[107], _07920_, _06514_);
  xor g_12392_(out[105], out[233], _06515_);
  xor g_12393_(out[96], out[224], _06516_);
  xor g_12394_(out[110], out[238], _06517_);
  xor g_12395_(out[100], out[228], _06518_);
  or g_12396_(_06517_, _06518_, _06519_);
  xor g_12397_(out[109], out[237], _06520_);
  xor g_12398_(out[99], out[227], _06521_);
  and g_12399_(_07832_, out[235], _06522_);
  xor g_12400_(out[102], out[230], _06523_);
  xor g_12401_(out[106], out[234], _06524_);
  xor g_12402_(out[101], out[229], _06525_);
  xor g_12403_(out[111], out[239], _06526_);
  xor g_12404_(out[104], out[232], _06527_);
  or g_12405_(_06520_, _06527_, _06528_);
  xor g_12406_(out[98], out[226], _06529_);
  or g_12407_(_06524_, _06529_, _06530_);
  or g_12408_(_06528_, _06530_, _06531_);
  or g_12409_(_06515_, _06521_, _06532_);
  or g_12410_(_06525_, _06532_, _06533_);
  or g_12411_(_06531_, _06533_, _06534_);
  or g_12412_(_06519_, _06534_, _06535_);
  xor g_12413_(out[108], out[236], _06536_);
  or g_12414_(_06522_, _06536_, _06537_);
  xor g_12415_(out[103], out[231], _06538_);
  or g_12416_(_06523_, _06538_, _06539_);
  or g_12417_(_06537_, _06539_, _06540_);
  or g_12418_(_06513_, _06514_, _06541_);
  or g_12419_(_06526_, _06541_, _06542_);
  or g_12420_(_06540_, _06542_, _06543_);
  or g_12421_(_06516_, _06543_, _06544_);
  or g_12422_(_06535_, _06544_, _06545_);
  xor g_12423_(out[87], out[231], _06546_);
  and g_12424_(_07821_, out[235], _06547_);
  xor g_12425_(out[94], out[238], _06548_);
  xor g_12426_(out[88], out[232], _06549_);
  xor g_12427_(out[81], out[225], _06550_);
  xor g_12428_(out[93], out[237], _06551_);
  xor g_12429_(out[89], out[233], _06552_);
  xor g_12430_(out[84], out[228], _06553_);
  xor g_12431_(out[82], out[226], _06554_);
  and g_12432_(out[91], _07920_, _06555_);
  xor g_12433_(out[83], out[227], _06556_);
  xor g_12434_(out[86], out[230], _06557_);
  xor g_12435_(out[95], out[239], _06558_);
  xor g_12436_(out[90], out[234], _06559_);
  xor g_12437_(out[85], out[229], _06560_);
  xor g_12438_(out[80], out[224], _06561_);
  or g_12439_(_06548_, _06553_, _06562_);
  or g_12440_(_06549_, _06551_, _06563_);
  or g_12441_(_06554_, _06559_, _06564_);
  or g_12442_(_06563_, _06564_, _06565_);
  or g_12443_(_06552_, _06556_, _06566_);
  or g_12444_(_06560_, _06561_, _06567_);
  or g_12445_(_06566_, _06567_, _06568_);
  or g_12446_(_06565_, _06568_, _06569_);
  xor g_12447_(out[92], out[236], _06570_);
  or g_12448_(_06547_, _06570_, _06571_);
  or g_12449_(_06546_, _06557_, _06572_);
  or g_12450_(_06571_, _06572_, _06573_);
  or g_12451_(_06550_, _06555_, _06574_);
  or g_12452_(_06558_, _06574_, _06575_);
  or g_12453_(_06573_, _06575_, _06576_);
  or g_12454_(_06569_, _06576_, _06577_);
  or g_12455_(_06562_, _06577_, _06578_);
  and g_12456_(out[75], _07920_, _06579_);
  xor g_12457_(out[68], out[228], _06580_);
  xor g_12458_(out[78], out[238], _06581_);
  or g_12459_(_06580_, _06581_, _06582_);
  xor g_12460_(out[77], out[237], _06583_);
  xor g_12461_(out[67], out[227], _06584_);
  xor g_12462_(out[64], out[224], _06585_);
  and g_12463_(_07810_, out[235], _06586_);
  xor g_12464_(out[74], out[234], _06587_);
  xor g_12465_(out[79], out[239], _06588_);
  xor g_12466_(out[70], out[230], _06589_);
  xor g_12467_(out[69], out[229], _06590_);
  xor g_12468_(out[72], out[232], _06591_);
  or g_12469_(_06583_, _06591_, _06592_);
  xor g_12470_(out[66], out[226], _06593_);
  xor g_12471_(out[73], out[233], _06594_);
  xor g_12472_(out[65], out[225], _06595_);
  or g_12473_(_06587_, _06593_, _06596_);
  or g_12474_(_06592_, _06596_, _06597_);
  or g_12475_(_06584_, _06594_, _06598_);
  or g_12476_(_06590_, _06598_, _06599_);
  or g_12477_(_06597_, _06599_, _06600_);
  or g_12478_(_06582_, _06600_, _06601_);
  xor g_12479_(out[76], out[236], _06602_);
  or g_12480_(_06586_, _06602_, _06603_);
  xor g_12481_(out[71], out[231], _06604_);
  or g_12482_(_06589_, _06604_, _06605_);
  or g_12483_(_06603_, _06605_, _06606_);
  or g_12484_(_06579_, _06595_, _06607_);
  or g_12485_(_06588_, _06607_, _06608_);
  or g_12486_(_06606_, _06608_, _06609_);
  or g_12487_(_06585_, _06609_, _06610_);
  or g_12488_(_06601_, _06610_, _06611_);
  not g_12489_(_06611_, _06612_);
  xor g_12490_(out[55], out[231], _06613_);
  and g_12491_(_07799_, out[235], _06614_);
  xor g_12492_(out[62], out[238], _06615_);
  xor g_12493_(out[56], out[232], _06616_);
  xor g_12494_(out[49], out[225], _06617_);
  xor g_12495_(out[61], out[237], _06618_);
  xor g_12496_(out[57], out[233], _06619_);
  xor g_12497_(out[52], out[228], _06620_);
  xor g_12498_(out[50], out[226], _06621_);
  and g_12499_(out[59], _07920_, _06622_);
  xor g_12500_(out[51], out[227], _06623_);
  xor g_12501_(out[54], out[230], _06624_);
  xor g_12502_(out[63], out[239], _06625_);
  xor g_12503_(out[58], out[234], _06626_);
  xor g_12504_(out[53], out[229], _06627_);
  xor g_12505_(out[48], out[224], _06628_);
  or g_12506_(_06615_, _06620_, _06629_);
  or g_12507_(_06616_, _06618_, _06630_);
  or g_12508_(_06621_, _06626_, _06631_);
  or g_12509_(_06630_, _06631_, _06632_);
  or g_12510_(_06619_, _06623_, _06633_);
  or g_12511_(_06627_, _06628_, _06634_);
  or g_12512_(_06633_, _06634_, _06635_);
  or g_12513_(_06632_, _06635_, _06636_);
  xor g_12514_(out[60], out[236], _06637_);
  or g_12515_(_06614_, _06637_, _06638_);
  or g_12516_(_06613_, _06624_, _06639_);
  or g_12517_(_06638_, _06639_, _06640_);
  or g_12518_(_06617_, _06622_, _06641_);
  or g_12519_(_06625_, _06641_, _06642_);
  or g_12520_(_06640_, _06642_, _06643_);
  or g_12521_(_06636_, _06643_, _06644_);
  or g_12522_(_06629_, _06644_, _06645_);
  xor g_12523_(out[44], out[236], _06646_);
  and g_12524_(_07788_, out[235], _06647_);
  xor g_12525_(out[45], out[237], _06648_);
  xor g_12526_(out[38], out[230], _06649_);
  xor g_12527_(out[40], out[232], _06650_);
  xor g_12528_(out[41], out[233], _06651_);
  xor g_12529_(out[46], out[238], _06652_);
  xor g_12530_(out[36], out[228], _06653_);
  or g_12531_(_06652_, _06653_, _06654_);
  xor g_12532_(out[37], out[229], _06655_);
  xor g_12533_(out[33], out[225], _06656_);
  and g_12534_(out[43], _07920_, _06657_);
  xor g_12535_(out[47], out[239], _06658_);
  xor g_12536_(out[42], out[234], _06659_);
  xor g_12537_(out[32], out[224], _06660_);
  xor g_12538_(out[34], out[226], _06661_);
  xor g_12539_(out[35], out[227], _06662_);
  or g_12540_(_06648_, _06650_, _06663_);
  or g_12541_(_06659_, _06661_, _06664_);
  or g_12542_(_06663_, _06664_, _06665_);
  or g_12543_(_06651_, _06662_, _06666_);
  or g_12544_(_06655_, _06660_, _06667_);
  or g_12545_(_06666_, _06667_, _06668_);
  or g_12546_(_06665_, _06668_, _06669_);
  or g_12547_(_06646_, _06647_, _06670_);
  xor g_12548_(out[39], out[231], _06671_);
  or g_12549_(_06649_, _06671_, _06672_);
  or g_12550_(_06670_, _06672_, _06673_);
  or g_12551_(_06656_, _06657_, _06674_);
  or g_12552_(_06658_, _06674_, _06675_);
  or g_12553_(_06673_, _06675_, _06676_);
  or g_12554_(_06669_, _06676_, _06677_);
  or g_12555_(_06654_, _06677_, _06678_);
  not g_12556_(_06678_, _06679_);
  xor g_12557_(out[23], out[231], _06680_);
  and g_12558_(_07755_, out[235], _06681_);
  xor g_12559_(out[30], out[238], _06682_);
  xor g_12560_(out[24], out[232], _06683_);
  xor g_12561_(out[17], out[225], _06684_);
  xor g_12562_(out[29], out[237], _06685_);
  xor g_12563_(out[25], out[233], _06686_);
  xor g_12564_(out[20], out[228], _06687_);
  xor g_12565_(out[18], out[226], _06688_);
  and g_12566_(out[27], _07920_, _06689_);
  xor g_12567_(out[19], out[227], _06690_);
  xor g_12568_(out[22], out[230], _06691_);
  xor g_12569_(out[31], out[239], _06692_);
  xor g_12570_(out[26], out[234], _06693_);
  xor g_12571_(out[21], out[229], _06694_);
  xor g_12572_(out[16], out[224], _06695_);
  or g_12573_(_06682_, _06687_, _06696_);
  or g_12574_(_06683_, _06685_, _06697_);
  or g_12575_(_06688_, _06693_, _06698_);
  or g_12576_(_06697_, _06698_, _06699_);
  or g_12577_(_06686_, _06690_, _06700_);
  or g_12578_(_06694_, _06695_, _06701_);
  or g_12579_(_06700_, _06701_, _06702_);
  or g_12580_(_06699_, _06702_, _06703_);
  xor g_12581_(out[28], out[236], _06704_);
  or g_12582_(_06681_, _06704_, _06705_);
  or g_12583_(_06680_, _06691_, _06706_);
  or g_12584_(_06705_, _06706_, _06707_);
  or g_12585_(_06684_, _06689_, _06708_);
  or g_12586_(_06692_, _06708_, _06709_);
  or g_12587_(_06707_, _06709_, _06710_);
  or g_12588_(_06703_, _06710_, _06711_);
  or g_12589_(_06696_, _06711_, _06712_);
  not g_12590_(_06712_, _06713_);
  and g_12591_(out[11], _07920_, _06714_);
  and g_12592_(_07722_, out[235], _06715_);
  xor g_12593_(out[3], out[227], _06716_);
  xor g_12594_(out[1], out[225], _06717_);
  xor g_12595_(out[14], out[238], _06718_);
  xor g_12596_(out[5], out[229], _06719_);
  xor g_12597_(out[8], out[232], _06720_);
  xor g_12598_(out[10], out[234], _06721_);
  xor g_12599_(out[6], out[230], _06722_);
  xor g_12600_(out[4], out[228], _06723_);
  xor g_12601_(out[13], out[237], _06724_);
  xor g_12602_(out[15], out[239], _06725_);
  xor g_12603_(out[0], out[224], _06726_);
  xor g_12604_(out[2], out[226], _06727_);
  xor g_12605_(out[9], out[233], _06728_);
  or g_12606_(_06718_, _06723_, _06729_);
  or g_12607_(_06720_, _06724_, _06730_);
  or g_12608_(_06721_, _06727_, _06731_);
  or g_12609_(_06730_, _06731_, _06732_);
  or g_12610_(_06716_, _06728_, _06733_);
  or g_12611_(_06719_, _06726_, _06734_);
  or g_12612_(_06733_, _06734_, _06735_);
  or g_12613_(_06732_, _06735_, _06736_);
  xor g_12614_(out[12], out[236], _06737_);
  or g_12615_(_06715_, _06737_, _06738_);
  xor g_12616_(out[7], out[231], _06739_);
  or g_12617_(_06722_, _06739_, _06740_);
  or g_12618_(_06738_, _06740_, _06741_);
  or g_12619_(_06714_, _06717_, _06742_);
  or g_12620_(_06725_, _06742_, _06743_);
  or g_12621_(_06741_, _06743_, _06744_);
  or g_12622_(_06736_, _06744_, _06745_);
  or g_12623_(_06729_, _06745_, _06746_);
  xor g_12624_(out[145], out[209], _06747_);
  and g_12625_(out[155], _07909_, _06748_);
  xor g_12626_(out[153], out[217], _06749_);
  xor g_12627_(out[144], out[208], _06750_);
  xor g_12628_(out[158], out[222], _06751_);
  xor g_12629_(out[148], out[212], _06752_);
  or g_12630_(_06751_, _06752_, _06753_);
  xor g_12631_(out[157], out[221], _06754_);
  xor g_12632_(out[147], out[211], _06755_);
  and g_12633_(_07876_, out[219], _06756_);
  xor g_12634_(out[150], out[214], _06757_);
  xor g_12635_(out[154], out[218], _06758_);
  xor g_12636_(out[149], out[213], _06759_);
  xor g_12637_(out[159], out[223], _06760_);
  xor g_12638_(out[152], out[216], _06761_);
  or g_12639_(_06754_, _06761_, _06762_);
  xor g_12640_(out[146], out[210], _06763_);
  or g_12641_(_06758_, _06763_, _06764_);
  or g_12642_(_06762_, _06764_, _06765_);
  or g_12643_(_06749_, _06755_, _06766_);
  or g_12644_(_06759_, _06766_, _06767_);
  or g_12645_(_06765_, _06767_, _06768_);
  or g_12646_(_06753_, _06768_, _06769_);
  xor g_12647_(out[156], out[220], _06770_);
  or g_12648_(_06756_, _06770_, _06771_);
  xor g_12649_(out[151], out[215], _06772_);
  or g_12650_(_06757_, _06772_, _06773_);
  or g_12651_(_06771_, _06773_, _06774_);
  or g_12652_(_06747_, _06748_, _06775_);
  or g_12653_(_06760_, _06775_, _06776_);
  or g_12654_(_06774_, _06776_, _06777_);
  or g_12655_(_06750_, _06777_, _06778_);
  or g_12656_(_06769_, _06778_, _06779_);
  xor g_12657_(out[135], out[215], _06780_);
  and g_12658_(_07854_, out[219], _06781_);
  xor g_12659_(out[142], out[222], _06782_);
  xor g_12660_(out[136], out[216], _06783_);
  xor g_12661_(out[129], out[209], _06784_);
  xor g_12662_(out[141], out[221], _06785_);
  xor g_12663_(out[137], out[217], _06786_);
  xor g_12664_(out[132], out[212], _06787_);
  xor g_12665_(out[130], out[210], _06788_);
  and g_12666_(out[139], _07909_, _06789_);
  xor g_12667_(out[131], out[211], _06790_);
  xor g_12668_(out[134], out[214], _06791_);
  xor g_12669_(out[143], out[223], _06792_);
  xor g_12670_(out[138], out[218], _06793_);
  xor g_12671_(out[133], out[213], _06794_);
  xor g_12672_(out[128], out[208], _06795_);
  or g_12673_(_06782_, _06787_, _06796_);
  or g_12674_(_06783_, _06785_, _06797_);
  or g_12675_(_06788_, _06793_, _06798_);
  or g_12676_(_06797_, _06798_, _06799_);
  or g_12677_(_06786_, _06790_, _06800_);
  or g_12678_(_06794_, _06795_, _06801_);
  or g_12679_(_06800_, _06801_, _06802_);
  or g_12680_(_06799_, _06802_, _06803_);
  xor g_12681_(out[140], out[220], _06804_);
  or g_12682_(_06781_, _06804_, _06805_);
  or g_12683_(_06780_, _06791_, _06806_);
  or g_12684_(_06805_, _06806_, _06807_);
  or g_12685_(_06784_, _06789_, _06808_);
  or g_12686_(_06792_, _06808_, _06809_);
  or g_12687_(_06807_, _06809_, _06810_);
  or g_12688_(_06803_, _06810_, _06811_);
  or g_12689_(_06796_, _06811_, _06812_);
  not g_12690_(_06812_, _06813_);
  xor g_12691_(out[120], out[216], _06814_);
  xor g_12692_(out[117], out[213], _06815_);
  xor g_12693_(out[115], out[211], _06816_);
  xor g_12694_(out[126], out[222], _06817_);
  xor g_12695_(out[125], out[221], _06818_);
  xor g_12696_(out[114], out[210], _06819_);
  xor g_12697_(out[121], out[217], _06820_);
  xor g_12698_(out[118], out[214], _06821_);
  xor g_12699_(out[127], out[223], _06822_);
  xor g_12700_(out[122], out[218], _06823_);
  xor g_12701_(out[116], out[212], _06824_);
  xor g_12702_(out[112], out[208], _06825_);
  and g_12703_(_07843_, out[219], _06826_);
  and g_12704_(out[123], _07909_, _06827_);
  or g_12705_(_06814_, _06818_, _06828_);
  xor g_12706_(out[113], out[209], _06829_);
  or g_12707_(_06819_, _06823_, _06830_);
  or g_12708_(_06828_, _06830_, _06831_);
  or g_12709_(_06816_, _06820_, _06832_);
  or g_12710_(_06815_, _06832_, _06833_);
  or g_12711_(_06831_, _06833_, _06834_);
  or g_12712_(_06817_, _06824_, _06835_);
  or g_12713_(_06834_, _06835_, _06836_);
  xor g_12714_(out[124], out[220], _06837_);
  or g_12715_(_06826_, _06837_, _06838_);
  xor g_12716_(out[119], out[215], _06839_);
  or g_12717_(_06821_, _06839_, _06840_);
  or g_12718_(_06838_, _06840_, _06841_);
  or g_12719_(_06827_, _06829_, _06842_);
  or g_12720_(_06822_, _06842_, _06843_);
  or g_12721_(_06841_, _06843_, _06844_);
  or g_12722_(_06825_, _06844_, _06845_);
  or g_12723_(_06836_, _06845_, _06846_);
  not g_12724_(_06846_, _06847_);
  xor g_12725_(out[103], out[215], _06848_);
  and g_12726_(_07832_, out[219], _06849_);
  xor g_12727_(out[110], out[222], _06850_);
  xor g_12728_(out[104], out[216], _06851_);
  xor g_12729_(out[97], out[209], _06852_);
  xor g_12730_(out[109], out[221], _06853_);
  xor g_12731_(out[105], out[217], _06854_);
  xor g_12732_(out[100], out[212], _06855_);
  xor g_12733_(out[98], out[210], _06856_);
  and g_12734_(out[107], _07909_, _06857_);
  xor g_12735_(out[99], out[211], _06858_);
  xor g_12736_(out[102], out[214], _06859_);
  xor g_12737_(out[111], out[223], _06860_);
  xor g_12738_(out[106], out[218], _06861_);
  xor g_12739_(out[101], out[213], _06862_);
  xor g_12740_(out[96], out[208], _06863_);
  or g_12741_(_06850_, _06855_, _06864_);
  or g_12742_(_06851_, _06853_, _06865_);
  or g_12743_(_06856_, _06861_, _06866_);
  or g_12744_(_06865_, _06866_, _06867_);
  or g_12745_(_06854_, _06858_, _06868_);
  or g_12746_(_06862_, _06863_, _06869_);
  or g_12747_(_06868_, _06869_, _06870_);
  or g_12748_(_06867_, _06870_, _06871_);
  xor g_12749_(out[108], out[220], _06872_);
  or g_12750_(_06849_, _06872_, _06873_);
  or g_12751_(_06848_, _06859_, _06874_);
  or g_12752_(_06873_, _06874_, _06875_);
  or g_12753_(_06852_, _06857_, _06876_);
  or g_12754_(_06860_, _06876_, _06877_);
  or g_12755_(_06875_, _06877_, _06878_);
  or g_12756_(_06871_, _06878_, _06879_);
  or g_12757_(_06864_, _06879_, _06880_);
  not g_12758_(_06880_, _06881_);
  xor g_12759_(out[81], out[209], _06882_);
  and g_12760_(out[91], _07909_, _06883_);
  xor g_12761_(out[89], out[217], _06884_);
  xor g_12762_(out[80], out[208], _06885_);
  xor g_12763_(out[94], out[222], _06886_);
  xor g_12764_(out[84], out[212], _06887_);
  or g_12765_(_06886_, _06887_, _06888_);
  xor g_12766_(out[93], out[221], _06889_);
  xor g_12767_(out[83], out[211], _06890_);
  and g_12768_(_07821_, out[219], _06891_);
  xor g_12769_(out[86], out[214], _06892_);
  xor g_12770_(out[90], out[218], _06893_);
  xor g_12771_(out[85], out[213], _06894_);
  xor g_12772_(out[95], out[223], _06895_);
  xor g_12773_(out[88], out[216], _06896_);
  or g_12774_(_06889_, _06896_, _06897_);
  xor g_12775_(out[82], out[210], _06898_);
  or g_12776_(_06893_, _06898_, _06899_);
  or g_12777_(_06897_, _06899_, _06900_);
  or g_12778_(_06884_, _06890_, _06901_);
  or g_12779_(_06894_, _06901_, _06902_);
  or g_12780_(_06900_, _06902_, _06903_);
  or g_12781_(_06888_, _06903_, _06904_);
  xor g_12782_(out[92], out[220], _06905_);
  or g_12783_(_06891_, _06905_, _06906_);
  xor g_12784_(out[87], out[215], _06907_);
  or g_12785_(_06892_, _06907_, _06908_);
  or g_12786_(_06906_, _06908_, _06909_);
  or g_12787_(_06882_, _06883_, _06910_);
  or g_12788_(_06895_, _06910_, _06911_);
  or g_12789_(_06909_, _06911_, _06912_);
  or g_12790_(_06885_, _06912_, _06913_);
  or g_12791_(_06904_, _06913_, _06914_);
  not g_12792_(_06914_, _06915_);
  xor g_12793_(out[71], out[215], _06916_);
  and g_12794_(_07810_, out[219], _06917_);
  xor g_12795_(out[78], out[222], _06918_);
  xor g_12796_(out[72], out[216], _06919_);
  xor g_12797_(out[65], out[209], _06920_);
  xor g_12798_(out[77], out[221], _06921_);
  xor g_12799_(out[73], out[217], _06922_);
  xor g_12800_(out[68], out[212], _06923_);
  xor g_12801_(out[66], out[210], _06924_);
  and g_12802_(out[75], _07909_, _06925_);
  xor g_12803_(out[67], out[211], _06926_);
  xor g_12804_(out[70], out[214], _06927_);
  xor g_12805_(out[79], out[223], _06928_);
  xor g_12806_(out[74], out[218], _06929_);
  xor g_12807_(out[69], out[213], _06930_);
  xor g_12808_(out[64], out[208], _06931_);
  or g_12809_(_06918_, _06923_, _06932_);
  or g_12810_(_06919_, _06921_, _06933_);
  or g_12811_(_06924_, _06929_, _06934_);
  or g_12812_(_06933_, _06934_, _06935_);
  or g_12813_(_06922_, _06926_, _06936_);
  or g_12814_(_06930_, _06931_, _06937_);
  or g_12815_(_06936_, _06937_, _06938_);
  or g_12816_(_06935_, _06938_, _06939_);
  xor g_12817_(out[76], out[220], _06940_);
  or g_12818_(_06917_, _06940_, _06941_);
  or g_12819_(_06916_, _06927_, _06942_);
  or g_12820_(_06941_, _06942_, _06943_);
  or g_12821_(_06920_, _06925_, _06944_);
  or g_12822_(_06928_, _06944_, _06945_);
  or g_12823_(_06943_, _06945_, _06946_);
  or g_12824_(_06939_, _06946_, _06947_);
  or g_12825_(_06932_, _06947_, _06948_);
  and g_12826_(out[59], _07909_, _06949_);
  xor g_12827_(out[52], out[212], _06950_);
  xor g_12828_(out[50], out[210], _06951_);
  xor g_12829_(out[57], out[217], _06952_);
  xor g_12830_(out[48], out[208], _06953_);
  xor g_12831_(out[51], out[211], _06954_);
  and g_12832_(_07799_, out[219], _06955_);
  xor g_12833_(out[58], out[218], _06956_);
  xor g_12834_(out[63], out[223], _06957_);
  xor g_12835_(out[54], out[214], _06958_);
  xor g_12836_(out[53], out[213], _06959_);
  xor g_12837_(out[61], out[221], _06960_);
  xor g_12838_(out[62], out[222], _06961_);
  xor g_12839_(out[56], out[216], _06962_);
  xor g_12840_(out[49], out[209], _06963_);
  or g_12841_(_06950_, _06961_, _06964_);
  or g_12842_(_06960_, _06962_, _06965_);
  or g_12843_(_06951_, _06956_, _06966_);
  or g_12844_(_06965_, _06966_, _06967_);
  or g_12845_(_06952_, _06954_, _06968_);
  or g_12846_(_06953_, _06959_, _06969_);
  or g_12847_(_06968_, _06969_, _06970_);
  or g_12848_(_06967_, _06970_, _06971_);
  xor g_12849_(out[60], out[220], _06972_);
  or g_12850_(_06955_, _06972_, _06973_);
  xor g_12851_(out[55], out[215], _06974_);
  or g_12852_(_06958_, _06974_, _06975_);
  or g_12853_(_06973_, _06975_, _06976_);
  or g_12854_(_06949_, _06963_, _06977_);
  or g_12855_(_06957_, _06977_, _06978_);
  or g_12856_(_06976_, _06978_, _06979_);
  or g_12857_(_06971_, _06979_, _06980_);
  or g_12858_(_06964_, _06980_, _06981_);
  xor g_12859_(out[39], out[215], _06982_);
  and g_12860_(_07788_, out[219], _06983_);
  xor g_12861_(out[46], out[222], _06984_);
  xor g_12862_(out[40], out[216], _06985_);
  xor g_12863_(out[33], out[209], _06986_);
  xor g_12864_(out[45], out[221], _06987_);
  xor g_12865_(out[41], out[217], _06988_);
  xor g_12866_(out[36], out[212], _06989_);
  xor g_12867_(out[34], out[210], _06990_);
  and g_12868_(out[43], _07909_, _06991_);
  xor g_12869_(out[35], out[211], _06992_);
  xor g_12870_(out[38], out[214], _06993_);
  xor g_12871_(out[47], out[223], _06994_);
  xor g_12872_(out[42], out[218], _06995_);
  xor g_12873_(out[37], out[213], _06996_);
  xor g_12874_(out[32], out[208], _06997_);
  or g_12875_(_06984_, _06989_, _06998_);
  or g_12876_(_06985_, _06987_, _06999_);
  or g_12877_(_06990_, _06995_, _07000_);
  or g_12878_(_06999_, _07000_, _07001_);
  or g_12879_(_06988_, _06992_, _07002_);
  or g_12880_(_06996_, _06997_, _07003_);
  or g_12881_(_07002_, _07003_, _07004_);
  or g_12882_(_07001_, _07004_, _07005_);
  xor g_12883_(out[44], out[220], _07006_);
  or g_12884_(_06983_, _07006_, _07007_);
  or g_12885_(_06982_, _06993_, _07008_);
  or g_12886_(_07007_, _07008_, _07009_);
  or g_12887_(_06986_, _06991_, _07010_);
  or g_12888_(_06994_, _07010_, _07011_);
  or g_12889_(_07009_, _07011_, _07012_);
  or g_12890_(_07005_, _07012_, _07013_);
  or g_12891_(_06998_, _07013_, _07014_);
  xor g_12892_(out[17], out[209], _07015_);
  and g_12893_(out[27], _07909_, _07016_);
  xor g_12894_(out[30], out[222], _07017_);
  xor g_12895_(out[19], out[211], _07018_);
  xor g_12896_(out[20], out[212], _07019_);
  xor g_12897_(out[18], out[210], _07020_);
  xor g_12898_(out[25], out[217], _07021_);
  xor g_12899_(out[16], out[208], _07022_);
  and g_12900_(_07755_, out[219], _07023_);
  xor g_12901_(out[22], out[214], _07024_);
  xor g_12902_(out[26], out[218], _07025_);
  xor g_12903_(out[21], out[213], _07026_);
  xor g_12904_(out[31], out[223], _07027_);
  xor g_12905_(out[29], out[221], _07028_);
  xor g_12906_(out[24], out[216], _07029_);
  or g_12907_(_07017_, _07019_, _07030_);
  or g_12908_(_07028_, _07029_, _07031_);
  or g_12909_(_07020_, _07025_, _07032_);
  or g_12910_(_07031_, _07032_, _07033_);
  or g_12911_(_07018_, _07021_, _07034_);
  or g_12912_(_07022_, _07026_, _07035_);
  or g_12913_(_07034_, _07035_, _07036_);
  or g_12914_(_07033_, _07036_, _07037_);
  xor g_12915_(out[28], out[220], _07038_);
  or g_12916_(_07023_, _07038_, _07039_);
  xor g_12917_(out[23], out[215], _07040_);
  or g_12918_(_07024_, _07040_, _07041_);
  or g_12919_(_07039_, _07041_, _07042_);
  or g_12920_(_07015_, _07016_, _07043_);
  or g_12921_(_07027_, _07043_, _07044_);
  or g_12922_(_07042_, _07044_, _07045_);
  or g_12923_(_07037_, _07045_, _07046_);
  or g_12924_(_07030_, _07046_, _07047_);
  not g_12925_(_07047_, _07048_);
  xor g_12926_(out[1], out[209], _07049_);
  and g_12927_(_07722_, out[219], _07050_);
  and g_12928_(out[11], _07909_, _07051_);
  xor g_12929_(out[9], out[217], _07052_);
  xor g_12930_(out[0], out[208], _07053_);
  xor g_12931_(out[14], out[222], _07054_);
  xor g_12932_(out[4], out[212], _07055_);
  or g_12933_(_07054_, _07055_, _07056_);
  xor g_12934_(out[13], out[221], _07057_);
  xor g_12935_(out[3], out[211], _07058_);
  xor g_12936_(out[12], out[220], _07059_);
  xor g_12937_(out[6], out[214], _07060_);
  xor g_12938_(out[10], out[218], _07061_);
  xor g_12939_(out[5], out[213], _07062_);
  xor g_12940_(out[15], out[223], _07063_);
  xor g_12941_(out[8], out[216], _07064_);
  or g_12942_(_07057_, _07064_, _07065_);
  xor g_12943_(out[2], out[210], _07066_);
  or g_12944_(_07061_, _07066_, _07067_);
  or g_12945_(_07065_, _07067_, _07068_);
  or g_12946_(_07052_, _07058_, _07069_);
  or g_12947_(_07062_, _07069_, _07070_);
  or g_12948_(_07068_, _07070_, _07071_);
  or g_12949_(_07056_, _07071_, _07072_);
  or g_12950_(_07050_, _07059_, _07073_);
  xor g_12951_(out[7], out[215], _07074_);
  or g_12952_(_07060_, _07074_, _07075_);
  or g_12953_(_07073_, _07075_, _07076_);
  or g_12954_(_07049_, _07051_, _07077_);
  or g_12955_(_07063_, _07077_, _07078_);
  or g_12956_(_07076_, _07078_, _07079_);
  or g_12957_(_07053_, _07079_, _07080_);
  or g_12958_(_07072_, _07080_, _07081_);
  not g_12959_(_07081_, _07082_);
  xor g_12960_(out[151], out[199], _07083_);
  and g_12961_(_07876_, out[203], _07084_);
  xor g_12962_(out[158], out[206], _07085_);
  xor g_12963_(out[152], out[200], _07086_);
  xor g_12964_(out[145], out[193], _07087_);
  xor g_12965_(out[157], out[205], _07088_);
  xor g_12966_(out[153], out[201], _07089_);
  xor g_12967_(out[148], out[196], _07090_);
  xor g_12968_(out[146], out[194], _07091_);
  and g_12969_(out[155], _07898_, _07092_);
  xor g_12970_(out[147], out[195], _07093_);
  xor g_12971_(out[150], out[198], _07094_);
  xor g_12972_(out[159], out[207], _07095_);
  xor g_12973_(out[154], out[202], _07096_);
  xor g_12974_(out[149], out[197], _07097_);
  xor g_12975_(out[144], out[192], _07098_);
  or g_12976_(_07085_, _07090_, _07099_);
  or g_12977_(_07086_, _07088_, _07100_);
  or g_12978_(_07091_, _07096_, _07101_);
  or g_12979_(_07100_, _07101_, _07102_);
  or g_12980_(_07089_, _07093_, _07103_);
  or g_12981_(_07097_, _07098_, _07104_);
  or g_12982_(_07103_, _07104_, _07105_);
  or g_12983_(_07102_, _07105_, _07106_);
  xor g_12984_(out[156], out[204], _07107_);
  or g_12985_(_07084_, _07107_, _07108_);
  or g_12986_(_07083_, _07094_, _07109_);
  or g_12987_(_07108_, _07109_, _07110_);
  or g_12988_(_07087_, _07092_, _07111_);
  or g_12989_(_07095_, _07111_, _07112_);
  or g_12990_(_07110_, _07112_, _07113_);
  or g_12991_(_07106_, _07113_, _07114_);
  or g_12992_(_07099_, _07114_, _07115_);
  xor g_12993_(out[140], out[204], _07116_);
  and g_12994_(_07854_, out[203], _07117_);
  xor g_12995_(out[136], out[200], _07118_);
  xor g_12996_(out[134], out[198], _07119_);
  xor g_12997_(out[141], out[205], _07120_);
  xor g_12998_(out[142], out[206], _07121_);
  xor g_12999_(out[130], out[194], _07122_);
  xor g_13000_(out[137], out[201], _07123_);
  xor g_13001_(out[133], out[197], _07124_);
  xor g_13002_(out[129], out[193], _07125_);
  and g_13003_(out[139], _07898_, _07126_);
  or g_13004_(_07118_, _07120_, _07127_);
  xor g_13005_(out[143], out[207], _07128_);
  xor g_13006_(out[138], out[202], _07129_);
  xor g_13007_(out[132], out[196], _07130_);
  xor g_13008_(out[131], out[195], _07131_);
  xor g_13009_(out[128], out[192], _07132_);
  or g_13010_(_07122_, _07129_, _07133_);
  or g_13011_(_07127_, _07133_, _07134_);
  or g_13012_(_07123_, _07131_, _07135_);
  or g_13013_(_07124_, _07135_, _07136_);
  or g_13014_(_07134_, _07136_, _07137_);
  or g_13015_(_07121_, _07130_, _07138_);
  or g_13016_(_07137_, _07138_, _07139_);
  or g_13017_(_07116_, _07117_, _07140_);
  xor g_13018_(out[135], out[199], _07141_);
  or g_13019_(_07119_, _07141_, _07142_);
  or g_13020_(_07140_, _07142_, _07143_);
  or g_13021_(_07125_, _07126_, _07144_);
  or g_13022_(_07128_, _07144_, _07145_);
  or g_13023_(_07143_, _07145_, _07146_);
  or g_13024_(_07132_, _07146_, _07147_);
  or g_13025_(_07139_, _07147_, _07148_);
  xor g_13026_(out[119], out[199], _07149_);
  and g_13027_(_07843_, out[203], _07150_);
  xor g_13028_(out[126], out[206], _07151_);
  xor g_13029_(out[120], out[200], _07152_);
  xor g_13030_(out[113], out[193], _07153_);
  xor g_13031_(out[125], out[205], _07154_);
  xor g_13032_(out[121], out[201], _07155_);
  xor g_13033_(out[116], out[196], _07156_);
  xor g_13034_(out[114], out[194], _07157_);
  and g_13035_(out[123], _07898_, _07158_);
  xor g_13036_(out[115], out[195], _07159_);
  xor g_13037_(out[118], out[198], _07160_);
  xor g_13038_(out[127], out[207], _07161_);
  xor g_13039_(out[122], out[202], _07162_);
  xor g_13040_(out[117], out[197], _07163_);
  xor g_13041_(out[112], out[192], _07164_);
  or g_13042_(_07151_, _07156_, _07165_);
  or g_13043_(_07152_, _07154_, _07166_);
  or g_13044_(_07157_, _07162_, _07167_);
  or g_13045_(_07166_, _07167_, _07168_);
  or g_13046_(_07155_, _07159_, _07169_);
  or g_13047_(_07163_, _07164_, _07170_);
  or g_13048_(_07169_, _07170_, _07171_);
  or g_13049_(_07168_, _07171_, _07172_);
  xor g_13050_(out[124], out[204], _07173_);
  or g_13051_(_07150_, _07173_, _07174_);
  or g_13052_(_07149_, _07160_, _07175_);
  or g_13053_(_07174_, _07175_, _07176_);
  or g_13054_(_07153_, _07158_, _07177_);
  or g_13055_(_07161_, _07177_, _07178_);
  or g_13056_(_07176_, _07178_, _07179_);
  or g_13057_(_07172_, _07179_, _07180_);
  or g_13058_(_07165_, _07180_, _07181_);
  not g_13059_(_07181_, _07182_);
  xor g_13060_(out[97], out[193], _07183_);
  and g_13061_(out[107], _07898_, _07184_);
  xor g_13062_(out[105], out[201], _07185_);
  xor g_13063_(out[96], out[192], _07186_);
  xor g_13064_(out[110], out[206], _07187_);
  xor g_13065_(out[100], out[196], _07188_);
  or g_13066_(_07187_, _07188_, _07189_);
  xor g_13067_(out[109], out[205], _07190_);
  xor g_13068_(out[99], out[195], _07191_);
  and g_13069_(_07832_, out[203], _07192_);
  xor g_13070_(out[102], out[198], _07193_);
  xor g_13071_(out[106], out[202], _07194_);
  xor g_13072_(out[101], out[197], _07195_);
  xor g_13073_(out[111], out[207], _07196_);
  xor g_13074_(out[104], out[200], _07197_);
  or g_13075_(_07190_, _07197_, _07198_);
  xor g_13076_(out[98], out[194], _07199_);
  or g_13077_(_07194_, _07199_, _07200_);
  or g_13078_(_07198_, _07200_, _07201_);
  or g_13079_(_07185_, _07191_, _07202_);
  or g_13080_(_07195_, _07202_, _07203_);
  or g_13081_(_07201_, _07203_, _07204_);
  or g_13082_(_07189_, _07204_, _07205_);
  xor g_13083_(out[108], out[204], _07206_);
  or g_13084_(_07192_, _07206_, _07207_);
  xor g_13085_(out[103], out[199], _07208_);
  or g_13086_(_07193_, _07208_, _07209_);
  or g_13087_(_07207_, _07209_, _07210_);
  or g_13088_(_07183_, _07184_, _07211_);
  or g_13089_(_07196_, _07211_, _07212_);
  or g_13090_(_07210_, _07212_, _07213_);
  or g_13091_(_07186_, _07213_, _07214_);
  or g_13092_(_07205_, _07214_, _07215_);
  xor g_13093_(out[87], out[199], _07216_);
  and g_13094_(_07821_, out[203], _07217_);
  xor g_13095_(out[94], out[206], _07218_);
  xor g_13096_(out[88], out[200], _07219_);
  xor g_13097_(out[81], out[193], _07220_);
  xor g_13098_(out[93], out[205], _07221_);
  xor g_13099_(out[89], out[201], _07222_);
  xor g_13100_(out[84], out[196], _07223_);
  xor g_13101_(out[82], out[194], _07224_);
  and g_13102_(out[91], _07898_, _07225_);
  xor g_13103_(out[83], out[195], _07226_);
  xor g_13104_(out[86], out[198], _07227_);
  xor g_13105_(out[95], out[207], _07228_);
  xor g_13106_(out[90], out[202], _07229_);
  xor g_13107_(out[85], out[197], _07230_);
  xor g_13108_(out[80], out[192], _07231_);
  or g_13109_(_07218_, _07223_, _07232_);
  or g_13110_(_07219_, _07221_, _07233_);
  or g_13111_(_07224_, _07229_, _07234_);
  or g_13112_(_07233_, _07234_, _07235_);
  or g_13113_(_07222_, _07226_, _07236_);
  or g_13114_(_07230_, _07231_, _07237_);
  or g_13115_(_07236_, _07237_, _07238_);
  or g_13116_(_07235_, _07238_, _07239_);
  xor g_13117_(out[92], out[204], _07240_);
  or g_13118_(_07217_, _07240_, _07241_);
  or g_13119_(_07216_, _07227_, _07242_);
  or g_13120_(_07241_, _07242_, _07243_);
  or g_13121_(_07220_, _07225_, _07244_);
  or g_13122_(_07228_, _07244_, _07245_);
  or g_13123_(_07243_, _07245_, _07246_);
  or g_13124_(_07239_, _07246_, _07247_);
  or g_13125_(_07232_, _07247_, _07248_);
  xor g_13126_(out[74], out[202], _07249_);
  xor g_13127_(out[72], out[200], _07250_);
  xor g_13128_(out[65], out[193], _07251_);
  and g_13129_(_07810_, out[203], _07252_);
  and g_13130_(out[75], _07898_, _07253_);
  xor g_13131_(out[66], out[194], _07254_);
  xor g_13132_(out[69], out[197], _07255_);
  xor g_13133_(out[73], out[201], _07256_);
  xor g_13134_(out[76], out[204], _07257_);
  xor g_13135_(out[77], out[205], _07258_);
  xor g_13136_(out[79], out[207], _07259_);
  xor g_13137_(out[68], out[196], _07260_);
  xor g_13138_(out[70], out[198], _07261_);
  xor g_13139_(out[67], out[195], _07262_);
  xor g_13140_(out[64], out[192], _07263_);
  xor g_13141_(out[78], out[206], _07264_);
  or g_13142_(_07260_, _07264_, _07265_);
  or g_13143_(_07250_, _07258_, _07266_);
  or g_13144_(_07249_, _07254_, _07267_);
  or g_13145_(_07266_, _07267_, _07268_);
  or g_13146_(_07256_, _07262_, _07269_);
  or g_13147_(_07255_, _07263_, _07270_);
  or g_13148_(_07269_, _07270_, _07271_);
  or g_13149_(_07268_, _07271_, _07272_);
  or g_13150_(_07252_, _07257_, _07273_);
  xor g_13151_(out[71], out[199], _07274_);
  or g_13152_(_07261_, _07274_, _07275_);
  or g_13153_(_07273_, _07275_, _07276_);
  or g_13154_(_07251_, _07253_, _07277_);
  or g_13155_(_07259_, _07277_, _07278_);
  or g_13156_(_07276_, _07278_, _07279_);
  or g_13157_(_07272_, _07279_, _07280_);
  or g_13158_(_07265_, _07280_, _07281_);
  not g_13159_(_07281_, _07282_);
  xor g_13160_(out[55], out[199], _07283_);
  and g_13161_(_07799_, out[203], _07284_);
  xor g_13162_(out[62], out[206], _07285_);
  xor g_13163_(out[56], out[200], _07286_);
  xor g_13164_(out[49], out[193], _07287_);
  xor g_13165_(out[61], out[205], _07288_);
  xor g_13166_(out[57], out[201], _07289_);
  xor g_13167_(out[52], out[196], _07290_);
  xor g_13168_(out[50], out[194], _07291_);
  and g_13169_(out[59], _07898_, _07292_);
  xor g_13170_(out[51], out[195], _07293_);
  xor g_13171_(out[54], out[198], _07294_);
  xor g_13172_(out[63], out[207], _07295_);
  xor g_13173_(out[58], out[202], _07296_);
  xor g_13174_(out[53], out[197], _07297_);
  xor g_13175_(out[48], out[192], _07298_);
  or g_13176_(_07285_, _07290_, _07299_);
  or g_13177_(_07286_, _07288_, _07300_);
  or g_13178_(_07291_, _07296_, _07301_);
  or g_13179_(_07300_, _07301_, _07302_);
  or g_13180_(_07289_, _07293_, _07303_);
  or g_13181_(_07297_, _07298_, _07304_);
  or g_13182_(_07303_, _07304_, _07305_);
  or g_13183_(_07302_, _07305_, _07306_);
  xor g_13184_(out[60], out[204], _07307_);
  or g_13185_(_07284_, _07307_, _07308_);
  or g_13186_(_07283_, _07294_, _07309_);
  or g_13187_(_07308_, _07309_, _07310_);
  or g_13188_(_07287_, _07292_, _07311_);
  or g_13189_(_07295_, _07311_, _07312_);
  or g_13190_(_07310_, _07312_, _07313_);
  or g_13191_(_07306_, _07313_, _07314_);
  or g_13192_(_07299_, _07314_, _07315_);
  not g_13193_(_07315_, _07316_);
  xor g_13194_(out[33], out[193], _07317_);
  and g_13195_(out[43], _07898_, _07318_);
  xor g_13196_(out[41], out[201], _07319_);
  xor g_13197_(out[32], out[192], _07320_);
  xor g_13198_(out[46], out[206], _07321_);
  xor g_13199_(out[36], out[196], _07322_);
  or g_13200_(_07321_, _07322_, _07323_);
  xor g_13201_(out[45], out[205], _07324_);
  xor g_13202_(out[35], out[195], _07325_);
  and g_13203_(_07788_, out[203], _07326_);
  xor g_13204_(out[38], out[198], _07327_);
  xor g_13205_(out[42], out[202], _07328_);
  xor g_13206_(out[37], out[197], _07329_);
  xor g_13207_(out[47], out[207], _07330_);
  xor g_13208_(out[40], out[200], _07331_);
  or g_13209_(_07324_, _07331_, _07332_);
  xor g_13210_(out[34], out[194], _07333_);
  or g_13211_(_07328_, _07333_, _07334_);
  or g_13212_(_07332_, _07334_, _07335_);
  or g_13213_(_07319_, _07325_, _07336_);
  or g_13214_(_07329_, _07336_, _07337_);
  or g_13215_(_07335_, _07337_, _07338_);
  or g_13216_(_07323_, _07338_, _07339_);
  xor g_13217_(out[44], out[204], _07340_);
  or g_13218_(_07326_, _07340_, _07341_);
  xor g_13219_(out[39], out[199], _07342_);
  or g_13220_(_07327_, _07342_, _07343_);
  or g_13221_(_07341_, _07343_, _07344_);
  or g_13222_(_07317_, _07318_, _07345_);
  or g_13223_(_07330_, _07345_, _07346_);
  or g_13224_(_07344_, _07346_, _07347_);
  or g_13225_(_07320_, _07347_, _07348_);
  or g_13226_(_07339_, _07348_, _07349_);
  xor g_13227_(out[23], out[199], _07350_);
  and g_13228_(_07755_, out[203], _07351_);
  xor g_13229_(out[30], out[206], _07352_);
  xor g_13230_(out[24], out[200], _07353_);
  xor g_13231_(out[17], out[193], _07354_);
  xor g_13232_(out[29], out[205], _07355_);
  xor g_13233_(out[25], out[201], _07356_);
  xor g_13234_(out[20], out[196], _07357_);
  xor g_13235_(out[18], out[194], _07358_);
  and g_13236_(out[27], _07898_, _07359_);
  xor g_13237_(out[19], out[195], _07360_);
  xor g_13238_(out[22], out[198], _07361_);
  xor g_13239_(out[31], out[207], _07362_);
  xor g_13240_(out[26], out[202], _07363_);
  xor g_13241_(out[21], out[197], _07364_);
  xor g_13242_(out[16], out[192], _07365_);
  or g_13243_(_07352_, _07357_, _07366_);
  or g_13244_(_07353_, _07355_, _07367_);
  or g_13245_(_07358_, _07363_, _07368_);
  or g_13246_(_07367_, _07368_, _07369_);
  or g_13247_(_07356_, _07360_, _07370_);
  or g_13248_(_07364_, _07365_, _07371_);
  or g_13249_(_07370_, _07371_, _07372_);
  or g_13250_(_07369_, _07372_, _07373_);
  xor g_13251_(out[28], out[204], _07374_);
  or g_13252_(_07351_, _07374_, _07375_);
  or g_13253_(_07350_, _07361_, _07376_);
  or g_13254_(_07375_, _07376_, _07377_);
  or g_13255_(_07354_, _07359_, _07378_);
  or g_13256_(_07362_, _07378_, _07379_);
  or g_13257_(_07377_, _07379_, _07380_);
  or g_13258_(_07373_, _07380_, _07381_);
  or g_13259_(_07366_, _07381_, _07382_);
  xor g_13260_(out[1], out[193], _07383_);
  and g_13261_(out[11], _07898_, _07384_);
  xor g_13262_(out[9], out[201], _07385_);
  xor g_13263_(out[0], out[192], _07386_);
  xor g_13264_(out[14], out[206], _07387_);
  xor g_13265_(out[4], out[196], _07388_);
  or g_13266_(_07387_, _07388_, _07389_);
  xor g_13267_(out[13], out[205], _07390_);
  xor g_13268_(out[3], out[195], _07391_);
  and g_13269_(_07722_, out[203], _07392_);
  xor g_13270_(out[6], out[198], _07393_);
  xor g_13271_(out[10], out[202], _07394_);
  xor g_13272_(out[5], out[197], _07395_);
  xor g_13273_(out[15], out[207], _07396_);
  xor g_13274_(out[8], out[200], _07397_);
  or g_13275_(_07390_, _07397_, _07398_);
  xor g_13276_(out[2], out[194], _07399_);
  or g_13277_(_07394_, _07399_, _07400_);
  or g_13278_(_07398_, _07400_, _07401_);
  or g_13279_(_07385_, _07391_, _07402_);
  or g_13280_(_07395_, _07402_, _07403_);
  or g_13281_(_07401_, _07403_, _07404_);
  or g_13282_(_07389_, _07404_, _07405_);
  xor g_13283_(out[12], out[204], _07406_);
  or g_13284_(_07392_, _07406_, _07407_);
  xor g_13285_(out[7], out[199], _07408_);
  or g_13286_(_07393_, _07408_, _07409_);
  or g_13287_(_07407_, _07409_, _07410_);
  or g_13288_(_07383_, _07384_, _07411_);
  or g_13289_(_07396_, _07411_, _07412_);
  or g_13290_(_07410_, _07412_, _07413_);
  or g_13291_(_07386_, _07413_, _07414_);
  or g_13292_(_07405_, _07414_, _07415_);
  not g_13293_(_07415_, _07416_);
  xor g_13294_(out[145], out[177], _07417_);
  and g_13295_(out[155], _07887_, _07418_);
  xor g_13296_(out[153], out[185], _07419_);
  xor g_13297_(out[144], out[176], _07420_);
  xor g_13298_(out[158], out[190], _07421_);
  xor g_13299_(out[148], out[180], _07422_);
  or g_13300_(_07421_, _07422_, _07423_);
  xor g_13301_(out[157], out[189], _07424_);
  xor g_13302_(out[147], out[179], _07425_);
  and g_13303_(_07876_, out[187], _07426_);
  xor g_13304_(out[150], out[182], _07427_);
  xor g_13305_(out[154], out[186], _07428_);
  xor g_13306_(out[149], out[181], _07429_);
  xor g_13307_(out[159], out[191], _07430_);
  xor g_13308_(out[152], out[184], _07431_);
  or g_13309_(_07424_, _07431_, _07432_);
  xor g_13310_(out[146], out[178], _07433_);
  or g_13311_(_07428_, _07433_, _07434_);
  or g_13312_(_07432_, _07434_, _07435_);
  or g_13313_(_07419_, _07425_, _07436_);
  or g_13314_(_07429_, _07436_, _07437_);
  or g_13315_(_07435_, _07437_, _07438_);
  or g_13316_(_07423_, _07438_, _07439_);
  xor g_13317_(out[156], out[188], _07440_);
  or g_13318_(_07426_, _07440_, _07441_);
  xor g_13319_(out[151], out[183], _07442_);
  or g_13320_(_07427_, _07442_, _07443_);
  or g_13321_(_07441_, _07443_, _07444_);
  or g_13322_(_07417_, _07418_, _07445_);
  or g_13323_(_07430_, _07445_, _07446_);
  or g_13324_(_07444_, _07446_, _07447_);
  or g_13325_(_07420_, _07447_, _07448_);
  or g_13326_(_07439_, _07448_, _07449_);
  xor g_13327_(out[135], out[183], _07450_);
  and g_13328_(_07854_, out[187], _07451_);
  xor g_13329_(out[142], out[190], _07452_);
  xor g_13330_(out[136], out[184], _07453_);
  xor g_13331_(out[129], out[177], _07454_);
  xor g_13332_(out[141], out[189], _07455_);
  xor g_13333_(out[137], out[185], _07456_);
  xor g_13334_(out[132], out[180], _07457_);
  xor g_13335_(out[130], out[178], _07458_);
  and g_13336_(out[139], _07887_, _07459_);
  xor g_13337_(out[131], out[179], _07460_);
  xor g_13338_(out[134], out[182], _07461_);
  xor g_13339_(out[143], out[191], _07462_);
  xor g_13340_(out[138], out[186], _07463_);
  xor g_13341_(out[133], out[181], _07464_);
  xor g_13342_(out[128], out[176], _07465_);
  or g_13343_(_07452_, _07457_, _07466_);
  or g_13344_(_07453_, _07455_, _07467_);
  or g_13345_(_07458_, _07463_, _07468_);
  or g_13346_(_07467_, _07468_, _07469_);
  or g_13347_(_07456_, _07460_, _07470_);
  or g_13348_(_07464_, _07465_, _07471_);
  or g_13349_(_07470_, _07471_, _07472_);
  or g_13350_(_07469_, _07472_, _07473_);
  xor g_13351_(out[140], out[188], _07474_);
  or g_13352_(_07451_, _07474_, _07475_);
  or g_13353_(_07450_, _07461_, _07476_);
  or g_13354_(_07475_, _07476_, _07477_);
  or g_13355_(_07454_, _07459_, _07478_);
  or g_13356_(_07462_, _07478_, _07479_);
  or g_13357_(_07477_, _07479_, _07480_);
  or g_13358_(_07473_, _07480_, _07481_);
  or g_13359_(_07466_, _07481_, _07482_);
  xor g_13360_(out[113], out[177], _07483_);
  and g_13361_(out[123], _07887_, _07484_);
  xor g_13362_(out[126], out[190], _07485_);
  xor g_13363_(out[115], out[179], _07486_);
  xor g_13364_(out[116], out[180], _07487_);
  xor g_13365_(out[114], out[178], _07488_);
  xor g_13366_(out[121], out[185], _07489_);
  xor g_13367_(out[112], out[176], _07490_);
  and g_13368_(_07843_, out[187], _07491_);
  xor g_13369_(out[118], out[182], _07492_);
  xor g_13370_(out[122], out[186], _07493_);
  xor g_13371_(out[117], out[181], _07494_);
  xor g_13372_(out[127], out[191], _07495_);
  xor g_13373_(out[125], out[189], _07496_);
  xor g_13374_(out[120], out[184], _07497_);
  or g_13375_(_07485_, _07487_, _07498_);
  or g_13376_(_07496_, _07497_, _07499_);
  or g_13377_(_07488_, _07493_, _07500_);
  or g_13378_(_07499_, _07500_, _07501_);
  or g_13379_(_07486_, _07489_, _07502_);
  or g_13380_(_07490_, _07494_, _07503_);
  or g_13381_(_07502_, _07503_, _07504_);
  or g_13382_(_07501_, _07504_, _07505_);
  xor g_13383_(out[124], out[188], _07506_);
  or g_13384_(_07491_, _07506_, _07507_);
  xor g_13385_(out[119], out[183], _07508_);
  or g_13386_(_07492_, _07508_, _07509_);
  or g_13387_(_07507_, _07509_, _07510_);
  or g_13388_(_07483_, _07484_, _07511_);
  or g_13389_(_07495_, _07511_, _07512_);
  or g_13390_(_07510_, _07512_, _07513_);
  or g_13391_(_07505_, _07513_, _07514_);
  or g_13392_(_07498_, _07514_, _07515_);
  xor g_13393_(out[103], out[183], _07516_);
  and g_13394_(_07832_, out[187], _07517_);
  xor g_13395_(out[110], out[190], _07518_);
  xor g_13396_(out[104], out[184], _07519_);
  xor g_13397_(out[97], out[177], _07520_);
  xor g_13398_(out[109], out[189], _07521_);
  xor g_13399_(out[105], out[185], _07522_);
  xor g_13400_(out[100], out[180], _07523_);
  xor g_13401_(out[98], out[178], _07524_);
  and g_13402_(out[107], _07887_, _07525_);
  xor g_13403_(out[99], out[179], _07526_);
  xor g_13404_(out[102], out[182], _07527_);
  xor g_13405_(out[111], out[191], _07528_);
  xor g_13406_(out[106], out[186], _07529_);
  xor g_13407_(out[101], out[181], _07530_);
  xor g_13408_(out[96], out[176], _07531_);
  or g_13409_(_07518_, _07523_, _07532_);
  or g_13410_(_07519_, _07521_, _07533_);
  or g_13411_(_07524_, _07529_, _07534_);
  or g_13412_(_07533_, _07534_, _07535_);
  or g_13413_(_07522_, _07526_, _07536_);
  or g_13414_(_07530_, _07531_, _07537_);
  or g_13415_(_07536_, _07537_, _07538_);
  or g_13416_(_07535_, _07538_, _07539_);
  xor g_13417_(out[108], out[188], _07540_);
  or g_13418_(_07517_, _07540_, _07541_);
  or g_13419_(_07516_, _07527_, _07542_);
  or g_13420_(_07541_, _07542_, _07543_);
  or g_13421_(_07520_, _07525_, _07544_);
  or g_13422_(_07528_, _07544_, _07545_);
  or g_13423_(_07543_, _07545_, _07546_);
  or g_13424_(_07539_, _07546_, _07547_);
  or g_13425_(_07532_, _07547_, _07548_);
  xor g_13426_(out[88], out[184], _07549_);
  xor g_13427_(out[85], out[181], _07550_);
  xor g_13428_(out[83], out[179], _07551_);
  xor g_13429_(out[94], out[190], _07552_);
  xor g_13430_(out[93], out[189], _07553_);
  xor g_13431_(out[82], out[178], _07554_);
  xor g_13432_(out[89], out[185], _07555_);
  xor g_13433_(out[86], out[182], _07556_);
  xor g_13434_(out[95], out[191], _07557_);
  xor g_13435_(out[90], out[186], _07558_);
  xor g_13436_(out[84], out[180], _07559_);
  xor g_13437_(out[80], out[176], _07560_);
  and g_13438_(_07821_, out[187], _07561_);
  and g_13439_(out[91], _07887_, _07562_);
  or g_13440_(_07549_, _07553_, _07563_);
  xor g_13441_(out[81], out[177], _07564_);
  or g_13442_(_07554_, _07558_, _07565_);
  or g_13443_(_07563_, _07565_, _07566_);
  or g_13444_(_07551_, _07555_, _07567_);
  or g_13445_(_07550_, _07567_, _07568_);
  or g_13446_(_07566_, _07568_, _07569_);
  or g_13447_(_07552_, _07559_, _07570_);
  or g_13448_(_07569_, _07570_, _07571_);
  xor g_13449_(out[92], out[188], _07572_);
  or g_13450_(_07561_, _07572_, _07573_);
  xor g_13451_(out[87], out[183], _07574_);
  or g_13452_(_07556_, _07574_, _07575_);
  or g_13453_(_07573_, _07575_, _07576_);
  or g_13454_(_07562_, _07564_, _07577_);
  or g_13455_(_07557_, _07577_, _07578_);
  or g_13456_(_07576_, _07578_, _07579_);
  or g_13457_(_07560_, _07579_, _07580_);
  or g_13458_(_07571_, _07580_, _07581_);
  not g_13459_(_07581_, _07582_);
  xor g_13460_(out[71], out[183], _07583_);
  and g_13461_(_07810_, out[187], _07584_);
  xor g_13462_(out[78], out[190], _07585_);
  xor g_13463_(out[72], out[184], _07586_);
  xor g_13464_(out[65], out[177], _07587_);
  xor g_13465_(out[77], out[189], _07588_);
  xor g_13466_(out[73], out[185], _07589_);
  xor g_13467_(out[68], out[180], _07590_);
  xor g_13468_(out[66], out[178], _07591_);
  and g_13469_(out[75], _07887_, _07592_);
  xor g_13470_(out[67], out[179], _07593_);
  xor g_13471_(out[70], out[182], _07594_);
  xor g_13472_(out[79], out[191], _07595_);
  xor g_13473_(out[74], out[186], _07596_);
  xor g_13474_(out[69], out[181], _07597_);
  xor g_13475_(out[64], out[176], _07598_);
  or g_13476_(_07585_, _07590_, _07599_);
  or g_13477_(_07586_, _07588_, _07600_);
  or g_13478_(_07591_, _07596_, _07601_);
  or g_13479_(_07600_, _07601_, _07602_);
  or g_13480_(_07589_, _07593_, _07603_);
  or g_13481_(_07597_, _07598_, _07604_);
  or g_13482_(_07603_, _07604_, _07605_);
  or g_13483_(_07602_, _07605_, _07606_);
  xor g_13484_(out[76], out[188], _07607_);
  or g_13485_(_07584_, _07607_, _07608_);
  or g_13486_(_07583_, _07594_, _07609_);
  or g_13487_(_07608_, _07609_, _07610_);
  or g_13488_(_07587_, _07592_, _07611_);
  or g_13489_(_07595_, _07611_, _07612_);
  or g_13490_(_07610_, _07612_, _07613_);
  or g_13491_(_07606_, _07613_, _07614_);
  or g_13492_(_07599_, _07614_, _07615_);
  not g_13493_(_07615_, _07616_);
  xor g_13494_(out[49], out[177], _07617_);
  and g_13495_(out[59], _07887_, _07618_);
  xor g_13496_(out[57], out[185], _07619_);
  xor g_13497_(out[48], out[176], _07620_);
  xor g_13498_(out[62], out[190], _07621_);
  xor g_13499_(out[52], out[180], _07622_);
  or g_13500_(_07621_, _07622_, _07623_);
  xor g_13501_(out[61], out[189], _07624_);
  xor g_13502_(out[51], out[179], _07625_);
  and g_13503_(_07799_, out[187], _07626_);
  xor g_13504_(out[54], out[182], _07627_);
  xor g_13505_(out[58], out[186], _07628_);
  xor g_13506_(out[53], out[181], _07629_);
  xor g_13507_(out[63], out[191], _07630_);
  xor g_13508_(out[56], out[184], _07631_);
  or g_13509_(_07624_, _07631_, _07632_);
  xor g_13510_(out[50], out[178], _07633_);
  or g_13511_(_07628_, _07633_, _07634_);
  or g_13512_(_07632_, _07634_, _07635_);
  or g_13513_(_07619_, _07625_, _07636_);
  or g_13514_(_07629_, _07636_, _07637_);
  or g_13515_(_07635_, _07637_, _07638_);
  or g_13516_(_07623_, _07638_, _07639_);
  xor g_13517_(out[60], out[188], _07640_);
  or g_13518_(_07626_, _07640_, _07641_);
  xor g_13519_(out[55], out[183], _07642_);
  or g_13520_(_07627_, _07642_, _07643_);
  or g_13521_(_07641_, _07643_, _07644_);
  or g_13522_(_07617_, _07618_, _07645_);
  or g_13523_(_07630_, _07645_, _07646_);
  or g_13524_(_07644_, _07646_, _07647_);
  or g_13525_(_07620_, _07647_, _07648_);
  or g_13526_(_07639_, _07648_, _07649_);
  xor g_13527_(out[39], out[183], _07650_);
  and g_13528_(_07788_, out[187], _07651_);
  xor g_13529_(out[46], out[190], _07652_);
  xor g_13530_(out[40], out[184], _07653_);
  xor g_13531_(out[33], out[177], _07654_);
  xor g_13532_(out[45], out[189], _07655_);
  xor g_13533_(out[41], out[185], _07656_);
  xor g_13534_(out[36], out[180], _07657_);
  xor g_13535_(out[34], out[178], _07658_);
  and g_13536_(out[43], _07887_, _07659_);
  xor g_13537_(out[35], out[179], _07660_);
  xor g_13538_(out[38], out[182], _07661_);
  xor g_13539_(out[47], out[191], _07662_);
  xor g_13540_(out[42], out[186], _07663_);
  xor g_13541_(out[37], out[181], _07664_);
  xor g_13542_(out[32], out[176], _07665_);
  or g_13543_(_07652_, _07657_, _07666_);
  or g_13544_(_07653_, _07655_, _07667_);
  or g_13545_(_07658_, _07663_, _07668_);
  or g_13546_(_07667_, _07668_, _07669_);
  or g_13547_(_07656_, _07660_, _07670_);
  or g_13548_(_07664_, _07665_, _07671_);
  or g_13549_(_07670_, _07671_, _07672_);
  or g_13550_(_07669_, _07672_, _07673_);
  xor g_13551_(out[44], out[188], _07674_);
  or g_13552_(_07651_, _07674_, _07675_);
  or g_13553_(_07650_, _07661_, _07676_);
  or g_13554_(_07675_, _07676_, _07677_);
  or g_13555_(_07654_, _07659_, _07678_);
  or g_13556_(_07662_, _07678_, _07679_);
  or g_13557_(_07677_, _07679_, _07680_);
  or g_13558_(_07673_, _07680_, _07681_);
  or g_13559_(_07666_, _07681_, _07682_);
  xor g_13560_(out[17], out[177], _07683_);
  and g_13561_(_07755_, out[187], _07684_);
  and g_13562_(out[27], _07887_, _07685_);
  xor g_13563_(out[24], out[184], _07686_);
  xor g_13564_(out[26], out[186], _07687_);
  xor g_13565_(out[18], out[178], _07688_);
  xor g_13566_(out[20], out[180], _07689_);
  xor g_13567_(out[21], out[181], _07690_);
  xor g_13568_(out[25], out[185], _07691_);
  xor g_13569_(out[19], out[179], _07692_);
  xor g_13570_(out[30], out[190], _07693_);
  xor g_13571_(out[16], out[176], _07694_);
  xor g_13572_(out[31], out[191], _07695_);
  xor g_13573_(out[29], out[189], _07696_);
  or g_13574_(_07686_, _07696_, _07697_);
  xor g_13575_(out[22], out[182], _07698_);
  or g_13576_(_07687_, _07688_, _07699_);
  or g_13577_(_07697_, _07699_, _07701_);
  or g_13578_(_07691_, _07692_, _07702_);
  or g_13579_(_07690_, _07702_, _07703_);
  or g_13580_(_07701_, _07703_, _07704_);
  or g_13581_(_07689_, _07693_, _07705_);
  or g_13582_(_07704_, _07705_, _07706_);
  xor g_13583_(out[28], out[188], _07707_);
  or g_13584_(_07684_, _07707_, _07708_);
  xor g_13585_(out[23], out[183], _07709_);
  or g_13586_(_07698_, _07709_, _07710_);
  or g_13587_(_07708_, _07710_, _07712_);
  or g_13588_(_07683_, _07685_, _07713_);
  or g_13589_(_07695_, _07713_, _07714_);
  or g_13590_(_07712_, _07714_, _07715_);
  or g_13591_(_07694_, _07715_, _07716_);
  or g_13592_(_07706_, _07716_, _07717_);
  xor g_13593_(out[1], out[177], _07718_);
  and g_13594_(out[11], _07887_, _07719_);
  xor g_13595_(out[9], out[185], _07720_);
  xor g_13596_(out[0], out[176], _07721_);
  xor g_13597_(out[14], out[190], _07723_);
  xor g_13598_(out[4], out[180], _07724_);
  or g_13599_(_07723_, _07724_, _07725_);
  xor g_13600_(out[13], out[189], _07726_);
  xor g_13601_(out[3], out[179], _07727_);
  and g_13602_(_07722_, out[187], _07728_);
  xor g_13603_(out[6], out[182], _07729_);
  xor g_13604_(out[10], out[186], _07730_);
  xor g_13605_(out[5], out[181], _07731_);
  xor g_13606_(out[15], out[191], _07732_);
  xor g_13607_(out[8], out[184], _07734_);
  or g_13608_(_07726_, _07734_, _07735_);
  xor g_13609_(out[2], out[178], _07736_);
  or g_13610_(_07730_, _07736_, _07737_);
  or g_13611_(_07735_, _07737_, _07738_);
  or g_13612_(_07720_, _07727_, _07739_);
  or g_13613_(_07731_, _07739_, _07740_);
  or g_13614_(_07738_, _07740_, _07741_);
  or g_13615_(_07725_, _07741_, _07742_);
  xor g_13616_(out[12], out[188], _07743_);
  or g_13617_(_07728_, _07743_, _07745_);
  xor g_13618_(out[7], out[183], _07746_);
  or g_13619_(_07729_, _07746_, _07747_);
  or g_13620_(_07745_, _07747_, _07748_);
  or g_13621_(_07718_, _07719_, _07749_);
  or g_13622_(_07732_, _07749_, _07750_);
  or g_13623_(_07748_, _07750_, _07751_);
  or g_13624_(_07721_, _07751_, _07752_);
  or g_13625_(_07742_, _07752_, _07753_);
  xor g_13626_(out[172], out[156], _07754_);
  and g_13627_(_07733_, out[155], _07756_);
  xor g_13628_(out[168], out[152], _07757_);
  xor g_13629_(out[166], out[150], _07758_);
  xor g_13630_(out[173], out[157], _07759_);
  xor g_13631_(out[174], out[158], _07760_);
  xor g_13632_(out[162], out[146], _07761_);
  xor g_13633_(out[169], out[153], _07762_);
  xor g_13634_(out[165], out[149], _07763_);
  xor g_13635_(out[161], out[145], _07764_);
  and g_13636_(out[171], _07876_, _07765_);
  or g_13637_(_07757_, _07759_, _07767_);
  xor g_13638_(out[175], out[159], _07768_);
  xor g_13639_(out[170], out[154], _07769_);
  xor g_13640_(out[164], out[148], _07770_);
  xor g_13641_(out[163], out[147], _07771_);
  xor g_13642_(out[160], out[144], _07772_);
  or g_13643_(_07761_, _07769_, _07773_);
  or g_13644_(_07767_, _07773_, _07774_);
  or g_13645_(_07762_, _07771_, _07775_);
  or g_13646_(_07763_, _07775_, _07776_);
  or g_13647_(_07774_, _07776_, _07778_);
  or g_13648_(_07760_, _07770_, _07779_);
  or g_13649_(_07778_, _07779_, _07780_);
  or g_13650_(_07754_, _07756_, _07781_);
  xor g_13651_(out[167], out[151], _07782_);
  or g_13652_(_07758_, _07782_, _07783_);
  or g_13653_(_07781_, _07783_, _07784_);
  or g_13654_(_07764_, _07765_, _07785_);
  or g_13655_(_07768_, _07785_, _07786_);
  or g_13656_(_07784_, _07786_, _07787_);
  or g_13657_(_07772_, _07787_, _07789_);
  or g_13658_(_07780_, _07789_, _07790_);
  not g_13659_(_07790_, _07791_);
  xor g_13660_(out[161], out[129], _07792_);
  and g_13661_(out[171], _07854_, _07793_);
  xor g_13662_(out[169], out[137], _07794_);
  xor g_13663_(out[160], out[128], _07795_);
  xor g_13664_(out[174], out[142], _07796_);
  xor g_13665_(out[164], out[132], _07797_);
  or g_13666_(_07796_, _07797_, _07798_);
  xor g_13667_(out[173], out[141], _07800_);
  xor g_13668_(out[163], out[131], _07801_);
  and g_13669_(_07733_, out[139], _07802_);
  xor g_13670_(out[166], out[134], _07803_);
  xor g_13671_(out[170], out[138], _07804_);
  xor g_13672_(out[165], out[133], _07805_);
  xor g_13673_(out[175], out[143], _07806_);
  xor g_13674_(out[168], out[136], _07807_);
  or g_13675_(_07800_, _07807_, _07808_);
  xor g_13676_(out[162], out[130], _07809_);
  or g_13677_(_07804_, _07809_, _07811_);
  or g_13678_(_07808_, _07811_, _07812_);
  or g_13679_(_07794_, _07801_, _07813_);
  or g_13680_(_07805_, _07813_, _07814_);
  or g_13681_(_07812_, _07814_, _07815_);
  or g_13682_(_07798_, _07815_, _07816_);
  xor g_13683_(out[172], out[140], _07817_);
  or g_13684_(_07802_, _07817_, _07818_);
  xor g_13685_(out[167], out[135], _07819_);
  or g_13686_(_07803_, _07819_, _07820_);
  or g_13687_(_07818_, _07820_, _07822_);
  or g_13688_(_07792_, _07793_, _07823_);
  or g_13689_(_07806_, _07823_, _07824_);
  or g_13690_(_07822_, _07824_, _07825_);
  or g_13691_(_07795_, _07825_, _07826_);
  or g_13692_(_07816_, _07826_, _07827_);
  not g_13693_(_07827_, _07828_);
  xor g_13694_(out[170], out[122], _07829_);
  xor g_13695_(out[162], out[114], _07830_);
  xor g_13696_(out[161], out[113], _07831_);
  and g_13697_(_07733_, out[123], _07833_);
  and g_13698_(out[171], _07843_, _07834_);
  xor g_13699_(out[173], out[125], _07835_);
  xor g_13700_(out[163], out[115], _07836_);
  xor g_13701_(out[174], out[126], _07837_);
  xor g_13702_(out[172], out[124], _07838_);
  xor g_13703_(out[168], out[120], _07839_);
  xor g_13704_(out[175], out[127], _07840_);
  xor g_13705_(out[165], out[117], _07841_);
  xor g_13706_(out[166], out[118], _07842_);
  xor g_13707_(out[160], out[112], _07844_);
  xor g_13708_(out[164], out[116], _07845_);
  or g_13709_(_07835_, _07839_, _07846_);
  xor g_13710_(out[169], out[121], _07847_);
  or g_13711_(_07829_, _07830_, _07848_);
  or g_13712_(_07846_, _07848_, _07849_);
  or g_13713_(_07836_, _07847_, _07850_);
  or g_13714_(_07841_, _07850_, _07851_);
  or g_13715_(_07849_, _07851_, _07852_);
  or g_13716_(_07837_, _07845_, _07853_);
  or g_13717_(_07852_, _07853_, _07855_);
  or g_13718_(_07833_, _07838_, _07856_);
  xor g_13719_(out[167], out[119], _07857_);
  or g_13720_(_07842_, _07857_, _07858_);
  or g_13721_(_07856_, _07858_, _07859_);
  or g_13722_(_07831_, _07834_, _07860_);
  or g_13723_(_07840_, _07860_, _07861_);
  or g_13724_(_07859_, _07861_, _07862_);
  or g_13725_(_07844_, _07862_, _07863_);
  or g_13726_(_07855_, _07863_, _07864_);
  not g_13727_(_07864_, _07866_);
  xor g_13728_(out[161], out[97], _07867_);
  and g_13729_(out[171], _07832_, _07868_);
  xor g_13730_(out[169], out[105], _07869_);
  xor g_13731_(out[160], out[96], _07870_);
  xor g_13732_(out[174], out[110], _07871_);
  xor g_13733_(out[164], out[100], _07872_);
  or g_13734_(_07871_, _07872_, _07873_);
  xor g_13735_(out[173], out[109], _07874_);
  xor g_13736_(out[163], out[99], _07875_);
  and g_13737_(_07733_, out[107], _07877_);
  xor g_13738_(out[166], out[102], _07878_);
  xor g_13739_(out[170], out[106], _07879_);
  xor g_13740_(out[165], out[101], _07880_);
  xor g_13741_(out[175], out[111], _07881_);
  xor g_13742_(out[168], out[104], _07882_);
  or g_13743_(_07874_, _07882_, _07883_);
  xor g_13744_(out[162], out[98], _07884_);
  or g_13745_(_07879_, _07884_, _07885_);
  or g_13746_(_07883_, _07885_, _07886_);
  or g_13747_(_07869_, _07875_, _07888_);
  or g_13748_(_07880_, _07888_, _07889_);
  or g_13749_(_07886_, _07889_, _07890_);
  or g_13750_(_07873_, _07890_, _07891_);
  xor g_13751_(out[172], out[108], _07892_);
  or g_13752_(_07877_, _07892_, _07893_);
  xor g_13753_(out[167], out[103], _07894_);
  or g_13754_(_07878_, _07894_, _07895_);
  or g_13755_(_07893_, _07895_, _07896_);
  or g_13756_(_07867_, _07868_, _07897_);
  or g_13757_(_07881_, _07897_, _07899_);
  or g_13758_(_07896_, _07899_, _07900_);
  or g_13759_(_07870_, _07900_, _07901_);
  or g_13760_(_07891_, _07901_, _07902_);
  not g_13761_(_07902_, _07903_);
  xor g_13762_(out[172], out[92], _07904_);
  and g_13763_(_07733_, out[91], _07905_);
  xor g_13764_(out[173], out[93], _07906_);
  xor g_13765_(out[166], out[86], _07907_);
  xor g_13766_(out[168], out[88], _07908_);
  xor g_13767_(out[169], out[89], _07910_);
  xor g_13768_(out[174], out[94], _07911_);
  xor g_13769_(out[164], out[84], _07912_);
  or g_13770_(_07911_, _07912_, _07913_);
  xor g_13771_(out[165], out[85], _07914_);
  xor g_13772_(out[161], out[81], _07915_);
  and g_13773_(out[171], _07821_, _07916_);
  xor g_13774_(out[175], out[95], _07917_);
  xor g_13775_(out[170], out[90], _07918_);
  xor g_13776_(out[160], out[80], _07919_);
  xor g_13777_(out[162], out[82], _07921_);
  xor g_13778_(out[163], out[83], _07922_);
  or g_13779_(_07906_, _07908_, _07923_);
  or g_13780_(_07918_, _07921_, _07924_);
  or g_13781_(_07923_, _07924_, _07925_);
  or g_13782_(_07910_, _07922_, _07926_);
  or g_13783_(_07914_, _07919_, _07927_);
  or g_13784_(_07926_, _07927_, _07928_);
  or g_13785_(_07925_, _07928_, _07929_);
  or g_13786_(_07904_, _07905_, _07930_);
  xor g_13787_(out[167], out[87], _07932_);
  or g_13788_(_07907_, _07932_, _07933_);
  or g_13789_(_07930_, _07933_, _07934_);
  or g_13790_(_07915_, _07916_, _07935_);
  or g_13791_(_07917_, _07935_, _07936_);
  or g_13792_(_07934_, _07936_, _07937_);
  or g_13793_(_07929_, _07937_, _07938_);
  or g_13794_(_07913_, _07938_, _07939_);
  not g_13795_(_07939_, _07940_);
  xor g_13796_(out[172], out[76], _07941_);
  and g_13797_(_07733_, out[75], _07943_);
  xor g_13798_(out[168], out[72], _07944_);
  xor g_13799_(out[166], out[70], _07945_);
  xor g_13800_(out[173], out[77], _07946_);
  xor g_13801_(out[174], out[78], _07947_);
  xor g_13802_(out[162], out[66], _07948_);
  xor g_13803_(out[169], out[73], _07949_);
  xor g_13804_(out[165], out[69], _07950_);
  xor g_13805_(out[161], out[65], _07951_);
  and g_13806_(out[171], _07810_, _07952_);
  or g_13807_(_07944_, _07946_, _07954_);
  xor g_13808_(out[175], out[79], _07955_);
  xor g_13809_(out[170], out[74], _07956_);
  xor g_13810_(out[164], out[68], _07957_);
  xor g_13811_(out[163], out[67], _07958_);
  xor g_13812_(out[160], out[64], _07959_);
  or g_13813_(_07948_, _07956_, _07960_);
  or g_13814_(_07954_, _07960_, _07961_);
  or g_13815_(_07949_, _07958_, _07962_);
  or g_13816_(_07950_, _07962_, _07963_);
  or g_13817_(_07961_, _07963_, _07965_);
  or g_13818_(_07947_, _07957_, _07966_);
  or g_13819_(_07965_, _07966_, _07967_);
  or g_13820_(_07941_, _07943_, _07968_);
  xor g_13821_(out[167], out[71], _07969_);
  or g_13822_(_07945_, _07969_, _07970_);
  or g_13823_(_07968_, _07970_, _07971_);
  or g_13824_(_07951_, _07952_, _07972_);
  or g_13825_(_07955_, _07972_, _07973_);
  or g_13826_(_07971_, _07973_, _07974_);
  or g_13827_(_07959_, _07974_, _07976_);
  or g_13828_(_07967_, _07976_, _07977_);
  not g_13829_(_07977_, _07978_);
  xor g_13830_(out[166], out[54], _07979_);
  xor g_13831_(out[161], out[49], _07980_);
  xor g_13832_(out[160], out[48], _07981_);
  xor g_13833_(out[162], out[50], _07982_);
  xor g_13834_(out[163], out[51], _07983_);
  xor g_13835_(out[169], out[57], _07984_);
  xor g_13836_(out[174], out[62], _07985_);
  and g_13837_(_07733_, out[59], _07987_);
  xor g_13838_(out[167], out[55], _07988_);
  and g_13839_(out[171], _07799_, _07989_);
  xor g_13840_(out[173], out[61], _07990_);
  xor g_13841_(out[168], out[56], _07991_);
  or g_13842_(_07990_, _07991_, _07992_);
  xor g_13843_(out[175], out[63], _07993_);
  xor g_13844_(out[170], out[58], _07994_);
  xor g_13845_(out[165], out[53], _07995_);
  xor g_13846_(out[164], out[52], _07996_);
  or g_13847_(_07982_, _07994_, _07998_);
  or g_13848_(_07992_, _07998_, _07999_);
  or g_13849_(_07983_, _07984_, _08000_);
  or g_13850_(_07995_, _08000_, _08001_);
  or g_13851_(_07999_, _08001_, _08002_);
  or g_13852_(_07985_, _07996_, _08003_);
  or g_13853_(_08002_, _08003_, _08004_);
  xor g_13854_(out[172], out[60], _08005_);
  or g_13855_(_07987_, _08005_, _08006_);
  or g_13856_(_07979_, _07988_, _08007_);
  or g_13857_(_08006_, _08007_, _08009_);
  or g_13858_(_07980_, _07989_, _08010_);
  or g_13859_(_07993_, _08010_, _08011_);
  or g_13860_(_08009_, _08011_, _08012_);
  or g_13861_(_07981_, _08012_, _08013_);
  or g_13862_(_08004_, _08013_, _08014_);
  and g_13863_(out[167], _07777_, _08015_);
  and g_13864_(_07711_, out[39], _08016_);
  xor g_13865_(out[163], out[35], _08017_);
  xor g_13866_(out[172], out[44], _08018_);
  xor g_13867_(out[169], out[41], _08020_);
  xor g_13868_(out[166], out[38], _08021_);
  xor g_13869_(out[170], out[42], _08022_);
  or g_13870_(_08021_, _08022_, _08023_);
  xor g_13871_(out[165], out[37], _08024_);
  xor g_13872_(out[161], out[33], _08025_);
  xor g_13873_(out[171], out[43], _08026_);
  xor g_13874_(out[160], out[32], _08027_);
  xor g_13875_(out[168], out[40], _08028_);
  xor g_13876_(out[173], out[45], _08029_);
  xor g_13877_(out[164], out[36], _08031_);
  or g_13878_(_08017_, _08031_, _08032_);
  xor g_13879_(out[174], out[46], _08033_);
  or g_13880_(_08023_, _08032_, _08034_);
  or g_13881_(_08024_, _08026_, _08035_);
  or g_13882_(_08029_, _08035_, _08036_);
  or g_13883_(_08034_, _08036_, _08037_);
  or g_13884_(_08018_, _08027_, _08038_);
  or g_13885_(_08037_, _08038_, _08039_);
  xor g_13886_(out[162], out[34], _08040_);
  or g_13887_(_08016_, _08040_, _08042_);
  xor g_13888_(out[175], out[47], _08043_);
  or g_13889_(_08033_, _08043_, _08044_);
  or g_13890_(_08042_, _08044_, _08045_);
  or g_13891_(_08015_, _08020_, _08046_);
  or g_13892_(_08025_, _08046_, _08047_);
  or g_13893_(_08045_, _08047_, _08048_);
  or g_13894_(_08028_, _08048_, _08049_);
  or g_13895_(_08039_, _08049_, _08050_);
  not g_13896_(_08050_, _08051_);
  xor g_13897_(out[166], out[22], _08053_);
  xor g_13898_(out[170], out[26], _08054_);
  xor g_13899_(out[174], out[30], _08055_);
  xor g_13900_(out[164], out[20], _08056_);
  xor g_13901_(out[163], out[19], _08057_);
  xor g_13902_(out[175], out[31], _08058_);
  xor g_13903_(out[173], out[29], _08059_);
  and g_13904_(_07744_, out[28], _08060_);
  xor g_13905_(out[165], out[21], _08061_);
  and g_13906_(out[172], _07766_, _08062_);
  xor g_13907_(out[167], out[23], _08064_);
  xor g_13908_(out[160], out[16], _08065_);
  xor g_13909_(out[169], out[25], _08066_);
  xor g_13910_(out[171], out[27], _08067_);
  xor g_13911_(out[162], out[18], _08068_);
  xor g_13912_(out[161], out[17], _08069_);
  or g_13913_(_08055_, _08066_, _08070_);
  or g_13914_(_08053_, _08067_, _08071_);
  or g_13915_(_08070_, _08071_, _08072_);
  or g_13916_(_08054_, _08064_, _08073_);
  or g_13917_(_08056_, _08073_, _08075_);
  or g_13918_(_08072_, _08075_, _08076_);
  or g_13919_(_08065_, _08068_, _08077_);
  or g_13920_(_08076_, _08077_, _08078_);
  or g_13921_(_08059_, _08060_, _08079_);
  xor g_13922_(out[168], out[24], _08080_);
  or g_13923_(_08069_, _08080_, _08081_);
  or g_13924_(_08079_, _08081_, _08082_);
  or g_13925_(_08061_, _08062_, _08083_);
  or g_13926_(_08058_, _08083_, _08084_);
  or g_13927_(_08082_, _08084_, _08086_);
  or g_13928_(_08057_, _08086_, _08087_);
  or g_13929_(_08078_, _08087_, _08088_);
  xor g_13930_(out[10], out[170], _08089_);
  xor g_13931_(out[5], out[165], _08090_);
  xor g_13932_(out[9], out[169], _08091_);
  and g_13933_(out[7], _07711_, _08092_);
  xor g_13934_(out[12], out[172], _08093_);
  xor g_13935_(out[8], out[168], _08094_);
  xor g_13936_(out[2], out[162], _08095_);
  and g_13937_(_07700_, out[167], _08097_);
  xor g_13938_(out[11], out[171], _08098_);
  xor g_13939_(out[0], out[160], _08099_);
  xor g_13940_(out[4], out[164], _08100_);
  xor g_13941_(out[6], out[166], _08101_);
  xor g_13942_(out[3], out[163], _08102_);
  xor g_13943_(out[13], out[173], _08103_);
  xor g_13944_(out[14], out[174], _08104_);
  xor g_13945_(out[1], out[161], _08105_);
  or g_13946_(_08100_, _08102_, _08106_);
  or g_13947_(_08089_, _08101_, _08108_);
  or g_13948_(_08106_, _08108_, _08109_);
  or g_13949_(_08090_, _08098_, _08110_);
  or g_13950_(_08103_, _08110_, _08111_);
  or g_13951_(_08109_, _08111_, _08112_);
  or g_13952_(_08093_, _08099_, _08113_);
  or g_13953_(_08112_, _08113_, _08114_);
  or g_13954_(_08095_, _08097_, _08115_);
  xor g_13955_(out[15], out[175], _08116_);
  or g_13956_(_08104_, _08116_, _08117_);
  or g_13957_(_08115_, _08117_, _08119_);
  or g_13958_(_08091_, _08092_, _08120_);
  or g_13959_(_08105_, _08120_, _08121_);
  or g_13960_(_08119_, _08121_, _08122_);
  or g_13961_(_08094_, _08122_, _08123_);
  or g_13962_(_08114_, _08123_, _08124_);
  or g_13963_(_08088_, _08124_, _08125_);
  and g_13964_(_08088_, _08124_, _08126_);
  xor g_13965_(_08088_, _08124_, _08127_);
  xor g_13966_(_08051_, _08127_, _08128_);
  not g_13967_(_08128_, _08130_);
  or g_13968_(_08014_, _08130_, _08131_);
  xor g_13969_(_08014_, _08128_, _08132_);
  or g_13970_(_07977_, _08132_, _08133_);
  xor g_13971_(_07978_, _08132_, _08134_);
  or g_13972_(_07939_, _08134_, _08135_);
  xor g_13973_(_07940_, _08134_, _08136_);
  or g_13974_(_07902_, _08136_, _08137_);
  xor g_13975_(_07903_, _08136_, _08138_);
  or g_13976_(_07864_, _08138_, _08139_);
  xor g_13977_(_07866_, _08138_, _08141_);
  or g_13978_(_07827_, _08141_, _08142_);
  xor g_13979_(_07828_, _08141_, _08143_);
  or g_13980_(_07790_, _08143_, _08144_);
  xor g_13981_(_07791_, _08143_, _08145_);
  or g_13982_(_07753_, _08145_, _08146_);
  xor g_13983_(_07753_, _08145_, _08147_);
  not g_13984_(_08147_, _08148_);
  or g_13985_(_07717_, _08148_, _08149_);
  xor g_13986_(_07717_, _08147_, _08150_);
  not g_13987_(_08150_, _08152_);
  or g_13988_(_07682_, _08150_, _08153_);
  xor g_13989_(_07682_, _08150_, _08154_);
  xor g_13990_(_07682_, _08152_, _08155_);
  or g_13991_(_07649_, _08155_, _08156_);
  xor g_13992_(_07649_, _08154_, _08157_);
  or g_13993_(_07615_, _08157_, _08158_);
  xor g_13994_(_07616_, _08157_, _08159_);
  or g_13995_(_07581_, _08159_, _08160_);
  xor g_13996_(_07582_, _08159_, _08161_);
  or g_13997_(_07548_, _08161_, _08163_);
  xor g_13998_(_07548_, _08161_, _08164_);
  not g_13999_(_08164_, _08165_);
  or g_14000_(_07515_, _08165_, _08166_);
  xor g_14001_(_07515_, _08164_, _08167_);
  not g_14002_(_08167_, _08168_);
  or g_14003_(_07482_, _08167_, _08169_);
  xor g_14004_(_07482_, _08167_, _08170_);
  xor g_14005_(_07482_, _08168_, _08171_);
  or g_14006_(_07449_, _08171_, _08172_);
  xor g_14007_(_07449_, _08170_, _08174_);
  or g_14008_(_07415_, _08174_, _08175_);
  xor g_14009_(_07416_, _08174_, _08176_);
  or g_14010_(_07382_, _08176_, _08177_);
  xor g_14011_(_07382_, _08176_, _08178_);
  not g_14012_(_08178_, _08179_);
  or g_14013_(_07349_, _08179_, _08180_);
  xor g_14014_(_07349_, _08178_, _08181_);
  or g_14015_(_07315_, _08181_, _08182_);
  xor g_14016_(_07316_, _08181_, _08183_);
  or g_14017_(_07281_, _08183_, _08185_);
  xor g_14018_(_07282_, _08183_, _08186_);
  or g_14019_(_07248_, _08186_, _08187_);
  xor g_14020_(_07248_, _08186_, _08188_);
  not g_14021_(_08188_, _08189_);
  or g_14022_(_07215_, _08189_, _08190_);
  not g_14023_(_08190_, _08191_);
  xor g_14024_(_07215_, _08188_, _08192_);
  or g_14025_(_07181_, _08192_, _08193_);
  not g_14026_(_08193_, _08194_);
  xor g_14027_(_07182_, _08192_, _08196_);
  or g_14028_(_07148_, _08196_, _08197_);
  not g_14029_(_08197_, _08198_);
  and g_14030_(_07148_, _08196_, _08199_);
  xor g_14031_(_07148_, _08196_, _08200_);
  or g_14032_(_08198_, _08199_, _08201_);
  or g_14033_(_07115_, _08201_, _08202_);
  xor g_14034_(_07115_, _08200_, _08203_);
  or g_14035_(_07081_, _08203_, _08204_);
  xor g_14036_(_07082_, _08203_, _08205_);
  or g_14037_(_07047_, _08205_, _08207_);
  xor g_14038_(_07048_, _08205_, _08208_);
  not g_14039_(_08208_, _08209_);
  or g_14040_(_07014_, _08208_, _08210_);
  xor g_14041_(_07014_, _08208_, _08211_);
  xor g_14042_(_07014_, _08209_, _08212_);
  or g_14043_(_06981_, _08212_, _08213_);
  xor g_14044_(_06981_, _08211_, _08214_);
  or g_14045_(_06948_, _08214_, _08215_);
  not g_14046_(_08215_, _08216_);
  xor g_14047_(_06948_, _08214_, _08218_);
  not g_14048_(_08218_, _08219_);
  and g_14049_(_06915_, _08218_, _08220_);
  or g_14050_(_06914_, _08219_, _08221_);
  xor g_14051_(_06914_, _08218_, _08222_);
  or g_14052_(_06880_, _08222_, _08223_);
  xor g_14053_(_06881_, _08222_, _08224_);
  or g_14054_(_06846_, _08224_, _08225_);
  xor g_14055_(_06847_, _08224_, _08226_);
  or g_14056_(_06812_, _08226_, _08227_);
  xor g_14057_(_06813_, _08226_, _08229_);
  or g_14058_(_06779_, _08229_, _08230_);
  not g_14059_(_08230_, _08231_);
  and g_14060_(_06779_, _08229_, _08232_);
  xor g_14061_(_06779_, _08229_, _08233_);
  or g_14062_(_08231_, _08232_, _08234_);
  or g_14063_(_06746_, _08234_, _08235_);
  xor g_14064_(_06746_, _08233_, _08236_);
  or g_14065_(_06712_, _08236_, _08237_);
  not g_14066_(_08237_, _08238_);
  xor g_14067_(_06713_, _08236_, _08240_);
  or g_14068_(_06678_, _08240_, _08241_);
  xor g_14069_(_06678_, _08240_, _08242_);
  xor g_14070_(_06679_, _08240_, _08243_);
  or g_14071_(_06645_, _08243_, _08244_);
  xor g_14072_(_06645_, _08242_, _08245_);
  or g_14073_(_06611_, _08245_, _08246_);
  xor g_14074_(_06612_, _08245_, _08247_);
  not g_14075_(_08247_, _08248_);
  or g_14076_(_06578_, _08247_, _08249_);
  not g_14077_(_08249_, _08251_);
  xor g_14078_(_06578_, _08247_, _08252_);
  xor g_14079_(_06578_, _08248_, _08253_);
  or g_14080_(_06545_, _08253_, _08254_);
  xor g_14081_(_06545_, _08252_, _08255_);
  or g_14082_(_06511_, _08255_, _08256_);
  xor g_14083_(_06512_, _08255_, _08257_);
  or g_14084_(_06477_, _08257_, _08258_);
  xor g_14085_(_06478_, _08257_, _08259_);
  or g_14086_(_06443_, _08259_, _08260_);
  xor g_14087_(_06443_, _08259_, _08262_);
  xor g_14088_(_06444_, _08259_, _08263_);
  and g_14089_(_06410_, _08262_, _08264_);
  or g_14090_(_06409_, _08263_, _08265_);
  xor g_14091_(_06410_, _08262_, _08266_);
  xor g_14092_(_06409_, _08262_, _08267_);
  or g_14093_(_06376_, _08267_, _08268_);
  xor g_14094_(_06376_, _08266_, _08269_);
  or g_14095_(_06342_, _08269_, _08270_);
  xor g_14096_(_06343_, _08269_, _08271_);
  not g_14097_(_08271_, _08273_);
  or g_14098_(_06309_, _08271_, _08274_);
  xor g_14099_(_06309_, _08271_, _08275_);
  xor g_14100_(_06309_, _08273_, _08276_);
  or g_14101_(_06276_, _08276_, _08277_);
  xor g_14102_(_06276_, _08275_, _08278_);
  or g_14103_(_06242_, _08278_, _08279_);
  xor g_14104_(_06243_, _08278_, _08280_);
  or g_14105_(_06208_, _08280_, _08281_);
  xor g_14106_(_06209_, _08280_, _08282_);
  or g_14107_(_06174_, _08282_, _08284_);
  xor g_14108_(_06175_, _08282_, _08285_);
  or g_14109_(_06140_, _08285_, _08286_);
  not g_14110_(_08286_, _08287_);
  xor g_14111_(_06141_, _08285_, _08288_);
  not g_14112_(_08288_, _08289_);
  or g_14113_(_06107_, _08288_, _08290_);
  xor g_14114_(_06107_, _08288_, _08291_);
  xor g_14115_(_06107_, _08289_, _08292_);
  or g_14116_(_06074_, _08292_, _08293_);
  xor g_14117_(_06074_, _08291_, _08295_);
  not g_14118_(_08295_, _08296_);
  or g_14119_(_06041_, _08295_, _08297_);
  not g_14120_(_08297_, _08298_);
  xor g_14121_(_06041_, _08296_, _08299_);
  not g_14122_(_08299_, _08300_);
  or g_14123_(_06008_, _08299_, _08301_);
  not g_14124_(_08301_, _08302_);
  xor g_14125_(_06008_, _08300_, _08303_);
  not g_14126_(_08303_, _08304_);
  and g_14127_(_05975_, _08304_, _08306_);
  or g_14128_(_05974_, _08303_, _08307_);
  xor g_14129_(_05974_, _08303_, _08308_);
  xor g_14130_(_05975_, _08303_, _08309_);
  and g_14131_(_05941_, _08308_, _08310_);
  or g_14132_(_05940_, _08309_, _08311_);
  xor g_14133_(_05941_, _08308_, _08312_);
  xor g_14134_(_05940_, _08308_, _08313_);
  or g_14135_(_05907_, _08313_, _08314_);
  xor g_14136_(_05907_, _08312_, _08315_);
  not g_14137_(_08315_, _08317_);
  or g_14138_(_05874_, _08315_, _08318_);
  xor g_14139_(_05874_, _08317_, _08319_);
  not g_14140_(_08319_, _08320_);
  or g_14141_(_05841_, _08319_, _08321_);
  xor g_14142_(_05841_, _08319_, _08322_);
  xor g_14143_(_05841_, _08320_, _08323_);
  or g_14144_(_05808_, _08323_, _08324_);
  xor g_14145_(_05808_, _08322_, _08325_);
  not g_14146_(_08325_, _08326_);
  or g_14147_(_05775_, _08325_, _08328_);
  not g_14148_(_08328_, _08329_);
  xor g_14149_(_05775_, _08326_, _08330_);
  or g_14150_(_05742_, _08330_, _08331_);
  xor g_14151_(_05742_, _08330_, _08332_);
  not g_14152_(_08332_, _08333_);
  or g_14153_(_05709_, _08333_, _08334_);
  xor g_14154_(_05709_, _08332_, _08335_);
  or g_14155_(_05675_, _08335_, _08336_);
  xor g_14156_(_05676_, _08335_, _08337_);
  not g_14157_(_08337_, _08339_);
  or g_14158_(_05642_, _08337_, _08340_);
  xor g_14159_(_05642_, _08337_, _08341_);
  xor g_14160_(_05642_, _08339_, _08342_);
  or g_14161_(_05609_, _08342_, _08343_);
  not g_14162_(_08343_, _08344_);
  xor g_14163_(_05609_, _08341_, _08345_);
  or g_14164_(_05575_, _08345_, _08346_);
  xor g_14165_(_05576_, _08345_, _08347_);
  not g_14166_(_08347_, _08348_);
  or g_14167_(_05542_, _08347_, _08350_);
  xor g_14168_(_05542_, _08347_, _08351_);
  xor g_14169_(_05542_, _08348_, _08352_);
  or g_14170_(_05509_, _08352_, _08353_);
  xor g_14171_(_05509_, _08351_, _08354_);
  or g_14172_(_05475_, _08354_, _08355_);
  xor g_14173_(_05475_, _08354_, _08356_);
  xor g_14174_(_05476_, _08354_, _08357_);
  or g_14175_(_05442_, _08357_, _08358_);
  xor g_14176_(_05442_, _08356_, _08359_);
  or g_14177_(_05408_, _08359_, _08361_);
  xor g_14178_(_05409_, _08359_, _08362_);
  or g_14179_(_10254_, _08362_, _08363_);
  xor g_14180_(_10254_, _08362_, _08364_);
  not g_14181_(_08364_, _08365_);
  or g_14182_(_10221_, _08365_, _08366_);
  xor g_14183_(_10221_, _08364_, _08367_);
  not g_14184_(_08367_, _08368_);
  or g_14185_(_10188_, _08367_, _08369_);
  xor g_14186_(_10188_, _08367_, _08370_);
  xor g_14187_(_10188_, _08368_, _08372_);
  or g_14188_(_10155_, _08372_, _08373_);
  xor g_14189_(_10155_, _08370_, _08374_);
  not g_14190_(_08374_, _08375_);
  or g_14191_(_10122_, _08374_, _08376_);
  xor g_14192_(_10122_, _08374_, _08377_);
  xor g_14193_(_10122_, _08375_, _08378_);
  or g_14194_(_10089_, _08378_, _08379_);
  xor g_14195_(_10089_, _08377_, _08380_);
  not g_14196_(_08380_, _08381_);
  or g_14197_(_10056_, _08380_, _08383_);
  not g_14198_(_08383_, _08384_);
  xor g_14199_(_10056_, _08381_, _08385_);
  or g_14200_(_10023_, _08385_, _08386_);
  not g_14201_(_08386_, _08387_);
  xor g_14202_(_10023_, _08385_, _08388_);
  not g_14203_(_08388_, _08389_);
  or g_14204_(_09990_, _08389_, _08390_);
  not g_14205_(_08390_, _08391_);
  xor g_14206_(_09990_, _08388_, _08392_);
  or g_14207_(_09957_, _08392_, _08394_);
  not g_14208_(_08394_, _08395_);
  xor g_14209_(_09957_, _08392_, _08396_);
  not g_14210_(_08396_, _08397_);
  or g_14211_(_09924_, _08397_, _08398_);
  xor g_14212_(_09924_, _08396_, _08399_);
  not g_14213_(_08399_, _08400_);
  or g_14214_(_09891_, _08399_, _08401_);
  not g_14215_(_08401_, _08402_);
  xor g_14216_(_09891_, _08400_, _08403_);
  or g_14217_(_09857_, _08403_, _08405_);
  xor g_14218_(_09858_, _08403_, _08406_);
  or g_14219_(_09823_, _08406_, _08407_);
  xor g_14220_(_09823_, _08406_, _08408_);
  xor g_14221_(_09824_, _08406_, _08409_);
  or g_14222_(_09790_, _08409_, _08410_);
  xor g_14223_(_09790_, _08408_, _08411_);
  not g_14224_(_08411_, _08412_);
  or g_14225_(_09434_, _08411_, _08413_);
  xor g_14226_(_09434_, _08412_, _08414_);
  not g_14227_(_08414_, _08416_);
  or g_14228_(_09072_, _08414_, _08417_);
  xor g_14229_(_09072_, _08414_, _08418_);
  xor g_14230_(_09072_, _08416_, _08419_);
  or g_14231_(_08711_, _08419_, _08420_);
  xor g_14232_(_08711_, _08418_, _08421_);
  or g_14233_(_08349_, _08421_, _08422_);
  xor g_14234_(_08349_, _08421_, out[320]);
  and g_14235_(_08420_, _08422_, _08423_);
  and g_14236_(_08413_, _08417_, _08424_);
  not g_14237_(_08424_, _08426_);
  and g_14238_(_08366_, _08369_, _08427_);
  and g_14239_(_08361_, _08363_, _08428_);
  and g_14240_(_08355_, _08358_, _08429_);
  and g_14241_(_08350_, _08353_, _08430_);
  and g_14242_(_08281_, _08284_, _08431_);
  and g_14243_(_08270_, _08274_, _08432_);
  and g_14244_(_08139_, _08142_, _08433_);
  not g_14245_(_08433_, _08434_);
  and g_14246_(_08050_, _08125_, _08435_);
  or g_14247_(_08126_, _08435_, _08437_);
  not g_14248_(_08437_, _08438_);
  or g_14249_(_08131_, _08437_, _08439_);
  not g_14250_(_08439_, _08440_);
  or g_14251_(_08133_, _08437_, _08441_);
  xor g_14252_(_08133_, _08438_, _08442_);
  and g_14253_(_08131_, _08442_, _08443_);
  or g_14254_(_08440_, _08443_, _08444_);
  not g_14255_(_08444_, _08445_);
  and g_14256_(_08135_, _08137_, _08446_);
  xor g_14257_(_08445_, _08446_, _08448_);
  xor g_14258_(_08434_, _08448_, _08449_);
  xor g_14259_(_08433_, _08448_, _08450_);
  or g_14260_(_08144_, _08449_, _08451_);
  xor g_14261_(_08144_, _08450_, _08452_);
  or g_14262_(_08146_, _08452_, _08453_);
  not g_14263_(_08453_, _08454_);
  and g_14264_(_08146_, _08452_, _08455_);
  or g_14265_(_08454_, _08455_, _08456_);
  not g_14266_(_08456_, _08457_);
  and g_14267_(_08149_, _08153_, _08459_);
  xor g_14268_(_08457_, _08459_, _08460_);
  xor g_14269_(_08456_, _08459_, _08461_);
  and g_14270_(_08156_, _08158_, _08462_);
  or g_14271_(_08460_, _08462_, _08463_);
  xor g_14272_(_08461_, _08462_, _08464_);
  not g_14273_(_08464_, _08465_);
  and g_14274_(_08160_, _08163_, _08466_);
  xor g_14275_(_08465_, _08466_, _08467_);
  or g_14276_(_08160_, _08464_, _08468_);
  or g_14277_(_08163_, _08464_, _08470_);
  or g_14278_(_08166_, _08467_, _08471_);
  xor g_14279_(_08166_, _08467_, _08472_);
  not g_14280_(_08472_, _08473_);
  or g_14281_(_08169_, _08473_, _08474_);
  xor g_14282_(_08169_, _08472_, _08475_);
  not g_14283_(_08475_, _08476_);
  or g_14284_(_08172_, _08475_, _08477_);
  xor g_14285_(_08172_, _08475_, _08478_);
  xor g_14286_(_08172_, _08476_, _08479_);
  or g_14287_(_08175_, _08479_, _08481_);
  xor g_14288_(_08175_, _08478_, _08482_);
  not g_14289_(_08482_, _08483_);
  or g_14290_(_08177_, _08482_, _08484_);
  xor g_14291_(_08177_, _08483_, _08485_);
  not g_14292_(_08485_, _08486_);
  or g_14293_(_08180_, _08485_, _08487_);
  xor g_14294_(_08180_, _08485_, _08488_);
  xor g_14295_(_08180_, _08486_, _08489_);
  or g_14296_(_08182_, _08489_, _08490_);
  xor g_14297_(_08182_, _08488_, _08492_);
  not g_14298_(_08492_, _08493_);
  or g_14299_(_08185_, _08492_, _08494_);
  xor g_14300_(_08185_, _08492_, _08495_);
  xor g_14301_(_08185_, _08493_, _08496_);
  or g_14302_(_08187_, _08496_, _08497_);
  xor g_14303_(_08187_, _08495_, _08498_);
  or g_14304_(_08190_, _08498_, _08499_);
  xor g_14305_(_08191_, _08498_, _08500_);
  or g_14306_(_08193_, _08500_, _08501_);
  xor g_14307_(_08194_, _08500_, _08503_);
  or g_14308_(_08197_, _08503_, _08504_);
  xor g_14309_(_08197_, _08503_, _08505_);
  xor g_14310_(_08198_, _08503_, _08506_);
  or g_14311_(_08202_, _08506_, _08507_);
  xor g_14312_(_08202_, _08505_, _08508_);
  not g_14313_(_08508_, _08509_);
  or g_14314_(_08207_, _08508_, _08510_);
  not g_14315_(_08510_, _08511_);
  or g_14316_(_08204_, _08508_, _08512_);
  and g_14317_(_08204_, _08207_, _08514_);
  or g_14318_(_08508_, _08514_, _08515_);
  xor g_14319_(_08508_, _08514_, _08516_);
  not g_14320_(_08516_, _08517_);
  or g_14321_(_08210_, _08517_, _08518_);
  xor g_14322_(_08210_, _08516_, _08519_);
  xor g_14323_(_08509_, _08514_, _08520_);
  xor g_14324_(_08508_, _08514_, _08521_);
  or g_14325_(_08210_, _08520_, _08522_);
  xor g_14326_(_08210_, _08520_, _08523_);
  xor g_14327_(_08210_, _08521_, _08525_);
  or g_14328_(_08213_, _08519_, _08526_);
  or g_14329_(_08213_, _08525_, _08527_);
  xor g_14330_(_08213_, _08523_, _08528_);
  or g_14331_(_08215_, _08528_, _08529_);
  xor g_14332_(_08216_, _08528_, _08530_);
  or g_14333_(_08221_, _08530_, _08531_);
  xor g_14334_(_08220_, _08530_, _08532_);
  not g_14335_(_08532_, _08533_);
  or g_14336_(_08223_, _08532_, _08534_);
  xor g_14337_(_08223_, _08533_, _08536_);
  and g_14338_(_08225_, _08227_, _08537_);
  xor g_14339_(_08536_, _08537_, _08538_);
  not g_14340_(_08538_, _08539_);
  and g_14341_(_08231_, _08538_, _08540_);
  or g_14342_(_08230_, _08539_, _08541_);
  xor g_14343_(_08231_, _08538_, _08542_);
  xor g_14344_(_08230_, _08538_, _08543_);
  or g_14345_(_08235_, _08543_, _08544_);
  xor g_14346_(_08235_, _08542_, _08545_);
  or g_14347_(_08237_, _08545_, _08547_);
  xor g_14348_(_08238_, _08545_, _08548_);
  not g_14349_(_08548_, _08549_);
  or g_14350_(_08241_, _08548_, _08550_);
  not g_14351_(_08550_, _08551_);
  xor g_14352_(_08241_, _08548_, _08552_);
  xor g_14353_(_08241_, _08549_, _08553_);
  and g_14354_(_08244_, _08246_, _08554_);
  xor g_14355_(_08552_, _08554_, _08555_);
  xor g_14356_(_08552_, _08554_, _08556_);
  or g_14357_(_08249_, _08555_, _08558_);
  xor g_14358_(_08249_, _08556_, _08559_);
  xor g_14359_(_08251_, _08556_, _08560_);
  or g_14360_(_08254_, _08560_, _08561_);
  xor g_14361_(_08254_, _08560_, _08562_);
  xor g_14362_(_08254_, _08559_, _08563_);
  or g_14363_(_08256_, _08563_, _08564_);
  xor g_14364_(_08256_, _08562_, _08565_);
  not g_14365_(_08565_, _08566_);
  and g_14366_(_08258_, _08260_, _08567_);
  xor g_14367_(_08566_, _08567_, _08569_);
  not g_14368_(_08569_, _08570_);
  or g_14369_(_08268_, _08569_, _08571_);
  not g_14370_(_08571_, _08572_);
  and g_14371_(_08265_, _08268_, _08573_);
  and g_14372_(_08569_, _08573_, _08574_);
  and g_14373_(_08264_, _08570_, _08575_);
  not g_14374_(_08575_, _08576_);
  or g_14375_(_08574_, _08575_, _08577_);
  or g_14376_(_08572_, _08577_, _08578_);
  not g_14377_(_08578_, _08580_);
  xor g_14378_(_08570_, _08573_, _08581_);
  or g_14379_(_08270_, _08581_, _08582_);
  xor g_14380_(_08432_, _08580_, _08583_);
  not g_14381_(_08583_, _08584_);
  and g_14382_(_08277_, _08279_, _08585_);
  xor g_14383_(_08584_, _08585_, _08586_);
  not g_14384_(_08586_, _08587_);
  or g_14385_(_08277_, _08583_, _08588_);
  or g_14386_(_08279_, _08583_, _08589_);
  not g_14387_(_08589_, _08591_);
  xor g_14388_(_08431_, _08587_, _08592_);
  xor g_14389_(_08431_, _08586_, _08593_);
  and g_14390_(_08286_, _08290_, _08594_);
  or g_14391_(_08290_, _08592_, _08595_);
  and g_14392_(_08287_, _08593_, _08596_);
  or g_14393_(_08286_, _08592_, _08597_);
  xor g_14394_(_08593_, _08594_, _08598_);
  not g_14395_(_08598_, _08599_);
  or g_14396_(_08293_, _08598_, _08600_);
  xor g_14397_(_08293_, _08598_, _08602_);
  xor g_14398_(_08293_, _08599_, _08603_);
  or g_14399_(_08301_, _08603_, _08604_);
  not g_14400_(_08604_, _08605_);
  or g_14401_(_08297_, _08598_, _08606_);
  not g_14402_(_08606_, _08607_);
  and g_14403_(_08297_, _08603_, _08608_);
  or g_14404_(_08298_, _08602_, _08609_);
  and g_14405_(_08606_, _08609_, _08610_);
  or g_14406_(_08607_, _08608_, _08611_);
  and g_14407_(_08301_, _08611_, _08613_);
  or g_14408_(_08302_, _08610_, _08614_);
  and g_14409_(_08604_, _08614_, _08615_);
  or g_14410_(_08605_, _08613_, _08616_);
  and g_14411_(_08310_, _08615_, _08617_);
  and g_14412_(_08307_, _08616_, _08618_);
  or g_14413_(_08303_, _08611_, _08619_);
  and g_14414_(_08306_, _08610_, _08620_);
  or g_14415_(_08618_, _08620_, _08621_);
  and g_14416_(_08311_, _08621_, _08622_);
  or g_14417_(_08617_, _08622_, _08624_);
  not g_14418_(_08624_, _08625_);
  or g_14419_(_08309_, _08616_, _08626_);
  or g_14420_(_08617_, _08620_, _08627_);
  or g_14421_(_08618_, _08627_, _08628_);
  or g_14422_(_08311_, _08615_, _08629_);
  and g_14423_(_08628_, _08629_, _08630_);
  or g_14424_(_08314_, _08624_, _08631_);
  xor g_14425_(_08314_, _08630_, _08632_);
  xor g_14426_(_08314_, _08625_, _08633_);
  or g_14427_(_08321_, _08633_, _08635_);
  xor g_14428_(_08321_, _08632_, _08636_);
  and g_14429_(_08318_, _08636_, _08637_);
  or g_14430_(_08318_, _08624_, _08638_);
  not g_14431_(_08638_, _08639_);
  or g_14432_(_08637_, _08639_, _08640_);
  not g_14433_(_08640_, _08641_);
  or g_14434_(_08324_, _08640_, _08642_);
  xor g_14435_(_08324_, _08640_, _08643_);
  xor g_14436_(_08324_, _08641_, _08644_);
  and g_14437_(_08329_, _08643_, _08646_);
  not g_14438_(_08646_, _08647_);
  xor g_14439_(_08328_, _08643_, _08648_);
  not g_14440_(_08648_, _08649_);
  or g_14441_(_08334_, _08648_, _08650_);
  not g_14442_(_08650_, _08651_);
  or g_14443_(_08331_, _08644_, _08652_);
  xor g_14444_(_08331_, _08649_, _08653_);
  and g_14445_(_08334_, _08653_, _08654_);
  or g_14446_(_08651_, _08654_, _08655_);
  and g_14447_(_08336_, _08340_, _08657_);
  xor g_14448_(_08655_, _08657_, _08658_);
  not g_14449_(_08658_, _08659_);
  and g_14450_(_08343_, _08346_, _08660_);
  and g_14451_(_08344_, _08658_, _08661_);
  or g_14452_(_08343_, _08659_, _08662_);
  or g_14453_(_08346_, _08659_, _08663_);
  xor g_14454_(_08658_, _08660_, _08664_);
  xor g_14455_(_08658_, _08660_, _08665_);
  not g_14456_(_08665_, _08666_);
  xor g_14457_(_08430_, _08666_, _08668_);
  xor g_14458_(_08430_, _08665_, _08669_);
  xor g_14459_(_08429_, _08669_, _08670_);
  not g_14460_(_08670_, _08671_);
  xor g_14461_(_08428_, _08671_, _08672_);
  not g_14462_(_08672_, _08673_);
  xor g_14463_(_08427_, _08673_, _08674_);
  and g_14464_(_08373_, _08376_, _08675_);
  xor g_14465_(_08427_, _08673_, _08676_);
  not g_14466_(_08676_, _08677_);
  or g_14467_(_08376_, _08674_, _08679_);
  or g_14468_(_08373_, _08674_, _08680_);
  xor g_14469_(_08675_, _08676_, _08681_);
  xor g_14470_(_08675_, _08677_, _08682_);
  or g_14471_(_08379_, _08682_, _08683_);
  xor g_14472_(_08379_, _08682_, _08684_);
  xor g_14473_(_08379_, _08681_, _08685_);
  and g_14474_(_08383_, _08685_, _08686_);
  or g_14475_(_08384_, _08684_, _08687_);
  or g_14476_(_08383_, _08682_, _08688_);
  not g_14477_(_08688_, _08690_);
  and g_14478_(_08687_, _08688_, _08691_);
  or g_14479_(_08686_, _08690_, _08692_);
  or g_14480_(_08390_, _08692_, _08693_);
  not g_14481_(_08693_, _08694_);
  or g_14482_(_08386_, _08685_, _08695_);
  not g_14483_(_08695_, _08696_);
  and g_14484_(_08386_, _08692_, _08697_);
  or g_14485_(_08387_, _08691_, _08698_);
  and g_14486_(_08695_, _08698_, _08699_);
  or g_14487_(_08696_, _08697_, _08701_);
  and g_14488_(_08390_, _08701_, _08702_);
  or g_14489_(_08391_, _08699_, _08703_);
  and g_14490_(_08693_, _08703_, _08704_);
  or g_14491_(_08694_, _08702_, _08705_);
  and g_14492_(_08394_, _08398_, _08706_);
  xor g_14493_(_08704_, _08706_, _08707_);
  or g_14494_(_08401_, _08707_, _08708_);
  xor g_14495_(_08401_, _08707_, _08709_);
  xor g_14496_(_08402_, _08707_, _08710_);
  or g_14497_(_08405_, _08710_, _08712_);
  xor g_14498_(_08405_, _08710_, _08713_);
  xor g_14499_(_08405_, _08709_, _08714_);
  or g_14500_(_08407_, _08714_, _08715_);
  not g_14501_(_08715_, _08716_);
  or g_14502_(_08410_, _08714_, _08717_);
  not g_14503_(_08717_, _08718_);
  xor g_14504_(_08410_, _08713_, _08719_);
  and g_14505_(_08407_, _08719_, _08720_);
  or g_14506_(_08716_, _08720_, _08721_);
  xor g_14507_(_08426_, _08721_, _08723_);
  xor g_14508_(_08423_, _08723_, out[321]);
  or g_14509_(_08422_, _08723_, _08724_);
  or g_14510_(_08420_, _08723_, _08725_);
  not g_14511_(_08725_, _08726_);
  or g_14512_(_08417_, _08721_, _08727_);
  not g_14513_(_08727_, _08728_);
  or g_14514_(_08398_, _08705_, _08729_);
  not g_14515_(_08729_, _08730_);
  and g_14516_(_08395_, _08704_, _08731_);
  or g_14517_(_08369_, _08672_, _08733_);
  not g_14518_(_08733_, _08734_);
  or g_14519_(_08366_, _08672_, _08735_);
  or g_14520_(_08363_, _08670_, _08736_);
  or g_14521_(_08358_, _08668_, _08737_);
  or g_14522_(_08355_, _08668_, _08738_);
  or g_14523_(_08340_, _08655_, _08739_);
  or g_14524_(_08336_, _08653_, _08740_);
  and g_14525_(_08635_, _08642_, _08741_);
  or g_14526_(_08284_, _08586_, _08742_);
  or g_14527_(_08260_, _08565_, _08744_);
  or g_14528_(_08258_, _08565_, _08745_);
  not g_14529_(_08745_, _08746_);
  or g_14530_(_08246_, _08553_, _08747_);
  or g_14531_(_08244_, _08548_, _08748_);
  and g_14532_(_08518_, _08526_, _08749_);
  and g_14533_(_08504_, _08507_, _08750_);
  and g_14534_(_08499_, _08501_, _08751_);
  and g_14535_(_08494_, _08497_, _08752_);
  not g_14536_(_08752_, _08753_);
  or g_14537_(_08153_, _08456_, _08755_);
  or g_14538_(_08142_, _08448_, _08756_);
  or g_14539_(_08139_, _08448_, _08757_);
  not g_14540_(_08757_, _08758_);
  or g_14541_(_08137_, _08443_, _08759_);
  and g_14542_(_08439_, _08441_, _08760_);
  or g_14543_(_08135_, _08444_, _08761_);
  and g_14544_(_08760_, _08761_, _08762_);
  and g_14545_(_08759_, _08762_, _08763_);
  or g_14546_(_08757_, _08763_, _08764_);
  xor g_14547_(_08757_, _08763_, _08766_);
  xor g_14548_(_08758_, _08763_, _08767_);
  or g_14549_(_08756_, _08767_, _08768_);
  xor g_14550_(_08756_, _08766_, _08769_);
  not g_14551_(_08769_, _08770_);
  or g_14552_(_08451_, _08769_, _08771_);
  xor g_14553_(_08451_, _08770_, _08772_);
  and g_14554_(_08149_, _08453_, _08773_);
  or g_14555_(_08455_, _08773_, _08774_);
  not g_14556_(_08774_, _08775_);
  or g_14557_(_08772_, _08774_, _08777_);
  xor g_14558_(_08772_, _08774_, _08778_);
  xor g_14559_(_08772_, _08775_, _08779_);
  or g_14560_(_08755_, _08779_, _08780_);
  xor g_14561_(_08755_, _08778_, _08781_);
  not g_14562_(_08781_, _08782_);
  or g_14563_(_08463_, _08781_, _08783_);
  xor g_14564_(_08463_, _08781_, _08784_);
  xor g_14565_(_08463_, _08782_, _08785_);
  or g_14566_(_08468_, _08785_, _08786_);
  not g_14567_(_08786_, _08788_);
  xor g_14568_(_08468_, _08784_, _08789_);
  not g_14569_(_08789_, _08790_);
  or g_14570_(_08470_, _08789_, _08791_);
  xor g_14571_(_08470_, _08789_, _08792_);
  xor g_14572_(_08470_, _08790_, _08793_);
  and g_14573_(_08471_, _08474_, _08794_);
  or g_14574_(_08793_, _08794_, _08795_);
  xor g_14575_(_08793_, _08794_, _08796_);
  xor g_14576_(_08792_, _08794_, _08797_);
  or g_14577_(_08477_, _08797_, _08799_);
  xor g_14578_(_08477_, _08796_, _08800_);
  not g_14579_(_08800_, _08801_);
  and g_14580_(_08481_, _08484_, _08802_);
  or g_14581_(_08484_, _08800_, _08803_);
  or g_14582_(_08481_, _08800_, _08804_);
  xor g_14583_(_08801_, _08802_, _08805_);
  not g_14584_(_08805_, _08806_);
  and g_14585_(_08487_, _08490_, _08807_);
  xor g_14586_(_08806_, _08807_, _08808_);
  xor g_14587_(_08753_, _08808_, _08810_);
  not g_14588_(_08810_, _08811_);
  or g_14589_(_08490_, _08805_, _08812_);
  or g_14590_(_08487_, _08805_, _08813_);
  xor g_14591_(_08751_, _08811_, _08814_);
  xor g_14592_(_08750_, _08814_, _08815_);
  not g_14593_(_08815_, _08816_);
  xor g_14594_(_08515_, _08815_, _08817_);
  not g_14595_(_08817_, _08818_);
  or g_14596_(_08749_, _08817_, _08819_);
  xor g_14597_(_08749_, _08818_, _08821_);
  not g_14598_(_08821_, _08822_);
  or g_14599_(_08529_, _08821_, _08823_);
  xor g_14600_(_08529_, _08821_, _08824_);
  xor g_14601_(_08529_, _08822_, _08825_);
  and g_14602_(_08522_, _08527_, _08826_);
  xor g_14603_(_08817_, _08826_, _08827_);
  xor g_14604_(_08529_, _08827_, _08828_);
  or g_14605_(_08512_, _08816_, _08829_);
  and g_14606_(_08511_, _08815_, _08830_);
  not g_14607_(_08830_, _08832_);
  or g_14608_(_08531_, _08825_, _08833_);
  xor g_14609_(_08531_, _08828_, _08834_);
  xor g_14610_(_08531_, _08824_, _08835_);
  or g_14611_(_08534_, _08835_, _08836_);
  not g_14612_(_08836_, _08837_);
  xor g_14613_(_08534_, _08834_, _08838_);
  or g_14614_(_08225_, _08532_, _08839_);
  not g_14615_(_08839_, _08840_);
  or g_14616_(_08838_, _08839_, _08841_);
  xor g_14617_(_08838_, _08839_, _08843_);
  xor g_14618_(_08838_, _08840_, _08844_);
  or g_14619_(_08227_, _08536_, _08845_);
  or g_14620_(_08844_, _08845_, _08846_);
  xor g_14621_(_08843_, _08845_, _08847_);
  or g_14622_(_08541_, _08847_, _08848_);
  not g_14623_(_08848_, _08849_);
  xor g_14624_(_08540_, _08847_, _08850_);
  not g_14625_(_08850_, _08851_);
  and g_14626_(_08544_, _08547_, _08852_);
  xor g_14627_(_08850_, _08852_, _08854_);
  xor g_14628_(_08851_, _08852_, _08855_);
  and g_14629_(_08551_, _08854_, _08856_);
  or g_14630_(_08550_, _08855_, _08857_);
  xor g_14631_(_08550_, _08854_, _08858_);
  or g_14632_(_08544_, _08850_, _08859_);
  xor g_14633_(_08544_, _08850_, _08860_);
  xor g_14634_(_08547_, _08860_, _08861_);
  xor g_14635_(_08550_, _08861_, _08862_);
  or g_14636_(_08748_, _08858_, _08863_);
  not g_14637_(_08863_, _08865_);
  xor g_14638_(_08748_, _08862_, _08866_);
  or g_14639_(_08747_, _08866_, _08867_);
  not g_14640_(_08867_, _08868_);
  xor g_14641_(_08747_, _08866_, _08869_);
  not g_14642_(_08869_, _08870_);
  or g_14643_(_08558_, _08870_, _08871_);
  xor g_14644_(_08558_, _08869_, _08872_);
  not g_14645_(_08872_, _08873_);
  and g_14646_(_08561_, _08564_, _08874_);
  or g_14647_(_08561_, _08872_, _08876_);
  or g_14648_(_08564_, _08872_, _08877_);
  not g_14649_(_08877_, _08878_);
  xor g_14650_(_08872_, _08874_, _08879_);
  xor g_14651_(_08873_, _08874_, _08880_);
  and g_14652_(_08746_, _08879_, _08881_);
  or g_14653_(_08745_, _08880_, _08882_);
  xor g_14654_(_08746_, _08879_, _08883_);
  xor g_14655_(_08745_, _08879_, _08884_);
  or g_14656_(_08744_, _08884_, _08885_);
  xor g_14657_(_08744_, _08883_, _08887_);
  or g_14658_(_08576_, _08887_, _08888_);
  xor g_14659_(_08575_, _08887_, _08889_);
  or g_14660_(_08571_, _08889_, _08890_);
  xor g_14661_(_08571_, _08889_, _08891_);
  not g_14662_(_08891_, _08892_);
  or g_14663_(_08270_, _08578_, _08893_);
  or g_14664_(_08892_, _08893_, _08894_);
  xor g_14665_(_08582_, _08892_, _08895_);
  xor g_14666_(_08582_, _08891_, _08896_);
  or g_14667_(_08274_, _08578_, _08898_);
  or g_14668_(_08896_, _08898_, _08899_);
  not g_14669_(_08899_, _08900_);
  xor g_14670_(_08895_, _08898_, _08901_);
  and g_14671_(_08588_, _08901_, _08902_);
  or g_14672_(_08588_, _08901_, _08903_);
  not g_14673_(_08903_, _08904_);
  or g_14674_(_08902_, _08904_, _08905_);
  not g_14675_(_08905_, _08906_);
  or g_14676_(_08281_, _08586_, _08907_);
  and g_14677_(_08589_, _08907_, _08909_);
  xor g_14678_(_08905_, _08909_, _08910_);
  xor g_14679_(_08906_, _08909_, _08911_);
  or g_14680_(_08742_, _08911_, _08912_);
  not g_14681_(_08912_, _08913_);
  xor g_14682_(_08742_, _08910_, _08914_);
  or g_14683_(_08597_, _08914_, _08915_);
  not g_14684_(_08915_, _08916_);
  xor g_14685_(_08596_, _08914_, _08917_);
  and g_14686_(_08591_, _08906_, _08918_);
  and g_14687_(_08595_, _08917_, _08920_);
  or g_14688_(_08595_, _08917_, _08921_);
  not g_14689_(_08921_, _08922_);
  or g_14690_(_08920_, _08922_, _08923_);
  not g_14691_(_08923_, _08924_);
  or g_14692_(_08600_, _08923_, _08925_);
  xor g_14693_(_08600_, _08924_, _08926_);
  or g_14694_(_08606_, _08926_, _08927_);
  xor g_14695_(_08607_, _08926_, _08928_);
  or g_14696_(_08604_, _08928_, _08929_);
  not g_14697_(_08929_, _08931_);
  xor g_14698_(_08605_, _08928_, _08932_);
  xor g_14699_(_08627_, _08932_, _08933_);
  not g_14700_(_08933_, _08934_);
  or g_14701_(_08631_, _08933_, _08935_);
  xor g_14702_(_08631_, _08934_, _08936_);
  or g_14703_(_08638_, _08936_, _08937_);
  xor g_14704_(_08639_, _08936_, _08938_);
  xor g_14705_(_08741_, _08938_, _08939_);
  not g_14706_(_08939_, _08940_);
  or g_14707_(_08647_, _08940_, _08942_);
  not g_14708_(_08942_, _08943_);
  xor g_14709_(_08646_, _08939_, _08944_);
  not g_14710_(_08944_, _08945_);
  or g_14711_(_08652_, _08945_, _08946_);
  not g_14712_(_08946_, _08947_);
  xor g_14713_(_08652_, _08944_, _08948_);
  or g_14714_(_08650_, _08948_, _08949_);
  xor g_14715_(_08650_, _08948_, _08950_);
  xor g_14716_(_08651_, _08948_, _08951_);
  or g_14717_(_08740_, _08951_, _08953_);
  xor g_14718_(_08740_, _08950_, _08954_);
  not g_14719_(_08954_, _08955_);
  or g_14720_(_08739_, _08954_, _08956_);
  xor g_14721_(_08739_, _08955_, _08957_);
  or g_14722_(_08662_, _08957_, _08958_);
  not g_14723_(_08958_, _08959_);
  xor g_14724_(_08661_, _08957_, _08960_);
  not g_14725_(_08960_, _08961_);
  or g_14726_(_08350_, _08664_, _08962_);
  and g_14727_(_08663_, _08962_, _08964_);
  or g_14728_(_08663_, _08960_, _08965_);
  not g_14729_(_08965_, _08966_);
  xor g_14730_(_08961_, _08964_, _08967_);
  or g_14731_(_08353_, _08664_, _08968_);
  or g_14732_(_08353_, _08665_, _08969_);
  not g_14733_(_08969_, _08970_);
  or g_14734_(_08967_, _08968_, _08971_);
  not g_14735_(_08971_, _08972_);
  xor g_14736_(_08967_, _08970_, _08973_);
  not g_14737_(_08973_, _08975_);
  or g_14738_(_08738_, _08973_, _08976_);
  xor g_14739_(_08738_, _08975_, _08977_);
  not g_14740_(_08977_, _08978_);
  or g_14741_(_08737_, _08977_, _08979_);
  xor g_14742_(_08737_, _08977_, _08980_);
  xor g_14743_(_08737_, _08978_, _08981_);
  or g_14744_(_08361_, _08670_, _08982_);
  or g_14745_(_08981_, _08982_, _08983_);
  xor g_14746_(_08980_, _08982_, _08984_);
  or g_14747_(_08736_, _08984_, _08986_);
  xor g_14748_(_08736_, _08984_, _08987_);
  not g_14749_(_08987_, _08988_);
  or g_14750_(_08735_, _08988_, _08989_);
  xor g_14751_(_08735_, _08987_, _08990_);
  or g_14752_(_08733_, _08990_, _08991_);
  xor g_14753_(_08734_, _08990_, _08992_);
  or g_14754_(_08373_, _08676_, _08993_);
  not g_14755_(_08993_, _08994_);
  or g_14756_(_08680_, _08992_, _08995_);
  xor g_14757_(_08992_, _08994_, _08997_);
  or g_14758_(_08376_, _08676_, _08998_);
  not g_14759_(_08998_, _08999_);
  or g_14760_(_08679_, _08997_, _09000_);
  xor g_14761_(_08997_, _08999_, _09001_);
  and g_14762_(_08683_, _08688_, _09002_);
  not g_14763_(_09002_, _09003_);
  or g_14764_(_08688_, _09001_, _09004_);
  or g_14765_(_08683_, _09001_, _09005_);
  xor g_14766_(_09001_, _09003_, _09006_);
  or g_14767_(_08695_, _09006_, _09008_);
  xor g_14768_(_08696_, _09006_, _09009_);
  or g_14769_(_08693_, _09009_, _09010_);
  xor g_14770_(_08693_, _09009_, _09011_);
  xor g_14771_(_08694_, _09009_, _09012_);
  or g_14772_(_08731_, _09011_, _09013_);
  or g_14773_(_08394_, _08701_, _09014_);
  or g_14774_(_09012_, _09014_, _09015_);
  and g_14775_(_09013_, _09015_, _09016_);
  not g_14776_(_09016_, _09017_);
  and g_14777_(_08730_, _09016_, _09019_);
  or g_14778_(_08729_, _09017_, _09020_);
  xor g_14779_(_08729_, _09016_, _09021_);
  not g_14780_(_09021_, _09022_);
  and g_14781_(_08708_, _08712_, _09023_);
  xor g_14782_(_09022_, _09023_, _09024_);
  or g_14783_(_08715_, _09024_, _09025_);
  xor g_14784_(_08715_, _09024_, _09026_);
  xor g_14785_(_08716_, _09024_, _09027_);
  or g_14786_(_08413_, _08721_, _09028_);
  not g_14787_(_09028_, _09030_);
  or g_14788_(_09027_, _09028_, _09031_);
  not g_14789_(_09031_, _09032_);
  and g_14790_(_08718_, _09026_, _09033_);
  not g_14791_(_09033_, _09034_);
  xor g_14792_(_08718_, _09026_, _09035_);
  xor g_14793_(_08717_, _09026_, _09036_);
  and g_14794_(_09028_, _09036_, _09037_);
  or g_14795_(_09030_, _09035_, _09038_);
  and g_14796_(_09031_, _09038_, _09039_);
  or g_14797_(_09032_, _09037_, _09041_);
  and g_14798_(_08728_, _09039_, _09042_);
  or g_14799_(_08727_, _09041_, _09043_);
  xor g_14800_(_08727_, _09039_, _09044_);
  not g_14801_(_09044_, _09045_);
  and g_14802_(_08726_, _09045_, _09046_);
  or g_14803_(_08725_, _09044_, _09047_);
  xor g_14804_(_08726_, _09044_, _09048_);
  or g_14805_(_08724_, _09048_, _09049_);
  xor g_14806_(_08724_, _09048_, out[322]);
  or g_14807_(_08712_, _09021_, _09051_);
  not g_14808_(_09051_, _09052_);
  or g_14809_(_08708_, _09021_, _09053_);
  not g_14810_(_09053_, _09054_);
  or g_14811_(_08960_, _08962_, _09055_);
  or g_14812_(_08642_, _08936_, _09056_);
  not g_14813_(_09056_, _09057_);
  or g_14814_(_08635_, _08938_, _09058_);
  or g_14815_(_08626_, _08932_, _09059_);
  not g_14816_(_09059_, _09060_);
  or g_14817_(_05940_, _09059_, _09062_);
  or g_14818_(_08619_, _08932_, _09063_);
  not g_14819_(_09063_, _09064_);
  or g_14820_(_08905_, _08907_, _09065_);
  not g_14821_(_09065_, _09066_);
  or g_14822_(_08547_, _08850_, _09067_);
  not g_14823_(_09067_, _09068_);
  or g_14824_(_08856_, _09068_, _09069_);
  or g_14825_(_08507_, _08814_, _09070_);
  not g_14826_(_09070_, _09071_);
  or g_14827_(_08504_, _08814_, _09073_);
  not g_14828_(_09073_, _09074_);
  or g_14829_(_08501_, _08810_, _09075_);
  or g_14830_(_08499_, _08810_, _09076_);
  or g_14831_(_08497_, _08808_, _09077_);
  or g_14832_(_08494_, _08808_, _09078_);
  and g_14833_(_08799_, _08804_, _09079_);
  not g_14834_(_09079_, _09080_);
  and g_14835_(_08764_, _08768_, _09081_);
  and g_14836_(_08771_, _09081_, _09082_);
  and g_14837_(_08777_, _09082_, _09084_);
  and g_14838_(_08780_, _09084_, _09085_);
  and g_14839_(_08783_, _09085_, _09086_);
  or g_14840_(_08786_, _09086_, _09087_);
  xor g_14841_(_08786_, _09086_, _09088_);
  xor g_14842_(_08788_, _09086_, _09089_);
  or g_14843_(_08791_, _09089_, _09090_);
  xor g_14844_(_08791_, _09088_, _09091_);
  not g_14845_(_09091_, _09092_);
  xor g_14846_(_08795_, _09092_, _09093_);
  or g_14847_(_09079_, _09093_, _09095_);
  xor g_14848_(_09079_, _09093_, _09096_);
  xor g_14849_(_09080_, _09093_, _09097_);
  or g_14850_(_08803_, _09097_, _09098_);
  xor g_14851_(_08803_, _09096_, _09099_);
  not g_14852_(_09099_, _09100_);
  or g_14853_(_08813_, _09099_, _09101_);
  xor g_14854_(_08813_, _09100_, _09102_);
  not g_14855_(_09102_, _09103_);
  or g_14856_(_08812_, _09102_, _09104_);
  xor g_14857_(_08812_, _09102_, _09106_);
  xor g_14858_(_08812_, _09103_, _09107_);
  or g_14859_(_09078_, _09107_, _09108_);
  xor g_14860_(_09078_, _09106_, _09109_);
  not g_14861_(_09109_, _09110_);
  or g_14862_(_09077_, _09109_, _09111_);
  xor g_14863_(_09077_, _09110_, _09112_);
  not g_14864_(_09112_, _09113_);
  or g_14865_(_09076_, _09112_, _09114_);
  xor g_14866_(_09076_, _09113_, _09115_);
  or g_14867_(_09075_, _09115_, _09117_);
  xor g_14868_(_09075_, _09115_, _09118_);
  and g_14869_(_09074_, _09118_, _09119_);
  xor g_14870_(_09073_, _09118_, _09120_);
  or g_14871_(_09070_, _09120_, _09121_);
  xor g_14872_(_09071_, _09120_, _09122_);
  not g_14873_(_09122_, _09123_);
  or g_14874_(_08829_, _09122_, _09124_);
  xor g_14875_(_08829_, _09123_, _09125_);
  or g_14876_(_08832_, _09125_, _09126_);
  xor g_14877_(_08832_, _09125_, _09128_);
  xor g_14878_(_08819_, _09128_, _09129_);
  and g_14879_(_08823_, _08833_, _09130_);
  not g_14880_(_09130_, _09131_);
  or g_14881_(_09129_, _09130_, _09132_);
  xor g_14882_(_09129_, _09131_, _09133_);
  or g_14883_(_08836_, _09133_, _09134_);
  xor g_14884_(_08837_, _09133_, _09135_);
  and g_14885_(_08841_, _08846_, _09136_);
  not g_14886_(_09136_, _09137_);
  xor g_14887_(_09135_, _09137_, _09139_);
  xor g_14888_(_09135_, _09136_, _09140_);
  and g_14889_(_08848_, _08859_, _09141_);
  xor g_14890_(_09140_, _09141_, _09142_);
  xor g_14891_(_09069_, _09142_, _09143_);
  or g_14892_(_08863_, _09143_, _09144_);
  xor g_14893_(_08865_, _09143_, _09145_);
  or g_14894_(_08867_, _09145_, _09146_);
  xor g_14895_(_08868_, _09145_, _09147_);
  not g_14896_(_09147_, _09148_);
  and g_14897_(_08871_, _08876_, _09150_);
  xor g_14898_(_09148_, _09150_, _09151_);
  xor g_14899_(_09147_, _09150_, _09152_);
  or g_14900_(_08882_, _09151_, _09153_);
  or g_14901_(_08878_, _09152_, _09154_);
  or g_14902_(_08881_, _09154_, _09155_);
  or g_14903_(_08877_, _09151_, _09156_);
  and g_14904_(_09155_, _09156_, _09157_);
  and g_14905_(_09153_, _09157_, _09158_);
  not g_14906_(_09158_, _09159_);
  or g_14907_(_08885_, _09159_, _09161_);
  xor g_14908_(_08885_, _09158_, _09162_);
  not g_14909_(_09162_, _09163_);
  or g_14910_(_08888_, _09162_, _09164_);
  xor g_14911_(_08888_, _09162_, _09165_);
  xor g_14912_(_08888_, _09163_, _09166_);
  and g_14913_(_08890_, _08894_, _09167_);
  xor g_14914_(_09166_, _09167_, _09168_);
  xor g_14915_(_09165_, _09167_, _09169_);
  and g_14916_(_08904_, _09168_, _09170_);
  and g_14917_(_08899_, _09169_, _09172_);
  and g_14918_(_08903_, _09172_, _09173_);
  and g_14919_(_08900_, _09168_, _09174_);
  or g_14920_(_09173_, _09174_, _09175_);
  or g_14921_(_09170_, _09175_, _09176_);
  not g_14922_(_09176_, _09177_);
  and g_14923_(_08918_, _09177_, _09178_);
  xor g_14924_(_08918_, _09176_, _09179_);
  or g_14925_(_09065_, _09179_, _09180_);
  not g_14926_(_09180_, _09181_);
  xor g_14927_(_09066_, _09179_, _09183_);
  or g_14928_(_08915_, _09183_, _09184_);
  not g_14929_(_09184_, _09185_);
  or g_14930_(_08912_, _09183_, _09186_);
  xor g_14931_(_08912_, _09183_, _09187_);
  xor g_14932_(_08913_, _09183_, _09188_);
  and g_14933_(_08915_, _09188_, _09189_);
  or g_14934_(_08916_, _09187_, _09190_);
  and g_14935_(_09184_, _09190_, _09191_);
  or g_14936_(_09185_, _09189_, _09192_);
  and g_14937_(_08922_, _09191_, _09194_);
  xor g_14938_(_08921_, _09191_, _09195_);
  or g_14939_(_08927_, _09195_, _09196_);
  not g_14940_(_09196_, _09197_);
  and g_14941_(_08925_, _09195_, _09198_);
  or g_14942_(_08925_, _09192_, _09199_);
  not g_14943_(_09199_, _09200_);
  or g_14944_(_09198_, _09200_, _09201_);
  and g_14945_(_08927_, _09201_, _09202_);
  or g_14946_(_09197_, _09202_, _09203_);
  xor g_14947_(_08931_, _09203_, _09205_);
  xor g_14948_(_08929_, _09203_, _09206_);
  and g_14949_(_09064_, _09206_, _09207_);
  or g_14950_(_09063_, _09205_, _09208_);
  and g_14951_(_05975_, _09207_, _09209_);
  or g_14952_(_05974_, _09208_, _09210_);
  or g_14953_(_05974_, _09063_, _09211_);
  not g_14954_(_09211_, _09212_);
  and g_14955_(_09205_, _09211_, _09213_);
  or g_14956_(_09206_, _09212_, _09214_);
  and g_14957_(_09210_, _09214_, _09216_);
  or g_14958_(_09209_, _09213_, _09217_);
  and g_14959_(_09062_, _09217_, _09218_);
  and g_14960_(_09060_, _09216_, _09219_);
  or g_14961_(_09059_, _09217_, _09220_);
  and g_14962_(_05941_, _09219_, _09221_);
  or g_14963_(_05940_, _09220_, _09222_);
  or g_14964_(_09218_, _09221_, _09223_);
  and g_14965_(_08935_, _08937_, _09224_);
  not g_14966_(_09224_, _09225_);
  xor g_14967_(_09223_, _09224_, _09227_);
  xor g_14968_(_09223_, _09225_, _09228_);
  or g_14969_(_09058_, _09228_, _09229_);
  not g_14970_(_09229_, _09230_);
  xor g_14971_(_09058_, _09227_, _09231_);
  or g_14972_(_09056_, _09231_, _09232_);
  not g_14973_(_09232_, _09233_);
  xor g_14974_(_09056_, _09231_, _09234_);
  xor g_14975_(_09057_, _09231_, _09235_);
  and g_14976_(_08942_, _09235_, _09236_);
  and g_14977_(_08946_, _09236_, _09238_);
  and g_14978_(_08947_, _09234_, _09239_);
  or g_14979_(_08946_, _09235_, _09240_);
  and g_14980_(_08943_, _09234_, _09241_);
  or g_14981_(_08942_, _09235_, _09242_);
  or g_14982_(_09239_, _09241_, _09243_);
  or g_14983_(_09238_, _09243_, _09244_);
  not g_14984_(_09244_, _09245_);
  and g_14985_(_08949_, _08953_, _09246_);
  xor g_14986_(_09244_, _09246_, _09247_);
  xor g_14987_(_09245_, _09246_, _09249_);
  or g_14988_(_08956_, _09249_, _09250_);
  xor g_14989_(_08956_, _09247_, _09251_);
  or g_14990_(_08958_, _09251_, _09252_);
  xor g_14991_(_08959_, _09251_, _09253_);
  or g_14992_(_08965_, _09253_, _09254_);
  xor g_14993_(_08966_, _09253_, _09255_);
  or g_14994_(_09055_, _09255_, _09256_);
  not g_14995_(_09256_, _09257_);
  xor g_14996_(_09055_, _09255_, _09258_);
  and g_14997_(_08972_, _09258_, _09260_);
  not g_14998_(_09260_, _09261_);
  xor g_14999_(_08972_, _09258_, _09262_);
  xor g_15000_(_08971_, _09258_, _09263_);
  or g_15001_(_08976_, _09263_, _09264_);
  not g_15002_(_09264_, _09265_);
  xor g_15003_(_08976_, _09262_, _09266_);
  not g_15004_(_09266_, _09267_);
  and g_15005_(_08979_, _08983_, _09268_);
  xor g_15006_(_09266_, _09268_, _09269_);
  xor g_15007_(_09267_, _09268_, _09271_);
  or g_15008_(_08986_, _09271_, _09272_);
  xor g_15009_(_08986_, _09269_, _09273_);
  not g_15010_(_09273_, _09274_);
  or g_15011_(_08989_, _09273_, _09275_);
  xor g_15012_(_08989_, _09273_, _09276_);
  xor g_15013_(_08989_, _09274_, _09277_);
  or g_15014_(_08991_, _09277_, _09278_);
  xor g_15015_(_08991_, _09276_, _09279_);
  not g_15016_(_09279_, _09280_);
  or g_15017_(_08995_, _09279_, _09282_);
  and g_15018_(_08995_, _09279_, _09283_);
  xor g_15019_(_08995_, _09279_, _09284_);
  xor g_15020_(_08995_, _09280_, _09285_);
  and g_15021_(_09000_, _09005_, _09286_);
  xor g_15022_(_09284_, _09286_, _09287_);
  not g_15023_(_09287_, _09288_);
  or g_15024_(_09004_, _09287_, _09289_);
  xor g_15025_(_09004_, _09288_, _09290_);
  and g_15026_(_09008_, _09010_, _09291_);
  xor g_15027_(_09290_, _09291_, _09293_);
  not g_15028_(_09293_, _09294_);
  or g_15029_(_09015_, _09294_, _09295_);
  xor g_15030_(_09015_, _09293_, _09296_);
  or g_15031_(_09020_, _09296_, _09297_);
  xor g_15032_(_09019_, _09296_, _09298_);
  or g_15033_(_09053_, _09298_, _09299_);
  xor g_15034_(_09054_, _09298_, _09300_);
  or g_15035_(_09051_, _09300_, _09301_);
  xor g_15036_(_09052_, _09300_, _09302_);
  and g_15037_(_09025_, _09302_, _09304_);
  or g_15038_(_09025_, _09302_, _09305_);
  not g_15039_(_09305_, _09306_);
  xor g_15040_(_09025_, _09302_, _09307_);
  or g_15041_(_09304_, _09306_, _09308_);
  and g_15042_(_09033_, _09307_, _09309_);
  or g_15043_(_09034_, _09308_, _09310_);
  xor g_15044_(_09034_, _09307_, _09311_);
  not g_15045_(_09311_, _09312_);
  or g_15046_(_09031_, _09311_, _09313_);
  not g_15047_(_09313_, _09315_);
  xor g_15048_(_09031_, _09311_, _09316_);
  xor g_15049_(_09032_, _09311_, _09317_);
  and g_15050_(_09043_, _09317_, _09318_);
  or g_15051_(_09042_, _09316_, _09319_);
  and g_15052_(_09042_, _09312_, _09320_);
  or g_15053_(_09043_, _09311_, _09321_);
  and g_15054_(_09319_, _09321_, _09322_);
  or g_15055_(_09318_, _09320_, _09323_);
  and g_15056_(_09046_, _09322_, _09324_);
  or g_15057_(_09047_, _09323_, _09326_);
  xor g_15058_(_09047_, _09322_, _09327_);
  or g_15059_(_09049_, _09327_, _09328_);
  not g_15060_(_09328_, _09329_);
  xor g_15061_(_09049_, _09327_, out[323]);
  or g_15062_(_09010_, _09290_, _09330_);
  not g_15063_(_09330_, _09331_);
  or g_15064_(_09008_, _09290_, _09332_);
  not g_15065_(_09332_, _09333_);
  or g_15066_(_09000_, _09283_, _09334_);
  and g_15067_(_09282_, _09334_, _09336_);
  and g_15068_(_09275_, _09278_, _09337_);
  or g_15069_(_08979_, _09266_, _09338_);
  not g_15070_(_09338_, _09339_);
  or g_15071_(_08953_, _09244_, _09340_);
  not g_15072_(_09340_, _09341_);
  or g_15073_(_08949_, _09244_, _09342_);
  not g_15074_(_09342_, _09343_);
  or g_15075_(_08937_, _09223_, _09344_);
  not g_15076_(_09344_, _09345_);
  and g_15077_(_09229_, _09344_, _09347_);
  or g_15078_(_08929_, _09201_, _09348_);
  and g_15079_(_09196_, _09199_, _09349_);
  not g_15080_(_09349_, _09350_);
  or g_15081_(_08894_, _09166_, _09351_);
  or g_15082_(_08876_, _09147_, _09352_);
  or g_15083_(_08857_, _09142_, _09353_);
  or g_15084_(_09067_, _09142_, _09354_);
  or g_15085_(_08859_, _09139_, _09355_);
  and g_15086_(_08849_, _09140_, _09356_);
  not g_15087_(_09356_, _09358_);
  or g_15088_(_08846_, _09135_, _09359_);
  or g_15089_(_08817_, _09125_, _09360_);
  or g_15090_(_08526_, _09360_, _09361_);
  not g_15091_(_09361_, _09362_);
  or g_15092_(_08795_, _09091_, _09363_);
  and g_15093_(_09087_, _09090_, _09364_);
  and g_15094_(_09363_, _09364_, _09365_);
  and g_15095_(_09095_, _09365_, _09366_);
  and g_15096_(_09098_, _09366_, _09367_);
  and g_15097_(_09101_, _09367_, _09369_);
  and g_15098_(_09104_, _09369_, _09370_);
  and g_15099_(_09108_, _09370_, _09371_);
  and g_15100_(_09111_, _09371_, _09372_);
  and g_15101_(_09114_, _09372_, _09373_);
  and g_15102_(_09117_, _09373_, _09374_);
  xor g_15103_(_09119_, _09374_, _09375_);
  and g_15104_(_09121_, _09375_, _09376_);
  and g_15105_(_09124_, _09376_, _09377_);
  not g_15106_(_09377_, _09378_);
  or g_15107_(_08518_, _09360_, _09380_);
  and g_15108_(_09126_, _09380_, _09381_);
  xor g_15109_(_09378_, _09381_, _09382_);
  or g_15110_(_09361_, _09382_, _09383_);
  xor g_15111_(_09362_, _09382_, _09384_);
  not g_15112_(_09384_, _09385_);
  or g_15113_(_09132_, _09384_, _09386_);
  xor g_15114_(_09132_, _09385_, _09387_);
  not g_15115_(_09387_, _09388_);
  or g_15116_(_08841_, _09135_, _09389_);
  and g_15117_(_09134_, _09389_, _09391_);
  or g_15118_(_09387_, _09391_, _09392_);
  xor g_15119_(_09387_, _09391_, _09393_);
  xor g_15120_(_09388_, _09391_, _09394_);
  or g_15121_(_09359_, _09394_, _09395_);
  xor g_15122_(_09359_, _09393_, _09396_);
  or g_15123_(_09358_, _09396_, _09397_);
  xor g_15124_(_09356_, _09396_, _09398_);
  not g_15125_(_09398_, _09399_);
  or g_15126_(_09355_, _09398_, _09400_);
  xor g_15127_(_09355_, _09398_, _09402_);
  xor g_15128_(_09355_, _09399_, _09403_);
  or g_15129_(_09354_, _09403_, _09404_);
  xor g_15130_(_09354_, _09402_, _09405_);
  not g_15131_(_09405_, _09406_);
  or g_15132_(_09353_, _09405_, _09407_);
  xor g_15133_(_09353_, _09406_, _09408_);
  not g_15134_(_09408_, _09409_);
  or g_15135_(_09144_, _09408_, _09410_);
  and g_15136_(_09144_, _09408_, _09411_);
  xor g_15137_(_09144_, _09409_, _09413_);
  not g_15138_(_09413_, _09414_);
  or g_15139_(_08871_, _09147_, _09415_);
  and g_15140_(_09146_, _09415_, _09416_);
  xor g_15141_(_09413_, _09416_, _09417_);
  xor g_15142_(_09414_, _09416_, _09418_);
  or g_15143_(_09352_, _09418_, _09419_);
  xor g_15144_(_09352_, _09417_, _09420_);
  not g_15145_(_09420_, _09421_);
  or g_15146_(_09156_, _09420_, _09422_);
  xor g_15147_(_09156_, _09421_, _09424_);
  not g_15148_(_09424_, _09425_);
  or g_15149_(_09161_, _09424_, _09426_);
  not g_15150_(_09426_, _09427_);
  or g_15151_(_09153_, _09424_, _09428_);
  xor g_15152_(_09153_, _09425_, _09429_);
  and g_15153_(_09161_, _09429_, _09430_);
  or g_15154_(_09427_, _09430_, _09431_);
  not g_15155_(_09431_, _09432_);
  or g_15156_(_08890_, _09166_, _09433_);
  and g_15157_(_09164_, _09433_, _09435_);
  xor g_15158_(_09432_, _09435_, _09436_);
  or g_15159_(_09351_, _09436_, _09437_);
  xor g_15160_(_09351_, _09436_, _09438_);
  and g_15161_(_09174_, _09438_, _09439_);
  or g_15162_(_09174_, _09438_, _09440_);
  xor g_15163_(_09174_, _09438_, _09441_);
  or g_15164_(_09170_, _09178_, _09442_);
  xor g_15165_(_09441_, _09442_, _09443_);
  not g_15166_(_09443_, _09444_);
  or g_15167_(_09186_, _09444_, _09446_);
  and g_15168_(_09181_, _09443_, _09447_);
  xor g_15169_(_09180_, _09443_, _09448_);
  and g_15170_(_09186_, _09448_, _09449_);
  not g_15171_(_09449_, _09450_);
  and g_15172_(_09446_, _09450_, _09451_);
  or g_15173_(_08921_, _09189_, _09452_);
  and g_15174_(_09184_, _09452_, _09453_);
  xor g_15175_(_09451_, _09453_, _09454_);
  or g_15176_(_09349_, _09454_, _09455_);
  xor g_15177_(_09350_, _09454_, _09457_);
  not g_15178_(_09457_, _09458_);
  or g_15179_(_09348_, _09457_, _09459_);
  xor g_15180_(_09348_, _09457_, _09460_);
  xor g_15181_(_09348_, _09458_, _09461_);
  and g_15182_(_09207_, _09460_, _09462_);
  or g_15183_(_09208_, _09461_, _09463_);
  and g_15184_(_05975_, _09462_, _09464_);
  or g_15185_(_05974_, _09463_, _09465_);
  and g_15186_(_09210_, _09461_, _09466_);
  not g_15187_(_09466_, _09468_);
  and g_15188_(_09465_, _09468_, _09469_);
  or g_15189_(_09464_, _09466_, _09470_);
  or g_15190_(_08935_, _09223_, _09471_);
  not g_15191_(_09471_, _09472_);
  and g_15192_(_09222_, _09471_, _09473_);
  xor g_15193_(_09470_, _09473_, _09474_);
  xor g_15194_(_09469_, _09473_, _09475_);
  xor g_15195_(_09347_, _09474_, _09476_);
  xor g_15196_(_09347_, _09475_, _09477_);
  or g_15197_(_09233_, _09477_, _09479_);
  or g_15198_(_09241_, _09479_, _09480_);
  not g_15199_(_09480_, _09481_);
  and g_15200_(_09241_, _09477_, _09482_);
  or g_15201_(_09242_, _09476_, _09483_);
  or g_15202_(_09232_, _09476_, _09484_);
  not g_15203_(_09484_, _09485_);
  and g_15204_(_09483_, _09484_, _09486_);
  or g_15205_(_09482_, _09485_, _09487_);
  and g_15206_(_09480_, _09486_, _09488_);
  or g_15207_(_09481_, _09487_, _09490_);
  or g_15208_(_09240_, _09490_, _09491_);
  not g_15209_(_09491_, _09492_);
  xor g_15210_(_09240_, _09488_, _09493_);
  or g_15211_(_09342_, _09493_, _09494_);
  not g_15212_(_09494_, _09495_);
  xor g_15213_(_09343_, _09493_, _09496_);
  or g_15214_(_09340_, _09496_, _09497_);
  xor g_15215_(_09341_, _09496_, _09498_);
  not g_15216_(_09498_, _09499_);
  and g_15217_(_09250_, _09252_, _09501_);
  or g_15218_(_09498_, _09501_, _09502_);
  xor g_15219_(_09498_, _09501_, _09503_);
  xor g_15220_(_09499_, _09501_, _09504_);
  or g_15221_(_09254_, _09504_, _09505_);
  xor g_15222_(_09254_, _09503_, _09506_);
  not g_15223_(_09506_, _09507_);
  and g_15224_(_09260_, _09507_, _09508_);
  not g_15225_(_09508_, _09509_);
  or g_15226_(_09256_, _09506_, _09510_);
  xor g_15227_(_09256_, _09506_, _09512_);
  xor g_15228_(_09257_, _09506_, _09513_);
  and g_15229_(_09265_, _09512_, _09514_);
  or g_15230_(_09264_, _09513_, _09515_);
  xor g_15231_(_09264_, _09513_, _09516_);
  xor g_15232_(_09264_, _09512_, _09517_);
  and g_15233_(_09261_, _09517_, _09518_);
  or g_15234_(_09260_, _09516_, _09519_);
  and g_15235_(_09509_, _09519_, _09520_);
  or g_15236_(_09508_, _09518_, _09521_);
  and g_15237_(_09339_, _09520_, _09523_);
  or g_15238_(_09338_, _09521_, _09524_);
  xor g_15239_(_09338_, _09520_, _09525_);
  not g_15240_(_09525_, _09526_);
  or g_15241_(_08983_, _09266_, _09527_);
  and g_15242_(_09272_, _09527_, _09528_);
  xor g_15243_(_09526_, _09528_, _09529_);
  not g_15244_(_09529_, _09530_);
  xor g_15245_(_09337_, _09530_, _09531_);
  or g_15246_(_09336_, _09531_, _09532_);
  xor g_15247_(_09336_, _09531_, _09534_);
  not g_15248_(_09534_, _09535_);
  or g_15249_(_09005_, _09285_, _09536_);
  and g_15250_(_09289_, _09536_, _09537_);
  xor g_15251_(_09534_, _09537_, _09538_);
  or g_15252_(_09332_, _09538_, _09539_);
  xor g_15253_(_09333_, _09538_, _09540_);
  or g_15254_(_09330_, _09540_, _09541_);
  xor g_15255_(_09330_, _09540_, _09542_);
  xor g_15256_(_09331_, _09540_, _09543_);
  and g_15257_(_09295_, _09297_, _09545_);
  xor g_15258_(_09542_, _09545_, _09546_);
  or g_15259_(_09299_, _09546_, _09547_);
  xor g_15260_(_09299_, _09546_, _09548_);
  not g_15261_(_09548_, _09549_);
  and g_15262_(_09306_, _09548_, _09550_);
  not g_15263_(_09550_, _09551_);
  or g_15264_(_09301_, _09549_, _09552_);
  xor g_15265_(_09301_, _09548_, _09553_);
  or g_15266_(_09310_, _09553_, _09554_);
  xor g_15267_(_09309_, _09553_, _09556_);
  and g_15268_(_09305_, _09556_, _09557_);
  or g_15269_(_09550_, _09557_, _09558_);
  or g_15270_(_09313_, _09558_, _09559_);
  xor g_15271_(_09313_, _09558_, _09560_);
  xor g_15272_(_09315_, _09558_, _09561_);
  or g_15273_(_09320_, _09324_, _09562_);
  or g_15274_(_09560_, _09562_, _09563_);
  and g_15275_(_09320_, _09560_, _09564_);
  or g_15276_(_09321_, _09561_, _09565_);
  or g_15277_(_09326_, _09561_, _09567_);
  and g_15278_(_09565_, _09567_, _09568_);
  and g_15279_(_09563_, _09568_, _09569_);
  and g_15280_(_09329_, _09569_, _09570_);
  xor g_15281_(_09329_, _09569_, out[324]);
  or g_15282_(_09295_, _09543_, _09571_);
  not g_15283_(_09571_, _09572_);
  and g_15284_(_09539_, _09541_, _09573_);
  not g_15285_(_09573_, _09574_);
  or g_15286_(_09289_, _09535_, _09575_);
  not g_15287_(_09575_, _09577_);
  or g_15288_(_09535_, _09536_, _09578_);
  or g_15289_(_09278_, _09529_, _09579_);
  or g_15290_(_09275_, _09529_, _09580_);
  not g_15291_(_09580_, _09581_);
  or g_15292_(_09272_, _09525_, _09582_);
  not g_15293_(_09582_, _09583_);
  or g_15294_(_09525_, _09527_, _09584_);
  and g_15295_(_09497_, _09502_, _09585_);
  and g_15296_(_09230_, _09474_, _09586_);
  or g_15297_(_09229_, _09475_, _09588_);
  and g_15298_(_09469_, _09472_, _09589_);
  or g_15299_(_09470_, _09471_, _09590_);
  or g_15300_(_09222_, _09470_, _09591_);
  and g_15301_(_09465_, _09591_, _09592_);
  and g_15302_(_09455_, _09459_, _09593_);
  and g_15303_(_09194_, _09451_, _09594_);
  and g_15304_(_09184_, _09446_, _09595_);
  or g_15305_(_09449_, _09595_, _09596_);
  and g_15306_(_09178_, _09438_, _09597_);
  or g_15307_(_09431_, _09433_, _09599_);
  or g_15308_(_09164_, _09430_, _09600_);
  or g_15309_(_09413_, _09415_, _09601_);
  or g_15310_(_09146_, _09411_, _09602_);
  or g_15311_(_07014_, _08205_, _09603_);
  or g_15312_(_08508_, _09603_, _09604_);
  or g_15313_(_08816_, _09604_, _09605_);
  or g_15314_(_09125_, _09605_, _09606_);
  and g_15315_(_09380_, _09606_, _09607_);
  or g_15316_(_09377_, _09607_, _09608_);
  and g_15317_(_09383_, _09608_, _09610_);
  and g_15318_(_09386_, _09610_, _09611_);
  and g_15319_(_09392_, _09611_, _09612_);
  and g_15320_(_09395_, _09612_, _09613_);
  and g_15321_(_09397_, _09613_, _09614_);
  and g_15322_(_09400_, _09614_, _09615_);
  and g_15323_(_09404_, _09615_, _09616_);
  and g_15324_(_09407_, _09616_, _09617_);
  and g_15325_(_09410_, _09617_, _09618_);
  and g_15326_(_09602_, _09618_, _09619_);
  and g_15327_(_09601_, _09619_, _09621_);
  and g_15328_(_09419_, _09621_, _09622_);
  and g_15329_(_09422_, _09622_, _09623_);
  and g_15330_(_09428_, _09623_, _09624_);
  and g_15331_(_09426_, _09624_, _09625_);
  and g_15332_(_09600_, _09625_, _09626_);
  and g_15333_(_09599_, _09626_, _09627_);
  and g_15334_(_09437_, _09627_, _09628_);
  or g_15335_(_09170_, _09439_, _09629_);
  and g_15336_(_09440_, _09629_, _09630_);
  xor g_15337_(_09628_, _09630_, _09632_);
  xor g_15338_(_09597_, _09632_, _09633_);
  xor g_15339_(_09447_, _09633_, _09634_);
  xor g_15340_(_09596_, _09634_, _09635_);
  xor g_15341_(_09594_, _09635_, _09636_);
  xor g_15342_(_09593_, _09636_, _09637_);
  not g_15343_(_09637_, _09638_);
  xor g_15344_(_09592_, _09638_, _09639_);
  xor g_15345_(_09592_, _09637_, _09640_);
  and g_15346_(_09589_, _09640_, _09641_);
  or g_15347_(_09590_, _09639_, _09643_);
  or g_15348_(_09589_, _09640_, _09644_);
  xor g_15349_(_09589_, _09639_, _09645_);
  and g_15350_(_09345_, _09474_, _09646_);
  or g_15351_(_09344_, _09475_, _09647_);
  and g_15352_(_09645_, _09647_, _09648_);
  and g_15353_(_09644_, _09646_, _09649_);
  and g_15354_(_09643_, _09649_, _09650_);
  or g_15355_(_09648_, _09650_, _09651_);
  or g_15356_(_09588_, _09651_, _09652_);
  xor g_15357_(_09586_, _09651_, _09654_);
  or g_15358_(_09484_, _09654_, _09655_);
  xor g_15359_(_09484_, _09654_, _09656_);
  xor g_15360_(_09485_, _09654_, _09657_);
  and g_15361_(_09482_, _09656_, _09658_);
  or g_15362_(_09483_, _09657_, _09659_);
  and g_15363_(_09483_, _09657_, _09660_);
  or g_15364_(_09482_, _09656_, _09661_);
  and g_15365_(_09659_, _09661_, _09662_);
  or g_15366_(_09658_, _09660_, _09663_);
  and g_15367_(_09491_, _09494_, _09665_);
  or g_15368_(_09492_, _09495_, _09666_);
  and g_15369_(_09663_, _09665_, _09667_);
  or g_15370_(_09662_, _09666_, _09668_);
  and g_15371_(_09661_, _09666_, _09669_);
  or g_15372_(_09660_, _09665_, _09670_);
  and g_15373_(_09659_, _09669_, _09671_);
  or g_15374_(_09658_, _09670_, _09672_);
  and g_15375_(_09668_, _09672_, _09673_);
  or g_15376_(_09667_, _09671_, _09674_);
  xor g_15377_(_09585_, _09673_, _09676_);
  and g_15378_(_09505_, _09510_, _09677_);
  or g_15379_(_09676_, _09677_, _09678_);
  xor g_15380_(_09676_, _09677_, _09679_);
  and g_15381_(_09508_, _09679_, _09680_);
  or g_15382_(_09508_, _09679_, _09681_);
  xor g_15383_(_09508_, _09679_, _09682_);
  not g_15384_(_09682_, _09683_);
  and g_15385_(_09523_, _09682_, _09684_);
  or g_15386_(_09524_, _09683_, _09685_);
  xor g_15387_(_09515_, _09682_, _09687_);
  and g_15388_(_09524_, _09687_, _09688_);
  or g_15389_(_09684_, _09688_, _09689_);
  xor g_15390_(_09584_, _09689_, _09690_);
  and g_15391_(_09583_, _09690_, _09691_);
  xor g_15392_(_09582_, _09690_, _09692_);
  or g_15393_(_09580_, _09692_, _09693_);
  xor g_15394_(_09581_, _09692_, _09694_);
  not g_15395_(_09694_, _09695_);
  or g_15396_(_09579_, _09694_, _09696_);
  xor g_15397_(_09579_, _09694_, _09698_);
  xor g_15398_(_09579_, _09695_, _09699_);
  or g_15399_(_09532_, _09699_, _09700_);
  xor g_15400_(_09532_, _09698_, _09701_);
  or g_15401_(_09578_, _09701_, _09702_);
  and g_15402_(_09578_, _09701_, _09703_);
  xor g_15403_(_09578_, _09701_, _09704_);
  xor g_15404_(_09577_, _09704_, _09705_);
  and g_15405_(_09574_, _09705_, _09706_);
  xor g_15406_(_09573_, _09705_, _09707_);
  or g_15407_(_09571_, _09707_, _09709_);
  and g_15408_(_09571_, _09707_, _09710_);
  xor g_15409_(_09572_, _09707_, _09711_);
  not g_15410_(_09711_, _09712_);
  or g_15411_(_09297_, _09543_, _09713_);
  and g_15412_(_09547_, _09713_, _09714_);
  xor g_15413_(_09711_, _09714_, _09715_);
  xor g_15414_(_09712_, _09714_, _09716_);
  or g_15415_(_09552_, _09716_, _09717_);
  and g_15416_(_09552_, _09716_, _09718_);
  xor g_15417_(_09552_, _09715_, _09720_);
  xor g_15418_(_09550_, _09720_, _09721_);
  or g_15419_(_09554_, _09721_, _09722_);
  and g_15420_(_09554_, _09721_, _09723_);
  xor g_15421_(_09554_, _09721_, _09724_);
  not g_15422_(_09724_, _09725_);
  and g_15423_(_09564_, _09724_, _09726_);
  or g_15424_(_09565_, _09725_, _09727_);
  xor g_15425_(_09559_, _09724_, _09728_);
  and g_15426_(_09565_, _09728_, _09729_);
  or g_15427_(_09726_, _09729_, _09731_);
  xor g_15428_(_09567_, _09731_, _09732_);
  and g_15429_(_09570_, _09732_, _09733_);
  xor g_15430_(_09570_, _09732_, out[325]);
  or g_15431_(_09567_, _09729_, _09734_);
  and g_15432_(_09727_, _09734_, _09735_);
  or g_15433_(_09551_, _09718_, _09736_);
  and g_15434_(_09717_, _09736_, _09737_);
  or g_15435_(_09710_, _09713_, _09738_);
  and g_15436_(_09709_, _09738_, _09739_);
  and g_15437_(_09693_, _09696_, _09741_);
  and g_15438_(_09584_, _09685_, _09742_);
  or g_15439_(_09688_, _09742_, _09743_);
  or g_15440_(_09514_, _09680_, _09744_);
  and g_15441_(_09681_, _09744_, _09745_);
  or g_15442_(_09498_, _09674_, _09746_);
  or g_15443_(_09252_, _09746_, _09747_);
  or g_15444_(_09250_, _09746_, _09748_);
  or g_15445_(_09497_, _09674_, _09749_);
  and g_15446_(_09652_, _09655_, _09750_);
  not g_15447_(_09750_, _09752_);
  and g_15448_(_09220_, _09463_, _09753_);
  or g_15449_(_05940_, _09466_, _09754_);
  or g_15450_(_09637_, _09754_, _09755_);
  or g_15451_(_09753_, _09755_, _09756_);
  or g_15452_(_09641_, _09649_, _09757_);
  not g_15453_(_09757_, _09758_);
  xor g_15454_(_09756_, _09758_, _09759_);
  xor g_15455_(_09756_, _09757_, _09760_);
  and g_15456_(_09752_, _09760_, _09761_);
  and g_15457_(_09750_, _09759_, _09763_);
  or g_15458_(_09658_, _09763_, _09764_);
  or g_15459_(_09761_, _09764_, _09765_);
  or g_15460_(_09669_, _09765_, _09766_);
  xor g_15461_(_09749_, _09766_, _09767_);
  and g_15462_(_09748_, _09767_, _09768_);
  xor g_15463_(_09747_, _09768_, _09769_);
  xor g_15464_(_09678_, _09769_, _09770_);
  xor g_15465_(_09745_, _09770_, _09771_);
  xor g_15466_(_09743_, _09771_, _09772_);
  xor g_15467_(_09691_, _09772_, _09774_);
  xor g_15468_(_09741_, _09774_, _09775_);
  xor g_15469_(_09700_, _09775_, _09776_);
  or g_15470_(_09575_, _09703_, _09777_);
  and g_15471_(_09702_, _09777_, _09778_);
  xor g_15472_(_09776_, _09778_, _09779_);
  xor g_15473_(_09739_, _09779_, _09780_);
  or g_15474_(_09547_, _09711_, _09781_);
  xor g_15475_(_09706_, _09781_, _09782_);
  xor g_15476_(_09780_, _09782_, _09783_);
  xor g_15477_(_09737_, _09783_, _09785_);
  and g_15478_(_09559_, _09722_, _09786_);
  or g_15479_(_09723_, _09786_, _09787_);
  xor g_15480_(_09785_, _09787_, _09788_);
  xor g_15481_(_09735_, _09788_, _09789_);
  xor g_15482_(_09733_, _09789_, out[326]);
  buf b_0_(set1[83], out[243]);
  buf b_1_(set1[98], out[258]);
  buf b_2_(set2[155], out[155]);
  buf b_3_(set1[124], out[284]);
  buf b_4_(set2[129], out[129]);
  buf b_5_(set2[54], out[54]);
  buf b_6_(set1[17], out[177]);
  buf b_7_(set2[141], out[141]);
  buf b_8_(set2[57], out[57]);
  buf b_9_(set2[28], out[28]);
  buf b_10_(set1[62], out[222]);
  buf b_11_(set2[97], out[97]);
  buf b_12_(set1[93], out[253]);
  buf b_13_(set1[0], out[160]);
  buf b_14_(set1[127], out[287]);
  buf b_15_(set2[31], out[31]);
  buf b_16_(set1[57], out[217]);
  buf b_17_(set1[48], out[208]);
  buf b_18_(set1[141], out[301]);
  buf b_19_(set1[66], out[226]);
  buf b_20_(set2[3], out[3]);
  buf b_21_(set1[43], out[203]);
  buf b_22_(set2[127], out[127]);
  buf b_23_(set2[46], out[46]);
  buf b_24_(set2[98], out[98]);
  buf b_25_(set1[130], out[290]);
  buf b_26_(set2[35], out[35]);
  buf b_27_(set2[89], out[89]);
  buf b_28_(set2[29], out[29]);
  buf b_29_(set1[51], out[211]);
  buf b_30_(set2[88], out[88]);
  buf b_31_(set1[69], out[229]);
  buf b_32_(set1[46], out[206]);
  buf b_33_(set1[41], out[201]);
  buf b_34_(set2[83], out[83]);
  buf b_35_(set2[53], out[53]);
  buf b_36_(set1[80], out[240]);
  buf b_37_(set1[145], out[305]);
  buf b_38_(set1[27], out[187]);
  buf b_39_(set1[5], out[165]);
  buf b_40_(set2[69], out[69]);
  buf b_41_(set2[133], out[133]);
  buf b_42_(set2[104], out[104]);
  buf b_43_(set2[123], out[123]);
  buf b_44_(set2[138], out[138]);
  buf b_45_(set2[148], out[148]);
  buf b_46_(set1[37], out[197]);
  buf b_47_(set2[87], out[87]);
  buf b_48_(set1[25], out[185]);
  buf b_49_(set1[20], out[180]);
  buf b_50_(set1[144], out[304]);
  buf b_51_(set2[78], out[78]);
  buf b_52_(set2[84], out[84]);
  buf b_53_(set1[103], out[263]);
  buf b_54_(set2[59], out[59]);
  buf b_55_(set2[153], out[153]);
  buf b_56_(set2[44], out[44]);
  buf b_57_(set1[49], out[209]);
  buf b_58_(set1[95], out[255]);
  buf b_59_(set1[10], out[170]);
  buf b_60_(set1[122], out[282]);
  buf b_61_(set2[18], out[18]);
  buf b_62_(set2[6], out[6]);
  buf b_63_(set1[131], out[291]);
  buf b_64_(set1[11], out[171]);
  buf b_65_(set1[28], out[188]);
  buf b_66_(set1[142], out[302]);
  buf b_67_(set2[149], out[149]);
  buf b_68_(set2[157], out[157]);
  buf b_69_(set1[32], out[192]);
  buf b_70_(set2[76], out[76]);
  buf b_71_(set1[107], out[267]);
  buf b_72_(set1[139], out[299]);
  buf b_73_(set1[143], out[303]);
  buf b_74_(set1[94], out[254]);
  czero b_75_(_10276_);
  buf b_76_(set1[75], out[235]);
  buf b_77_(set2[56], out[56]);
  buf b_78_(set2[85], out[85]);
  buf b_79_(set1[132], out[292]);
  buf b_80_(set2[64], out[64]);
  buf b_81_(set1[74], out[234]);
  buf b_82_(set1[13], out[173]);
  buf b_83_(set1[87], out[247]);
  buf b_84_(set2[119], out[119]);
  buf b_85_(set2[82], out[82]);
  buf b_86_(set1[159], out[319]);
  buf b_87_(set2[118], out[118]);
  buf b_88_(set2[109], out[109]);
  buf b_89_(set1[34], out[194]);
  buf b_90_(set2[121], out[121]);
  buf b_91_(set2[134], out[134]);
  buf b_92_(set1[78], out[238]);
  buf b_93_(set1[105], out[265]);
  buf b_94_(set2[126], out[126]);
  buf b_95_(set2[12], out[12]);
  buf b_96_(set1[86], out[246]);
  buf b_97_(set2[86], out[86]);
  buf b_98_(set1[2], out[162]);
  buf b_99_(set2[19], out[19]);
  buf b_100_(set2[1], out[1]);
  buf b_101_(set1[152], out[312]);
  buf b_102_(set1[134], out[294]);
  buf b_103_(set1[101], out[261]);
  buf b_104_(set2[140], out[140]);
  buf b_105_(set2[92], out[92]);
  buf b_106_(set1[26], out[186]);
  buf b_107_(set2[23], out[23]);
  buf b_108_(set1[155], out[315]);
  buf b_109_(set2[130], out[130]);
  buf b_110_(set2[101], out[101]);
  buf b_111_(set2[80], out[80]);
  buf b_112_(set2[9], out[9]);
  buf b_113_(set2[96], out[96]);
  buf b_114_(set1[110], out[270]);
  buf b_115_(set2[156], out[156]);
  buf b_116_(set2[0], out[0]);
  buf b_117_(set2[105], out[105]);
  buf b_118_(set1[53], out[213]);
  buf b_119_(set2[142], out[142]);
  buf b_120_(set1[50], out[210]);
  buf b_121_(set1[114], out[274]);
  buf b_122_(set1[55], out[215]);
  buf b_123_(set1[82], out[242]);
  buf b_124_(set2[95], out[95]);
  buf b_125_(set1[44], out[204]);
  buf b_126_(set1[111], out[271]);
  buf b_127_(set1[7], out[167]);
  buf b_128_(set1[85], out[245]);
  buf b_129_(set2[75], out[75]);
  buf b_130_(set2[91], out[91]);
  buf b_131_(set1[45], out[205]);
  buf b_132_(set1[18], out[178]);
  buf b_133_(set2[24], out[24]);
  buf b_134_(set2[34], out[34]);
  buf b_135_(set2[137], out[137]);
  buf b_136_(set2[70], out[70]);
  buf b_137_(set1[118], out[278]);
  buf b_138_(set2[51], out[51]);
  buf b_139_(set2[15], out[15]);
  buf b_140_(set1[138], out[298]);
  buf b_141_(set1[126], out[286]);
  buf b_142_(set2[90], out[90]);
  buf b_143_(set2[116], out[116]);
  buf b_144_(set2[39], out[39]);
  buf b_145_(set2[159], out[159]);
  buf b_146_(set1[19], out[179]);
  buf b_147_(set1[30], out[190]);
  buf b_148_(set2[72], out[72]);
  buf b_149_(set1[123], out[283]);
  buf b_150_(set1[135], out[295]);
  buf b_151_(set1[47], out[207]);
  buf b_152_(set2[131], out[131]);
  buf b_153_(set2[79], out[79]);
  buf b_154_(set2[68], out[68]);
  buf b_155_(set1[70], out[230]);
  buf b_156_(set2[66], out[66]);
  buf b_157_(set2[147], out[147]);
  buf b_158_(set2[37], out[37]);
  buf b_159_(set1[154], out[314]);
  buf b_160_(set1[102], out[262]);
  buf b_161_(set1[113], out[273]);
  buf b_162_(set2[40], out[40]);
  buf b_163_(set2[47], out[47]);
  buf b_164_(set2[36], out[36]);
  buf b_165_(set2[77], out[77]);
  buf b_166_(set2[65], out[65]);
  buf b_167_(set2[10], out[10]);
  buf b_168_(set1[42], out[202]);
  buf b_169_(set2[108], out[108]);
  buf b_170_(set1[153], out[313]);
  buf b_171_(set1[8], out[168]);
  buf b_172_(set1[73], out[233]);
  buf b_173_(set1[108], out[268]);
  buf b_174_(set1[151], out[311]);
  buf b_175_(set1[58], out[218]);
  buf b_176_(set1[64], out[224]);
  buf b_177_(set2[106], out[106]);
  buf b_178_(set1[40], out[200]);
  buf b_179_(set1[121], out[281]);
  buf b_180_(set1[52], out[212]);
  buf b_181_(set1[84], out[244]);
  buf b_182_(set2[120], out[120]);
  buf b_183_(set1[116], out[276]);
  czero b_184_(out[327]);
  buf b_185_(set1[136], out[296]);
  buf b_186_(set1[65], out[225]);
  buf b_187_(set2[52], out[52]);
  buf b_188_(set1[96], out[256]);
  buf b_189_(set1[23], out[183]);
  buf b_190_(set2[11], out[11]);
  buf b_191_(set2[128], out[128]);
  buf b_192_(set2[26], out[26]);
  buf b_193_(set2[21], out[21]);
  buf b_194_(set1[150], out[310]);
  buf b_195_(set1[60], out[220]);
  buf b_196_(set2[17], out[17]);
  buf b_197_(set1[140], out[300]);
  buf b_198_(set1[71], out[231]);
  buf b_199_(set2[48], out[48]);
  buf b_200_(set1[67], out[227]);
  buf b_201_(set1[3], out[163]);
  buf b_202_(set1[90], out[250]);
  buf b_203_(set2[13], out[13]);
  buf b_204_(set2[71], out[71]);
  buf b_205_(set1[115], out[275]);
  buf b_206_(set2[58], out[58]);
  buf b_207_(set2[152], out[152]);
  buf b_208_(set1[104], out[264]);
  buf b_209_(set2[102], out[102]);
  buf b_210_(set2[100], out[100]);
  buf b_211_(set2[154], out[154]);
  buf b_212_(set2[103], out[103]);
  buf b_213_(set1[12], out[172]);
  buf b_214_(set2[55], out[55]);
  buf b_215_(set2[93], out[93]);
  buf b_216_(set2[143], out[143]);
  buf b_217_(set2[94], out[94]);
  buf b_218_(set1[61], out[221]);
  buf b_219_(set2[30], out[30]);
  buf b_220_(set1[156], out[316]);
  buf b_221_(set1[133], out[293]);
  buf b_222_(set1[128], out[288]);
  buf b_223_(set1[72], out[232]);
  buf b_224_(set2[5], out[5]);
  czero b_225_(out[327]);
  buf b_226_(set1[16], out[176]);
  buf b_227_(set2[25], out[25]);
  buf b_228_(set2[22], out[22]);
  buf b_229_(set2[112], out[112]);
  buf b_230_(set1[6], out[166]);
  buf b_231_(set2[135], out[135]);
  buf b_232_(set2[114], out[114]);
  buf b_233_(set1[129], out[289]);
  buf b_234_(set1[14], out[174]);
  buf b_235_(set1[38], out[198]);
  buf b_236_(set2[145], out[145]);
  buf b_237_(set2[117], out[117]);
  buf b_238_(set1[120], out[280]);
  buf b_239_(set1[92], out[252]);
  buf b_240_(set2[33], out[33]);
  buf b_241_(set1[109], out[269]);
  buf b_242_(set2[144], out[144]);
  buf b_243_(set2[14], out[14]);
  buf b_244_(set1[149], out[309]);
  buf b_245_(set2[2], out[2]);
  buf b_246_(set2[16], out[16]);
  buf b_247_(set1[63], out[223]);
  buf b_248_(set2[63], out[63]);
  buf b_249_(set2[32], out[32]);
  buf b_250_(set2[139], out[139]);
  buf b_251_(set1[81], out[241]);
  buf b_252_(set1[146], out[306]);
  buf b_253_(set2[42], out[42]);
  buf b_254_(set1[21], out[181]);
  buf b_255_(set2[132], out[132]);
  buf b_256_(set2[27], out[27]);
  buf b_257_(set1[158], out[318]);
  buf b_258_(set1[77], out[237]);
  buf b_259_(set1[35], out[195]);
  buf b_260_(set2[67], out[67]);
  buf b_261_(set2[8], out[8]);
  buf b_262_(set1[39], out[199]);
  buf b_263_(set2[136], out[136]);
  buf b_264_(set1[157], out[317]);
  buf b_265_(set2[124], out[124]);
  buf b_266_(set2[99], out[99]);
  buf b_267_(set2[146], out[146]);
  buf b_268_(set1[91], out[251]);
  buf b_269_(set1[76], out[236]);
  buf b_270_(set1[117], out[277]);
  buf b_271_(set2[115], out[115]);
  buf b_272_(set1[97], out[257]);
  buf b_273_(set2[38], out[38]);
  buf b_274_(set1[36], out[196]);
  buf b_275_(set2[7], out[7]);
  buf b_276_(set1[137], out[297]);
  buf b_277_(set1[148], out[308]);
  buf b_278_(set2[74], out[74]);
  buf b_279_(set2[61], out[61]);
  buf b_280_(set2[158], out[158]);
  buf b_281_(set2[125], out[125]);
  buf b_282_(set1[22], out[182]);
  buf b_283_(set1[56], out[216]);
  buf b_284_(set1[88], out[248]);
  buf b_285_(set1[31], out[191]);
  buf b_286_(set1[15], out[175]);
  buf b_287_(set2[111], out[111]);
  buf b_288_(set2[73], out[73]);
  buf b_289_(set2[151], out[151]);
  buf b_290_(set2[107], out[107]);
  buf b_291_(set2[113], out[113]);
  buf b_292_(set2[60], out[60]);
  buf b_293_(set1[119], out[279]);
  buf b_294_(set2[81], out[81]);
  buf b_295_(set1[112], out[272]);
  buf b_296_(set1[59], out[219]);
  buf b_297_(set1[100], out[260]);
  buf b_298_(set2[110], out[110]);
  buf b_299_(set1[1], out[161]);
  buf b_300_(set2[4], out[4]);
  buf b_301_(set1[68], out[228]);
  buf b_302_(set1[99], out[259]);
  buf b_303_(set1[89], out[249]);
  buf b_304_(set1[9], out[169]);
  buf b_305_(set1[24], out[184]);
  buf b_306_(set2[20], out[20]);
  buf b_307_(set2[150], out[150]);
  buf b_308_(set2[49], out[49]);
  buf b_309_(set1[4], out[164]);
  buf b_310_(set2[41], out[41]);
  buf b_311_(set2[50], out[50]);
  buf b_312_(set1[54], out[214]);
  buf b_313_(set2[62], out[62]);
  buf b_314_(set1[29], out[189]);
  buf b_315_(set2[45], out[45]);
  buf b_316_(set1[33], out[193]);
  buf b_317_(set1[147], out[307]);
  buf b_318_(set1[106], out[266]);
  buf b_319_(set2[43], out[43]);
  buf b_320_(set1[125], out[285]);
  buf b_321_(set1[79], out[239]);
  buf b_322_(set2[122], out[122]);

endmodule
