module min_hash(
  input wire [159:0] set1,
  input wire [159:0] set2,
  output wire [335:0] out
);
  wire [15:0] set1_unflattened[10];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  wire [15:0] set2_unflattened[10];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  wire [15:0] array_index_21426;
  wire [11:0] add_21430;
  wire [12:0] concat_21434;
  wire [10:0] add_21437;
  wire eq_21440;
  wire [12:0] concat_21443;
  wire [15:0] array_index_21445;
  wire ne_21457;
  wire [11:0] sel_21458;
  wire [8:0] add_21461;
  wire [11:0] concat_21464;
  wire [11:0] add_21469;
  wire [11:0] sel_21471;
  wire [12:0] concat_21472;
  wire [11:0] sel_21476;
  wire [12:0] concat_21479;
  wire [12:0] concat_21480;
  wire [10:0] add_21485;
  wire [11:0] sel_21488;
  wire eq_21490;
  wire [10:0] add_21493;
  wire [11:0] concat_21495;
  wire [12:0] concat_21499;
  wire [12:0] concat_21500;
  wire [15:0] array_index_21501;
  wire [12:0] concat_21504;
  wire [11:0] sel_21508;
  wire nor_21513;
  wire [11:0] sel_21514;
  wire [11:0] sel_21515;
  wire [8:0] add_21520;
  wire [11:0] sel_21523;
  wire [11:0] concat_21525;
  wire [11:0] add_21528;
  wire [11:0] sel_21530;
  wire [10:0] add_21532;
  wire [11:0] concat_21534;
  wire [12:0] concat_21538;
  wire [12:0] concat_21539;
  wire [11:0] sel_21542;
  wire [11:0] sel_21543;
  wire [12:0] concat_21545;
  wire [12:0] concat_21546;
  wire [12:0] concat_21547;
  wire [11:0] sel_21550;
  wire [10:0] add_21554;
  wire [11:0] sel_21557;
  wire eq_21559;
  wire [10:0] add_21564;
  wire [11:0] sel_21566;
  wire [11:0] concat_21568;
  wire [12:0] concat_21570;
  wire [12:0] concat_21571;
  wire [15:0] array_index_21572;
  wire [11:0] concat_21576;
  wire [12:0] concat_21580;
  wire [12:0] concat_21581;
  wire [11:0] sel_21584;
  wire [11:0] sel_21585;
  wire or_21589;
  wire [11:0] sel_21590;
  wire [11:0] sel_21594;
  wire [8:0] add_21598;
  wire [11:0] sel_21601;
  wire [11:0] concat_21603;
  wire [11:0] add_21607;
  wire [11:0] sel_21609;
  wire [15:0] array_index_21610;
  wire [10:0] add_21612;
  wire [11:0] sel_21614;
  wire [11:0] concat_21616;
  wire [12:0] concat_21618;
  wire [12:0] concat_21619;
  wire [11:0] sel_21622;
  wire eq_21624;
  wire [12:0] concat_21625;
  wire [12:0] concat_21626;
  wire [12:0] concat_21629;
  wire [12:0] concat_21630;
  wire [11:0] sel_21632;
  wire [11:0] sel_21633;
  wire [10:0] add_21636;
  wire [11:0] sel_21639;
  wire or_21642;
  wire [11:0] add_21646;
  wire [10:0] add_21649;
  wire [11:0] sel_21651;
  wire [11:0] concat_21653;
  wire [12:0] concat_21655;
  wire [12:0] concat_21656;
  wire [15:0] array_index_21659;
  wire [15:0] array_index_21664;
  wire [11:0] concat_21668;
  wire [12:0] concat_21670;
  wire [12:0] concat_21671;
  wire [11:0] sel_21674;
  wire [10:0] add_21678;
  wire nor_21680;
  wire and_21683;
  wire [11:0] sel_21691;
  wire [11:0] sel_21692;
  wire [8:0] add_21695;
  wire [11:0] sel_21698;
  wire [11:0] concat_21700;
  wire [11:0] add_21707;
  wire [11:0] sel_21709;
  wire [11:0] add_21712;
  wire [11:0] sel_21714;
  wire [10:0] add_21716;
  wire [11:0] sel_21718;
  wire [11:0] concat_21720;
  wire [12:0] concat_21722;
  wire [12:0] concat_21723;
  wire or_21735;
  wire eq_21736;
  wire [12:0] concat_21737;
  wire [12:0] concat_21738;
  wire [15:0] array_index_21739;
  wire [12:0] concat_21742;
  wire [12:0] concat_21743;
  wire [11:0] sel_21745;
  wire [8:0] add_21749;
  wire [10:0] add_21752;
  wire [11:0] sel_21755;
  wire [10:0] add_21757;
  wire [11:0] sel_21760;
  wire or_21763;
  wire [10:0] add_21770;
  wire [11:0] sel_21772;
  wire [11:0] concat_21774;
  wire [12:0] concat_21778;
  wire [12:0] concat_21779;
  wire [15:0] array_index_21782;
  wire [11:0] add_21789;
  wire [11:0] sel_21791;
  wire [11:0] concat_21793;
  wire [12:0] concat_21795;
  wire [12:0] concat_21796;
  wire and_21812;
  wire and_21815;
  wire [15:0] array_index_21818;
  wire [11:0] sel_21822;
  wire [10:0] add_21826;
  wire [8:0] add_21828;
  wire [11:0] sel_21831;
  wire [8:0] add_21833;
  wire [11:0] sel_21836;
  wire [11:0] concat_21838;
  wire [10:0] add_21841;
  wire [11:0] sel_21844;
  wire [11:0] add_21848;
  wire [11:0] sel_21850;
  wire [10:0] add_21855;
  wire [11:0] sel_21857;
  wire [11:0] concat_21859;
  wire [12:0] concat_21863;
  wire [12:0] concat_21864;
  wire or_21873;
  wire eq_21874;
  wire [12:0] concat_21875;
  wire [12:0] concat_21876;
  wire [11:0] add_21879;
  wire [11:0] sel_21881;
  wire [12:0] concat_21882;
  wire [12:0] concat_21883;
  wire [10:0] add_21898;
  wire [11:0] sel_21901;
  wire or_21908;
  wire [15:0] array_index_21910;
  wire [10:0] add_21915;
  wire [10:0] add_21917;
  wire [11:0] sel_21919;
  wire [10:0] add_21921;
  wire [11:0] sel_21923;
  wire [11:0] concat_21925;
  wire [8:0] add_21928;
  wire [11:0] sel_21931;
  wire [12:0] concat_21932;
  wire [12:0] concat_21933;
  wire [10:0] add_21935;
  wire [11:0] sel_21938;
  wire [15:0] array_index_21939;
  wire [11:0] concat_21948;
  wire [12:0] concat_21952;
  wire [12:0] concat_21953;
  wire and_21967;
  wire [11:0] add_21972;
  wire [11:0] sel_21974;
  wire [8:0] add_21987;
  wire [11:0] sel_21990;
  wire [11:0] concat_21996;
  wire [11:0] add_22003;
  wire [11:0] sel_22005;
  wire [15:0] array_index_22006;
  wire [10:0] add_22010;
  wire [11:0] sel_22012;
  wire [10:0] add_22014;
  wire [11:0] sel_22016;
  wire [11:0] concat_22018;
  wire [10:0] add_22021;
  wire [11:0] sel_22023;
  wire [12:0] concat_22024;
  wire [12:0] concat_22025;
  wire [8:0] add_22027;
  wire [11:0] sel_22030;
  wire [10:0] add_22036;
  wire [11:0] sel_22039;
  wire and_22040;
  wire [12:0] concat_22042;
  wire [12:0] concat_22043;
  wire [12:0] concat_22047;
  wire [12:0] concat_22048;
  wire [10:0] add_22060;
  wire [11:0] sel_22063;
  wire eq_22068;
  wire [11:0] add_22072;
  wire [11:0] sel_22074;
  wire [10:0] add_22080;
  wire [11:0] sel_22082;
  wire [11:0] concat_22087;
  wire [12:0] concat_22093;
  wire [12:0] concat_22094;
  wire [15:0] array_index_22099;
  wire or_22100;
  wire [15:0] array_index_22103;
  wire [11:0] concat_22107;
  wire [10:0] add_22110;
  wire [11:0] sel_22112;
  wire [12:0] concat_22113;
  wire [12:0] concat_22114;
  wire [10:0] add_22116;
  wire [11:0] sel_22118;
  wire [8:0] add_22124;
  wire [11:0] sel_22127;
  wire [10:0] add_22130;
  wire [11:0] sel_22133;
  wire or_22136;
  wire [11:0] sel_22137;
  wire [8:0] add_22151;
  wire [11:0] sel_22154;
  wire [11:0] concat_22158;
  wire [11:0] add_22164;
  wire [11:0] add_22169;
  wire [11:0] sel_22171;
  wire [10:0] add_22173;
  wire [11:0] sel_22175;
  wire [11:0] concat_22180;
  wire [12:0] concat_22185;
  wire [12:0] concat_22186;
  wire [11:0] sel_22193;
  wire [15:0] array_index_22199;
  wire [15:0] array_index_22202;
  wire [12:0] concat_22205;
  wire [12:0] concat_22206;
  wire [10:0] add_22208;
  wire [11:0] sel_22210;
  wire [10:0] add_22215;
  wire [11:0] sel_22217;
  wire [8:0] add_22220;
  wire [11:0] sel_22223;
  wire [10:0] add_22225;
  wire [10:0] add_22230;
  wire [11:0] sel_22233;
  wire [10:0] add_22244;
  wire [11:0] sel_22246;
  wire [11:0] concat_22250;
  wire [11:0] add_22260;
  wire [11:0] sel_22262;
  wire [11:0] add_22265;
  wire [11:0] sel_22267;
  wire [11:0] concat_22269;
  wire [12:0] concat_22274;
  wire [12:0] concat_22275;
  wire [11:0] sel_22281;
  wire and_22295;
  wire [15:0] array_index_22297;
  wire [15:0] array_index_22300;
  wire [10:0] add_22307;
  wire [11:0] sel_22309;
  wire [10:0] add_22312;
  wire [11:0] sel_22314;
  wire [8:0] add_22316;
  wire [8:0] add_22321;
  wire [11:0] sel_22324;
  wire [10:0] add_22326;
  wire [11:0] sel_22329;
  wire [10:0] add_22331;
  wire [11:0] sel_22334;
  wire [10:0] add_22345;
  wire [11:0] sel_22347;
  wire [11:0] concat_22351;
  wire or_22364;
  wire [11:0] add_22369;
  wire [11:0] sel_22371;
  wire [11:0] add_22374;
  wire [11:0] sel_22376;
  wire [12:0] concat_22377;
  wire [12:0] concat_22378;
  wire [11:0] sel_22383;
  wire or_22405;
  wire and_22406;
  wire [12:0] concat_22410;
  wire [12:0] concat_22411;
  wire [15:0] array_index_22412;
  wire [10:0] add_22417;
  wire [11:0] sel_22419;
  wire [10:0] add_22421;
  wire [10:0] add_22425;
  wire [11:0] sel_22427;
  wire [8:0] add_22429;
  wire [11:0] sel_22432;
  wire [8:0] add_22434;
  wire [11:0] sel_22437;
  wire [10:0] add_22440;
  wire [11:0] sel_22443;
  wire [10:0] add_22445;
  wire [11:0] sel_22448;
  wire eq_22452;
  wire [11:0] concat_22458;
  wire [12:0] concat_22472;
  wire [12:0] concat_22473;
  wire [11:0] add_22483;
  wire [11:0] sel_22485;
  wire [11:0] sel_22487;
  wire and_22513;
  wire ne_22516;
  wire [10:0] add_22522;
  wire [10:0] add_22526;
  wire [11:0] sel_22528;
  wire [10:0] add_22530;
  wire [11:0] sel_22532;
  wire [10:0] add_22534;
  wire [11:0] sel_22536;
  wire [8:0] add_22539;
  wire [11:0] sel_22542;
  wire [8:0] add_22544;
  wire [11:0] sel_22547;
  wire [11:0] concat_22550;
  wire [10:0] add_22553;
  wire [11:0] sel_22556;
  wire and_22557;
  wire [12:0] concat_22571;
  wire [12:0] concat_22572;
  wire [10:0] add_22608;
  wire [11:0] sel_22610;
  wire [10:0] add_22612;
  wire [11:0] sel_22614;
  wire [10:0] add_22617;
  wire [11:0] sel_22619;
  wire [10:0] add_22621;
  wire [11:0] sel_22623;
  wire [11:0] concat_22626;
  wire [8:0] add_22629;
  wire [11:0] sel_22632;
  wire [1:0] concat_22635;
  wire [12:0] concat_22643;
  wire [12:0] concat_22644;
  wire [1:0] add_22653;
  wire [10:0] add_22674;
  wire [11:0] sel_22676;
  wire [10:0] add_22678;
  wire [11:0] sel_22680;
  wire [11:0] concat_22683;
  wire [10:0] add_22686;
  wire [11:0] sel_22688;
  wire [2:0] concat_22691;
  wire [12:0] concat_22694;
  wire [12:0] concat_22695;
  wire [2:0] add_22704;
  wire [11:0] concat_22718;
  wire [10:0] add_22721;
  wire [11:0] sel_22723;
  wire [3:0] concat_22726;
  wire [3:0] add_22734;
  wire [4:0] concat_22743;
  wire [4:0] add_22746;
  assign array_index_21426 = set1_unflattened[4'h0];
  assign add_21430 = array_index_21426[11:0] + 12'h247;
  assign concat_21434 = {1'h0, add_21430};
  assign add_21437 = array_index_21426[11:1] + 11'h247;
  assign eq_21440 = array_index_21426 == 16'h0000;
  assign concat_21443 = {1'h0, add_21437, array_index_21426[0]};
  assign array_index_21445 = set1_unflattened[4'h1];
  assign ne_21457 = array_index_21426 != 16'h0000;
  assign sel_21458 = eq_21440 | $signed(concat_21434) >= $signed(13'h0fff) ? 12'hfff : add_21430;
  assign add_21461 = array_index_21426[11:3] + 9'h0bd;
  assign concat_21464 = {add_21437, array_index_21426[0]};
  assign add_21469 = array_index_21445[11:0] + 12'h247;
  assign sel_21471 = ne_21457 ? ($signed(concat_21434) < $signed(13'h0fff) ? add_21430 : 12'hfff) : sel_21458;
  assign concat_21472 = {1'h0, add_21461, array_index_21426[2:0]};
  assign sel_21476 = eq_21440 | $signed(concat_21443) >= $signed(13'h0fff) ? 12'hfff : concat_21464;
  assign concat_21479 = {1'h0, add_21469};
  assign concat_21480 = {1'h0, sel_21471};
  assign add_21485 = array_index_21445[11:1] + 11'h247;
  assign sel_21488 = ne_21457 ? ($signed(concat_21443) < $signed(13'h0fff) ? concat_21464 : 12'hfff) : sel_21476;
  assign eq_21490 = array_index_21445 == 16'h0000;
  assign add_21493 = array_index_21426[11:1] + 11'h347;
  assign concat_21495 = {add_21461, array_index_21426[2:0]};
  assign concat_21499 = {1'h0, add_21485, array_index_21445[0]};
  assign concat_21500 = {1'h0, sel_21488};
  assign array_index_21501 = set1_unflattened[4'h2];
  assign concat_21504 = {1'h0, add_21493, array_index_21426[0]};
  assign sel_21508 = eq_21440 | $signed(concat_21472) >= $signed(13'h0fff) ? 12'hfff : concat_21495;
  assign nor_21513 = ~(eq_21490 | eq_21440);
  assign sel_21514 = eq_21490 | $signed(concat_21479) >= $signed(concat_21480) ? sel_21471 : add_21469;
  assign sel_21515 = $signed(concat_21479) < $signed(concat_21480) ? add_21469 : sel_21471;
  assign add_21520 = array_index_21445[11:3] + 9'h0bd;
  assign sel_21523 = ne_21457 ? ($signed(concat_21472) < $signed(13'h0fff) ? concat_21495 : 12'hfff) : sel_21508;
  assign concat_21525 = {add_21485, array_index_21445[0]};
  assign add_21528 = array_index_21501[11:0] + 12'h247;
  assign sel_21530 = nor_21513 ? sel_21515 : sel_21514;
  assign add_21532 = array_index_21426[11:1] + 11'h79d;
  assign concat_21534 = {add_21493, array_index_21426[0]};
  assign concat_21538 = {1'h0, add_21520, array_index_21445[2:0]};
  assign concat_21539 = {1'h0, sel_21523};
  assign sel_21542 = eq_21490 | $signed(concat_21499) >= $signed(concat_21500) ? sel_21488 : concat_21525;
  assign sel_21543 = $signed(concat_21499) < $signed(concat_21500) ? concat_21525 : sel_21488;
  assign concat_21545 = {1'h0, add_21528};
  assign concat_21546 = {1'h0, sel_21530};
  assign concat_21547 = {1'h0, add_21532, array_index_21426[0]};
  assign sel_21550 = eq_21440 | $signed(concat_21504) >= $signed(13'h0fff) ? 12'hfff : concat_21534;
  assign add_21554 = array_index_21501[11:1] + 11'h247;
  assign sel_21557 = nor_21513 ? sel_21543 : sel_21542;
  assign eq_21559 = array_index_21501 == 16'h0000;
  assign add_21564 = array_index_21445[11:1] + 11'h347;
  assign sel_21566 = ne_21457 ? ($signed(concat_21504) < $signed(13'h0fff) ? concat_21534 : 12'hfff) : sel_21550;
  assign concat_21568 = {add_21520, array_index_21445[2:0]};
  assign concat_21570 = {1'h0, add_21554, array_index_21501[0]};
  assign concat_21571 = {1'h0, sel_21557};
  assign array_index_21572 = set1_unflattened[4'h3];
  assign concat_21576 = {add_21532, array_index_21426[0]};
  assign concat_21580 = {1'h0, add_21564, array_index_21445[0]};
  assign concat_21581 = {1'h0, sel_21566};
  assign sel_21584 = eq_21490 | $signed(concat_21538) >= $signed(concat_21539) ? sel_21523 : concat_21568;
  assign sel_21585 = $signed(concat_21538) < $signed(concat_21539) ? concat_21568 : sel_21523;
  assign or_21589 = eq_21440 | eq_21490 | eq_21559;
  assign sel_21590 = $signed(concat_21545) < $signed(concat_21546) ? add_21528 : sel_21530;
  assign sel_21594 = eq_21440 | $signed(concat_21547) >= $signed(13'h0fff) ? 12'hfff : concat_21576;
  assign add_21598 = array_index_21501[11:3] + 9'h0bd;
  assign sel_21601 = nor_21513 ? sel_21585 : sel_21584;
  assign concat_21603 = {add_21554, array_index_21501[0]};
  assign add_21607 = array_index_21572[11:0] + 12'h247;
  assign sel_21609 = or_21589 ? (eq_21559 | $signed(concat_21545) >= $signed(concat_21546) ? sel_21530 : add_21528) : sel_21590;
  assign array_index_21610 = set2_unflattened[4'h0];
  assign add_21612 = array_index_21445[11:1] + 11'h79d;
  assign sel_21614 = ne_21457 ? ($signed(concat_21547) < $signed(13'h0fff) ? concat_21576 : 12'hfff) : sel_21594;
  assign concat_21616 = {add_21564, array_index_21445[0]};
  assign concat_21618 = {1'h0, add_21598, array_index_21501[2:0]};
  assign concat_21619 = {1'h0, sel_21601};
  assign sel_21622 = $signed(concat_21570) < $signed(concat_21571) ? concat_21603 : sel_21557;
  assign eq_21624 = array_index_21572 == 16'h0000;
  assign concat_21625 = {1'h0, add_21607};
  assign concat_21626 = {1'h0, sel_21609};
  assign concat_21629 = {1'h0, add_21612, array_index_21445[0]};
  assign concat_21630 = {1'h0, sel_21614};
  assign sel_21632 = eq_21490 | $signed(concat_21580) >= $signed(concat_21581) ? sel_21566 : concat_21616;
  assign sel_21633 = $signed(concat_21580) < $signed(concat_21581) ? concat_21616 : sel_21566;
  assign add_21636 = array_index_21572[11:1] + 11'h247;
  assign sel_21639 = or_21589 ? (eq_21559 | $signed(concat_21570) >= $signed(concat_21571) ? sel_21557 : concat_21603) : sel_21622;
  assign or_21642 = or_21589 | eq_21624;
  assign add_21646 = array_index_21610[11:0] + 12'h247;
  assign add_21649 = array_index_21501[11:1] + 11'h347;
  assign sel_21651 = nor_21513 ? sel_21633 : sel_21632;
  assign concat_21653 = {add_21598, array_index_21501[2:0]};
  assign concat_21655 = {1'h0, add_21636, array_index_21572[0]};
  assign concat_21656 = {1'h0, sel_21639};
  assign array_index_21659 = set1_unflattened[4'h4];
  assign array_index_21664 = set2_unflattened[4'h1];
  assign concat_21668 = {add_21612, array_index_21445[0]};
  assign concat_21670 = {1'h0, add_21649, array_index_21501[0]};
  assign concat_21671 = {1'h0, sel_21651};
  assign sel_21674 = $signed(concat_21618) < $signed(concat_21619) ? concat_21653 : sel_21601;
  assign add_21678 = array_index_21610[11:1] + 11'h247;
  assign nor_21680 = ~(eq_21440 | eq_21490 | eq_21559);
  assign and_21683 = array_index_21572 != 16'h0000 & ~or_21642;
  assign sel_21691 = eq_21490 | $signed(concat_21629) >= $signed(concat_21630) ? sel_21614 : concat_21668;
  assign sel_21692 = $signed(concat_21629) < $signed(concat_21630) ? concat_21668 : sel_21614;
  assign add_21695 = array_index_21572[11:3] + 9'h0bd;
  assign sel_21698 = or_21589 ? (eq_21559 | $signed(concat_21618) >= $signed(concat_21619) ? sel_21601 : concat_21653) : sel_21674;
  assign concat_21700 = {add_21636, array_index_21572[0]};
  assign add_21707 = array_index_21659[11:0] + 12'h247;
  assign sel_21709 = and_21683 ? ($signed(concat_21625) < $signed(concat_21626) ? add_21607 : sel_21590) : (eq_21624 | $signed(concat_21625) >= $signed(concat_21626) ? sel_21609 : add_21607);
  assign add_21712 = array_index_21664[11:0] + 12'h247;
  assign sel_21714 = $signed({1'h0, add_21646}) < $signed(13'h0fff) ? add_21646 : 12'hfff;
  assign add_21716 = array_index_21501[11:1] + 11'h79d;
  assign sel_21718 = nor_21513 ? sel_21692 : sel_21691;
  assign concat_21720 = {add_21649, array_index_21501[0]};
  assign concat_21722 = {1'h0, add_21695, array_index_21572[2:0]};
  assign concat_21723 = {1'h0, sel_21698};
  assign or_21735 = or_21589 | or_21642 & nor_21680;
  assign eq_21736 = array_index_21659 == 16'h0000;
  assign concat_21737 = {1'h0, add_21707};
  assign concat_21738 = {1'h0, sel_21709};
  assign array_index_21739 = set2_unflattened[4'h2];
  assign concat_21742 = {1'h0, add_21716, array_index_21501[0]};
  assign concat_21743 = {1'h0, sel_21718};
  assign sel_21745 = $signed(concat_21670) < $signed(concat_21671) ? concat_21720 : sel_21651;
  assign add_21749 = array_index_21610[11:3] + 9'h0bd;
  assign add_21752 = array_index_21659[11:1] + 11'h247;
  assign sel_21755 = and_21683 ? ($signed(concat_21655) < $signed(concat_21656) ? concat_21700 : sel_21622) : (eq_21624 | $signed(concat_21655) >= $signed(concat_21656) ? sel_21639 : concat_21700);
  assign add_21757 = array_index_21664[11:1] + 11'h247;
  assign sel_21760 = $signed({1'h0, add_21678, array_index_21610[0]}) < $signed(13'h0fff) ? {add_21678, array_index_21610[0]} : 12'hfff;
  assign or_21763 = or_21735 | eq_21736;
  assign add_21770 = array_index_21572[11:1] + 11'h347;
  assign sel_21772 = or_21589 ? (eq_21559 | $signed(concat_21670) >= $signed(concat_21671) ? sel_21651 : concat_21720) : sel_21745;
  assign concat_21774 = {add_21695, array_index_21572[2:0]};
  assign concat_21778 = {1'h0, add_21752, array_index_21659[0]};
  assign concat_21779 = {1'h0, sel_21755};
  assign array_index_21782 = set1_unflattened[4'h5];
  assign add_21789 = array_index_21739[11:0] + 12'h247;
  assign sel_21791 = $signed({1'h0, add_21712}) < $signed({1'h0, sel_21714}) ? add_21712 : sel_21714;
  assign concat_21793 = {add_21716, array_index_21501[0]};
  assign concat_21795 = {1'h0, add_21770, array_index_21572[0]};
  assign concat_21796 = {1'h0, sel_21772};
  assign and_21812 = nor_21680 & ~or_21642;
  assign and_21815 = array_index_21659 != 16'h0000 & ~or_21763;
  assign array_index_21818 = set2_unflattened[4'h3];
  assign sel_21822 = $signed(concat_21742) < $signed(concat_21743) ? concat_21793 : sel_21718;
  assign add_21826 = array_index_21610[11:1] + 11'h347;
  assign add_21828 = array_index_21659[11:3] + 9'h0bd;
  assign sel_21831 = and_21683 ? ($signed(concat_21722) < $signed(concat_21723) ? concat_21774 : sel_21674) : (eq_21624 | $signed(concat_21722) >= $signed(concat_21723) ? sel_21698 : concat_21774);
  assign add_21833 = array_index_21664[11:3] + 9'h0bd;
  assign sel_21836 = $signed({1'h0, add_21749, array_index_21610[2:0]}) < $signed(13'h0fff) ? {add_21749, array_index_21610[2:0]} : 12'hfff;
  assign concat_21838 = {add_21752, array_index_21659[0]};
  assign add_21841 = array_index_21739[11:1] + 11'h247;
  assign sel_21844 = $signed({1'h0, add_21757, array_index_21664[0]}) < $signed({1'h0, sel_21760}) ? {add_21757, array_index_21664[0]} : sel_21760;
  assign add_21848 = array_index_21782[11:0] + 12'h247;
  assign sel_21850 = and_21815 ? ($signed(concat_21737) < $signed(concat_21738) ? add_21707 : sel_21709) : (eq_21736 | $signed(concat_21737) >= $signed(concat_21738) ? sel_21709 : add_21707);
  assign add_21855 = array_index_21572[11:1] + 11'h79d;
  assign sel_21857 = or_21589 ? (eq_21559 | $signed(concat_21742) >= $signed(concat_21743) ? sel_21718 : concat_21793) : sel_21822;
  assign concat_21859 = {add_21770, array_index_21572[0]};
  assign concat_21863 = {1'h0, add_21828, array_index_21659[2:0]};
  assign concat_21864 = {1'h0, sel_21831};
  assign or_21873 = or_21735 | or_21763 & and_21812;
  assign eq_21874 = array_index_21782 == 16'h0000;
  assign concat_21875 = {1'h0, add_21848};
  assign concat_21876 = {1'h0, sel_21850};
  assign add_21879 = array_index_21818[11:0] + 12'h247;
  assign sel_21881 = $signed({1'h0, add_21789}) < $signed({1'h0, sel_21791}) ? add_21789 : sel_21791;
  assign concat_21882 = {1'h0, add_21855, array_index_21572[0]};
  assign concat_21883 = {1'h0, sel_21857};
  assign add_21898 = array_index_21782[11:1] + 11'h247;
  assign sel_21901 = and_21815 ? ($signed(concat_21778) < $signed(concat_21779) ? concat_21838 : sel_21755) : (eq_21736 | $signed(concat_21778) >= $signed(concat_21779) ? sel_21755 : concat_21838);
  assign or_21908 = or_21873 | eq_21874;
  assign array_index_21910 = set2_unflattened[4'h4];
  assign add_21915 = array_index_21610[11:1] + 11'h79d;
  assign add_21917 = array_index_21659[11:1] + 11'h347;
  assign sel_21919 = and_21683 ? ($signed(concat_21795) < $signed(concat_21796) ? concat_21859 : sel_21745) : (eq_21624 | $signed(concat_21795) >= $signed(concat_21796) ? sel_21772 : concat_21859);
  assign add_21921 = array_index_21664[11:1] + 11'h347;
  assign sel_21923 = $signed({1'h0, add_21826, array_index_21610[0]}) < $signed(13'h0fff) ? {add_21826, array_index_21610[0]} : 12'hfff;
  assign concat_21925 = {add_21828, array_index_21659[2:0]};
  assign add_21928 = array_index_21739[11:3] + 9'h0bd;
  assign sel_21931 = $signed({1'h0, add_21833, array_index_21664[2:0]}) < $signed({1'h0, sel_21836}) ? {add_21833, array_index_21664[2:0]} : sel_21836;
  assign concat_21932 = {1'h0, add_21898, array_index_21782[0]};
  assign concat_21933 = {1'h0, sel_21901};
  assign add_21935 = array_index_21818[11:1] + 11'h247;
  assign sel_21938 = $signed({1'h0, add_21841, array_index_21739[0]}) < $signed({1'h0, sel_21844}) ? {add_21841, array_index_21739[0]} : sel_21844;
  assign array_index_21939 = set1_unflattened[4'h6];
  assign concat_21948 = {add_21855, array_index_21572[0]};
  assign concat_21952 = {1'h0, add_21917, array_index_21659[0]};
  assign concat_21953 = {1'h0, sel_21919};
  assign and_21967 = array_index_21782 != 16'h0000 & ~or_21908;
  assign add_21972 = array_index_21910[11:0] + 12'h247;
  assign sel_21974 = $signed({1'h0, add_21879}) < $signed({1'h0, sel_21881}) ? add_21879 : sel_21881;
  assign add_21987 = array_index_21782[11:3] + 9'h0bd;
  assign sel_21990 = and_21815 ? ($signed(concat_21863) < $signed(concat_21864) ? concat_21925 : sel_21831) : (eq_21736 | $signed(concat_21863) >= $signed(concat_21864) ? sel_21831 : concat_21925);
  assign concat_21996 = {add_21898, array_index_21782[0]};
  assign add_22003 = array_index_21939[11:0] + 12'h247;
  assign sel_22005 = and_21967 ? ($signed(concat_21875) < $signed(concat_21876) ? add_21848 : sel_21850) : (eq_21874 | $signed(concat_21875) >= $signed(concat_21876) ? sel_21850 : add_21848);
  assign array_index_22006 = set2_unflattened[4'h5];
  assign add_22010 = array_index_21659[11:1] + 11'h79d;
  assign sel_22012 = and_21683 ? ($signed(concat_21882) < $signed(concat_21883) ? concat_21948 : sel_21822) : (eq_21624 | $signed(concat_21882) >= $signed(concat_21883) ? sel_21857 : concat_21948);
  assign add_22014 = array_index_21664[11:1] + 11'h79d;
  assign sel_22016 = $signed({1'h0, add_21915, array_index_21610[0]}) < $signed(13'h0fff) ? {add_21915, array_index_21610[0]} : 12'hfff;
  assign concat_22018 = {add_21917, array_index_21659[0]};
  assign add_22021 = array_index_21739[11:1] + 11'h347;
  assign sel_22023 = $signed({1'h0, add_21921, array_index_21664[0]}) < $signed({1'h0, sel_21923}) ? {add_21921, array_index_21664[0]} : sel_21923;
  assign concat_22024 = {1'h0, add_21987, array_index_21782[2:0]};
  assign concat_22025 = {1'h0, sel_21990};
  assign add_22027 = array_index_21818[11:3] + 9'h0bd;
  assign sel_22030 = $signed({1'h0, add_21928, array_index_21739[2:0]}) < $signed({1'h0, sel_21931}) ? {add_21928, array_index_21739[2:0]} : sel_21931;
  assign add_22036 = array_index_21910[11:1] + 11'h247;
  assign sel_22039 = $signed({1'h0, add_21935, array_index_21818[0]}) < $signed({1'h0, sel_21938}) ? {add_21935, array_index_21818[0]} : sel_21938;
  assign and_22040 = and_21812 & ~or_21763;
  assign concat_22042 = {1'h0, add_22003};
  assign concat_22043 = {1'h0, sel_22005};
  assign concat_22047 = {1'h0, add_22010, array_index_21659[0]};
  assign concat_22048 = {1'h0, sel_22012};
  assign add_22060 = array_index_21939[11:1] + 11'h247;
  assign sel_22063 = and_21967 ? ($signed(concat_21932) < $signed(concat_21933) ? concat_21996 : sel_21901) : (eq_21874 | $signed(concat_21932) >= $signed(concat_21933) ? sel_21901 : concat_21996);
  assign eq_22068 = array_index_21939 == 16'h0000;
  assign add_22072 = array_index_22006[11:0] + 12'h247;
  assign sel_22074 = $signed({1'h0, add_21972}) < $signed({1'h0, sel_21974}) ? add_21972 : sel_21974;
  assign add_22080 = array_index_21782[11:1] + 11'h347;
  assign sel_22082 = and_21815 ? ($signed(concat_21952) < $signed(concat_21953) ? concat_22018 : sel_21919) : (eq_21736 | $signed(concat_21952) >= $signed(concat_21953) ? sel_21919 : concat_22018);
  assign concat_22087 = {add_21987, array_index_21782[2:0]};
  assign concat_22093 = {1'h0, add_22060, array_index_21939[0]};
  assign concat_22094 = {1'h0, sel_22063};
  assign array_index_22099 = set1_unflattened[4'h7];
  assign or_22100 = or_21873 | or_21908 & and_22040;
  assign array_index_22103 = set2_unflattened[4'h6];
  assign concat_22107 = {add_22010, array_index_21659[0]};
  assign add_22110 = array_index_21739[11:1] + 11'h79d;
  assign sel_22112 = $signed({1'h0, add_22014, array_index_21664[0]}) < $signed({1'h0, sel_22016}) ? {add_22014, array_index_21664[0]} : sel_22016;
  assign concat_22113 = {1'h0, add_22080, array_index_21782[0]};
  assign concat_22114 = {1'h0, sel_22082};
  assign add_22116 = array_index_21818[11:1] + 11'h347;
  assign sel_22118 = $signed({1'h0, add_22021, array_index_21739[0]}) < $signed({1'h0, sel_22023}) ? {add_22021, array_index_21739[0]} : sel_22023;
  assign add_22124 = array_index_21910[11:3] + 9'h0bd;
  assign sel_22127 = $signed({1'h0, add_22027, array_index_21818[2:0]}) < $signed({1'h0, sel_22030}) ? {add_22027, array_index_21818[2:0]} : sel_22030;
  assign add_22130 = array_index_22006[11:1] + 11'h247;
  assign sel_22133 = $signed({1'h0, add_22036, array_index_21910[0]}) < $signed({1'h0, sel_22039}) ? {add_22036, array_index_21910[0]} : sel_22039;
  assign or_22136 = or_22100 | eq_22068;
  assign sel_22137 = $signed(concat_22042) < $signed(concat_22043) ? add_22003 : sel_22005;
  assign add_22151 = array_index_21939[11:3] + 9'h0bd;
  assign sel_22154 = and_21967 ? ($signed(concat_22024) < $signed(concat_22025) ? concat_22087 : sel_21990) : (eq_21874 | $signed(concat_22024) >= $signed(concat_22025) ? sel_21990 : concat_22087);
  assign concat_22158 = {add_22060, array_index_21939[0]};
  assign add_22164 = array_index_22099[11:0] + 12'h247;
  assign add_22169 = array_index_22103[11:0] + 12'h247;
  assign sel_22171 = $signed({1'h0, add_22072}) < $signed({1'h0, sel_22074}) ? add_22072 : sel_22074;
  assign add_22173 = array_index_21782[11:1] + 11'h79d;
  assign sel_22175 = and_21815 ? ($signed(concat_22047) < $signed(concat_22048) ? concat_22107 : sel_22012) : (eq_21736 | $signed(concat_22047) >= $signed(concat_22048) ? sel_22012 : concat_22107);
  assign concat_22180 = {add_22080, array_index_21782[0]};
  assign concat_22185 = {1'h0, add_22151, array_index_21939[2:0]};
  assign concat_22186 = {1'h0, sel_22154};
  assign sel_22193 = $signed(concat_22093) < $signed(concat_22094) ? concat_22158 : sel_22063;
  assign array_index_22199 = set1_unflattened[4'h8];
  assign array_index_22202 = set2_unflattened[4'h7];
  assign concat_22205 = {1'h0, add_22173, array_index_21782[0]};
  assign concat_22206 = {1'h0, sel_22175};
  assign add_22208 = array_index_21818[11:1] + 11'h79d;
  assign sel_22210 = $signed({1'h0, add_22110, array_index_21739[0]}) < $signed({1'h0, sel_22112}) ? {add_22110, array_index_21739[0]} : sel_22112;
  assign add_22215 = array_index_21910[11:1] + 11'h347;
  assign sel_22217 = $signed({1'h0, add_22116, array_index_21818[0]}) < $signed({1'h0, sel_22118}) ? {add_22116, array_index_21818[0]} : sel_22118;
  assign add_22220 = array_index_22006[11:3] + 9'h0bd;
  assign sel_22223 = $signed({1'h0, add_22124, array_index_21910[2:0]}) < $signed({1'h0, sel_22127}) ? {add_22124, array_index_21910[2:0]} : sel_22127;
  assign add_22225 = array_index_22099[11:1] + 11'h247;
  assign add_22230 = array_index_22103[11:1] + 11'h247;
  assign sel_22233 = $signed({1'h0, add_22130, array_index_22006[0]}) < $signed({1'h0, sel_22133}) ? {add_22130, array_index_22006[0]} : sel_22133;
  assign add_22244 = array_index_21939[11:1] + 11'h347;
  assign sel_22246 = and_21967 ? ($signed(concat_22113) < $signed(concat_22114) ? concat_22180 : sel_22082) : (eq_21874 | $signed(concat_22113) >= $signed(concat_22114) ? sel_22082 : concat_22180);
  assign concat_22250 = {add_22151, array_index_21939[2:0]};
  assign add_22260 = array_index_22199[11:0] + 12'h247;
  assign sel_22262 = $signed({1'h0, add_22164}) < $signed({1'h0, or_22136 ? (eq_22068 | $signed(concat_22042) >= $signed(concat_22043) ? sel_22005 : add_22003) : sel_22137}) ? add_22164 : sel_22137;
  assign add_22265 = array_index_22202[11:0] + 12'h247;
  assign sel_22267 = $signed({1'h0, add_22169}) < $signed({1'h0, sel_22171}) ? add_22169 : sel_22171;
  assign concat_22269 = {add_22173, array_index_21782[0]};
  assign concat_22274 = {1'h0, add_22244, array_index_21939[0]};
  assign concat_22275 = {1'h0, sel_22246};
  assign sel_22281 = $signed(concat_22185) < $signed(concat_22186) ? concat_22250 : sel_22154;
  assign and_22295 = and_22040 & ~or_21908;
  assign array_index_22297 = set1_unflattened[4'h9];
  assign array_index_22300 = set2_unflattened[4'h8];
  assign add_22307 = array_index_21910[11:1] + 11'h79d;
  assign sel_22309 = $signed({1'h0, add_22208, array_index_21818[0]}) < $signed({1'h0, sel_22210}) ? {add_22208, array_index_21818[0]} : sel_22210;
  assign add_22312 = array_index_22006[11:1] + 11'h347;
  assign sel_22314 = $signed({1'h0, add_22215, array_index_21910[0]}) < $signed({1'h0, sel_22217}) ? {add_22215, array_index_21910[0]} : sel_22217;
  assign add_22316 = array_index_22099[11:3] + 9'h0bd;
  assign add_22321 = array_index_22103[11:3] + 9'h0bd;
  assign sel_22324 = $signed({1'h0, add_22220, array_index_22006[2:0]}) < $signed({1'h0, sel_22223}) ? {add_22220, array_index_22006[2:0]} : sel_22223;
  assign add_22326 = array_index_22199[11:1] + 11'h247;
  assign sel_22329 = $signed({1'h0, add_22225, array_index_22099[0]}) < $signed({1'h0, or_22136 ? (eq_22068 | $signed(concat_22093) >= $signed(concat_22094) ? sel_22063 : concat_22158) : sel_22193}) ? {add_22225, array_index_22099[0]} : sel_22193;
  assign add_22331 = array_index_22202[11:1] + 11'h247;
  assign sel_22334 = $signed({1'h0, add_22230, array_index_22103[0]}) < $signed({1'h0, sel_22233}) ? {add_22230, array_index_22103[0]} : sel_22233;
  assign add_22345 = array_index_21939[11:1] + 11'h79d;
  assign sel_22347 = and_21967 ? ($signed(concat_22205) < $signed(concat_22206) ? concat_22269 : sel_22175) : (eq_21874 | $signed(concat_22205) >= $signed(concat_22206) ? sel_22175 : concat_22269);
  assign concat_22351 = {add_22244, array_index_21939[0]};
  assign or_22364 = or_22100 | or_22136 & and_22295;
  assign add_22369 = array_index_22297[11:0] + 12'h247;
  assign sel_22371 = $signed({1'h0, add_22260}) < $signed({1'h0, sel_22262}) ? add_22260 : sel_22262;
  assign add_22374 = array_index_22300[11:0] + 12'h247;
  assign sel_22376 = $signed({1'h0, add_22265}) < $signed({1'h0, sel_22267}) ? add_22265 : sel_22267;
  assign concat_22377 = {1'h0, add_22345, array_index_21939[0]};
  assign concat_22378 = {1'h0, sel_22347};
  assign sel_22383 = $signed(concat_22274) < $signed(concat_22275) ? concat_22351 : sel_22246;
  assign or_22405 = or_22364 | array_index_22099 == 16'h0000;
  assign and_22406 = and_22295 & ~or_22136;
  assign concat_22410 = {1'h0, add_22369};
  assign concat_22411 = {1'h0, sel_22371};
  assign array_index_22412 = set2_unflattened[4'h9];
  assign add_22417 = array_index_22006[11:1] + 11'h79d;
  assign sel_22419 = $signed({1'h0, add_22307, array_index_21910[0]}) < $signed({1'h0, sel_22309}) ? {add_22307, array_index_21910[0]} : sel_22309;
  assign add_22421 = array_index_22099[11:1] + 11'h347;
  assign add_22425 = array_index_22103[11:1] + 11'h347;
  assign sel_22427 = $signed({1'h0, add_22312, array_index_22006[0]}) < $signed({1'h0, sel_22314}) ? {add_22312, array_index_22006[0]} : sel_22314;
  assign add_22429 = array_index_22199[11:3] + 9'h0bd;
  assign sel_22432 = $signed({1'h0, add_22316, array_index_22099[2:0]}) < $signed({1'h0, or_22136 ? (eq_22068 | $signed(concat_22185) >= $signed(concat_22186) ? sel_22154 : concat_22250) : sel_22281}) ? {add_22316, array_index_22099[2:0]} : sel_22281;
  assign add_22434 = array_index_22202[11:3] + 9'h0bd;
  assign sel_22437 = $signed({1'h0, add_22321, array_index_22103[2:0]}) < $signed({1'h0, sel_22324}) ? {add_22321, array_index_22103[2:0]} : sel_22324;
  assign add_22440 = array_index_22297[11:1] + 11'h247;
  assign sel_22443 = $signed({1'h0, add_22326, array_index_22199[0]}) < $signed({1'h0, sel_22329}) ? {add_22326, array_index_22199[0]} : sel_22329;
  assign add_22445 = array_index_22300[11:1] + 11'h247;
  assign sel_22448 = $signed({1'h0, add_22331, array_index_22202[0]}) < $signed({1'h0, sel_22334}) ? {add_22331, array_index_22202[0]} : sel_22334;
  assign eq_22452 = array_index_22297 == 16'h0000;
  assign concat_22458 = {add_22345, array_index_21939[0]};
  assign concat_22472 = {1'h0, add_22440, array_index_22297[0]};
  assign concat_22473 = {1'h0, sel_22443};
  assign add_22483 = array_index_22412[11:0] + 12'h247;
  assign sel_22485 = $signed({1'h0, add_22374}) < $signed({1'h0, sel_22376}) ? add_22374 : sel_22376;
  assign sel_22487 = $signed(concat_22377) < $signed(concat_22378) ? concat_22458 : sel_22347;
  assign and_22513 = and_22406 & ~or_22405;
  assign ne_22516 = array_index_22297 != 16'h0000;
  assign add_22522 = array_index_22099[11:1] + 11'h79d;
  assign add_22526 = array_index_22103[11:1] + 11'h79d;
  assign sel_22528 = $signed({1'h0, add_22417, array_index_22006[0]}) < $signed({1'h0, sel_22419}) ? {add_22417, array_index_22006[0]} : sel_22419;
  assign add_22530 = array_index_22199[11:1] + 11'h347;
  assign sel_22532 = $signed({1'h0, add_22421, array_index_22099[0]}) < $signed({1'h0, or_22136 ? (eq_22068 | $signed(concat_22274) >= $signed(concat_22275) ? sel_22246 : concat_22351) : sel_22383}) ? {add_22421, array_index_22099[0]} : sel_22383;
  assign add_22534 = array_index_22202[11:1] + 11'h347;
  assign sel_22536 = $signed({1'h0, add_22425, array_index_22103[0]}) < $signed({1'h0, sel_22427}) ? {add_22425, array_index_22103[0]} : sel_22427;
  assign add_22539 = array_index_22297[11:3] + 9'h0bd;
  assign sel_22542 = $signed({1'h0, add_22429, array_index_22199[2:0]}) < $signed({1'h0, sel_22432}) ? {add_22429, array_index_22199[2:0]} : sel_22432;
  assign add_22544 = array_index_22300[11:3] + 9'h0bd;
  assign sel_22547 = $signed({1'h0, add_22434, array_index_22202[2:0]}) < $signed({1'h0, sel_22437}) ? {add_22434, array_index_22202[2:0]} : sel_22437;
  assign concat_22550 = {add_22440, array_index_22297[0]};
  assign add_22553 = array_index_22412[11:1] + 11'h247;
  assign sel_22556 = $signed({1'h0, add_22445, array_index_22300[0]}) < $signed({1'h0, sel_22448}) ? {add_22445, array_index_22300[0]} : sel_22448;
  assign and_22557 = and_22513 & ~(or_22364 | or_22405 & and_22406 | array_index_22199 == 16'h0000);
  assign concat_22571 = {1'h0, add_22539, array_index_22297[2:0]};
  assign concat_22572 = {1'h0, sel_22542};
  assign add_22608 = array_index_22199[11:1] + 11'h79d;
  assign sel_22610 = $signed({1'h0, add_22522, array_index_22099[0]}) < $signed({1'h0, or_22136 ? (eq_22068 | $signed(concat_22377) >= $signed(concat_22378) ? sel_22347 : concat_22458) : sel_22487}) ? {add_22522, array_index_22099[0]} : sel_22487;
  assign add_22612 = array_index_22202[11:1] + 11'h79d;
  assign sel_22614 = $signed({1'h0, add_22526, array_index_22103[0]}) < $signed({1'h0, sel_22528}) ? {add_22526, array_index_22103[0]} : sel_22528;
  assign add_22617 = array_index_22297[11:1] + 11'h347;
  assign sel_22619 = $signed({1'h0, add_22530, array_index_22199[0]}) < $signed({1'h0, sel_22532}) ? {add_22530, array_index_22199[0]} : sel_22532;
  assign add_22621 = array_index_22300[11:1] + 11'h347;
  assign sel_22623 = $signed({1'h0, add_22534, array_index_22202[0]}) < $signed({1'h0, sel_22536}) ? {add_22534, array_index_22202[0]} : sel_22536;
  assign concat_22626 = {add_22539, array_index_22297[2:0]};
  assign add_22629 = array_index_22412[11:3] + 9'h0bd;
  assign sel_22632 = $signed({1'h0, add_22544, array_index_22300[2:0]}) < $signed({1'h0, sel_22547}) ? {add_22544, array_index_22300[2:0]} : sel_22547;
  assign concat_22635 = {1'h0, (and_22557 ? (ne_22516 ? ($signed(concat_22410) < $signed(concat_22411) ? add_22369 : sel_22371) : (eq_22452 | $signed(concat_22410) >= $signed(concat_22411) ? sel_22371 : add_22369)) : (and_22513 ? sel_22262 : (and_22406 ? sel_22137 : (and_22295 ? sel_22005 : (and_22040 ? sel_21850 : (and_21812 ? sel_21709 : (or_21589 ? (nor_21513 ? sel_21515 : (ne_21457 ? sel_21514 : sel_21458)) : sel_21590))))))) == ($signed({1'h0, add_22483}) < $signed({1'h0, sel_22485}) ? add_22483 : sel_22485)};
  assign concat_22643 = {1'h0, add_22617, array_index_22297[0]};
  assign concat_22644 = {1'h0, sel_22619};
  assign add_22653 = concat_22635 + 2'h1;
  assign add_22674 = array_index_22297[11:1] + 11'h79d;
  assign sel_22676 = $signed({1'h0, add_22608, array_index_22199[0]}) < $signed({1'h0, sel_22610}) ? {add_22608, array_index_22199[0]} : sel_22610;
  assign add_22678 = array_index_22300[11:1] + 11'h79d;
  assign sel_22680 = $signed({1'h0, add_22612, array_index_22202[0]}) < $signed({1'h0, sel_22614}) ? {add_22612, array_index_22202[0]} : sel_22614;
  assign concat_22683 = {add_22617, array_index_22297[0]};
  assign add_22686 = array_index_22412[11:1] + 11'h347;
  assign sel_22688 = $signed({1'h0, add_22621, array_index_22300[0]}) < $signed({1'h0, sel_22623}) ? {add_22621, array_index_22300[0]} : sel_22623;
  assign concat_22691 = {1'h0, (and_22557 ? (ne_22516 ? ($signed(concat_22472) < $signed(concat_22473) ? concat_22550 : sel_22443) : (eq_22452 | $signed(concat_22472) >= $signed(concat_22473) ? sel_22443 : concat_22550)) : (and_22513 ? sel_22329 : (and_22406 ? sel_22193 : (and_22295 ? sel_22063 : (and_22040 ? sel_21901 : (and_21812 ? sel_21755 : (or_21589 ? (nor_21513 ? sel_21543 : (ne_21457 ? sel_21542 : sel_21476)) : sel_21622))))))) == ($signed({1'h0, add_22553, array_index_22412[0]}) < $signed({1'h0, sel_22556}) ? {add_22553, array_index_22412[0]} : sel_22556) ? add_22653 : concat_22635};
  assign concat_22694 = {1'h0, add_22674, array_index_22297[0]};
  assign concat_22695 = {1'h0, sel_22676};
  assign add_22704 = concat_22691 + 3'h1;
  assign concat_22718 = {add_22674, array_index_22297[0]};
  assign add_22721 = array_index_22412[11:1] + 11'h79d;
  assign sel_22723 = $signed({1'h0, add_22678, array_index_22300[0]}) < $signed({1'h0, sel_22680}) ? {add_22678, array_index_22300[0]} : sel_22680;
  assign concat_22726 = {1'h0, (and_22557 ? (ne_22516 ? ($signed(concat_22571) < $signed(concat_22572) ? concat_22626 : sel_22542) : (eq_22452 | $signed(concat_22571) >= $signed(concat_22572) ? sel_22542 : concat_22626)) : (and_22513 ? sel_22432 : (and_22406 ? sel_22281 : (and_22295 ? sel_22154 : (and_22040 ? sel_21990 : (and_21812 ? sel_21831 : (or_21589 ? (nor_21513 ? sel_21585 : (ne_21457 ? sel_21584 : sel_21508)) : sel_21674))))))) == ($signed({1'h0, add_22629, array_index_22412[2:0]}) < $signed({1'h0, sel_22632}) ? {add_22629, array_index_22412[2:0]} : sel_22632) ? add_22704 : concat_22691};
  assign add_22734 = concat_22726 + 4'h1;
  assign concat_22743 = {1'h0, (and_22557 ? (ne_22516 ? ($signed(concat_22643) < $signed(concat_22644) ? concat_22683 : sel_22619) : (eq_22452 | $signed(concat_22643) >= $signed(concat_22644) ? sel_22619 : concat_22683)) : (and_22513 ? sel_22532 : (and_22406 ? sel_22383 : (and_22295 ? sel_22246 : (and_22040 ? sel_22082 : (and_21812 ? sel_21919 : (or_21589 ? (nor_21513 ? sel_21633 : (ne_21457 ? sel_21632 : sel_21550)) : sel_21745))))))) == ($signed({1'h0, add_22686, array_index_22412[0]}) < $signed({1'h0, sel_22688}) ? {add_22686, array_index_22412[0]} : sel_22688) ? add_22734 : concat_22726};
  assign add_22746 = concat_22743 + 5'h01;
  assign out = {{11'h000, (and_22557 ? (ne_22516 ? ($signed(concat_22694) < $signed(concat_22695) ? concat_22718 : sel_22676) : (eq_22452 | $signed(concat_22694) >= $signed(concat_22695) ? sel_22676 : concat_22718)) : (and_22513 ? sel_22610 : (and_22406 ? sel_22487 : (and_22295 ? sel_22347 : (and_22040 ? sel_22175 : (and_21812 ? sel_22012 : (or_21589 ? (nor_21513 ? sel_21692 : (ne_21457 ? sel_21691 : sel_21594)) : sel_21822))))))) == ($signed({1'h0, add_22721, array_index_22412[0]}) < $signed({1'h0, sel_22723}) ? {add_22721, array_index_22412[0]} : sel_22723) ? add_22746 : concat_22743}, {set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
