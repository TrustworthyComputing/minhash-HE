module min_hash(
  input wire [479:0] set1,
  input wire [479:0] set2,
  output wire [967:0] out
);
  wire [15:0] set1_unflattened[30];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  wire [15:0] set2_unflattened[30];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  wire [15:0] array_index_86651;
  wire [15:0] array_index_86652;
  wire [15:0] array_index_86656;
  wire [1:0] concat_86657;
  wire [1:0] add_86660;
  wire [15:0] array_index_86664;
  wire [2:0] concat_86665;
  wire [2:0] add_86668;
  wire [15:0] array_index_86672;
  wire [3:0] concat_86673;
  wire [3:0] add_86676;
  wire [15:0] array_index_86680;
  wire [4:0] concat_86681;
  wire [4:0] add_86684;
  wire [15:0] array_index_86688;
  wire [5:0] concat_86689;
  wire [5:0] add_86692;
  wire [15:0] array_index_86696;
  wire [6:0] concat_86697;
  wire [6:0] add_86700;
  wire [15:0] array_index_86704;
  wire [7:0] concat_86705;
  wire [7:0] add_86709;
  wire [15:0] array_index_86710;
  wire [7:0] sel_86711;
  wire [7:0] add_86715;
  wire [15:0] array_index_86716;
  wire [7:0] sel_86717;
  wire [7:0] add_86721;
  wire [15:0] array_index_86722;
  wire [7:0] sel_86723;
  wire [7:0] add_86727;
  wire [15:0] array_index_86728;
  wire [7:0] sel_86729;
  wire [7:0] add_86733;
  wire [15:0] array_index_86734;
  wire [7:0] sel_86735;
  wire [7:0] add_86739;
  wire [15:0] array_index_86740;
  wire [7:0] sel_86741;
  wire [7:0] add_86745;
  wire [15:0] array_index_86746;
  wire [7:0] sel_86747;
  wire [7:0] add_86751;
  wire [15:0] array_index_86752;
  wire [7:0] sel_86753;
  wire [7:0] add_86757;
  wire [15:0] array_index_86758;
  wire [7:0] sel_86759;
  wire [7:0] add_86763;
  wire [15:0] array_index_86764;
  wire [7:0] sel_86765;
  wire [7:0] add_86769;
  wire [15:0] array_index_86770;
  wire [7:0] sel_86771;
  wire [7:0] add_86775;
  wire [15:0] array_index_86776;
  wire [7:0] sel_86777;
  wire [7:0] add_86781;
  wire [15:0] array_index_86782;
  wire [7:0] sel_86783;
  wire [7:0] add_86787;
  wire [15:0] array_index_86788;
  wire [7:0] sel_86789;
  wire [7:0] add_86793;
  wire [15:0] array_index_86794;
  wire [7:0] sel_86795;
  wire [7:0] add_86799;
  wire [15:0] array_index_86800;
  wire [7:0] sel_86801;
  wire [7:0] add_86805;
  wire [15:0] array_index_86806;
  wire [7:0] sel_86807;
  wire [7:0] add_86811;
  wire [15:0] array_index_86812;
  wire [7:0] sel_86813;
  wire [7:0] add_86817;
  wire [15:0] array_index_86818;
  wire [7:0] sel_86819;
  wire [7:0] add_86823;
  wire [15:0] array_index_86824;
  wire [7:0] sel_86825;
  wire [7:0] add_86829;
  wire [15:0] array_index_86830;
  wire [7:0] sel_86831;
  wire [7:0] add_86835;
  wire [15:0] array_index_86836;
  wire [7:0] sel_86837;
  wire [7:0] add_86841;
  wire [15:0] array_index_86842;
  wire [7:0] sel_86843;
  wire [7:0] add_86846;
  wire [7:0] sel_86847;
  wire [7:0] add_86850;
  wire [7:0] sel_86851;
  wire [7:0] add_86854;
  wire [7:0] sel_86855;
  wire [7:0] add_86858;
  wire [7:0] sel_86859;
  wire [7:0] add_86862;
  wire [7:0] sel_86863;
  wire [7:0] add_86866;
  wire [7:0] sel_86867;
  wire [7:0] add_86870;
  wire [7:0] sel_86871;
  wire [7:0] add_86874;
  wire [7:0] sel_86875;
  wire [7:0] add_86878;
  wire [7:0] sel_86879;
  wire [7:0] add_86882;
  wire [7:0] sel_86883;
  wire [7:0] add_86886;
  wire [7:0] sel_86887;
  wire [7:0] add_86890;
  wire [7:0] sel_86891;
  wire [7:0] add_86894;
  wire [7:0] sel_86895;
  wire [7:0] add_86898;
  wire [7:0] sel_86899;
  wire [7:0] add_86902;
  wire [7:0] sel_86903;
  wire [7:0] add_86906;
  wire [7:0] sel_86907;
  wire [7:0] add_86910;
  wire [7:0] sel_86911;
  wire [7:0] add_86914;
  wire [7:0] sel_86915;
  wire [7:0] add_86918;
  wire [7:0] sel_86919;
  wire [7:0] add_86922;
  wire [7:0] sel_86923;
  wire [7:0] add_86926;
  wire [7:0] sel_86927;
  wire [7:0] add_86930;
  wire [7:0] sel_86931;
  wire [7:0] add_86934;
  wire [7:0] sel_86935;
  wire [7:0] add_86938;
  wire [7:0] sel_86939;
  wire [7:0] add_86942;
  wire [7:0] sel_86943;
  wire [7:0] add_86946;
  wire [7:0] sel_86947;
  wire [7:0] add_86950;
  wire [7:0] sel_86951;
  wire [7:0] add_86954;
  wire [7:0] sel_86955;
  wire [7:0] add_86958;
  wire [7:0] sel_86959;
  wire [7:0] add_86963;
  wire [15:0] array_index_86964;
  wire [7:0] sel_86965;
  wire [7:0] add_86968;
  wire [7:0] sel_86969;
  wire [7:0] add_86972;
  wire [7:0] sel_86973;
  wire [7:0] add_86976;
  wire [7:0] sel_86977;
  wire [7:0] add_86980;
  wire [7:0] sel_86981;
  wire [7:0] add_86984;
  wire [7:0] sel_86985;
  wire [7:0] add_86988;
  wire [7:0] sel_86989;
  wire [7:0] add_86992;
  wire [7:0] sel_86993;
  wire [7:0] add_86996;
  wire [7:0] sel_86997;
  wire [7:0] add_87000;
  wire [7:0] sel_87001;
  wire [7:0] add_87004;
  wire [7:0] sel_87005;
  wire [7:0] add_87008;
  wire [7:0] sel_87009;
  wire [7:0] add_87012;
  wire [7:0] sel_87013;
  wire [7:0] add_87016;
  wire [7:0] sel_87017;
  wire [7:0] add_87020;
  wire [7:0] sel_87021;
  wire [7:0] add_87024;
  wire [7:0] sel_87025;
  wire [7:0] add_87028;
  wire [7:0] sel_87029;
  wire [7:0] add_87032;
  wire [7:0] sel_87033;
  wire [7:0] add_87036;
  wire [7:0] sel_87037;
  wire [7:0] add_87040;
  wire [7:0] sel_87041;
  wire [7:0] add_87044;
  wire [7:0] sel_87045;
  wire [7:0] add_87048;
  wire [7:0] sel_87049;
  wire [7:0] add_87052;
  wire [7:0] sel_87053;
  wire [7:0] add_87056;
  wire [7:0] sel_87057;
  wire [7:0] add_87060;
  wire [7:0] sel_87061;
  wire [7:0] add_87064;
  wire [7:0] sel_87065;
  wire [7:0] add_87068;
  wire [7:0] sel_87069;
  wire [7:0] add_87072;
  wire [7:0] sel_87073;
  wire [7:0] add_87076;
  wire [7:0] sel_87077;
  wire [7:0] add_87080;
  wire [7:0] sel_87081;
  wire [7:0] add_87085;
  wire [15:0] array_index_87086;
  wire [7:0] sel_87087;
  wire [7:0] add_87090;
  wire [7:0] sel_87091;
  wire [7:0] add_87094;
  wire [7:0] sel_87095;
  wire [7:0] add_87098;
  wire [7:0] sel_87099;
  wire [7:0] add_87102;
  wire [7:0] sel_87103;
  wire [7:0] add_87106;
  wire [7:0] sel_87107;
  wire [7:0] add_87110;
  wire [7:0] sel_87111;
  wire [7:0] add_87114;
  wire [7:0] sel_87115;
  wire [7:0] add_87118;
  wire [7:0] sel_87119;
  wire [7:0] add_87122;
  wire [7:0] sel_87123;
  wire [7:0] add_87126;
  wire [7:0] sel_87127;
  wire [7:0] add_87130;
  wire [7:0] sel_87131;
  wire [7:0] add_87134;
  wire [7:0] sel_87135;
  wire [7:0] add_87138;
  wire [7:0] sel_87139;
  wire [7:0] add_87142;
  wire [7:0] sel_87143;
  wire [7:0] add_87146;
  wire [7:0] sel_87147;
  wire [7:0] add_87150;
  wire [7:0] sel_87151;
  wire [7:0] add_87154;
  wire [7:0] sel_87155;
  wire [7:0] add_87158;
  wire [7:0] sel_87159;
  wire [7:0] add_87162;
  wire [7:0] sel_87163;
  wire [7:0] add_87166;
  wire [7:0] sel_87167;
  wire [7:0] add_87170;
  wire [7:0] sel_87171;
  wire [7:0] add_87174;
  wire [7:0] sel_87175;
  wire [7:0] add_87178;
  wire [7:0] sel_87179;
  wire [7:0] add_87182;
  wire [7:0] sel_87183;
  wire [7:0] add_87186;
  wire [7:0] sel_87187;
  wire [7:0] add_87190;
  wire [7:0] sel_87191;
  wire [7:0] add_87194;
  wire [7:0] sel_87195;
  wire [7:0] add_87198;
  wire [7:0] sel_87199;
  wire [7:0] add_87202;
  wire [7:0] sel_87203;
  wire [7:0] add_87207;
  wire [15:0] array_index_87208;
  wire [7:0] sel_87209;
  wire [7:0] add_87212;
  wire [7:0] sel_87213;
  wire [7:0] add_87216;
  wire [7:0] sel_87217;
  wire [7:0] add_87220;
  wire [7:0] sel_87221;
  wire [7:0] add_87224;
  wire [7:0] sel_87225;
  wire [7:0] add_87228;
  wire [7:0] sel_87229;
  wire [7:0] add_87232;
  wire [7:0] sel_87233;
  wire [7:0] add_87236;
  wire [7:0] sel_87237;
  wire [7:0] add_87240;
  wire [7:0] sel_87241;
  wire [7:0] add_87244;
  wire [7:0] sel_87245;
  wire [7:0] add_87248;
  wire [7:0] sel_87249;
  wire [7:0] add_87252;
  wire [7:0] sel_87253;
  wire [7:0] add_87256;
  wire [7:0] sel_87257;
  wire [7:0] add_87260;
  wire [7:0] sel_87261;
  wire [7:0] add_87264;
  wire [7:0] sel_87265;
  wire [7:0] add_87268;
  wire [7:0] sel_87269;
  wire [7:0] add_87272;
  wire [7:0] sel_87273;
  wire [7:0] add_87276;
  wire [7:0] sel_87277;
  wire [7:0] add_87280;
  wire [7:0] sel_87281;
  wire [7:0] add_87284;
  wire [7:0] sel_87285;
  wire [7:0] add_87288;
  wire [7:0] sel_87289;
  wire [7:0] add_87292;
  wire [7:0] sel_87293;
  wire [7:0] add_87296;
  wire [7:0] sel_87297;
  wire [7:0] add_87300;
  wire [7:0] sel_87301;
  wire [7:0] add_87304;
  wire [7:0] sel_87305;
  wire [7:0] add_87308;
  wire [7:0] sel_87309;
  wire [7:0] add_87312;
  wire [7:0] sel_87313;
  wire [7:0] add_87316;
  wire [7:0] sel_87317;
  wire [7:0] add_87320;
  wire [7:0] sel_87321;
  wire [7:0] add_87324;
  wire [7:0] sel_87325;
  wire [7:0] add_87329;
  wire [15:0] array_index_87330;
  wire [7:0] sel_87331;
  wire [7:0] add_87334;
  wire [7:0] sel_87335;
  wire [7:0] add_87338;
  wire [7:0] sel_87339;
  wire [7:0] add_87342;
  wire [7:0] sel_87343;
  wire [7:0] add_87346;
  wire [7:0] sel_87347;
  wire [7:0] add_87350;
  wire [7:0] sel_87351;
  wire [7:0] add_87354;
  wire [7:0] sel_87355;
  wire [7:0] add_87358;
  wire [7:0] sel_87359;
  wire [7:0] add_87362;
  wire [7:0] sel_87363;
  wire [7:0] add_87366;
  wire [7:0] sel_87367;
  wire [7:0] add_87370;
  wire [7:0] sel_87371;
  wire [7:0] add_87374;
  wire [7:0] sel_87375;
  wire [7:0] add_87378;
  wire [7:0] sel_87379;
  wire [7:0] add_87382;
  wire [7:0] sel_87383;
  wire [7:0] add_87386;
  wire [7:0] sel_87387;
  wire [7:0] add_87390;
  wire [7:0] sel_87391;
  wire [7:0] add_87394;
  wire [7:0] sel_87395;
  wire [7:0] add_87398;
  wire [7:0] sel_87399;
  wire [7:0] add_87402;
  wire [7:0] sel_87403;
  wire [7:0] add_87406;
  wire [7:0] sel_87407;
  wire [7:0] add_87410;
  wire [7:0] sel_87411;
  wire [7:0] add_87414;
  wire [7:0] sel_87415;
  wire [7:0] add_87418;
  wire [7:0] sel_87419;
  wire [7:0] add_87422;
  wire [7:0] sel_87423;
  wire [7:0] add_87426;
  wire [7:0] sel_87427;
  wire [7:0] add_87430;
  wire [7:0] sel_87431;
  wire [7:0] add_87434;
  wire [7:0] sel_87435;
  wire [7:0] add_87438;
  wire [7:0] sel_87439;
  wire [7:0] add_87442;
  wire [7:0] sel_87443;
  wire [7:0] add_87446;
  wire [7:0] sel_87447;
  wire [7:0] add_87451;
  wire [15:0] array_index_87452;
  wire [7:0] sel_87453;
  wire [7:0] add_87456;
  wire [7:0] sel_87457;
  wire [7:0] add_87460;
  wire [7:0] sel_87461;
  wire [7:0] add_87464;
  wire [7:0] sel_87465;
  wire [7:0] add_87468;
  wire [7:0] sel_87469;
  wire [7:0] add_87472;
  wire [7:0] sel_87473;
  wire [7:0] add_87476;
  wire [7:0] sel_87477;
  wire [7:0] add_87480;
  wire [7:0] sel_87481;
  wire [7:0] add_87484;
  wire [7:0] sel_87485;
  wire [7:0] add_87488;
  wire [7:0] sel_87489;
  wire [7:0] add_87492;
  wire [7:0] sel_87493;
  wire [7:0] add_87496;
  wire [7:0] sel_87497;
  wire [7:0] add_87500;
  wire [7:0] sel_87501;
  wire [7:0] add_87504;
  wire [7:0] sel_87505;
  wire [7:0] add_87508;
  wire [7:0] sel_87509;
  wire [7:0] add_87512;
  wire [7:0] sel_87513;
  wire [7:0] add_87516;
  wire [7:0] sel_87517;
  wire [7:0] add_87520;
  wire [7:0] sel_87521;
  wire [7:0] add_87524;
  wire [7:0] sel_87525;
  wire [7:0] add_87528;
  wire [7:0] sel_87529;
  wire [7:0] add_87532;
  wire [7:0] sel_87533;
  wire [7:0] add_87536;
  wire [7:0] sel_87537;
  wire [7:0] add_87540;
  wire [7:0] sel_87541;
  wire [7:0] add_87544;
  wire [7:0] sel_87545;
  wire [7:0] add_87548;
  wire [7:0] sel_87549;
  wire [7:0] add_87552;
  wire [7:0] sel_87553;
  wire [7:0] add_87556;
  wire [7:0] sel_87557;
  wire [7:0] add_87560;
  wire [7:0] sel_87561;
  wire [7:0] add_87564;
  wire [7:0] sel_87565;
  wire [7:0] add_87568;
  wire [7:0] sel_87569;
  wire [7:0] add_87573;
  wire [15:0] array_index_87574;
  wire [7:0] sel_87575;
  wire [7:0] add_87578;
  wire [7:0] sel_87579;
  wire [7:0] add_87582;
  wire [7:0] sel_87583;
  wire [7:0] add_87586;
  wire [7:0] sel_87587;
  wire [7:0] add_87590;
  wire [7:0] sel_87591;
  wire [7:0] add_87594;
  wire [7:0] sel_87595;
  wire [7:0] add_87598;
  wire [7:0] sel_87599;
  wire [7:0] add_87602;
  wire [7:0] sel_87603;
  wire [7:0] add_87606;
  wire [7:0] sel_87607;
  wire [7:0] add_87610;
  wire [7:0] sel_87611;
  wire [7:0] add_87614;
  wire [7:0] sel_87615;
  wire [7:0] add_87618;
  wire [7:0] sel_87619;
  wire [7:0] add_87622;
  wire [7:0] sel_87623;
  wire [7:0] add_87626;
  wire [7:0] sel_87627;
  wire [7:0] add_87630;
  wire [7:0] sel_87631;
  wire [7:0] add_87634;
  wire [7:0] sel_87635;
  wire [7:0] add_87638;
  wire [7:0] sel_87639;
  wire [7:0] add_87642;
  wire [7:0] sel_87643;
  wire [7:0] add_87646;
  wire [7:0] sel_87647;
  wire [7:0] add_87650;
  wire [7:0] sel_87651;
  wire [7:0] add_87654;
  wire [7:0] sel_87655;
  wire [7:0] add_87658;
  wire [7:0] sel_87659;
  wire [7:0] add_87662;
  wire [7:0] sel_87663;
  wire [7:0] add_87666;
  wire [7:0] sel_87667;
  wire [7:0] add_87670;
  wire [7:0] sel_87671;
  wire [7:0] add_87674;
  wire [7:0] sel_87675;
  wire [7:0] add_87678;
  wire [7:0] sel_87679;
  wire [7:0] add_87682;
  wire [7:0] sel_87683;
  wire [7:0] add_87686;
  wire [7:0] sel_87687;
  wire [7:0] add_87690;
  wire [7:0] sel_87691;
  wire [7:0] add_87695;
  wire [15:0] array_index_87696;
  wire [7:0] sel_87697;
  wire [7:0] add_87700;
  wire [7:0] sel_87701;
  wire [7:0] add_87704;
  wire [7:0] sel_87705;
  wire [7:0] add_87708;
  wire [7:0] sel_87709;
  wire [7:0] add_87712;
  wire [7:0] sel_87713;
  wire [7:0] add_87716;
  wire [7:0] sel_87717;
  wire [7:0] add_87720;
  wire [7:0] sel_87721;
  wire [7:0] add_87724;
  wire [7:0] sel_87725;
  wire [7:0] add_87728;
  wire [7:0] sel_87729;
  wire [7:0] add_87732;
  wire [7:0] sel_87733;
  wire [7:0] add_87736;
  wire [7:0] sel_87737;
  wire [7:0] add_87740;
  wire [7:0] sel_87741;
  wire [7:0] add_87744;
  wire [7:0] sel_87745;
  wire [7:0] add_87748;
  wire [7:0] sel_87749;
  wire [7:0] add_87752;
  wire [7:0] sel_87753;
  wire [7:0] add_87756;
  wire [7:0] sel_87757;
  wire [7:0] add_87760;
  wire [7:0] sel_87761;
  wire [7:0] add_87764;
  wire [7:0] sel_87765;
  wire [7:0] add_87768;
  wire [7:0] sel_87769;
  wire [7:0] add_87772;
  wire [7:0] sel_87773;
  wire [7:0] add_87776;
  wire [7:0] sel_87777;
  wire [7:0] add_87780;
  wire [7:0] sel_87781;
  wire [7:0] add_87784;
  wire [7:0] sel_87785;
  wire [7:0] add_87788;
  wire [7:0] sel_87789;
  wire [7:0] add_87792;
  wire [7:0] sel_87793;
  wire [7:0] add_87796;
  wire [7:0] sel_87797;
  wire [7:0] add_87800;
  wire [7:0] sel_87801;
  wire [7:0] add_87804;
  wire [7:0] sel_87805;
  wire [7:0] add_87808;
  wire [7:0] sel_87809;
  wire [7:0] add_87812;
  wire [7:0] sel_87813;
  wire [7:0] add_87817;
  wire [15:0] array_index_87818;
  wire [7:0] sel_87819;
  wire [7:0] add_87822;
  wire [7:0] sel_87823;
  wire [7:0] add_87826;
  wire [7:0] sel_87827;
  wire [7:0] add_87830;
  wire [7:0] sel_87831;
  wire [7:0] add_87834;
  wire [7:0] sel_87835;
  wire [7:0] add_87838;
  wire [7:0] sel_87839;
  wire [7:0] add_87842;
  wire [7:0] sel_87843;
  wire [7:0] add_87846;
  wire [7:0] sel_87847;
  wire [7:0] add_87850;
  wire [7:0] sel_87851;
  wire [7:0] add_87854;
  wire [7:0] sel_87855;
  wire [7:0] add_87858;
  wire [7:0] sel_87859;
  wire [7:0] add_87862;
  wire [7:0] sel_87863;
  wire [7:0] add_87866;
  wire [7:0] sel_87867;
  wire [7:0] add_87870;
  wire [7:0] sel_87871;
  wire [7:0] add_87874;
  wire [7:0] sel_87875;
  wire [7:0] add_87878;
  wire [7:0] sel_87879;
  wire [7:0] add_87882;
  wire [7:0] sel_87883;
  wire [7:0] add_87886;
  wire [7:0] sel_87887;
  wire [7:0] add_87890;
  wire [7:0] sel_87891;
  wire [7:0] add_87894;
  wire [7:0] sel_87895;
  wire [7:0] add_87898;
  wire [7:0] sel_87899;
  wire [7:0] add_87902;
  wire [7:0] sel_87903;
  wire [7:0] add_87906;
  wire [7:0] sel_87907;
  wire [7:0] add_87910;
  wire [7:0] sel_87911;
  wire [7:0] add_87914;
  wire [7:0] sel_87915;
  wire [7:0] add_87918;
  wire [7:0] sel_87919;
  wire [7:0] add_87922;
  wire [7:0] sel_87923;
  wire [7:0] add_87926;
  wire [7:0] sel_87927;
  wire [7:0] add_87930;
  wire [7:0] sel_87931;
  wire [7:0] add_87934;
  wire [7:0] sel_87935;
  wire [7:0] add_87939;
  wire [15:0] array_index_87940;
  wire [7:0] sel_87941;
  wire [7:0] add_87944;
  wire [7:0] sel_87945;
  wire [7:0] add_87948;
  wire [7:0] sel_87949;
  wire [7:0] add_87952;
  wire [7:0] sel_87953;
  wire [7:0] add_87956;
  wire [7:0] sel_87957;
  wire [7:0] add_87960;
  wire [7:0] sel_87961;
  wire [7:0] add_87964;
  wire [7:0] sel_87965;
  wire [7:0] add_87968;
  wire [7:0] sel_87969;
  wire [7:0] add_87972;
  wire [7:0] sel_87973;
  wire [7:0] add_87976;
  wire [7:0] sel_87977;
  wire [7:0] add_87980;
  wire [7:0] sel_87981;
  wire [7:0] add_87984;
  wire [7:0] sel_87985;
  wire [7:0] add_87988;
  wire [7:0] sel_87989;
  wire [7:0] add_87992;
  wire [7:0] sel_87993;
  wire [7:0] add_87996;
  wire [7:0] sel_87997;
  wire [7:0] add_88000;
  wire [7:0] sel_88001;
  wire [7:0] add_88004;
  wire [7:0] sel_88005;
  wire [7:0] add_88008;
  wire [7:0] sel_88009;
  wire [7:0] add_88012;
  wire [7:0] sel_88013;
  wire [7:0] add_88016;
  wire [7:0] sel_88017;
  wire [7:0] add_88020;
  wire [7:0] sel_88021;
  wire [7:0] add_88024;
  wire [7:0] sel_88025;
  wire [7:0] add_88028;
  wire [7:0] sel_88029;
  wire [7:0] add_88032;
  wire [7:0] sel_88033;
  wire [7:0] add_88036;
  wire [7:0] sel_88037;
  wire [7:0] add_88040;
  wire [7:0] sel_88041;
  wire [7:0] add_88044;
  wire [7:0] sel_88045;
  wire [7:0] add_88048;
  wire [7:0] sel_88049;
  wire [7:0] add_88052;
  wire [7:0] sel_88053;
  wire [7:0] add_88056;
  wire [7:0] sel_88057;
  wire [7:0] add_88061;
  wire [15:0] array_index_88062;
  wire [7:0] sel_88063;
  wire [7:0] add_88066;
  wire [7:0] sel_88067;
  wire [7:0] add_88070;
  wire [7:0] sel_88071;
  wire [7:0] add_88074;
  wire [7:0] sel_88075;
  wire [7:0] add_88078;
  wire [7:0] sel_88079;
  wire [7:0] add_88082;
  wire [7:0] sel_88083;
  wire [7:0] add_88086;
  wire [7:0] sel_88087;
  wire [7:0] add_88090;
  wire [7:0] sel_88091;
  wire [7:0] add_88094;
  wire [7:0] sel_88095;
  wire [7:0] add_88098;
  wire [7:0] sel_88099;
  wire [7:0] add_88102;
  wire [7:0] sel_88103;
  wire [7:0] add_88106;
  wire [7:0] sel_88107;
  wire [7:0] add_88110;
  wire [7:0] sel_88111;
  wire [7:0] add_88114;
  wire [7:0] sel_88115;
  wire [7:0] add_88118;
  wire [7:0] sel_88119;
  wire [7:0] add_88122;
  wire [7:0] sel_88123;
  wire [7:0] add_88126;
  wire [7:0] sel_88127;
  wire [7:0] add_88130;
  wire [7:0] sel_88131;
  wire [7:0] add_88134;
  wire [7:0] sel_88135;
  wire [7:0] add_88138;
  wire [7:0] sel_88139;
  wire [7:0] add_88142;
  wire [7:0] sel_88143;
  wire [7:0] add_88146;
  wire [7:0] sel_88147;
  wire [7:0] add_88150;
  wire [7:0] sel_88151;
  wire [7:0] add_88154;
  wire [7:0] sel_88155;
  wire [7:0] add_88158;
  wire [7:0] sel_88159;
  wire [7:0] add_88162;
  wire [7:0] sel_88163;
  wire [7:0] add_88166;
  wire [7:0] sel_88167;
  wire [7:0] add_88170;
  wire [7:0] sel_88171;
  wire [7:0] add_88174;
  wire [7:0] sel_88175;
  wire [7:0] add_88178;
  wire [7:0] sel_88179;
  wire [7:0] add_88183;
  wire [15:0] array_index_88184;
  wire [7:0] sel_88185;
  wire [7:0] add_88188;
  wire [7:0] sel_88189;
  wire [7:0] add_88192;
  wire [7:0] sel_88193;
  wire [7:0] add_88196;
  wire [7:0] sel_88197;
  wire [7:0] add_88200;
  wire [7:0] sel_88201;
  wire [7:0] add_88204;
  wire [7:0] sel_88205;
  wire [7:0] add_88208;
  wire [7:0] sel_88209;
  wire [7:0] add_88212;
  wire [7:0] sel_88213;
  wire [7:0] add_88216;
  wire [7:0] sel_88217;
  wire [7:0] add_88220;
  wire [7:0] sel_88221;
  wire [7:0] add_88224;
  wire [7:0] sel_88225;
  wire [7:0] add_88228;
  wire [7:0] sel_88229;
  wire [7:0] add_88232;
  wire [7:0] sel_88233;
  wire [7:0] add_88236;
  wire [7:0] sel_88237;
  wire [7:0] add_88240;
  wire [7:0] sel_88241;
  wire [7:0] add_88244;
  wire [7:0] sel_88245;
  wire [7:0] add_88248;
  wire [7:0] sel_88249;
  wire [7:0] add_88252;
  wire [7:0] sel_88253;
  wire [7:0] add_88256;
  wire [7:0] sel_88257;
  wire [7:0] add_88260;
  wire [7:0] sel_88261;
  wire [7:0] add_88264;
  wire [7:0] sel_88265;
  wire [7:0] add_88268;
  wire [7:0] sel_88269;
  wire [7:0] add_88272;
  wire [7:0] sel_88273;
  wire [7:0] add_88276;
  wire [7:0] sel_88277;
  wire [7:0] add_88280;
  wire [7:0] sel_88281;
  wire [7:0] add_88284;
  wire [7:0] sel_88285;
  wire [7:0] add_88288;
  wire [7:0] sel_88289;
  wire [7:0] add_88292;
  wire [7:0] sel_88293;
  wire [7:0] add_88296;
  wire [7:0] sel_88297;
  wire [7:0] add_88300;
  wire [7:0] sel_88301;
  wire [7:0] add_88305;
  wire [15:0] array_index_88306;
  wire [7:0] sel_88307;
  wire [7:0] add_88310;
  wire [7:0] sel_88311;
  wire [7:0] add_88314;
  wire [7:0] sel_88315;
  wire [7:0] add_88318;
  wire [7:0] sel_88319;
  wire [7:0] add_88322;
  wire [7:0] sel_88323;
  wire [7:0] add_88326;
  wire [7:0] sel_88327;
  wire [7:0] add_88330;
  wire [7:0] sel_88331;
  wire [7:0] add_88334;
  wire [7:0] sel_88335;
  wire [7:0] add_88338;
  wire [7:0] sel_88339;
  wire [7:0] add_88342;
  wire [7:0] sel_88343;
  wire [7:0] add_88346;
  wire [7:0] sel_88347;
  wire [7:0] add_88350;
  wire [7:0] sel_88351;
  wire [7:0] add_88354;
  wire [7:0] sel_88355;
  wire [7:0] add_88358;
  wire [7:0] sel_88359;
  wire [7:0] add_88362;
  wire [7:0] sel_88363;
  wire [7:0] add_88366;
  wire [7:0] sel_88367;
  wire [7:0] add_88370;
  wire [7:0] sel_88371;
  wire [7:0] add_88374;
  wire [7:0] sel_88375;
  wire [7:0] add_88378;
  wire [7:0] sel_88379;
  wire [7:0] add_88382;
  wire [7:0] sel_88383;
  wire [7:0] add_88386;
  wire [7:0] sel_88387;
  wire [7:0] add_88390;
  wire [7:0] sel_88391;
  wire [7:0] add_88394;
  wire [7:0] sel_88395;
  wire [7:0] add_88398;
  wire [7:0] sel_88399;
  wire [7:0] add_88402;
  wire [7:0] sel_88403;
  wire [7:0] add_88406;
  wire [7:0] sel_88407;
  wire [7:0] add_88410;
  wire [7:0] sel_88411;
  wire [7:0] add_88414;
  wire [7:0] sel_88415;
  wire [7:0] add_88418;
  wire [7:0] sel_88419;
  wire [7:0] add_88422;
  wire [7:0] sel_88423;
  wire [7:0] add_88427;
  wire [15:0] array_index_88428;
  wire [7:0] sel_88429;
  wire [7:0] add_88432;
  wire [7:0] sel_88433;
  wire [7:0] add_88436;
  wire [7:0] sel_88437;
  wire [7:0] add_88440;
  wire [7:0] sel_88441;
  wire [7:0] add_88444;
  wire [7:0] sel_88445;
  wire [7:0] add_88448;
  wire [7:0] sel_88449;
  wire [7:0] add_88452;
  wire [7:0] sel_88453;
  wire [7:0] add_88456;
  wire [7:0] sel_88457;
  wire [7:0] add_88460;
  wire [7:0] sel_88461;
  wire [7:0] add_88464;
  wire [7:0] sel_88465;
  wire [7:0] add_88468;
  wire [7:0] sel_88469;
  wire [7:0] add_88472;
  wire [7:0] sel_88473;
  wire [7:0] add_88476;
  wire [7:0] sel_88477;
  wire [7:0] add_88480;
  wire [7:0] sel_88481;
  wire [7:0] add_88484;
  wire [7:0] sel_88485;
  wire [7:0] add_88488;
  wire [7:0] sel_88489;
  wire [7:0] add_88492;
  wire [7:0] sel_88493;
  wire [7:0] add_88496;
  wire [7:0] sel_88497;
  wire [7:0] add_88500;
  wire [7:0] sel_88501;
  wire [7:0] add_88504;
  wire [7:0] sel_88505;
  wire [7:0] add_88508;
  wire [7:0] sel_88509;
  wire [7:0] add_88512;
  wire [7:0] sel_88513;
  wire [7:0] add_88516;
  wire [7:0] sel_88517;
  wire [7:0] add_88520;
  wire [7:0] sel_88521;
  wire [7:0] add_88524;
  wire [7:0] sel_88525;
  wire [7:0] add_88528;
  wire [7:0] sel_88529;
  wire [7:0] add_88532;
  wire [7:0] sel_88533;
  wire [7:0] add_88536;
  wire [7:0] sel_88537;
  wire [7:0] add_88540;
  wire [7:0] sel_88541;
  wire [7:0] add_88544;
  wire [7:0] sel_88545;
  wire [7:0] add_88549;
  wire [15:0] array_index_88550;
  wire [7:0] sel_88551;
  wire [7:0] add_88554;
  wire [7:0] sel_88555;
  wire [7:0] add_88558;
  wire [7:0] sel_88559;
  wire [7:0] add_88562;
  wire [7:0] sel_88563;
  wire [7:0] add_88566;
  wire [7:0] sel_88567;
  wire [7:0] add_88570;
  wire [7:0] sel_88571;
  wire [7:0] add_88574;
  wire [7:0] sel_88575;
  wire [7:0] add_88578;
  wire [7:0] sel_88579;
  wire [7:0] add_88582;
  wire [7:0] sel_88583;
  wire [7:0] add_88586;
  wire [7:0] sel_88587;
  wire [7:0] add_88590;
  wire [7:0] sel_88591;
  wire [7:0] add_88594;
  wire [7:0] sel_88595;
  wire [7:0] add_88598;
  wire [7:0] sel_88599;
  wire [7:0] add_88602;
  wire [7:0] sel_88603;
  wire [7:0] add_88606;
  wire [7:0] sel_88607;
  wire [7:0] add_88610;
  wire [7:0] sel_88611;
  wire [7:0] add_88614;
  wire [7:0] sel_88615;
  wire [7:0] add_88618;
  wire [7:0] sel_88619;
  wire [7:0] add_88622;
  wire [7:0] sel_88623;
  wire [7:0] add_88626;
  wire [7:0] sel_88627;
  wire [7:0] add_88630;
  wire [7:0] sel_88631;
  wire [7:0] add_88634;
  wire [7:0] sel_88635;
  wire [7:0] add_88638;
  wire [7:0] sel_88639;
  wire [7:0] add_88642;
  wire [7:0] sel_88643;
  wire [7:0] add_88646;
  wire [7:0] sel_88647;
  wire [7:0] add_88650;
  wire [7:0] sel_88651;
  wire [7:0] add_88654;
  wire [7:0] sel_88655;
  wire [7:0] add_88658;
  wire [7:0] sel_88659;
  wire [7:0] add_88662;
  wire [7:0] sel_88663;
  wire [7:0] add_88666;
  wire [7:0] sel_88667;
  wire [7:0] add_88671;
  wire [15:0] array_index_88672;
  wire [7:0] sel_88673;
  wire [7:0] add_88676;
  wire [7:0] sel_88677;
  wire [7:0] add_88680;
  wire [7:0] sel_88681;
  wire [7:0] add_88684;
  wire [7:0] sel_88685;
  wire [7:0] add_88688;
  wire [7:0] sel_88689;
  wire [7:0] add_88692;
  wire [7:0] sel_88693;
  wire [7:0] add_88696;
  wire [7:0] sel_88697;
  wire [7:0] add_88700;
  wire [7:0] sel_88701;
  wire [7:0] add_88704;
  wire [7:0] sel_88705;
  wire [7:0] add_88708;
  wire [7:0] sel_88709;
  wire [7:0] add_88712;
  wire [7:0] sel_88713;
  wire [7:0] add_88716;
  wire [7:0] sel_88717;
  wire [7:0] add_88720;
  wire [7:0] sel_88721;
  wire [7:0] add_88724;
  wire [7:0] sel_88725;
  wire [7:0] add_88728;
  wire [7:0] sel_88729;
  wire [7:0] add_88732;
  wire [7:0] sel_88733;
  wire [7:0] add_88736;
  wire [7:0] sel_88737;
  wire [7:0] add_88740;
  wire [7:0] sel_88741;
  wire [7:0] add_88744;
  wire [7:0] sel_88745;
  wire [7:0] add_88748;
  wire [7:0] sel_88749;
  wire [7:0] add_88752;
  wire [7:0] sel_88753;
  wire [7:0] add_88756;
  wire [7:0] sel_88757;
  wire [7:0] add_88760;
  wire [7:0] sel_88761;
  wire [7:0] add_88764;
  wire [7:0] sel_88765;
  wire [7:0] add_88768;
  wire [7:0] sel_88769;
  wire [7:0] add_88772;
  wire [7:0] sel_88773;
  wire [7:0] add_88776;
  wire [7:0] sel_88777;
  wire [7:0] add_88780;
  wire [7:0] sel_88781;
  wire [7:0] add_88784;
  wire [7:0] sel_88785;
  wire [7:0] add_88788;
  wire [7:0] sel_88789;
  wire [7:0] add_88793;
  wire [15:0] array_index_88794;
  wire [7:0] sel_88795;
  wire [7:0] add_88798;
  wire [7:0] sel_88799;
  wire [7:0] add_88802;
  wire [7:0] sel_88803;
  wire [7:0] add_88806;
  wire [7:0] sel_88807;
  wire [7:0] add_88810;
  wire [7:0] sel_88811;
  wire [7:0] add_88814;
  wire [7:0] sel_88815;
  wire [7:0] add_88818;
  wire [7:0] sel_88819;
  wire [7:0] add_88822;
  wire [7:0] sel_88823;
  wire [7:0] add_88826;
  wire [7:0] sel_88827;
  wire [7:0] add_88830;
  wire [7:0] sel_88831;
  wire [7:0] add_88834;
  wire [7:0] sel_88835;
  wire [7:0] add_88838;
  wire [7:0] sel_88839;
  wire [7:0] add_88842;
  wire [7:0] sel_88843;
  wire [7:0] add_88846;
  wire [7:0] sel_88847;
  wire [7:0] add_88850;
  wire [7:0] sel_88851;
  wire [7:0] add_88854;
  wire [7:0] sel_88855;
  wire [7:0] add_88858;
  wire [7:0] sel_88859;
  wire [7:0] add_88862;
  wire [7:0] sel_88863;
  wire [7:0] add_88866;
  wire [7:0] sel_88867;
  wire [7:0] add_88870;
  wire [7:0] sel_88871;
  wire [7:0] add_88874;
  wire [7:0] sel_88875;
  wire [7:0] add_88878;
  wire [7:0] sel_88879;
  wire [7:0] add_88882;
  wire [7:0] sel_88883;
  wire [7:0] add_88886;
  wire [7:0] sel_88887;
  wire [7:0] add_88890;
  wire [7:0] sel_88891;
  wire [7:0] add_88894;
  wire [7:0] sel_88895;
  wire [7:0] add_88898;
  wire [7:0] sel_88899;
  wire [7:0] add_88902;
  wire [7:0] sel_88903;
  wire [7:0] add_88906;
  wire [7:0] sel_88907;
  wire [7:0] add_88910;
  wire [7:0] sel_88911;
  wire [7:0] add_88915;
  wire [15:0] array_index_88916;
  wire [7:0] sel_88917;
  wire [7:0] add_88920;
  wire [7:0] sel_88921;
  wire [7:0] add_88924;
  wire [7:0] sel_88925;
  wire [7:0] add_88928;
  wire [7:0] sel_88929;
  wire [7:0] add_88932;
  wire [7:0] sel_88933;
  wire [7:0] add_88936;
  wire [7:0] sel_88937;
  wire [7:0] add_88940;
  wire [7:0] sel_88941;
  wire [7:0] add_88944;
  wire [7:0] sel_88945;
  wire [7:0] add_88948;
  wire [7:0] sel_88949;
  wire [7:0] add_88952;
  wire [7:0] sel_88953;
  wire [7:0] add_88956;
  wire [7:0] sel_88957;
  wire [7:0] add_88960;
  wire [7:0] sel_88961;
  wire [7:0] add_88964;
  wire [7:0] sel_88965;
  wire [7:0] add_88968;
  wire [7:0] sel_88969;
  wire [7:0] add_88972;
  wire [7:0] sel_88973;
  wire [7:0] add_88976;
  wire [7:0] sel_88977;
  wire [7:0] add_88980;
  wire [7:0] sel_88981;
  wire [7:0] add_88984;
  wire [7:0] sel_88985;
  wire [7:0] add_88988;
  wire [7:0] sel_88989;
  wire [7:0] add_88992;
  wire [7:0] sel_88993;
  wire [7:0] add_88996;
  wire [7:0] sel_88997;
  wire [7:0] add_89000;
  wire [7:0] sel_89001;
  wire [7:0] add_89004;
  wire [7:0] sel_89005;
  wire [7:0] add_89008;
  wire [7:0] sel_89009;
  wire [7:0] add_89012;
  wire [7:0] sel_89013;
  wire [7:0] add_89016;
  wire [7:0] sel_89017;
  wire [7:0] add_89020;
  wire [7:0] sel_89021;
  wire [7:0] add_89024;
  wire [7:0] sel_89025;
  wire [7:0] add_89028;
  wire [7:0] sel_89029;
  wire [7:0] add_89032;
  wire [7:0] sel_89033;
  wire [7:0] add_89037;
  wire [15:0] array_index_89038;
  wire [7:0] sel_89039;
  wire [7:0] add_89042;
  wire [7:0] sel_89043;
  wire [7:0] add_89046;
  wire [7:0] sel_89047;
  wire [7:0] add_89050;
  wire [7:0] sel_89051;
  wire [7:0] add_89054;
  wire [7:0] sel_89055;
  wire [7:0] add_89058;
  wire [7:0] sel_89059;
  wire [7:0] add_89062;
  wire [7:0] sel_89063;
  wire [7:0] add_89066;
  wire [7:0] sel_89067;
  wire [7:0] add_89070;
  wire [7:0] sel_89071;
  wire [7:0] add_89074;
  wire [7:0] sel_89075;
  wire [7:0] add_89078;
  wire [7:0] sel_89079;
  wire [7:0] add_89082;
  wire [7:0] sel_89083;
  wire [7:0] add_89086;
  wire [7:0] sel_89087;
  wire [7:0] add_89090;
  wire [7:0] sel_89091;
  wire [7:0] add_89094;
  wire [7:0] sel_89095;
  wire [7:0] add_89098;
  wire [7:0] sel_89099;
  wire [7:0] add_89102;
  wire [7:0] sel_89103;
  wire [7:0] add_89106;
  wire [7:0] sel_89107;
  wire [7:0] add_89110;
  wire [7:0] sel_89111;
  wire [7:0] add_89114;
  wire [7:0] sel_89115;
  wire [7:0] add_89118;
  wire [7:0] sel_89119;
  wire [7:0] add_89122;
  wire [7:0] sel_89123;
  wire [7:0] add_89126;
  wire [7:0] sel_89127;
  wire [7:0] add_89130;
  wire [7:0] sel_89131;
  wire [7:0] add_89134;
  wire [7:0] sel_89135;
  wire [7:0] add_89138;
  wire [7:0] sel_89139;
  wire [7:0] add_89142;
  wire [7:0] sel_89143;
  wire [7:0] add_89146;
  wire [7:0] sel_89147;
  wire [7:0] add_89150;
  wire [7:0] sel_89151;
  wire [7:0] add_89154;
  wire [7:0] sel_89155;
  wire [7:0] add_89159;
  wire [15:0] array_index_89160;
  wire [7:0] sel_89161;
  wire [7:0] add_89164;
  wire [7:0] sel_89165;
  wire [7:0] add_89168;
  wire [7:0] sel_89169;
  wire [7:0] add_89172;
  wire [7:0] sel_89173;
  wire [7:0] add_89176;
  wire [7:0] sel_89177;
  wire [7:0] add_89180;
  wire [7:0] sel_89181;
  wire [7:0] add_89184;
  wire [7:0] sel_89185;
  wire [7:0] add_89188;
  wire [7:0] sel_89189;
  wire [7:0] add_89192;
  wire [7:0] sel_89193;
  wire [7:0] add_89196;
  wire [7:0] sel_89197;
  wire [7:0] add_89200;
  wire [7:0] sel_89201;
  wire [7:0] add_89204;
  wire [7:0] sel_89205;
  wire [7:0] add_89208;
  wire [7:0] sel_89209;
  wire [7:0] add_89212;
  wire [7:0] sel_89213;
  wire [7:0] add_89216;
  wire [7:0] sel_89217;
  wire [7:0] add_89220;
  wire [7:0] sel_89221;
  wire [7:0] add_89224;
  wire [7:0] sel_89225;
  wire [7:0] add_89228;
  wire [7:0] sel_89229;
  wire [7:0] add_89232;
  wire [7:0] sel_89233;
  wire [7:0] add_89236;
  wire [7:0] sel_89237;
  wire [7:0] add_89240;
  wire [7:0] sel_89241;
  wire [7:0] add_89244;
  wire [7:0] sel_89245;
  wire [7:0] add_89248;
  wire [7:0] sel_89249;
  wire [7:0] add_89252;
  wire [7:0] sel_89253;
  wire [7:0] add_89256;
  wire [7:0] sel_89257;
  wire [7:0] add_89260;
  wire [7:0] sel_89261;
  wire [7:0] add_89264;
  wire [7:0] sel_89265;
  wire [7:0] add_89268;
  wire [7:0] sel_89269;
  wire [7:0] add_89272;
  wire [7:0] sel_89273;
  wire [7:0] add_89276;
  wire [7:0] sel_89277;
  wire [7:0] add_89281;
  wire [15:0] array_index_89282;
  wire [7:0] sel_89283;
  wire [7:0] add_89286;
  wire [7:0] sel_89287;
  wire [7:0] add_89290;
  wire [7:0] sel_89291;
  wire [7:0] add_89294;
  wire [7:0] sel_89295;
  wire [7:0] add_89298;
  wire [7:0] sel_89299;
  wire [7:0] add_89302;
  wire [7:0] sel_89303;
  wire [7:0] add_89306;
  wire [7:0] sel_89307;
  wire [7:0] add_89310;
  wire [7:0] sel_89311;
  wire [7:0] add_89314;
  wire [7:0] sel_89315;
  wire [7:0] add_89318;
  wire [7:0] sel_89319;
  wire [7:0] add_89322;
  wire [7:0] sel_89323;
  wire [7:0] add_89326;
  wire [7:0] sel_89327;
  wire [7:0] add_89330;
  wire [7:0] sel_89331;
  wire [7:0] add_89334;
  wire [7:0] sel_89335;
  wire [7:0] add_89338;
  wire [7:0] sel_89339;
  wire [7:0] add_89342;
  wire [7:0] sel_89343;
  wire [7:0] add_89346;
  wire [7:0] sel_89347;
  wire [7:0] add_89350;
  wire [7:0] sel_89351;
  wire [7:0] add_89354;
  wire [7:0] sel_89355;
  wire [7:0] add_89358;
  wire [7:0] sel_89359;
  wire [7:0] add_89362;
  wire [7:0] sel_89363;
  wire [7:0] add_89366;
  wire [7:0] sel_89367;
  wire [7:0] add_89370;
  wire [7:0] sel_89371;
  wire [7:0] add_89374;
  wire [7:0] sel_89375;
  wire [7:0] add_89378;
  wire [7:0] sel_89379;
  wire [7:0] add_89382;
  wire [7:0] sel_89383;
  wire [7:0] add_89386;
  wire [7:0] sel_89387;
  wire [7:0] add_89390;
  wire [7:0] sel_89391;
  wire [7:0] add_89394;
  wire [7:0] sel_89395;
  wire [7:0] add_89398;
  wire [7:0] sel_89399;
  wire [7:0] add_89403;
  wire [15:0] array_index_89404;
  wire [7:0] sel_89405;
  wire [7:0] add_89408;
  wire [7:0] sel_89409;
  wire [7:0] add_89412;
  wire [7:0] sel_89413;
  wire [7:0] add_89416;
  wire [7:0] sel_89417;
  wire [7:0] add_89420;
  wire [7:0] sel_89421;
  wire [7:0] add_89424;
  wire [7:0] sel_89425;
  wire [7:0] add_89428;
  wire [7:0] sel_89429;
  wire [7:0] add_89432;
  wire [7:0] sel_89433;
  wire [7:0] add_89436;
  wire [7:0] sel_89437;
  wire [7:0] add_89440;
  wire [7:0] sel_89441;
  wire [7:0] add_89444;
  wire [7:0] sel_89445;
  wire [7:0] add_89448;
  wire [7:0] sel_89449;
  wire [7:0] add_89452;
  wire [7:0] sel_89453;
  wire [7:0] add_89456;
  wire [7:0] sel_89457;
  wire [7:0] add_89460;
  wire [7:0] sel_89461;
  wire [7:0] add_89464;
  wire [7:0] sel_89465;
  wire [7:0] add_89468;
  wire [7:0] sel_89469;
  wire [7:0] add_89472;
  wire [7:0] sel_89473;
  wire [7:0] add_89476;
  wire [7:0] sel_89477;
  wire [7:0] add_89480;
  wire [7:0] sel_89481;
  wire [7:0] add_89484;
  wire [7:0] sel_89485;
  wire [7:0] add_89488;
  wire [7:0] sel_89489;
  wire [7:0] add_89492;
  wire [7:0] sel_89493;
  wire [7:0] add_89496;
  wire [7:0] sel_89497;
  wire [7:0] add_89500;
  wire [7:0] sel_89501;
  wire [7:0] add_89504;
  wire [7:0] sel_89505;
  wire [7:0] add_89508;
  wire [7:0] sel_89509;
  wire [7:0] add_89512;
  wire [7:0] sel_89513;
  wire [7:0] add_89516;
  wire [7:0] sel_89517;
  wire [7:0] add_89520;
  wire [7:0] sel_89521;
  wire [7:0] add_89525;
  wire [15:0] array_index_89526;
  wire [7:0] sel_89527;
  wire [7:0] add_89530;
  wire [7:0] sel_89531;
  wire [7:0] add_89534;
  wire [7:0] sel_89535;
  wire [7:0] add_89538;
  wire [7:0] sel_89539;
  wire [7:0] add_89542;
  wire [7:0] sel_89543;
  wire [7:0] add_89546;
  wire [7:0] sel_89547;
  wire [7:0] add_89550;
  wire [7:0] sel_89551;
  wire [7:0] add_89554;
  wire [7:0] sel_89555;
  wire [7:0] add_89558;
  wire [7:0] sel_89559;
  wire [7:0] add_89562;
  wire [7:0] sel_89563;
  wire [7:0] add_89566;
  wire [7:0] sel_89567;
  wire [7:0] add_89570;
  wire [7:0] sel_89571;
  wire [7:0] add_89574;
  wire [7:0] sel_89575;
  wire [7:0] add_89578;
  wire [7:0] sel_89579;
  wire [7:0] add_89582;
  wire [7:0] sel_89583;
  wire [7:0] add_89586;
  wire [7:0] sel_89587;
  wire [7:0] add_89590;
  wire [7:0] sel_89591;
  wire [7:0] add_89594;
  wire [7:0] sel_89595;
  wire [7:0] add_89598;
  wire [7:0] sel_89599;
  wire [7:0] add_89602;
  wire [7:0] sel_89603;
  wire [7:0] add_89606;
  wire [7:0] sel_89607;
  wire [7:0] add_89610;
  wire [7:0] sel_89611;
  wire [7:0] add_89614;
  wire [7:0] sel_89615;
  wire [7:0] add_89618;
  wire [7:0] sel_89619;
  wire [7:0] add_89622;
  wire [7:0] sel_89623;
  wire [7:0] add_89626;
  wire [7:0] sel_89627;
  wire [7:0] add_89630;
  wire [7:0] sel_89631;
  wire [7:0] add_89634;
  wire [7:0] sel_89635;
  wire [7:0] add_89638;
  wire [7:0] sel_89639;
  wire [7:0] add_89642;
  wire [7:0] sel_89643;
  wire [7:0] add_89647;
  wire [15:0] array_index_89648;
  wire [7:0] sel_89649;
  wire [7:0] add_89652;
  wire [7:0] sel_89653;
  wire [7:0] add_89656;
  wire [7:0] sel_89657;
  wire [7:0] add_89660;
  wire [7:0] sel_89661;
  wire [7:0] add_89664;
  wire [7:0] sel_89665;
  wire [7:0] add_89668;
  wire [7:0] sel_89669;
  wire [7:0] add_89672;
  wire [7:0] sel_89673;
  wire [7:0] add_89676;
  wire [7:0] sel_89677;
  wire [7:0] add_89680;
  wire [7:0] sel_89681;
  wire [7:0] add_89684;
  wire [7:0] sel_89685;
  wire [7:0] add_89688;
  wire [7:0] sel_89689;
  wire [7:0] add_89692;
  wire [7:0] sel_89693;
  wire [7:0] add_89696;
  wire [7:0] sel_89697;
  wire [7:0] add_89700;
  wire [7:0] sel_89701;
  wire [7:0] add_89704;
  wire [7:0] sel_89705;
  wire [7:0] add_89708;
  wire [7:0] sel_89709;
  wire [7:0] add_89712;
  wire [7:0] sel_89713;
  wire [7:0] add_89716;
  wire [7:0] sel_89717;
  wire [7:0] add_89720;
  wire [7:0] sel_89721;
  wire [7:0] add_89724;
  wire [7:0] sel_89725;
  wire [7:0] add_89728;
  wire [7:0] sel_89729;
  wire [7:0] add_89732;
  wire [7:0] sel_89733;
  wire [7:0] add_89736;
  wire [7:0] sel_89737;
  wire [7:0] add_89740;
  wire [7:0] sel_89741;
  wire [7:0] add_89744;
  wire [7:0] sel_89745;
  wire [7:0] add_89748;
  wire [7:0] sel_89749;
  wire [7:0] add_89752;
  wire [7:0] sel_89753;
  wire [7:0] add_89756;
  wire [7:0] sel_89757;
  wire [7:0] add_89760;
  wire [7:0] sel_89761;
  wire [7:0] add_89764;
  wire [7:0] sel_89765;
  wire [7:0] add_89769;
  wire [15:0] array_index_89770;
  wire [7:0] sel_89771;
  wire [7:0] add_89774;
  wire [7:0] sel_89775;
  wire [7:0] add_89778;
  wire [7:0] sel_89779;
  wire [7:0] add_89782;
  wire [7:0] sel_89783;
  wire [7:0] add_89786;
  wire [7:0] sel_89787;
  wire [7:0] add_89790;
  wire [7:0] sel_89791;
  wire [7:0] add_89794;
  wire [7:0] sel_89795;
  wire [7:0] add_89798;
  wire [7:0] sel_89799;
  wire [7:0] add_89802;
  wire [7:0] sel_89803;
  wire [7:0] add_89806;
  wire [7:0] sel_89807;
  wire [7:0] add_89810;
  wire [7:0] sel_89811;
  wire [7:0] add_89814;
  wire [7:0] sel_89815;
  wire [7:0] add_89818;
  wire [7:0] sel_89819;
  wire [7:0] add_89822;
  wire [7:0] sel_89823;
  wire [7:0] add_89826;
  wire [7:0] sel_89827;
  wire [7:0] add_89830;
  wire [7:0] sel_89831;
  wire [7:0] add_89834;
  wire [7:0] sel_89835;
  wire [7:0] add_89838;
  wire [7:0] sel_89839;
  wire [7:0] add_89842;
  wire [7:0] sel_89843;
  wire [7:0] add_89846;
  wire [7:0] sel_89847;
  wire [7:0] add_89850;
  wire [7:0] sel_89851;
  wire [7:0] add_89854;
  wire [7:0] sel_89855;
  wire [7:0] add_89858;
  wire [7:0] sel_89859;
  wire [7:0] add_89862;
  wire [7:0] sel_89863;
  wire [7:0] add_89866;
  wire [7:0] sel_89867;
  wire [7:0] add_89870;
  wire [7:0] sel_89871;
  wire [7:0] add_89874;
  wire [7:0] sel_89875;
  wire [7:0] add_89878;
  wire [7:0] sel_89879;
  wire [7:0] add_89882;
  wire [7:0] sel_89883;
  wire [7:0] add_89886;
  wire [7:0] sel_89887;
  wire [7:0] add_89891;
  wire [15:0] array_index_89892;
  wire [7:0] sel_89893;
  wire [7:0] add_89896;
  wire [7:0] sel_89897;
  wire [7:0] add_89900;
  wire [7:0] sel_89901;
  wire [7:0] add_89904;
  wire [7:0] sel_89905;
  wire [7:0] add_89908;
  wire [7:0] sel_89909;
  wire [7:0] add_89912;
  wire [7:0] sel_89913;
  wire [7:0] add_89916;
  wire [7:0] sel_89917;
  wire [7:0] add_89920;
  wire [7:0] sel_89921;
  wire [7:0] add_89924;
  wire [7:0] sel_89925;
  wire [7:0] add_89928;
  wire [7:0] sel_89929;
  wire [7:0] add_89932;
  wire [7:0] sel_89933;
  wire [7:0] add_89936;
  wire [7:0] sel_89937;
  wire [7:0] add_89940;
  wire [7:0] sel_89941;
  wire [7:0] add_89944;
  wire [7:0] sel_89945;
  wire [7:0] add_89948;
  wire [7:0] sel_89949;
  wire [7:0] add_89952;
  wire [7:0] sel_89953;
  wire [7:0] add_89956;
  wire [7:0] sel_89957;
  wire [7:0] add_89960;
  wire [7:0] sel_89961;
  wire [7:0] add_89964;
  wire [7:0] sel_89965;
  wire [7:0] add_89968;
  wire [7:0] sel_89969;
  wire [7:0] add_89972;
  wire [7:0] sel_89973;
  wire [7:0] add_89976;
  wire [7:0] sel_89977;
  wire [7:0] add_89980;
  wire [7:0] sel_89981;
  wire [7:0] add_89984;
  wire [7:0] sel_89985;
  wire [7:0] add_89988;
  wire [7:0] sel_89989;
  wire [7:0] add_89992;
  wire [7:0] sel_89993;
  wire [7:0] add_89996;
  wire [7:0] sel_89997;
  wire [7:0] add_90000;
  wire [7:0] sel_90001;
  wire [7:0] add_90004;
  wire [7:0] sel_90005;
  wire [7:0] add_90008;
  wire [7:0] sel_90009;
  wire [7:0] add_90013;
  wire [15:0] array_index_90014;
  wire [7:0] sel_90015;
  wire [7:0] add_90018;
  wire [7:0] sel_90019;
  wire [7:0] add_90022;
  wire [7:0] sel_90023;
  wire [7:0] add_90026;
  wire [7:0] sel_90027;
  wire [7:0] add_90030;
  wire [7:0] sel_90031;
  wire [7:0] add_90034;
  wire [7:0] sel_90035;
  wire [7:0] add_90038;
  wire [7:0] sel_90039;
  wire [7:0] add_90042;
  wire [7:0] sel_90043;
  wire [7:0] add_90046;
  wire [7:0] sel_90047;
  wire [7:0] add_90050;
  wire [7:0] sel_90051;
  wire [7:0] add_90054;
  wire [7:0] sel_90055;
  wire [7:0] add_90058;
  wire [7:0] sel_90059;
  wire [7:0] add_90062;
  wire [7:0] sel_90063;
  wire [7:0] add_90066;
  wire [7:0] sel_90067;
  wire [7:0] add_90070;
  wire [7:0] sel_90071;
  wire [7:0] add_90074;
  wire [7:0] sel_90075;
  wire [7:0] add_90078;
  wire [7:0] sel_90079;
  wire [7:0] add_90082;
  wire [7:0] sel_90083;
  wire [7:0] add_90086;
  wire [7:0] sel_90087;
  wire [7:0] add_90090;
  wire [7:0] sel_90091;
  wire [7:0] add_90094;
  wire [7:0] sel_90095;
  wire [7:0] add_90098;
  wire [7:0] sel_90099;
  wire [7:0] add_90102;
  wire [7:0] sel_90103;
  wire [7:0] add_90106;
  wire [7:0] sel_90107;
  wire [7:0] add_90110;
  wire [7:0] sel_90111;
  wire [7:0] add_90114;
  wire [7:0] sel_90115;
  wire [7:0] add_90118;
  wire [7:0] sel_90119;
  wire [7:0] add_90122;
  wire [7:0] sel_90123;
  wire [7:0] add_90126;
  wire [7:0] sel_90127;
  wire [7:0] add_90130;
  wire [7:0] sel_90131;
  wire [7:0] add_90135;
  wire [15:0] array_index_90136;
  wire [7:0] sel_90137;
  wire [7:0] add_90140;
  wire [7:0] sel_90141;
  wire [7:0] add_90144;
  wire [7:0] sel_90145;
  wire [7:0] add_90148;
  wire [7:0] sel_90149;
  wire [7:0] add_90152;
  wire [7:0] sel_90153;
  wire [7:0] add_90156;
  wire [7:0] sel_90157;
  wire [7:0] add_90160;
  wire [7:0] sel_90161;
  wire [7:0] add_90164;
  wire [7:0] sel_90165;
  wire [7:0] add_90168;
  wire [7:0] sel_90169;
  wire [7:0] add_90172;
  wire [7:0] sel_90173;
  wire [7:0] add_90176;
  wire [7:0] sel_90177;
  wire [7:0] add_90180;
  wire [7:0] sel_90181;
  wire [7:0] add_90184;
  wire [7:0] sel_90185;
  wire [7:0] add_90188;
  wire [7:0] sel_90189;
  wire [7:0] add_90192;
  wire [7:0] sel_90193;
  wire [7:0] add_90196;
  wire [7:0] sel_90197;
  wire [7:0] add_90200;
  wire [7:0] sel_90201;
  wire [7:0] add_90204;
  wire [7:0] sel_90205;
  wire [7:0] add_90208;
  wire [7:0] sel_90209;
  wire [7:0] add_90212;
  wire [7:0] sel_90213;
  wire [7:0] add_90216;
  wire [7:0] sel_90217;
  wire [7:0] add_90220;
  wire [7:0] sel_90221;
  wire [7:0] add_90224;
  wire [7:0] sel_90225;
  wire [7:0] add_90228;
  wire [7:0] sel_90229;
  wire [7:0] add_90232;
  wire [7:0] sel_90233;
  wire [7:0] add_90236;
  wire [7:0] sel_90237;
  wire [7:0] add_90240;
  wire [7:0] sel_90241;
  wire [7:0] add_90244;
  wire [7:0] sel_90245;
  wire [7:0] add_90248;
  wire [7:0] sel_90249;
  wire [7:0] add_90252;
  wire [7:0] sel_90253;
  wire [7:0] add_90257;
  wire [15:0] array_index_90258;
  wire [7:0] sel_90259;
  wire [7:0] add_90262;
  wire [7:0] sel_90263;
  wire [7:0] add_90266;
  wire [7:0] sel_90267;
  wire [7:0] add_90270;
  wire [7:0] sel_90271;
  wire [7:0] add_90274;
  wire [7:0] sel_90275;
  wire [7:0] add_90278;
  wire [7:0] sel_90279;
  wire [7:0] add_90282;
  wire [7:0] sel_90283;
  wire [7:0] add_90286;
  wire [7:0] sel_90287;
  wire [7:0] add_90290;
  wire [7:0] sel_90291;
  wire [7:0] add_90294;
  wire [7:0] sel_90295;
  wire [7:0] add_90298;
  wire [7:0] sel_90299;
  wire [7:0] add_90302;
  wire [7:0] sel_90303;
  wire [7:0] add_90306;
  wire [7:0] sel_90307;
  wire [7:0] add_90310;
  wire [7:0] sel_90311;
  wire [7:0] add_90314;
  wire [7:0] sel_90315;
  wire [7:0] add_90318;
  wire [7:0] sel_90319;
  wire [7:0] add_90322;
  wire [7:0] sel_90323;
  wire [7:0] add_90326;
  wire [7:0] sel_90327;
  wire [7:0] add_90330;
  wire [7:0] sel_90331;
  wire [7:0] add_90334;
  wire [7:0] sel_90335;
  wire [7:0] add_90338;
  wire [7:0] sel_90339;
  wire [7:0] add_90342;
  wire [7:0] sel_90343;
  wire [7:0] add_90346;
  wire [7:0] sel_90347;
  wire [7:0] add_90350;
  wire [7:0] sel_90351;
  wire [7:0] add_90354;
  wire [7:0] sel_90355;
  wire [7:0] add_90358;
  wire [7:0] sel_90359;
  wire [7:0] add_90362;
  wire [7:0] sel_90363;
  wire [7:0] add_90366;
  wire [7:0] sel_90367;
  wire [7:0] add_90370;
  wire [7:0] sel_90371;
  wire [7:0] add_90374;
  wire [7:0] sel_90375;
  wire [7:0] add_90378;
  assign array_index_86651 = set1_unflattened[5'h00];
  assign array_index_86652 = set2_unflattened[5'h00];
  assign array_index_86656 = set2_unflattened[5'h01];
  assign concat_86657 = {1'h0, array_index_86651 == array_index_86652};
  assign add_86660 = concat_86657 + 2'h1;
  assign array_index_86664 = set2_unflattened[5'h02];
  assign concat_86665 = {1'h0, array_index_86651 == array_index_86656 ? add_86660 : concat_86657};
  assign add_86668 = concat_86665 + 3'h1;
  assign array_index_86672 = set2_unflattened[5'h03];
  assign concat_86673 = {1'h0, array_index_86651 == array_index_86664 ? add_86668 : concat_86665};
  assign add_86676 = concat_86673 + 4'h1;
  assign array_index_86680 = set2_unflattened[5'h04];
  assign concat_86681 = {1'h0, array_index_86651 == array_index_86672 ? add_86676 : concat_86673};
  assign add_86684 = concat_86681 + 5'h01;
  assign array_index_86688 = set2_unflattened[5'h05];
  assign concat_86689 = {1'h0, array_index_86651 == array_index_86680 ? add_86684 : concat_86681};
  assign add_86692 = concat_86689 + 6'h01;
  assign array_index_86696 = set2_unflattened[5'h06];
  assign concat_86697 = {1'h0, array_index_86651 == array_index_86688 ? add_86692 : concat_86689};
  assign add_86700 = concat_86697 + 7'h01;
  assign array_index_86704 = set2_unflattened[5'h07];
  assign concat_86705 = {1'h0, array_index_86651 == array_index_86696 ? add_86700 : concat_86697};
  assign add_86709 = concat_86705 + 8'h01;
  assign array_index_86710 = set2_unflattened[5'h08];
  assign sel_86711 = array_index_86651 == array_index_86704 ? add_86709 : concat_86705;
  assign add_86715 = sel_86711 + 8'h01;
  assign array_index_86716 = set2_unflattened[5'h09];
  assign sel_86717 = array_index_86651 == array_index_86710 ? add_86715 : sel_86711;
  assign add_86721 = sel_86717 + 8'h01;
  assign array_index_86722 = set2_unflattened[5'h0a];
  assign sel_86723 = array_index_86651 == array_index_86716 ? add_86721 : sel_86717;
  assign add_86727 = sel_86723 + 8'h01;
  assign array_index_86728 = set2_unflattened[5'h0b];
  assign sel_86729 = array_index_86651 == array_index_86722 ? add_86727 : sel_86723;
  assign add_86733 = sel_86729 + 8'h01;
  assign array_index_86734 = set2_unflattened[5'h0c];
  assign sel_86735 = array_index_86651 == array_index_86728 ? add_86733 : sel_86729;
  assign add_86739 = sel_86735 + 8'h01;
  assign array_index_86740 = set2_unflattened[5'h0d];
  assign sel_86741 = array_index_86651 == array_index_86734 ? add_86739 : sel_86735;
  assign add_86745 = sel_86741 + 8'h01;
  assign array_index_86746 = set2_unflattened[5'h0e];
  assign sel_86747 = array_index_86651 == array_index_86740 ? add_86745 : sel_86741;
  assign add_86751 = sel_86747 + 8'h01;
  assign array_index_86752 = set2_unflattened[5'h0f];
  assign sel_86753 = array_index_86651 == array_index_86746 ? add_86751 : sel_86747;
  assign add_86757 = sel_86753 + 8'h01;
  assign array_index_86758 = set2_unflattened[5'h10];
  assign sel_86759 = array_index_86651 == array_index_86752 ? add_86757 : sel_86753;
  assign add_86763 = sel_86759 + 8'h01;
  assign array_index_86764 = set2_unflattened[5'h11];
  assign sel_86765 = array_index_86651 == array_index_86758 ? add_86763 : sel_86759;
  assign add_86769 = sel_86765 + 8'h01;
  assign array_index_86770 = set2_unflattened[5'h12];
  assign sel_86771 = array_index_86651 == array_index_86764 ? add_86769 : sel_86765;
  assign add_86775 = sel_86771 + 8'h01;
  assign array_index_86776 = set2_unflattened[5'h13];
  assign sel_86777 = array_index_86651 == array_index_86770 ? add_86775 : sel_86771;
  assign add_86781 = sel_86777 + 8'h01;
  assign array_index_86782 = set2_unflattened[5'h14];
  assign sel_86783 = array_index_86651 == array_index_86776 ? add_86781 : sel_86777;
  assign add_86787 = sel_86783 + 8'h01;
  assign array_index_86788 = set2_unflattened[5'h15];
  assign sel_86789 = array_index_86651 == array_index_86782 ? add_86787 : sel_86783;
  assign add_86793 = sel_86789 + 8'h01;
  assign array_index_86794 = set2_unflattened[5'h16];
  assign sel_86795 = array_index_86651 == array_index_86788 ? add_86793 : sel_86789;
  assign add_86799 = sel_86795 + 8'h01;
  assign array_index_86800 = set2_unflattened[5'h17];
  assign sel_86801 = array_index_86651 == array_index_86794 ? add_86799 : sel_86795;
  assign add_86805 = sel_86801 + 8'h01;
  assign array_index_86806 = set2_unflattened[5'h18];
  assign sel_86807 = array_index_86651 == array_index_86800 ? add_86805 : sel_86801;
  assign add_86811 = sel_86807 + 8'h01;
  assign array_index_86812 = set2_unflattened[5'h19];
  assign sel_86813 = array_index_86651 == array_index_86806 ? add_86811 : sel_86807;
  assign add_86817 = sel_86813 + 8'h01;
  assign array_index_86818 = set2_unflattened[5'h1a];
  assign sel_86819 = array_index_86651 == array_index_86812 ? add_86817 : sel_86813;
  assign add_86823 = sel_86819 + 8'h01;
  assign array_index_86824 = set2_unflattened[5'h1b];
  assign sel_86825 = array_index_86651 == array_index_86818 ? add_86823 : sel_86819;
  assign add_86829 = sel_86825 + 8'h01;
  assign array_index_86830 = set2_unflattened[5'h1c];
  assign sel_86831 = array_index_86651 == array_index_86824 ? add_86829 : sel_86825;
  assign add_86835 = sel_86831 + 8'h01;
  assign array_index_86836 = set2_unflattened[5'h1d];
  assign sel_86837 = array_index_86651 == array_index_86830 ? add_86835 : sel_86831;
  assign add_86841 = sel_86837 + 8'h01;
  assign array_index_86842 = set1_unflattened[5'h01];
  assign sel_86843 = array_index_86651 == array_index_86836 ? add_86841 : sel_86837;
  assign add_86846 = sel_86843 + 8'h01;
  assign sel_86847 = array_index_86842 == array_index_86652 ? add_86846 : sel_86843;
  assign add_86850 = sel_86847 + 8'h01;
  assign sel_86851 = array_index_86842 == array_index_86656 ? add_86850 : sel_86847;
  assign add_86854 = sel_86851 + 8'h01;
  assign sel_86855 = array_index_86842 == array_index_86664 ? add_86854 : sel_86851;
  assign add_86858 = sel_86855 + 8'h01;
  assign sel_86859 = array_index_86842 == array_index_86672 ? add_86858 : sel_86855;
  assign add_86862 = sel_86859 + 8'h01;
  assign sel_86863 = array_index_86842 == array_index_86680 ? add_86862 : sel_86859;
  assign add_86866 = sel_86863 + 8'h01;
  assign sel_86867 = array_index_86842 == array_index_86688 ? add_86866 : sel_86863;
  assign add_86870 = sel_86867 + 8'h01;
  assign sel_86871 = array_index_86842 == array_index_86696 ? add_86870 : sel_86867;
  assign add_86874 = sel_86871 + 8'h01;
  assign sel_86875 = array_index_86842 == array_index_86704 ? add_86874 : sel_86871;
  assign add_86878 = sel_86875 + 8'h01;
  assign sel_86879 = array_index_86842 == array_index_86710 ? add_86878 : sel_86875;
  assign add_86882 = sel_86879 + 8'h01;
  assign sel_86883 = array_index_86842 == array_index_86716 ? add_86882 : sel_86879;
  assign add_86886 = sel_86883 + 8'h01;
  assign sel_86887 = array_index_86842 == array_index_86722 ? add_86886 : sel_86883;
  assign add_86890 = sel_86887 + 8'h01;
  assign sel_86891 = array_index_86842 == array_index_86728 ? add_86890 : sel_86887;
  assign add_86894 = sel_86891 + 8'h01;
  assign sel_86895 = array_index_86842 == array_index_86734 ? add_86894 : sel_86891;
  assign add_86898 = sel_86895 + 8'h01;
  assign sel_86899 = array_index_86842 == array_index_86740 ? add_86898 : sel_86895;
  assign add_86902 = sel_86899 + 8'h01;
  assign sel_86903 = array_index_86842 == array_index_86746 ? add_86902 : sel_86899;
  assign add_86906 = sel_86903 + 8'h01;
  assign sel_86907 = array_index_86842 == array_index_86752 ? add_86906 : sel_86903;
  assign add_86910 = sel_86907 + 8'h01;
  assign sel_86911 = array_index_86842 == array_index_86758 ? add_86910 : sel_86907;
  assign add_86914 = sel_86911 + 8'h01;
  assign sel_86915 = array_index_86842 == array_index_86764 ? add_86914 : sel_86911;
  assign add_86918 = sel_86915 + 8'h01;
  assign sel_86919 = array_index_86842 == array_index_86770 ? add_86918 : sel_86915;
  assign add_86922 = sel_86919 + 8'h01;
  assign sel_86923 = array_index_86842 == array_index_86776 ? add_86922 : sel_86919;
  assign add_86926 = sel_86923 + 8'h01;
  assign sel_86927 = array_index_86842 == array_index_86782 ? add_86926 : sel_86923;
  assign add_86930 = sel_86927 + 8'h01;
  assign sel_86931 = array_index_86842 == array_index_86788 ? add_86930 : sel_86927;
  assign add_86934 = sel_86931 + 8'h01;
  assign sel_86935 = array_index_86842 == array_index_86794 ? add_86934 : sel_86931;
  assign add_86938 = sel_86935 + 8'h01;
  assign sel_86939 = array_index_86842 == array_index_86800 ? add_86938 : sel_86935;
  assign add_86942 = sel_86939 + 8'h01;
  assign sel_86943 = array_index_86842 == array_index_86806 ? add_86942 : sel_86939;
  assign add_86946 = sel_86943 + 8'h01;
  assign sel_86947 = array_index_86842 == array_index_86812 ? add_86946 : sel_86943;
  assign add_86950 = sel_86947 + 8'h01;
  assign sel_86951 = array_index_86842 == array_index_86818 ? add_86950 : sel_86947;
  assign add_86954 = sel_86951 + 8'h01;
  assign sel_86955 = array_index_86842 == array_index_86824 ? add_86954 : sel_86951;
  assign add_86958 = sel_86955 + 8'h01;
  assign sel_86959 = array_index_86842 == array_index_86830 ? add_86958 : sel_86955;
  assign add_86963 = sel_86959 + 8'h01;
  assign array_index_86964 = set1_unflattened[5'h02];
  assign sel_86965 = array_index_86842 == array_index_86836 ? add_86963 : sel_86959;
  assign add_86968 = sel_86965 + 8'h01;
  assign sel_86969 = array_index_86964 == array_index_86652 ? add_86968 : sel_86965;
  assign add_86972 = sel_86969 + 8'h01;
  assign sel_86973 = array_index_86964 == array_index_86656 ? add_86972 : sel_86969;
  assign add_86976 = sel_86973 + 8'h01;
  assign sel_86977 = array_index_86964 == array_index_86664 ? add_86976 : sel_86973;
  assign add_86980 = sel_86977 + 8'h01;
  assign sel_86981 = array_index_86964 == array_index_86672 ? add_86980 : sel_86977;
  assign add_86984 = sel_86981 + 8'h01;
  assign sel_86985 = array_index_86964 == array_index_86680 ? add_86984 : sel_86981;
  assign add_86988 = sel_86985 + 8'h01;
  assign sel_86989 = array_index_86964 == array_index_86688 ? add_86988 : sel_86985;
  assign add_86992 = sel_86989 + 8'h01;
  assign sel_86993 = array_index_86964 == array_index_86696 ? add_86992 : sel_86989;
  assign add_86996 = sel_86993 + 8'h01;
  assign sel_86997 = array_index_86964 == array_index_86704 ? add_86996 : sel_86993;
  assign add_87000 = sel_86997 + 8'h01;
  assign sel_87001 = array_index_86964 == array_index_86710 ? add_87000 : sel_86997;
  assign add_87004 = sel_87001 + 8'h01;
  assign sel_87005 = array_index_86964 == array_index_86716 ? add_87004 : sel_87001;
  assign add_87008 = sel_87005 + 8'h01;
  assign sel_87009 = array_index_86964 == array_index_86722 ? add_87008 : sel_87005;
  assign add_87012 = sel_87009 + 8'h01;
  assign sel_87013 = array_index_86964 == array_index_86728 ? add_87012 : sel_87009;
  assign add_87016 = sel_87013 + 8'h01;
  assign sel_87017 = array_index_86964 == array_index_86734 ? add_87016 : sel_87013;
  assign add_87020 = sel_87017 + 8'h01;
  assign sel_87021 = array_index_86964 == array_index_86740 ? add_87020 : sel_87017;
  assign add_87024 = sel_87021 + 8'h01;
  assign sel_87025 = array_index_86964 == array_index_86746 ? add_87024 : sel_87021;
  assign add_87028 = sel_87025 + 8'h01;
  assign sel_87029 = array_index_86964 == array_index_86752 ? add_87028 : sel_87025;
  assign add_87032 = sel_87029 + 8'h01;
  assign sel_87033 = array_index_86964 == array_index_86758 ? add_87032 : sel_87029;
  assign add_87036 = sel_87033 + 8'h01;
  assign sel_87037 = array_index_86964 == array_index_86764 ? add_87036 : sel_87033;
  assign add_87040 = sel_87037 + 8'h01;
  assign sel_87041 = array_index_86964 == array_index_86770 ? add_87040 : sel_87037;
  assign add_87044 = sel_87041 + 8'h01;
  assign sel_87045 = array_index_86964 == array_index_86776 ? add_87044 : sel_87041;
  assign add_87048 = sel_87045 + 8'h01;
  assign sel_87049 = array_index_86964 == array_index_86782 ? add_87048 : sel_87045;
  assign add_87052 = sel_87049 + 8'h01;
  assign sel_87053 = array_index_86964 == array_index_86788 ? add_87052 : sel_87049;
  assign add_87056 = sel_87053 + 8'h01;
  assign sel_87057 = array_index_86964 == array_index_86794 ? add_87056 : sel_87053;
  assign add_87060 = sel_87057 + 8'h01;
  assign sel_87061 = array_index_86964 == array_index_86800 ? add_87060 : sel_87057;
  assign add_87064 = sel_87061 + 8'h01;
  assign sel_87065 = array_index_86964 == array_index_86806 ? add_87064 : sel_87061;
  assign add_87068 = sel_87065 + 8'h01;
  assign sel_87069 = array_index_86964 == array_index_86812 ? add_87068 : sel_87065;
  assign add_87072 = sel_87069 + 8'h01;
  assign sel_87073 = array_index_86964 == array_index_86818 ? add_87072 : sel_87069;
  assign add_87076 = sel_87073 + 8'h01;
  assign sel_87077 = array_index_86964 == array_index_86824 ? add_87076 : sel_87073;
  assign add_87080 = sel_87077 + 8'h01;
  assign sel_87081 = array_index_86964 == array_index_86830 ? add_87080 : sel_87077;
  assign add_87085 = sel_87081 + 8'h01;
  assign array_index_87086 = set1_unflattened[5'h03];
  assign sel_87087 = array_index_86964 == array_index_86836 ? add_87085 : sel_87081;
  assign add_87090 = sel_87087 + 8'h01;
  assign sel_87091 = array_index_87086 == array_index_86652 ? add_87090 : sel_87087;
  assign add_87094 = sel_87091 + 8'h01;
  assign sel_87095 = array_index_87086 == array_index_86656 ? add_87094 : sel_87091;
  assign add_87098 = sel_87095 + 8'h01;
  assign sel_87099 = array_index_87086 == array_index_86664 ? add_87098 : sel_87095;
  assign add_87102 = sel_87099 + 8'h01;
  assign sel_87103 = array_index_87086 == array_index_86672 ? add_87102 : sel_87099;
  assign add_87106 = sel_87103 + 8'h01;
  assign sel_87107 = array_index_87086 == array_index_86680 ? add_87106 : sel_87103;
  assign add_87110 = sel_87107 + 8'h01;
  assign sel_87111 = array_index_87086 == array_index_86688 ? add_87110 : sel_87107;
  assign add_87114 = sel_87111 + 8'h01;
  assign sel_87115 = array_index_87086 == array_index_86696 ? add_87114 : sel_87111;
  assign add_87118 = sel_87115 + 8'h01;
  assign sel_87119 = array_index_87086 == array_index_86704 ? add_87118 : sel_87115;
  assign add_87122 = sel_87119 + 8'h01;
  assign sel_87123 = array_index_87086 == array_index_86710 ? add_87122 : sel_87119;
  assign add_87126 = sel_87123 + 8'h01;
  assign sel_87127 = array_index_87086 == array_index_86716 ? add_87126 : sel_87123;
  assign add_87130 = sel_87127 + 8'h01;
  assign sel_87131 = array_index_87086 == array_index_86722 ? add_87130 : sel_87127;
  assign add_87134 = sel_87131 + 8'h01;
  assign sel_87135 = array_index_87086 == array_index_86728 ? add_87134 : sel_87131;
  assign add_87138 = sel_87135 + 8'h01;
  assign sel_87139 = array_index_87086 == array_index_86734 ? add_87138 : sel_87135;
  assign add_87142 = sel_87139 + 8'h01;
  assign sel_87143 = array_index_87086 == array_index_86740 ? add_87142 : sel_87139;
  assign add_87146 = sel_87143 + 8'h01;
  assign sel_87147 = array_index_87086 == array_index_86746 ? add_87146 : sel_87143;
  assign add_87150 = sel_87147 + 8'h01;
  assign sel_87151 = array_index_87086 == array_index_86752 ? add_87150 : sel_87147;
  assign add_87154 = sel_87151 + 8'h01;
  assign sel_87155 = array_index_87086 == array_index_86758 ? add_87154 : sel_87151;
  assign add_87158 = sel_87155 + 8'h01;
  assign sel_87159 = array_index_87086 == array_index_86764 ? add_87158 : sel_87155;
  assign add_87162 = sel_87159 + 8'h01;
  assign sel_87163 = array_index_87086 == array_index_86770 ? add_87162 : sel_87159;
  assign add_87166 = sel_87163 + 8'h01;
  assign sel_87167 = array_index_87086 == array_index_86776 ? add_87166 : sel_87163;
  assign add_87170 = sel_87167 + 8'h01;
  assign sel_87171 = array_index_87086 == array_index_86782 ? add_87170 : sel_87167;
  assign add_87174 = sel_87171 + 8'h01;
  assign sel_87175 = array_index_87086 == array_index_86788 ? add_87174 : sel_87171;
  assign add_87178 = sel_87175 + 8'h01;
  assign sel_87179 = array_index_87086 == array_index_86794 ? add_87178 : sel_87175;
  assign add_87182 = sel_87179 + 8'h01;
  assign sel_87183 = array_index_87086 == array_index_86800 ? add_87182 : sel_87179;
  assign add_87186 = sel_87183 + 8'h01;
  assign sel_87187 = array_index_87086 == array_index_86806 ? add_87186 : sel_87183;
  assign add_87190 = sel_87187 + 8'h01;
  assign sel_87191 = array_index_87086 == array_index_86812 ? add_87190 : sel_87187;
  assign add_87194 = sel_87191 + 8'h01;
  assign sel_87195 = array_index_87086 == array_index_86818 ? add_87194 : sel_87191;
  assign add_87198 = sel_87195 + 8'h01;
  assign sel_87199 = array_index_87086 == array_index_86824 ? add_87198 : sel_87195;
  assign add_87202 = sel_87199 + 8'h01;
  assign sel_87203 = array_index_87086 == array_index_86830 ? add_87202 : sel_87199;
  assign add_87207 = sel_87203 + 8'h01;
  assign array_index_87208 = set1_unflattened[5'h04];
  assign sel_87209 = array_index_87086 == array_index_86836 ? add_87207 : sel_87203;
  assign add_87212 = sel_87209 + 8'h01;
  assign sel_87213 = array_index_87208 == array_index_86652 ? add_87212 : sel_87209;
  assign add_87216 = sel_87213 + 8'h01;
  assign sel_87217 = array_index_87208 == array_index_86656 ? add_87216 : sel_87213;
  assign add_87220 = sel_87217 + 8'h01;
  assign sel_87221 = array_index_87208 == array_index_86664 ? add_87220 : sel_87217;
  assign add_87224 = sel_87221 + 8'h01;
  assign sel_87225 = array_index_87208 == array_index_86672 ? add_87224 : sel_87221;
  assign add_87228 = sel_87225 + 8'h01;
  assign sel_87229 = array_index_87208 == array_index_86680 ? add_87228 : sel_87225;
  assign add_87232 = sel_87229 + 8'h01;
  assign sel_87233 = array_index_87208 == array_index_86688 ? add_87232 : sel_87229;
  assign add_87236 = sel_87233 + 8'h01;
  assign sel_87237 = array_index_87208 == array_index_86696 ? add_87236 : sel_87233;
  assign add_87240 = sel_87237 + 8'h01;
  assign sel_87241 = array_index_87208 == array_index_86704 ? add_87240 : sel_87237;
  assign add_87244 = sel_87241 + 8'h01;
  assign sel_87245 = array_index_87208 == array_index_86710 ? add_87244 : sel_87241;
  assign add_87248 = sel_87245 + 8'h01;
  assign sel_87249 = array_index_87208 == array_index_86716 ? add_87248 : sel_87245;
  assign add_87252 = sel_87249 + 8'h01;
  assign sel_87253 = array_index_87208 == array_index_86722 ? add_87252 : sel_87249;
  assign add_87256 = sel_87253 + 8'h01;
  assign sel_87257 = array_index_87208 == array_index_86728 ? add_87256 : sel_87253;
  assign add_87260 = sel_87257 + 8'h01;
  assign sel_87261 = array_index_87208 == array_index_86734 ? add_87260 : sel_87257;
  assign add_87264 = sel_87261 + 8'h01;
  assign sel_87265 = array_index_87208 == array_index_86740 ? add_87264 : sel_87261;
  assign add_87268 = sel_87265 + 8'h01;
  assign sel_87269 = array_index_87208 == array_index_86746 ? add_87268 : sel_87265;
  assign add_87272 = sel_87269 + 8'h01;
  assign sel_87273 = array_index_87208 == array_index_86752 ? add_87272 : sel_87269;
  assign add_87276 = sel_87273 + 8'h01;
  assign sel_87277 = array_index_87208 == array_index_86758 ? add_87276 : sel_87273;
  assign add_87280 = sel_87277 + 8'h01;
  assign sel_87281 = array_index_87208 == array_index_86764 ? add_87280 : sel_87277;
  assign add_87284 = sel_87281 + 8'h01;
  assign sel_87285 = array_index_87208 == array_index_86770 ? add_87284 : sel_87281;
  assign add_87288 = sel_87285 + 8'h01;
  assign sel_87289 = array_index_87208 == array_index_86776 ? add_87288 : sel_87285;
  assign add_87292 = sel_87289 + 8'h01;
  assign sel_87293 = array_index_87208 == array_index_86782 ? add_87292 : sel_87289;
  assign add_87296 = sel_87293 + 8'h01;
  assign sel_87297 = array_index_87208 == array_index_86788 ? add_87296 : sel_87293;
  assign add_87300 = sel_87297 + 8'h01;
  assign sel_87301 = array_index_87208 == array_index_86794 ? add_87300 : sel_87297;
  assign add_87304 = sel_87301 + 8'h01;
  assign sel_87305 = array_index_87208 == array_index_86800 ? add_87304 : sel_87301;
  assign add_87308 = sel_87305 + 8'h01;
  assign sel_87309 = array_index_87208 == array_index_86806 ? add_87308 : sel_87305;
  assign add_87312 = sel_87309 + 8'h01;
  assign sel_87313 = array_index_87208 == array_index_86812 ? add_87312 : sel_87309;
  assign add_87316 = sel_87313 + 8'h01;
  assign sel_87317 = array_index_87208 == array_index_86818 ? add_87316 : sel_87313;
  assign add_87320 = sel_87317 + 8'h01;
  assign sel_87321 = array_index_87208 == array_index_86824 ? add_87320 : sel_87317;
  assign add_87324 = sel_87321 + 8'h01;
  assign sel_87325 = array_index_87208 == array_index_86830 ? add_87324 : sel_87321;
  assign add_87329 = sel_87325 + 8'h01;
  assign array_index_87330 = set1_unflattened[5'h05];
  assign sel_87331 = array_index_87208 == array_index_86836 ? add_87329 : sel_87325;
  assign add_87334 = sel_87331 + 8'h01;
  assign sel_87335 = array_index_87330 == array_index_86652 ? add_87334 : sel_87331;
  assign add_87338 = sel_87335 + 8'h01;
  assign sel_87339 = array_index_87330 == array_index_86656 ? add_87338 : sel_87335;
  assign add_87342 = sel_87339 + 8'h01;
  assign sel_87343 = array_index_87330 == array_index_86664 ? add_87342 : sel_87339;
  assign add_87346 = sel_87343 + 8'h01;
  assign sel_87347 = array_index_87330 == array_index_86672 ? add_87346 : sel_87343;
  assign add_87350 = sel_87347 + 8'h01;
  assign sel_87351 = array_index_87330 == array_index_86680 ? add_87350 : sel_87347;
  assign add_87354 = sel_87351 + 8'h01;
  assign sel_87355 = array_index_87330 == array_index_86688 ? add_87354 : sel_87351;
  assign add_87358 = sel_87355 + 8'h01;
  assign sel_87359 = array_index_87330 == array_index_86696 ? add_87358 : sel_87355;
  assign add_87362 = sel_87359 + 8'h01;
  assign sel_87363 = array_index_87330 == array_index_86704 ? add_87362 : sel_87359;
  assign add_87366 = sel_87363 + 8'h01;
  assign sel_87367 = array_index_87330 == array_index_86710 ? add_87366 : sel_87363;
  assign add_87370 = sel_87367 + 8'h01;
  assign sel_87371 = array_index_87330 == array_index_86716 ? add_87370 : sel_87367;
  assign add_87374 = sel_87371 + 8'h01;
  assign sel_87375 = array_index_87330 == array_index_86722 ? add_87374 : sel_87371;
  assign add_87378 = sel_87375 + 8'h01;
  assign sel_87379 = array_index_87330 == array_index_86728 ? add_87378 : sel_87375;
  assign add_87382 = sel_87379 + 8'h01;
  assign sel_87383 = array_index_87330 == array_index_86734 ? add_87382 : sel_87379;
  assign add_87386 = sel_87383 + 8'h01;
  assign sel_87387 = array_index_87330 == array_index_86740 ? add_87386 : sel_87383;
  assign add_87390 = sel_87387 + 8'h01;
  assign sel_87391 = array_index_87330 == array_index_86746 ? add_87390 : sel_87387;
  assign add_87394 = sel_87391 + 8'h01;
  assign sel_87395 = array_index_87330 == array_index_86752 ? add_87394 : sel_87391;
  assign add_87398 = sel_87395 + 8'h01;
  assign sel_87399 = array_index_87330 == array_index_86758 ? add_87398 : sel_87395;
  assign add_87402 = sel_87399 + 8'h01;
  assign sel_87403 = array_index_87330 == array_index_86764 ? add_87402 : sel_87399;
  assign add_87406 = sel_87403 + 8'h01;
  assign sel_87407 = array_index_87330 == array_index_86770 ? add_87406 : sel_87403;
  assign add_87410 = sel_87407 + 8'h01;
  assign sel_87411 = array_index_87330 == array_index_86776 ? add_87410 : sel_87407;
  assign add_87414 = sel_87411 + 8'h01;
  assign sel_87415 = array_index_87330 == array_index_86782 ? add_87414 : sel_87411;
  assign add_87418 = sel_87415 + 8'h01;
  assign sel_87419 = array_index_87330 == array_index_86788 ? add_87418 : sel_87415;
  assign add_87422 = sel_87419 + 8'h01;
  assign sel_87423 = array_index_87330 == array_index_86794 ? add_87422 : sel_87419;
  assign add_87426 = sel_87423 + 8'h01;
  assign sel_87427 = array_index_87330 == array_index_86800 ? add_87426 : sel_87423;
  assign add_87430 = sel_87427 + 8'h01;
  assign sel_87431 = array_index_87330 == array_index_86806 ? add_87430 : sel_87427;
  assign add_87434 = sel_87431 + 8'h01;
  assign sel_87435 = array_index_87330 == array_index_86812 ? add_87434 : sel_87431;
  assign add_87438 = sel_87435 + 8'h01;
  assign sel_87439 = array_index_87330 == array_index_86818 ? add_87438 : sel_87435;
  assign add_87442 = sel_87439 + 8'h01;
  assign sel_87443 = array_index_87330 == array_index_86824 ? add_87442 : sel_87439;
  assign add_87446 = sel_87443 + 8'h01;
  assign sel_87447 = array_index_87330 == array_index_86830 ? add_87446 : sel_87443;
  assign add_87451 = sel_87447 + 8'h01;
  assign array_index_87452 = set1_unflattened[5'h06];
  assign sel_87453 = array_index_87330 == array_index_86836 ? add_87451 : sel_87447;
  assign add_87456 = sel_87453 + 8'h01;
  assign sel_87457 = array_index_87452 == array_index_86652 ? add_87456 : sel_87453;
  assign add_87460 = sel_87457 + 8'h01;
  assign sel_87461 = array_index_87452 == array_index_86656 ? add_87460 : sel_87457;
  assign add_87464 = sel_87461 + 8'h01;
  assign sel_87465 = array_index_87452 == array_index_86664 ? add_87464 : sel_87461;
  assign add_87468 = sel_87465 + 8'h01;
  assign sel_87469 = array_index_87452 == array_index_86672 ? add_87468 : sel_87465;
  assign add_87472 = sel_87469 + 8'h01;
  assign sel_87473 = array_index_87452 == array_index_86680 ? add_87472 : sel_87469;
  assign add_87476 = sel_87473 + 8'h01;
  assign sel_87477 = array_index_87452 == array_index_86688 ? add_87476 : sel_87473;
  assign add_87480 = sel_87477 + 8'h01;
  assign sel_87481 = array_index_87452 == array_index_86696 ? add_87480 : sel_87477;
  assign add_87484 = sel_87481 + 8'h01;
  assign sel_87485 = array_index_87452 == array_index_86704 ? add_87484 : sel_87481;
  assign add_87488 = sel_87485 + 8'h01;
  assign sel_87489 = array_index_87452 == array_index_86710 ? add_87488 : sel_87485;
  assign add_87492 = sel_87489 + 8'h01;
  assign sel_87493 = array_index_87452 == array_index_86716 ? add_87492 : sel_87489;
  assign add_87496 = sel_87493 + 8'h01;
  assign sel_87497 = array_index_87452 == array_index_86722 ? add_87496 : sel_87493;
  assign add_87500 = sel_87497 + 8'h01;
  assign sel_87501 = array_index_87452 == array_index_86728 ? add_87500 : sel_87497;
  assign add_87504 = sel_87501 + 8'h01;
  assign sel_87505 = array_index_87452 == array_index_86734 ? add_87504 : sel_87501;
  assign add_87508 = sel_87505 + 8'h01;
  assign sel_87509 = array_index_87452 == array_index_86740 ? add_87508 : sel_87505;
  assign add_87512 = sel_87509 + 8'h01;
  assign sel_87513 = array_index_87452 == array_index_86746 ? add_87512 : sel_87509;
  assign add_87516 = sel_87513 + 8'h01;
  assign sel_87517 = array_index_87452 == array_index_86752 ? add_87516 : sel_87513;
  assign add_87520 = sel_87517 + 8'h01;
  assign sel_87521 = array_index_87452 == array_index_86758 ? add_87520 : sel_87517;
  assign add_87524 = sel_87521 + 8'h01;
  assign sel_87525 = array_index_87452 == array_index_86764 ? add_87524 : sel_87521;
  assign add_87528 = sel_87525 + 8'h01;
  assign sel_87529 = array_index_87452 == array_index_86770 ? add_87528 : sel_87525;
  assign add_87532 = sel_87529 + 8'h01;
  assign sel_87533 = array_index_87452 == array_index_86776 ? add_87532 : sel_87529;
  assign add_87536 = sel_87533 + 8'h01;
  assign sel_87537 = array_index_87452 == array_index_86782 ? add_87536 : sel_87533;
  assign add_87540 = sel_87537 + 8'h01;
  assign sel_87541 = array_index_87452 == array_index_86788 ? add_87540 : sel_87537;
  assign add_87544 = sel_87541 + 8'h01;
  assign sel_87545 = array_index_87452 == array_index_86794 ? add_87544 : sel_87541;
  assign add_87548 = sel_87545 + 8'h01;
  assign sel_87549 = array_index_87452 == array_index_86800 ? add_87548 : sel_87545;
  assign add_87552 = sel_87549 + 8'h01;
  assign sel_87553 = array_index_87452 == array_index_86806 ? add_87552 : sel_87549;
  assign add_87556 = sel_87553 + 8'h01;
  assign sel_87557 = array_index_87452 == array_index_86812 ? add_87556 : sel_87553;
  assign add_87560 = sel_87557 + 8'h01;
  assign sel_87561 = array_index_87452 == array_index_86818 ? add_87560 : sel_87557;
  assign add_87564 = sel_87561 + 8'h01;
  assign sel_87565 = array_index_87452 == array_index_86824 ? add_87564 : sel_87561;
  assign add_87568 = sel_87565 + 8'h01;
  assign sel_87569 = array_index_87452 == array_index_86830 ? add_87568 : sel_87565;
  assign add_87573 = sel_87569 + 8'h01;
  assign array_index_87574 = set1_unflattened[5'h07];
  assign sel_87575 = array_index_87452 == array_index_86836 ? add_87573 : sel_87569;
  assign add_87578 = sel_87575 + 8'h01;
  assign sel_87579 = array_index_87574 == array_index_86652 ? add_87578 : sel_87575;
  assign add_87582 = sel_87579 + 8'h01;
  assign sel_87583 = array_index_87574 == array_index_86656 ? add_87582 : sel_87579;
  assign add_87586 = sel_87583 + 8'h01;
  assign sel_87587 = array_index_87574 == array_index_86664 ? add_87586 : sel_87583;
  assign add_87590 = sel_87587 + 8'h01;
  assign sel_87591 = array_index_87574 == array_index_86672 ? add_87590 : sel_87587;
  assign add_87594 = sel_87591 + 8'h01;
  assign sel_87595 = array_index_87574 == array_index_86680 ? add_87594 : sel_87591;
  assign add_87598 = sel_87595 + 8'h01;
  assign sel_87599 = array_index_87574 == array_index_86688 ? add_87598 : sel_87595;
  assign add_87602 = sel_87599 + 8'h01;
  assign sel_87603 = array_index_87574 == array_index_86696 ? add_87602 : sel_87599;
  assign add_87606 = sel_87603 + 8'h01;
  assign sel_87607 = array_index_87574 == array_index_86704 ? add_87606 : sel_87603;
  assign add_87610 = sel_87607 + 8'h01;
  assign sel_87611 = array_index_87574 == array_index_86710 ? add_87610 : sel_87607;
  assign add_87614 = sel_87611 + 8'h01;
  assign sel_87615 = array_index_87574 == array_index_86716 ? add_87614 : sel_87611;
  assign add_87618 = sel_87615 + 8'h01;
  assign sel_87619 = array_index_87574 == array_index_86722 ? add_87618 : sel_87615;
  assign add_87622 = sel_87619 + 8'h01;
  assign sel_87623 = array_index_87574 == array_index_86728 ? add_87622 : sel_87619;
  assign add_87626 = sel_87623 + 8'h01;
  assign sel_87627 = array_index_87574 == array_index_86734 ? add_87626 : sel_87623;
  assign add_87630 = sel_87627 + 8'h01;
  assign sel_87631 = array_index_87574 == array_index_86740 ? add_87630 : sel_87627;
  assign add_87634 = sel_87631 + 8'h01;
  assign sel_87635 = array_index_87574 == array_index_86746 ? add_87634 : sel_87631;
  assign add_87638 = sel_87635 + 8'h01;
  assign sel_87639 = array_index_87574 == array_index_86752 ? add_87638 : sel_87635;
  assign add_87642 = sel_87639 + 8'h01;
  assign sel_87643 = array_index_87574 == array_index_86758 ? add_87642 : sel_87639;
  assign add_87646 = sel_87643 + 8'h01;
  assign sel_87647 = array_index_87574 == array_index_86764 ? add_87646 : sel_87643;
  assign add_87650 = sel_87647 + 8'h01;
  assign sel_87651 = array_index_87574 == array_index_86770 ? add_87650 : sel_87647;
  assign add_87654 = sel_87651 + 8'h01;
  assign sel_87655 = array_index_87574 == array_index_86776 ? add_87654 : sel_87651;
  assign add_87658 = sel_87655 + 8'h01;
  assign sel_87659 = array_index_87574 == array_index_86782 ? add_87658 : sel_87655;
  assign add_87662 = sel_87659 + 8'h01;
  assign sel_87663 = array_index_87574 == array_index_86788 ? add_87662 : sel_87659;
  assign add_87666 = sel_87663 + 8'h01;
  assign sel_87667 = array_index_87574 == array_index_86794 ? add_87666 : sel_87663;
  assign add_87670 = sel_87667 + 8'h01;
  assign sel_87671 = array_index_87574 == array_index_86800 ? add_87670 : sel_87667;
  assign add_87674 = sel_87671 + 8'h01;
  assign sel_87675 = array_index_87574 == array_index_86806 ? add_87674 : sel_87671;
  assign add_87678 = sel_87675 + 8'h01;
  assign sel_87679 = array_index_87574 == array_index_86812 ? add_87678 : sel_87675;
  assign add_87682 = sel_87679 + 8'h01;
  assign sel_87683 = array_index_87574 == array_index_86818 ? add_87682 : sel_87679;
  assign add_87686 = sel_87683 + 8'h01;
  assign sel_87687 = array_index_87574 == array_index_86824 ? add_87686 : sel_87683;
  assign add_87690 = sel_87687 + 8'h01;
  assign sel_87691 = array_index_87574 == array_index_86830 ? add_87690 : sel_87687;
  assign add_87695 = sel_87691 + 8'h01;
  assign array_index_87696 = set1_unflattened[5'h08];
  assign sel_87697 = array_index_87574 == array_index_86836 ? add_87695 : sel_87691;
  assign add_87700 = sel_87697 + 8'h01;
  assign sel_87701 = array_index_87696 == array_index_86652 ? add_87700 : sel_87697;
  assign add_87704 = sel_87701 + 8'h01;
  assign sel_87705 = array_index_87696 == array_index_86656 ? add_87704 : sel_87701;
  assign add_87708 = sel_87705 + 8'h01;
  assign sel_87709 = array_index_87696 == array_index_86664 ? add_87708 : sel_87705;
  assign add_87712 = sel_87709 + 8'h01;
  assign sel_87713 = array_index_87696 == array_index_86672 ? add_87712 : sel_87709;
  assign add_87716 = sel_87713 + 8'h01;
  assign sel_87717 = array_index_87696 == array_index_86680 ? add_87716 : sel_87713;
  assign add_87720 = sel_87717 + 8'h01;
  assign sel_87721 = array_index_87696 == array_index_86688 ? add_87720 : sel_87717;
  assign add_87724 = sel_87721 + 8'h01;
  assign sel_87725 = array_index_87696 == array_index_86696 ? add_87724 : sel_87721;
  assign add_87728 = sel_87725 + 8'h01;
  assign sel_87729 = array_index_87696 == array_index_86704 ? add_87728 : sel_87725;
  assign add_87732 = sel_87729 + 8'h01;
  assign sel_87733 = array_index_87696 == array_index_86710 ? add_87732 : sel_87729;
  assign add_87736 = sel_87733 + 8'h01;
  assign sel_87737 = array_index_87696 == array_index_86716 ? add_87736 : sel_87733;
  assign add_87740 = sel_87737 + 8'h01;
  assign sel_87741 = array_index_87696 == array_index_86722 ? add_87740 : sel_87737;
  assign add_87744 = sel_87741 + 8'h01;
  assign sel_87745 = array_index_87696 == array_index_86728 ? add_87744 : sel_87741;
  assign add_87748 = sel_87745 + 8'h01;
  assign sel_87749 = array_index_87696 == array_index_86734 ? add_87748 : sel_87745;
  assign add_87752 = sel_87749 + 8'h01;
  assign sel_87753 = array_index_87696 == array_index_86740 ? add_87752 : sel_87749;
  assign add_87756 = sel_87753 + 8'h01;
  assign sel_87757 = array_index_87696 == array_index_86746 ? add_87756 : sel_87753;
  assign add_87760 = sel_87757 + 8'h01;
  assign sel_87761 = array_index_87696 == array_index_86752 ? add_87760 : sel_87757;
  assign add_87764 = sel_87761 + 8'h01;
  assign sel_87765 = array_index_87696 == array_index_86758 ? add_87764 : sel_87761;
  assign add_87768 = sel_87765 + 8'h01;
  assign sel_87769 = array_index_87696 == array_index_86764 ? add_87768 : sel_87765;
  assign add_87772 = sel_87769 + 8'h01;
  assign sel_87773 = array_index_87696 == array_index_86770 ? add_87772 : sel_87769;
  assign add_87776 = sel_87773 + 8'h01;
  assign sel_87777 = array_index_87696 == array_index_86776 ? add_87776 : sel_87773;
  assign add_87780 = sel_87777 + 8'h01;
  assign sel_87781 = array_index_87696 == array_index_86782 ? add_87780 : sel_87777;
  assign add_87784 = sel_87781 + 8'h01;
  assign sel_87785 = array_index_87696 == array_index_86788 ? add_87784 : sel_87781;
  assign add_87788 = sel_87785 + 8'h01;
  assign sel_87789 = array_index_87696 == array_index_86794 ? add_87788 : sel_87785;
  assign add_87792 = sel_87789 + 8'h01;
  assign sel_87793 = array_index_87696 == array_index_86800 ? add_87792 : sel_87789;
  assign add_87796 = sel_87793 + 8'h01;
  assign sel_87797 = array_index_87696 == array_index_86806 ? add_87796 : sel_87793;
  assign add_87800 = sel_87797 + 8'h01;
  assign sel_87801 = array_index_87696 == array_index_86812 ? add_87800 : sel_87797;
  assign add_87804 = sel_87801 + 8'h01;
  assign sel_87805 = array_index_87696 == array_index_86818 ? add_87804 : sel_87801;
  assign add_87808 = sel_87805 + 8'h01;
  assign sel_87809 = array_index_87696 == array_index_86824 ? add_87808 : sel_87805;
  assign add_87812 = sel_87809 + 8'h01;
  assign sel_87813 = array_index_87696 == array_index_86830 ? add_87812 : sel_87809;
  assign add_87817 = sel_87813 + 8'h01;
  assign array_index_87818 = set1_unflattened[5'h09];
  assign sel_87819 = array_index_87696 == array_index_86836 ? add_87817 : sel_87813;
  assign add_87822 = sel_87819 + 8'h01;
  assign sel_87823 = array_index_87818 == array_index_86652 ? add_87822 : sel_87819;
  assign add_87826 = sel_87823 + 8'h01;
  assign sel_87827 = array_index_87818 == array_index_86656 ? add_87826 : sel_87823;
  assign add_87830 = sel_87827 + 8'h01;
  assign sel_87831 = array_index_87818 == array_index_86664 ? add_87830 : sel_87827;
  assign add_87834 = sel_87831 + 8'h01;
  assign sel_87835 = array_index_87818 == array_index_86672 ? add_87834 : sel_87831;
  assign add_87838 = sel_87835 + 8'h01;
  assign sel_87839 = array_index_87818 == array_index_86680 ? add_87838 : sel_87835;
  assign add_87842 = sel_87839 + 8'h01;
  assign sel_87843 = array_index_87818 == array_index_86688 ? add_87842 : sel_87839;
  assign add_87846 = sel_87843 + 8'h01;
  assign sel_87847 = array_index_87818 == array_index_86696 ? add_87846 : sel_87843;
  assign add_87850 = sel_87847 + 8'h01;
  assign sel_87851 = array_index_87818 == array_index_86704 ? add_87850 : sel_87847;
  assign add_87854 = sel_87851 + 8'h01;
  assign sel_87855 = array_index_87818 == array_index_86710 ? add_87854 : sel_87851;
  assign add_87858 = sel_87855 + 8'h01;
  assign sel_87859 = array_index_87818 == array_index_86716 ? add_87858 : sel_87855;
  assign add_87862 = sel_87859 + 8'h01;
  assign sel_87863 = array_index_87818 == array_index_86722 ? add_87862 : sel_87859;
  assign add_87866 = sel_87863 + 8'h01;
  assign sel_87867 = array_index_87818 == array_index_86728 ? add_87866 : sel_87863;
  assign add_87870 = sel_87867 + 8'h01;
  assign sel_87871 = array_index_87818 == array_index_86734 ? add_87870 : sel_87867;
  assign add_87874 = sel_87871 + 8'h01;
  assign sel_87875 = array_index_87818 == array_index_86740 ? add_87874 : sel_87871;
  assign add_87878 = sel_87875 + 8'h01;
  assign sel_87879 = array_index_87818 == array_index_86746 ? add_87878 : sel_87875;
  assign add_87882 = sel_87879 + 8'h01;
  assign sel_87883 = array_index_87818 == array_index_86752 ? add_87882 : sel_87879;
  assign add_87886 = sel_87883 + 8'h01;
  assign sel_87887 = array_index_87818 == array_index_86758 ? add_87886 : sel_87883;
  assign add_87890 = sel_87887 + 8'h01;
  assign sel_87891 = array_index_87818 == array_index_86764 ? add_87890 : sel_87887;
  assign add_87894 = sel_87891 + 8'h01;
  assign sel_87895 = array_index_87818 == array_index_86770 ? add_87894 : sel_87891;
  assign add_87898 = sel_87895 + 8'h01;
  assign sel_87899 = array_index_87818 == array_index_86776 ? add_87898 : sel_87895;
  assign add_87902 = sel_87899 + 8'h01;
  assign sel_87903 = array_index_87818 == array_index_86782 ? add_87902 : sel_87899;
  assign add_87906 = sel_87903 + 8'h01;
  assign sel_87907 = array_index_87818 == array_index_86788 ? add_87906 : sel_87903;
  assign add_87910 = sel_87907 + 8'h01;
  assign sel_87911 = array_index_87818 == array_index_86794 ? add_87910 : sel_87907;
  assign add_87914 = sel_87911 + 8'h01;
  assign sel_87915 = array_index_87818 == array_index_86800 ? add_87914 : sel_87911;
  assign add_87918 = sel_87915 + 8'h01;
  assign sel_87919 = array_index_87818 == array_index_86806 ? add_87918 : sel_87915;
  assign add_87922 = sel_87919 + 8'h01;
  assign sel_87923 = array_index_87818 == array_index_86812 ? add_87922 : sel_87919;
  assign add_87926 = sel_87923 + 8'h01;
  assign sel_87927 = array_index_87818 == array_index_86818 ? add_87926 : sel_87923;
  assign add_87930 = sel_87927 + 8'h01;
  assign sel_87931 = array_index_87818 == array_index_86824 ? add_87930 : sel_87927;
  assign add_87934 = sel_87931 + 8'h01;
  assign sel_87935 = array_index_87818 == array_index_86830 ? add_87934 : sel_87931;
  assign add_87939 = sel_87935 + 8'h01;
  assign array_index_87940 = set1_unflattened[5'h0a];
  assign sel_87941 = array_index_87818 == array_index_86836 ? add_87939 : sel_87935;
  assign add_87944 = sel_87941 + 8'h01;
  assign sel_87945 = array_index_87940 == array_index_86652 ? add_87944 : sel_87941;
  assign add_87948 = sel_87945 + 8'h01;
  assign sel_87949 = array_index_87940 == array_index_86656 ? add_87948 : sel_87945;
  assign add_87952 = sel_87949 + 8'h01;
  assign sel_87953 = array_index_87940 == array_index_86664 ? add_87952 : sel_87949;
  assign add_87956 = sel_87953 + 8'h01;
  assign sel_87957 = array_index_87940 == array_index_86672 ? add_87956 : sel_87953;
  assign add_87960 = sel_87957 + 8'h01;
  assign sel_87961 = array_index_87940 == array_index_86680 ? add_87960 : sel_87957;
  assign add_87964 = sel_87961 + 8'h01;
  assign sel_87965 = array_index_87940 == array_index_86688 ? add_87964 : sel_87961;
  assign add_87968 = sel_87965 + 8'h01;
  assign sel_87969 = array_index_87940 == array_index_86696 ? add_87968 : sel_87965;
  assign add_87972 = sel_87969 + 8'h01;
  assign sel_87973 = array_index_87940 == array_index_86704 ? add_87972 : sel_87969;
  assign add_87976 = sel_87973 + 8'h01;
  assign sel_87977 = array_index_87940 == array_index_86710 ? add_87976 : sel_87973;
  assign add_87980 = sel_87977 + 8'h01;
  assign sel_87981 = array_index_87940 == array_index_86716 ? add_87980 : sel_87977;
  assign add_87984 = sel_87981 + 8'h01;
  assign sel_87985 = array_index_87940 == array_index_86722 ? add_87984 : sel_87981;
  assign add_87988 = sel_87985 + 8'h01;
  assign sel_87989 = array_index_87940 == array_index_86728 ? add_87988 : sel_87985;
  assign add_87992 = sel_87989 + 8'h01;
  assign sel_87993 = array_index_87940 == array_index_86734 ? add_87992 : sel_87989;
  assign add_87996 = sel_87993 + 8'h01;
  assign sel_87997 = array_index_87940 == array_index_86740 ? add_87996 : sel_87993;
  assign add_88000 = sel_87997 + 8'h01;
  assign sel_88001 = array_index_87940 == array_index_86746 ? add_88000 : sel_87997;
  assign add_88004 = sel_88001 + 8'h01;
  assign sel_88005 = array_index_87940 == array_index_86752 ? add_88004 : sel_88001;
  assign add_88008 = sel_88005 + 8'h01;
  assign sel_88009 = array_index_87940 == array_index_86758 ? add_88008 : sel_88005;
  assign add_88012 = sel_88009 + 8'h01;
  assign sel_88013 = array_index_87940 == array_index_86764 ? add_88012 : sel_88009;
  assign add_88016 = sel_88013 + 8'h01;
  assign sel_88017 = array_index_87940 == array_index_86770 ? add_88016 : sel_88013;
  assign add_88020 = sel_88017 + 8'h01;
  assign sel_88021 = array_index_87940 == array_index_86776 ? add_88020 : sel_88017;
  assign add_88024 = sel_88021 + 8'h01;
  assign sel_88025 = array_index_87940 == array_index_86782 ? add_88024 : sel_88021;
  assign add_88028 = sel_88025 + 8'h01;
  assign sel_88029 = array_index_87940 == array_index_86788 ? add_88028 : sel_88025;
  assign add_88032 = sel_88029 + 8'h01;
  assign sel_88033 = array_index_87940 == array_index_86794 ? add_88032 : sel_88029;
  assign add_88036 = sel_88033 + 8'h01;
  assign sel_88037 = array_index_87940 == array_index_86800 ? add_88036 : sel_88033;
  assign add_88040 = sel_88037 + 8'h01;
  assign sel_88041 = array_index_87940 == array_index_86806 ? add_88040 : sel_88037;
  assign add_88044 = sel_88041 + 8'h01;
  assign sel_88045 = array_index_87940 == array_index_86812 ? add_88044 : sel_88041;
  assign add_88048 = sel_88045 + 8'h01;
  assign sel_88049 = array_index_87940 == array_index_86818 ? add_88048 : sel_88045;
  assign add_88052 = sel_88049 + 8'h01;
  assign sel_88053 = array_index_87940 == array_index_86824 ? add_88052 : sel_88049;
  assign add_88056 = sel_88053 + 8'h01;
  assign sel_88057 = array_index_87940 == array_index_86830 ? add_88056 : sel_88053;
  assign add_88061 = sel_88057 + 8'h01;
  assign array_index_88062 = set1_unflattened[5'h0b];
  assign sel_88063 = array_index_87940 == array_index_86836 ? add_88061 : sel_88057;
  assign add_88066 = sel_88063 + 8'h01;
  assign sel_88067 = array_index_88062 == array_index_86652 ? add_88066 : sel_88063;
  assign add_88070 = sel_88067 + 8'h01;
  assign sel_88071 = array_index_88062 == array_index_86656 ? add_88070 : sel_88067;
  assign add_88074 = sel_88071 + 8'h01;
  assign sel_88075 = array_index_88062 == array_index_86664 ? add_88074 : sel_88071;
  assign add_88078 = sel_88075 + 8'h01;
  assign sel_88079 = array_index_88062 == array_index_86672 ? add_88078 : sel_88075;
  assign add_88082 = sel_88079 + 8'h01;
  assign sel_88083 = array_index_88062 == array_index_86680 ? add_88082 : sel_88079;
  assign add_88086 = sel_88083 + 8'h01;
  assign sel_88087 = array_index_88062 == array_index_86688 ? add_88086 : sel_88083;
  assign add_88090 = sel_88087 + 8'h01;
  assign sel_88091 = array_index_88062 == array_index_86696 ? add_88090 : sel_88087;
  assign add_88094 = sel_88091 + 8'h01;
  assign sel_88095 = array_index_88062 == array_index_86704 ? add_88094 : sel_88091;
  assign add_88098 = sel_88095 + 8'h01;
  assign sel_88099 = array_index_88062 == array_index_86710 ? add_88098 : sel_88095;
  assign add_88102 = sel_88099 + 8'h01;
  assign sel_88103 = array_index_88062 == array_index_86716 ? add_88102 : sel_88099;
  assign add_88106 = sel_88103 + 8'h01;
  assign sel_88107 = array_index_88062 == array_index_86722 ? add_88106 : sel_88103;
  assign add_88110 = sel_88107 + 8'h01;
  assign sel_88111 = array_index_88062 == array_index_86728 ? add_88110 : sel_88107;
  assign add_88114 = sel_88111 + 8'h01;
  assign sel_88115 = array_index_88062 == array_index_86734 ? add_88114 : sel_88111;
  assign add_88118 = sel_88115 + 8'h01;
  assign sel_88119 = array_index_88062 == array_index_86740 ? add_88118 : sel_88115;
  assign add_88122 = sel_88119 + 8'h01;
  assign sel_88123 = array_index_88062 == array_index_86746 ? add_88122 : sel_88119;
  assign add_88126 = sel_88123 + 8'h01;
  assign sel_88127 = array_index_88062 == array_index_86752 ? add_88126 : sel_88123;
  assign add_88130 = sel_88127 + 8'h01;
  assign sel_88131 = array_index_88062 == array_index_86758 ? add_88130 : sel_88127;
  assign add_88134 = sel_88131 + 8'h01;
  assign sel_88135 = array_index_88062 == array_index_86764 ? add_88134 : sel_88131;
  assign add_88138 = sel_88135 + 8'h01;
  assign sel_88139 = array_index_88062 == array_index_86770 ? add_88138 : sel_88135;
  assign add_88142 = sel_88139 + 8'h01;
  assign sel_88143 = array_index_88062 == array_index_86776 ? add_88142 : sel_88139;
  assign add_88146 = sel_88143 + 8'h01;
  assign sel_88147 = array_index_88062 == array_index_86782 ? add_88146 : sel_88143;
  assign add_88150 = sel_88147 + 8'h01;
  assign sel_88151 = array_index_88062 == array_index_86788 ? add_88150 : sel_88147;
  assign add_88154 = sel_88151 + 8'h01;
  assign sel_88155 = array_index_88062 == array_index_86794 ? add_88154 : sel_88151;
  assign add_88158 = sel_88155 + 8'h01;
  assign sel_88159 = array_index_88062 == array_index_86800 ? add_88158 : sel_88155;
  assign add_88162 = sel_88159 + 8'h01;
  assign sel_88163 = array_index_88062 == array_index_86806 ? add_88162 : sel_88159;
  assign add_88166 = sel_88163 + 8'h01;
  assign sel_88167 = array_index_88062 == array_index_86812 ? add_88166 : sel_88163;
  assign add_88170 = sel_88167 + 8'h01;
  assign sel_88171 = array_index_88062 == array_index_86818 ? add_88170 : sel_88167;
  assign add_88174 = sel_88171 + 8'h01;
  assign sel_88175 = array_index_88062 == array_index_86824 ? add_88174 : sel_88171;
  assign add_88178 = sel_88175 + 8'h01;
  assign sel_88179 = array_index_88062 == array_index_86830 ? add_88178 : sel_88175;
  assign add_88183 = sel_88179 + 8'h01;
  assign array_index_88184 = set1_unflattened[5'h0c];
  assign sel_88185 = array_index_88062 == array_index_86836 ? add_88183 : sel_88179;
  assign add_88188 = sel_88185 + 8'h01;
  assign sel_88189 = array_index_88184 == array_index_86652 ? add_88188 : sel_88185;
  assign add_88192 = sel_88189 + 8'h01;
  assign sel_88193 = array_index_88184 == array_index_86656 ? add_88192 : sel_88189;
  assign add_88196 = sel_88193 + 8'h01;
  assign sel_88197 = array_index_88184 == array_index_86664 ? add_88196 : sel_88193;
  assign add_88200 = sel_88197 + 8'h01;
  assign sel_88201 = array_index_88184 == array_index_86672 ? add_88200 : sel_88197;
  assign add_88204 = sel_88201 + 8'h01;
  assign sel_88205 = array_index_88184 == array_index_86680 ? add_88204 : sel_88201;
  assign add_88208 = sel_88205 + 8'h01;
  assign sel_88209 = array_index_88184 == array_index_86688 ? add_88208 : sel_88205;
  assign add_88212 = sel_88209 + 8'h01;
  assign sel_88213 = array_index_88184 == array_index_86696 ? add_88212 : sel_88209;
  assign add_88216 = sel_88213 + 8'h01;
  assign sel_88217 = array_index_88184 == array_index_86704 ? add_88216 : sel_88213;
  assign add_88220 = sel_88217 + 8'h01;
  assign sel_88221 = array_index_88184 == array_index_86710 ? add_88220 : sel_88217;
  assign add_88224 = sel_88221 + 8'h01;
  assign sel_88225 = array_index_88184 == array_index_86716 ? add_88224 : sel_88221;
  assign add_88228 = sel_88225 + 8'h01;
  assign sel_88229 = array_index_88184 == array_index_86722 ? add_88228 : sel_88225;
  assign add_88232 = sel_88229 + 8'h01;
  assign sel_88233 = array_index_88184 == array_index_86728 ? add_88232 : sel_88229;
  assign add_88236 = sel_88233 + 8'h01;
  assign sel_88237 = array_index_88184 == array_index_86734 ? add_88236 : sel_88233;
  assign add_88240 = sel_88237 + 8'h01;
  assign sel_88241 = array_index_88184 == array_index_86740 ? add_88240 : sel_88237;
  assign add_88244 = sel_88241 + 8'h01;
  assign sel_88245 = array_index_88184 == array_index_86746 ? add_88244 : sel_88241;
  assign add_88248 = sel_88245 + 8'h01;
  assign sel_88249 = array_index_88184 == array_index_86752 ? add_88248 : sel_88245;
  assign add_88252 = sel_88249 + 8'h01;
  assign sel_88253 = array_index_88184 == array_index_86758 ? add_88252 : sel_88249;
  assign add_88256 = sel_88253 + 8'h01;
  assign sel_88257 = array_index_88184 == array_index_86764 ? add_88256 : sel_88253;
  assign add_88260 = sel_88257 + 8'h01;
  assign sel_88261 = array_index_88184 == array_index_86770 ? add_88260 : sel_88257;
  assign add_88264 = sel_88261 + 8'h01;
  assign sel_88265 = array_index_88184 == array_index_86776 ? add_88264 : sel_88261;
  assign add_88268 = sel_88265 + 8'h01;
  assign sel_88269 = array_index_88184 == array_index_86782 ? add_88268 : sel_88265;
  assign add_88272 = sel_88269 + 8'h01;
  assign sel_88273 = array_index_88184 == array_index_86788 ? add_88272 : sel_88269;
  assign add_88276 = sel_88273 + 8'h01;
  assign sel_88277 = array_index_88184 == array_index_86794 ? add_88276 : sel_88273;
  assign add_88280 = sel_88277 + 8'h01;
  assign sel_88281 = array_index_88184 == array_index_86800 ? add_88280 : sel_88277;
  assign add_88284 = sel_88281 + 8'h01;
  assign sel_88285 = array_index_88184 == array_index_86806 ? add_88284 : sel_88281;
  assign add_88288 = sel_88285 + 8'h01;
  assign sel_88289 = array_index_88184 == array_index_86812 ? add_88288 : sel_88285;
  assign add_88292 = sel_88289 + 8'h01;
  assign sel_88293 = array_index_88184 == array_index_86818 ? add_88292 : sel_88289;
  assign add_88296 = sel_88293 + 8'h01;
  assign sel_88297 = array_index_88184 == array_index_86824 ? add_88296 : sel_88293;
  assign add_88300 = sel_88297 + 8'h01;
  assign sel_88301 = array_index_88184 == array_index_86830 ? add_88300 : sel_88297;
  assign add_88305 = sel_88301 + 8'h01;
  assign array_index_88306 = set1_unflattened[5'h0d];
  assign sel_88307 = array_index_88184 == array_index_86836 ? add_88305 : sel_88301;
  assign add_88310 = sel_88307 + 8'h01;
  assign sel_88311 = array_index_88306 == array_index_86652 ? add_88310 : sel_88307;
  assign add_88314 = sel_88311 + 8'h01;
  assign sel_88315 = array_index_88306 == array_index_86656 ? add_88314 : sel_88311;
  assign add_88318 = sel_88315 + 8'h01;
  assign sel_88319 = array_index_88306 == array_index_86664 ? add_88318 : sel_88315;
  assign add_88322 = sel_88319 + 8'h01;
  assign sel_88323 = array_index_88306 == array_index_86672 ? add_88322 : sel_88319;
  assign add_88326 = sel_88323 + 8'h01;
  assign sel_88327 = array_index_88306 == array_index_86680 ? add_88326 : sel_88323;
  assign add_88330 = sel_88327 + 8'h01;
  assign sel_88331 = array_index_88306 == array_index_86688 ? add_88330 : sel_88327;
  assign add_88334 = sel_88331 + 8'h01;
  assign sel_88335 = array_index_88306 == array_index_86696 ? add_88334 : sel_88331;
  assign add_88338 = sel_88335 + 8'h01;
  assign sel_88339 = array_index_88306 == array_index_86704 ? add_88338 : sel_88335;
  assign add_88342 = sel_88339 + 8'h01;
  assign sel_88343 = array_index_88306 == array_index_86710 ? add_88342 : sel_88339;
  assign add_88346 = sel_88343 + 8'h01;
  assign sel_88347 = array_index_88306 == array_index_86716 ? add_88346 : sel_88343;
  assign add_88350 = sel_88347 + 8'h01;
  assign sel_88351 = array_index_88306 == array_index_86722 ? add_88350 : sel_88347;
  assign add_88354 = sel_88351 + 8'h01;
  assign sel_88355 = array_index_88306 == array_index_86728 ? add_88354 : sel_88351;
  assign add_88358 = sel_88355 + 8'h01;
  assign sel_88359 = array_index_88306 == array_index_86734 ? add_88358 : sel_88355;
  assign add_88362 = sel_88359 + 8'h01;
  assign sel_88363 = array_index_88306 == array_index_86740 ? add_88362 : sel_88359;
  assign add_88366 = sel_88363 + 8'h01;
  assign sel_88367 = array_index_88306 == array_index_86746 ? add_88366 : sel_88363;
  assign add_88370 = sel_88367 + 8'h01;
  assign sel_88371 = array_index_88306 == array_index_86752 ? add_88370 : sel_88367;
  assign add_88374 = sel_88371 + 8'h01;
  assign sel_88375 = array_index_88306 == array_index_86758 ? add_88374 : sel_88371;
  assign add_88378 = sel_88375 + 8'h01;
  assign sel_88379 = array_index_88306 == array_index_86764 ? add_88378 : sel_88375;
  assign add_88382 = sel_88379 + 8'h01;
  assign sel_88383 = array_index_88306 == array_index_86770 ? add_88382 : sel_88379;
  assign add_88386 = sel_88383 + 8'h01;
  assign sel_88387 = array_index_88306 == array_index_86776 ? add_88386 : sel_88383;
  assign add_88390 = sel_88387 + 8'h01;
  assign sel_88391 = array_index_88306 == array_index_86782 ? add_88390 : sel_88387;
  assign add_88394 = sel_88391 + 8'h01;
  assign sel_88395 = array_index_88306 == array_index_86788 ? add_88394 : sel_88391;
  assign add_88398 = sel_88395 + 8'h01;
  assign sel_88399 = array_index_88306 == array_index_86794 ? add_88398 : sel_88395;
  assign add_88402 = sel_88399 + 8'h01;
  assign sel_88403 = array_index_88306 == array_index_86800 ? add_88402 : sel_88399;
  assign add_88406 = sel_88403 + 8'h01;
  assign sel_88407 = array_index_88306 == array_index_86806 ? add_88406 : sel_88403;
  assign add_88410 = sel_88407 + 8'h01;
  assign sel_88411 = array_index_88306 == array_index_86812 ? add_88410 : sel_88407;
  assign add_88414 = sel_88411 + 8'h01;
  assign sel_88415 = array_index_88306 == array_index_86818 ? add_88414 : sel_88411;
  assign add_88418 = sel_88415 + 8'h01;
  assign sel_88419 = array_index_88306 == array_index_86824 ? add_88418 : sel_88415;
  assign add_88422 = sel_88419 + 8'h01;
  assign sel_88423 = array_index_88306 == array_index_86830 ? add_88422 : sel_88419;
  assign add_88427 = sel_88423 + 8'h01;
  assign array_index_88428 = set1_unflattened[5'h0e];
  assign sel_88429 = array_index_88306 == array_index_86836 ? add_88427 : sel_88423;
  assign add_88432 = sel_88429 + 8'h01;
  assign sel_88433 = array_index_88428 == array_index_86652 ? add_88432 : sel_88429;
  assign add_88436 = sel_88433 + 8'h01;
  assign sel_88437 = array_index_88428 == array_index_86656 ? add_88436 : sel_88433;
  assign add_88440 = sel_88437 + 8'h01;
  assign sel_88441 = array_index_88428 == array_index_86664 ? add_88440 : sel_88437;
  assign add_88444 = sel_88441 + 8'h01;
  assign sel_88445 = array_index_88428 == array_index_86672 ? add_88444 : sel_88441;
  assign add_88448 = sel_88445 + 8'h01;
  assign sel_88449 = array_index_88428 == array_index_86680 ? add_88448 : sel_88445;
  assign add_88452 = sel_88449 + 8'h01;
  assign sel_88453 = array_index_88428 == array_index_86688 ? add_88452 : sel_88449;
  assign add_88456 = sel_88453 + 8'h01;
  assign sel_88457 = array_index_88428 == array_index_86696 ? add_88456 : sel_88453;
  assign add_88460 = sel_88457 + 8'h01;
  assign sel_88461 = array_index_88428 == array_index_86704 ? add_88460 : sel_88457;
  assign add_88464 = sel_88461 + 8'h01;
  assign sel_88465 = array_index_88428 == array_index_86710 ? add_88464 : sel_88461;
  assign add_88468 = sel_88465 + 8'h01;
  assign sel_88469 = array_index_88428 == array_index_86716 ? add_88468 : sel_88465;
  assign add_88472 = sel_88469 + 8'h01;
  assign sel_88473 = array_index_88428 == array_index_86722 ? add_88472 : sel_88469;
  assign add_88476 = sel_88473 + 8'h01;
  assign sel_88477 = array_index_88428 == array_index_86728 ? add_88476 : sel_88473;
  assign add_88480 = sel_88477 + 8'h01;
  assign sel_88481 = array_index_88428 == array_index_86734 ? add_88480 : sel_88477;
  assign add_88484 = sel_88481 + 8'h01;
  assign sel_88485 = array_index_88428 == array_index_86740 ? add_88484 : sel_88481;
  assign add_88488 = sel_88485 + 8'h01;
  assign sel_88489 = array_index_88428 == array_index_86746 ? add_88488 : sel_88485;
  assign add_88492 = sel_88489 + 8'h01;
  assign sel_88493 = array_index_88428 == array_index_86752 ? add_88492 : sel_88489;
  assign add_88496 = sel_88493 + 8'h01;
  assign sel_88497 = array_index_88428 == array_index_86758 ? add_88496 : sel_88493;
  assign add_88500 = sel_88497 + 8'h01;
  assign sel_88501 = array_index_88428 == array_index_86764 ? add_88500 : sel_88497;
  assign add_88504 = sel_88501 + 8'h01;
  assign sel_88505 = array_index_88428 == array_index_86770 ? add_88504 : sel_88501;
  assign add_88508 = sel_88505 + 8'h01;
  assign sel_88509 = array_index_88428 == array_index_86776 ? add_88508 : sel_88505;
  assign add_88512 = sel_88509 + 8'h01;
  assign sel_88513 = array_index_88428 == array_index_86782 ? add_88512 : sel_88509;
  assign add_88516 = sel_88513 + 8'h01;
  assign sel_88517 = array_index_88428 == array_index_86788 ? add_88516 : sel_88513;
  assign add_88520 = sel_88517 + 8'h01;
  assign sel_88521 = array_index_88428 == array_index_86794 ? add_88520 : sel_88517;
  assign add_88524 = sel_88521 + 8'h01;
  assign sel_88525 = array_index_88428 == array_index_86800 ? add_88524 : sel_88521;
  assign add_88528 = sel_88525 + 8'h01;
  assign sel_88529 = array_index_88428 == array_index_86806 ? add_88528 : sel_88525;
  assign add_88532 = sel_88529 + 8'h01;
  assign sel_88533 = array_index_88428 == array_index_86812 ? add_88532 : sel_88529;
  assign add_88536 = sel_88533 + 8'h01;
  assign sel_88537 = array_index_88428 == array_index_86818 ? add_88536 : sel_88533;
  assign add_88540 = sel_88537 + 8'h01;
  assign sel_88541 = array_index_88428 == array_index_86824 ? add_88540 : sel_88537;
  assign add_88544 = sel_88541 + 8'h01;
  assign sel_88545 = array_index_88428 == array_index_86830 ? add_88544 : sel_88541;
  assign add_88549 = sel_88545 + 8'h01;
  assign array_index_88550 = set1_unflattened[5'h0f];
  assign sel_88551 = array_index_88428 == array_index_86836 ? add_88549 : sel_88545;
  assign add_88554 = sel_88551 + 8'h01;
  assign sel_88555 = array_index_88550 == array_index_86652 ? add_88554 : sel_88551;
  assign add_88558 = sel_88555 + 8'h01;
  assign sel_88559 = array_index_88550 == array_index_86656 ? add_88558 : sel_88555;
  assign add_88562 = sel_88559 + 8'h01;
  assign sel_88563 = array_index_88550 == array_index_86664 ? add_88562 : sel_88559;
  assign add_88566 = sel_88563 + 8'h01;
  assign sel_88567 = array_index_88550 == array_index_86672 ? add_88566 : sel_88563;
  assign add_88570 = sel_88567 + 8'h01;
  assign sel_88571 = array_index_88550 == array_index_86680 ? add_88570 : sel_88567;
  assign add_88574 = sel_88571 + 8'h01;
  assign sel_88575 = array_index_88550 == array_index_86688 ? add_88574 : sel_88571;
  assign add_88578 = sel_88575 + 8'h01;
  assign sel_88579 = array_index_88550 == array_index_86696 ? add_88578 : sel_88575;
  assign add_88582 = sel_88579 + 8'h01;
  assign sel_88583 = array_index_88550 == array_index_86704 ? add_88582 : sel_88579;
  assign add_88586 = sel_88583 + 8'h01;
  assign sel_88587 = array_index_88550 == array_index_86710 ? add_88586 : sel_88583;
  assign add_88590 = sel_88587 + 8'h01;
  assign sel_88591 = array_index_88550 == array_index_86716 ? add_88590 : sel_88587;
  assign add_88594 = sel_88591 + 8'h01;
  assign sel_88595 = array_index_88550 == array_index_86722 ? add_88594 : sel_88591;
  assign add_88598 = sel_88595 + 8'h01;
  assign sel_88599 = array_index_88550 == array_index_86728 ? add_88598 : sel_88595;
  assign add_88602 = sel_88599 + 8'h01;
  assign sel_88603 = array_index_88550 == array_index_86734 ? add_88602 : sel_88599;
  assign add_88606 = sel_88603 + 8'h01;
  assign sel_88607 = array_index_88550 == array_index_86740 ? add_88606 : sel_88603;
  assign add_88610 = sel_88607 + 8'h01;
  assign sel_88611 = array_index_88550 == array_index_86746 ? add_88610 : sel_88607;
  assign add_88614 = sel_88611 + 8'h01;
  assign sel_88615 = array_index_88550 == array_index_86752 ? add_88614 : sel_88611;
  assign add_88618 = sel_88615 + 8'h01;
  assign sel_88619 = array_index_88550 == array_index_86758 ? add_88618 : sel_88615;
  assign add_88622 = sel_88619 + 8'h01;
  assign sel_88623 = array_index_88550 == array_index_86764 ? add_88622 : sel_88619;
  assign add_88626 = sel_88623 + 8'h01;
  assign sel_88627 = array_index_88550 == array_index_86770 ? add_88626 : sel_88623;
  assign add_88630 = sel_88627 + 8'h01;
  assign sel_88631 = array_index_88550 == array_index_86776 ? add_88630 : sel_88627;
  assign add_88634 = sel_88631 + 8'h01;
  assign sel_88635 = array_index_88550 == array_index_86782 ? add_88634 : sel_88631;
  assign add_88638 = sel_88635 + 8'h01;
  assign sel_88639 = array_index_88550 == array_index_86788 ? add_88638 : sel_88635;
  assign add_88642 = sel_88639 + 8'h01;
  assign sel_88643 = array_index_88550 == array_index_86794 ? add_88642 : sel_88639;
  assign add_88646 = sel_88643 + 8'h01;
  assign sel_88647 = array_index_88550 == array_index_86800 ? add_88646 : sel_88643;
  assign add_88650 = sel_88647 + 8'h01;
  assign sel_88651 = array_index_88550 == array_index_86806 ? add_88650 : sel_88647;
  assign add_88654 = sel_88651 + 8'h01;
  assign sel_88655 = array_index_88550 == array_index_86812 ? add_88654 : sel_88651;
  assign add_88658 = sel_88655 + 8'h01;
  assign sel_88659 = array_index_88550 == array_index_86818 ? add_88658 : sel_88655;
  assign add_88662 = sel_88659 + 8'h01;
  assign sel_88663 = array_index_88550 == array_index_86824 ? add_88662 : sel_88659;
  assign add_88666 = sel_88663 + 8'h01;
  assign sel_88667 = array_index_88550 == array_index_86830 ? add_88666 : sel_88663;
  assign add_88671 = sel_88667 + 8'h01;
  assign array_index_88672 = set1_unflattened[5'h10];
  assign sel_88673 = array_index_88550 == array_index_86836 ? add_88671 : sel_88667;
  assign add_88676 = sel_88673 + 8'h01;
  assign sel_88677 = array_index_88672 == array_index_86652 ? add_88676 : sel_88673;
  assign add_88680 = sel_88677 + 8'h01;
  assign sel_88681 = array_index_88672 == array_index_86656 ? add_88680 : sel_88677;
  assign add_88684 = sel_88681 + 8'h01;
  assign sel_88685 = array_index_88672 == array_index_86664 ? add_88684 : sel_88681;
  assign add_88688 = sel_88685 + 8'h01;
  assign sel_88689 = array_index_88672 == array_index_86672 ? add_88688 : sel_88685;
  assign add_88692 = sel_88689 + 8'h01;
  assign sel_88693 = array_index_88672 == array_index_86680 ? add_88692 : sel_88689;
  assign add_88696 = sel_88693 + 8'h01;
  assign sel_88697 = array_index_88672 == array_index_86688 ? add_88696 : sel_88693;
  assign add_88700 = sel_88697 + 8'h01;
  assign sel_88701 = array_index_88672 == array_index_86696 ? add_88700 : sel_88697;
  assign add_88704 = sel_88701 + 8'h01;
  assign sel_88705 = array_index_88672 == array_index_86704 ? add_88704 : sel_88701;
  assign add_88708 = sel_88705 + 8'h01;
  assign sel_88709 = array_index_88672 == array_index_86710 ? add_88708 : sel_88705;
  assign add_88712 = sel_88709 + 8'h01;
  assign sel_88713 = array_index_88672 == array_index_86716 ? add_88712 : sel_88709;
  assign add_88716 = sel_88713 + 8'h01;
  assign sel_88717 = array_index_88672 == array_index_86722 ? add_88716 : sel_88713;
  assign add_88720 = sel_88717 + 8'h01;
  assign sel_88721 = array_index_88672 == array_index_86728 ? add_88720 : sel_88717;
  assign add_88724 = sel_88721 + 8'h01;
  assign sel_88725 = array_index_88672 == array_index_86734 ? add_88724 : sel_88721;
  assign add_88728 = sel_88725 + 8'h01;
  assign sel_88729 = array_index_88672 == array_index_86740 ? add_88728 : sel_88725;
  assign add_88732 = sel_88729 + 8'h01;
  assign sel_88733 = array_index_88672 == array_index_86746 ? add_88732 : sel_88729;
  assign add_88736 = sel_88733 + 8'h01;
  assign sel_88737 = array_index_88672 == array_index_86752 ? add_88736 : sel_88733;
  assign add_88740 = sel_88737 + 8'h01;
  assign sel_88741 = array_index_88672 == array_index_86758 ? add_88740 : sel_88737;
  assign add_88744 = sel_88741 + 8'h01;
  assign sel_88745 = array_index_88672 == array_index_86764 ? add_88744 : sel_88741;
  assign add_88748 = sel_88745 + 8'h01;
  assign sel_88749 = array_index_88672 == array_index_86770 ? add_88748 : sel_88745;
  assign add_88752 = sel_88749 + 8'h01;
  assign sel_88753 = array_index_88672 == array_index_86776 ? add_88752 : sel_88749;
  assign add_88756 = sel_88753 + 8'h01;
  assign sel_88757 = array_index_88672 == array_index_86782 ? add_88756 : sel_88753;
  assign add_88760 = sel_88757 + 8'h01;
  assign sel_88761 = array_index_88672 == array_index_86788 ? add_88760 : sel_88757;
  assign add_88764 = sel_88761 + 8'h01;
  assign sel_88765 = array_index_88672 == array_index_86794 ? add_88764 : sel_88761;
  assign add_88768 = sel_88765 + 8'h01;
  assign sel_88769 = array_index_88672 == array_index_86800 ? add_88768 : sel_88765;
  assign add_88772 = sel_88769 + 8'h01;
  assign sel_88773 = array_index_88672 == array_index_86806 ? add_88772 : sel_88769;
  assign add_88776 = sel_88773 + 8'h01;
  assign sel_88777 = array_index_88672 == array_index_86812 ? add_88776 : sel_88773;
  assign add_88780 = sel_88777 + 8'h01;
  assign sel_88781 = array_index_88672 == array_index_86818 ? add_88780 : sel_88777;
  assign add_88784 = sel_88781 + 8'h01;
  assign sel_88785 = array_index_88672 == array_index_86824 ? add_88784 : sel_88781;
  assign add_88788 = sel_88785 + 8'h01;
  assign sel_88789 = array_index_88672 == array_index_86830 ? add_88788 : sel_88785;
  assign add_88793 = sel_88789 + 8'h01;
  assign array_index_88794 = set1_unflattened[5'h11];
  assign sel_88795 = array_index_88672 == array_index_86836 ? add_88793 : sel_88789;
  assign add_88798 = sel_88795 + 8'h01;
  assign sel_88799 = array_index_88794 == array_index_86652 ? add_88798 : sel_88795;
  assign add_88802 = sel_88799 + 8'h01;
  assign sel_88803 = array_index_88794 == array_index_86656 ? add_88802 : sel_88799;
  assign add_88806 = sel_88803 + 8'h01;
  assign sel_88807 = array_index_88794 == array_index_86664 ? add_88806 : sel_88803;
  assign add_88810 = sel_88807 + 8'h01;
  assign sel_88811 = array_index_88794 == array_index_86672 ? add_88810 : sel_88807;
  assign add_88814 = sel_88811 + 8'h01;
  assign sel_88815 = array_index_88794 == array_index_86680 ? add_88814 : sel_88811;
  assign add_88818 = sel_88815 + 8'h01;
  assign sel_88819 = array_index_88794 == array_index_86688 ? add_88818 : sel_88815;
  assign add_88822 = sel_88819 + 8'h01;
  assign sel_88823 = array_index_88794 == array_index_86696 ? add_88822 : sel_88819;
  assign add_88826 = sel_88823 + 8'h01;
  assign sel_88827 = array_index_88794 == array_index_86704 ? add_88826 : sel_88823;
  assign add_88830 = sel_88827 + 8'h01;
  assign sel_88831 = array_index_88794 == array_index_86710 ? add_88830 : sel_88827;
  assign add_88834 = sel_88831 + 8'h01;
  assign sel_88835 = array_index_88794 == array_index_86716 ? add_88834 : sel_88831;
  assign add_88838 = sel_88835 + 8'h01;
  assign sel_88839 = array_index_88794 == array_index_86722 ? add_88838 : sel_88835;
  assign add_88842 = sel_88839 + 8'h01;
  assign sel_88843 = array_index_88794 == array_index_86728 ? add_88842 : sel_88839;
  assign add_88846 = sel_88843 + 8'h01;
  assign sel_88847 = array_index_88794 == array_index_86734 ? add_88846 : sel_88843;
  assign add_88850 = sel_88847 + 8'h01;
  assign sel_88851 = array_index_88794 == array_index_86740 ? add_88850 : sel_88847;
  assign add_88854 = sel_88851 + 8'h01;
  assign sel_88855 = array_index_88794 == array_index_86746 ? add_88854 : sel_88851;
  assign add_88858 = sel_88855 + 8'h01;
  assign sel_88859 = array_index_88794 == array_index_86752 ? add_88858 : sel_88855;
  assign add_88862 = sel_88859 + 8'h01;
  assign sel_88863 = array_index_88794 == array_index_86758 ? add_88862 : sel_88859;
  assign add_88866 = sel_88863 + 8'h01;
  assign sel_88867 = array_index_88794 == array_index_86764 ? add_88866 : sel_88863;
  assign add_88870 = sel_88867 + 8'h01;
  assign sel_88871 = array_index_88794 == array_index_86770 ? add_88870 : sel_88867;
  assign add_88874 = sel_88871 + 8'h01;
  assign sel_88875 = array_index_88794 == array_index_86776 ? add_88874 : sel_88871;
  assign add_88878 = sel_88875 + 8'h01;
  assign sel_88879 = array_index_88794 == array_index_86782 ? add_88878 : sel_88875;
  assign add_88882 = sel_88879 + 8'h01;
  assign sel_88883 = array_index_88794 == array_index_86788 ? add_88882 : sel_88879;
  assign add_88886 = sel_88883 + 8'h01;
  assign sel_88887 = array_index_88794 == array_index_86794 ? add_88886 : sel_88883;
  assign add_88890 = sel_88887 + 8'h01;
  assign sel_88891 = array_index_88794 == array_index_86800 ? add_88890 : sel_88887;
  assign add_88894 = sel_88891 + 8'h01;
  assign sel_88895 = array_index_88794 == array_index_86806 ? add_88894 : sel_88891;
  assign add_88898 = sel_88895 + 8'h01;
  assign sel_88899 = array_index_88794 == array_index_86812 ? add_88898 : sel_88895;
  assign add_88902 = sel_88899 + 8'h01;
  assign sel_88903 = array_index_88794 == array_index_86818 ? add_88902 : sel_88899;
  assign add_88906 = sel_88903 + 8'h01;
  assign sel_88907 = array_index_88794 == array_index_86824 ? add_88906 : sel_88903;
  assign add_88910 = sel_88907 + 8'h01;
  assign sel_88911 = array_index_88794 == array_index_86830 ? add_88910 : sel_88907;
  assign add_88915 = sel_88911 + 8'h01;
  assign array_index_88916 = set1_unflattened[5'h12];
  assign sel_88917 = array_index_88794 == array_index_86836 ? add_88915 : sel_88911;
  assign add_88920 = sel_88917 + 8'h01;
  assign sel_88921 = array_index_88916 == array_index_86652 ? add_88920 : sel_88917;
  assign add_88924 = sel_88921 + 8'h01;
  assign sel_88925 = array_index_88916 == array_index_86656 ? add_88924 : sel_88921;
  assign add_88928 = sel_88925 + 8'h01;
  assign sel_88929 = array_index_88916 == array_index_86664 ? add_88928 : sel_88925;
  assign add_88932 = sel_88929 + 8'h01;
  assign sel_88933 = array_index_88916 == array_index_86672 ? add_88932 : sel_88929;
  assign add_88936 = sel_88933 + 8'h01;
  assign sel_88937 = array_index_88916 == array_index_86680 ? add_88936 : sel_88933;
  assign add_88940 = sel_88937 + 8'h01;
  assign sel_88941 = array_index_88916 == array_index_86688 ? add_88940 : sel_88937;
  assign add_88944 = sel_88941 + 8'h01;
  assign sel_88945 = array_index_88916 == array_index_86696 ? add_88944 : sel_88941;
  assign add_88948 = sel_88945 + 8'h01;
  assign sel_88949 = array_index_88916 == array_index_86704 ? add_88948 : sel_88945;
  assign add_88952 = sel_88949 + 8'h01;
  assign sel_88953 = array_index_88916 == array_index_86710 ? add_88952 : sel_88949;
  assign add_88956 = sel_88953 + 8'h01;
  assign sel_88957 = array_index_88916 == array_index_86716 ? add_88956 : sel_88953;
  assign add_88960 = sel_88957 + 8'h01;
  assign sel_88961 = array_index_88916 == array_index_86722 ? add_88960 : sel_88957;
  assign add_88964 = sel_88961 + 8'h01;
  assign sel_88965 = array_index_88916 == array_index_86728 ? add_88964 : sel_88961;
  assign add_88968 = sel_88965 + 8'h01;
  assign sel_88969 = array_index_88916 == array_index_86734 ? add_88968 : sel_88965;
  assign add_88972 = sel_88969 + 8'h01;
  assign sel_88973 = array_index_88916 == array_index_86740 ? add_88972 : sel_88969;
  assign add_88976 = sel_88973 + 8'h01;
  assign sel_88977 = array_index_88916 == array_index_86746 ? add_88976 : sel_88973;
  assign add_88980 = sel_88977 + 8'h01;
  assign sel_88981 = array_index_88916 == array_index_86752 ? add_88980 : sel_88977;
  assign add_88984 = sel_88981 + 8'h01;
  assign sel_88985 = array_index_88916 == array_index_86758 ? add_88984 : sel_88981;
  assign add_88988 = sel_88985 + 8'h01;
  assign sel_88989 = array_index_88916 == array_index_86764 ? add_88988 : sel_88985;
  assign add_88992 = sel_88989 + 8'h01;
  assign sel_88993 = array_index_88916 == array_index_86770 ? add_88992 : sel_88989;
  assign add_88996 = sel_88993 + 8'h01;
  assign sel_88997 = array_index_88916 == array_index_86776 ? add_88996 : sel_88993;
  assign add_89000 = sel_88997 + 8'h01;
  assign sel_89001 = array_index_88916 == array_index_86782 ? add_89000 : sel_88997;
  assign add_89004 = sel_89001 + 8'h01;
  assign sel_89005 = array_index_88916 == array_index_86788 ? add_89004 : sel_89001;
  assign add_89008 = sel_89005 + 8'h01;
  assign sel_89009 = array_index_88916 == array_index_86794 ? add_89008 : sel_89005;
  assign add_89012 = sel_89009 + 8'h01;
  assign sel_89013 = array_index_88916 == array_index_86800 ? add_89012 : sel_89009;
  assign add_89016 = sel_89013 + 8'h01;
  assign sel_89017 = array_index_88916 == array_index_86806 ? add_89016 : sel_89013;
  assign add_89020 = sel_89017 + 8'h01;
  assign sel_89021 = array_index_88916 == array_index_86812 ? add_89020 : sel_89017;
  assign add_89024 = sel_89021 + 8'h01;
  assign sel_89025 = array_index_88916 == array_index_86818 ? add_89024 : sel_89021;
  assign add_89028 = sel_89025 + 8'h01;
  assign sel_89029 = array_index_88916 == array_index_86824 ? add_89028 : sel_89025;
  assign add_89032 = sel_89029 + 8'h01;
  assign sel_89033 = array_index_88916 == array_index_86830 ? add_89032 : sel_89029;
  assign add_89037 = sel_89033 + 8'h01;
  assign array_index_89038 = set1_unflattened[5'h13];
  assign sel_89039 = array_index_88916 == array_index_86836 ? add_89037 : sel_89033;
  assign add_89042 = sel_89039 + 8'h01;
  assign sel_89043 = array_index_89038 == array_index_86652 ? add_89042 : sel_89039;
  assign add_89046 = sel_89043 + 8'h01;
  assign sel_89047 = array_index_89038 == array_index_86656 ? add_89046 : sel_89043;
  assign add_89050 = sel_89047 + 8'h01;
  assign sel_89051 = array_index_89038 == array_index_86664 ? add_89050 : sel_89047;
  assign add_89054 = sel_89051 + 8'h01;
  assign sel_89055 = array_index_89038 == array_index_86672 ? add_89054 : sel_89051;
  assign add_89058 = sel_89055 + 8'h01;
  assign sel_89059 = array_index_89038 == array_index_86680 ? add_89058 : sel_89055;
  assign add_89062 = sel_89059 + 8'h01;
  assign sel_89063 = array_index_89038 == array_index_86688 ? add_89062 : sel_89059;
  assign add_89066 = sel_89063 + 8'h01;
  assign sel_89067 = array_index_89038 == array_index_86696 ? add_89066 : sel_89063;
  assign add_89070 = sel_89067 + 8'h01;
  assign sel_89071 = array_index_89038 == array_index_86704 ? add_89070 : sel_89067;
  assign add_89074 = sel_89071 + 8'h01;
  assign sel_89075 = array_index_89038 == array_index_86710 ? add_89074 : sel_89071;
  assign add_89078 = sel_89075 + 8'h01;
  assign sel_89079 = array_index_89038 == array_index_86716 ? add_89078 : sel_89075;
  assign add_89082 = sel_89079 + 8'h01;
  assign sel_89083 = array_index_89038 == array_index_86722 ? add_89082 : sel_89079;
  assign add_89086 = sel_89083 + 8'h01;
  assign sel_89087 = array_index_89038 == array_index_86728 ? add_89086 : sel_89083;
  assign add_89090 = sel_89087 + 8'h01;
  assign sel_89091 = array_index_89038 == array_index_86734 ? add_89090 : sel_89087;
  assign add_89094 = sel_89091 + 8'h01;
  assign sel_89095 = array_index_89038 == array_index_86740 ? add_89094 : sel_89091;
  assign add_89098 = sel_89095 + 8'h01;
  assign sel_89099 = array_index_89038 == array_index_86746 ? add_89098 : sel_89095;
  assign add_89102 = sel_89099 + 8'h01;
  assign sel_89103 = array_index_89038 == array_index_86752 ? add_89102 : sel_89099;
  assign add_89106 = sel_89103 + 8'h01;
  assign sel_89107 = array_index_89038 == array_index_86758 ? add_89106 : sel_89103;
  assign add_89110 = sel_89107 + 8'h01;
  assign sel_89111 = array_index_89038 == array_index_86764 ? add_89110 : sel_89107;
  assign add_89114 = sel_89111 + 8'h01;
  assign sel_89115 = array_index_89038 == array_index_86770 ? add_89114 : sel_89111;
  assign add_89118 = sel_89115 + 8'h01;
  assign sel_89119 = array_index_89038 == array_index_86776 ? add_89118 : sel_89115;
  assign add_89122 = sel_89119 + 8'h01;
  assign sel_89123 = array_index_89038 == array_index_86782 ? add_89122 : sel_89119;
  assign add_89126 = sel_89123 + 8'h01;
  assign sel_89127 = array_index_89038 == array_index_86788 ? add_89126 : sel_89123;
  assign add_89130 = sel_89127 + 8'h01;
  assign sel_89131 = array_index_89038 == array_index_86794 ? add_89130 : sel_89127;
  assign add_89134 = sel_89131 + 8'h01;
  assign sel_89135 = array_index_89038 == array_index_86800 ? add_89134 : sel_89131;
  assign add_89138 = sel_89135 + 8'h01;
  assign sel_89139 = array_index_89038 == array_index_86806 ? add_89138 : sel_89135;
  assign add_89142 = sel_89139 + 8'h01;
  assign sel_89143 = array_index_89038 == array_index_86812 ? add_89142 : sel_89139;
  assign add_89146 = sel_89143 + 8'h01;
  assign sel_89147 = array_index_89038 == array_index_86818 ? add_89146 : sel_89143;
  assign add_89150 = sel_89147 + 8'h01;
  assign sel_89151 = array_index_89038 == array_index_86824 ? add_89150 : sel_89147;
  assign add_89154 = sel_89151 + 8'h01;
  assign sel_89155 = array_index_89038 == array_index_86830 ? add_89154 : sel_89151;
  assign add_89159 = sel_89155 + 8'h01;
  assign array_index_89160 = set1_unflattened[5'h14];
  assign sel_89161 = array_index_89038 == array_index_86836 ? add_89159 : sel_89155;
  assign add_89164 = sel_89161 + 8'h01;
  assign sel_89165 = array_index_89160 == array_index_86652 ? add_89164 : sel_89161;
  assign add_89168 = sel_89165 + 8'h01;
  assign sel_89169 = array_index_89160 == array_index_86656 ? add_89168 : sel_89165;
  assign add_89172 = sel_89169 + 8'h01;
  assign sel_89173 = array_index_89160 == array_index_86664 ? add_89172 : sel_89169;
  assign add_89176 = sel_89173 + 8'h01;
  assign sel_89177 = array_index_89160 == array_index_86672 ? add_89176 : sel_89173;
  assign add_89180 = sel_89177 + 8'h01;
  assign sel_89181 = array_index_89160 == array_index_86680 ? add_89180 : sel_89177;
  assign add_89184 = sel_89181 + 8'h01;
  assign sel_89185 = array_index_89160 == array_index_86688 ? add_89184 : sel_89181;
  assign add_89188 = sel_89185 + 8'h01;
  assign sel_89189 = array_index_89160 == array_index_86696 ? add_89188 : sel_89185;
  assign add_89192 = sel_89189 + 8'h01;
  assign sel_89193 = array_index_89160 == array_index_86704 ? add_89192 : sel_89189;
  assign add_89196 = sel_89193 + 8'h01;
  assign sel_89197 = array_index_89160 == array_index_86710 ? add_89196 : sel_89193;
  assign add_89200 = sel_89197 + 8'h01;
  assign sel_89201 = array_index_89160 == array_index_86716 ? add_89200 : sel_89197;
  assign add_89204 = sel_89201 + 8'h01;
  assign sel_89205 = array_index_89160 == array_index_86722 ? add_89204 : sel_89201;
  assign add_89208 = sel_89205 + 8'h01;
  assign sel_89209 = array_index_89160 == array_index_86728 ? add_89208 : sel_89205;
  assign add_89212 = sel_89209 + 8'h01;
  assign sel_89213 = array_index_89160 == array_index_86734 ? add_89212 : sel_89209;
  assign add_89216 = sel_89213 + 8'h01;
  assign sel_89217 = array_index_89160 == array_index_86740 ? add_89216 : sel_89213;
  assign add_89220 = sel_89217 + 8'h01;
  assign sel_89221 = array_index_89160 == array_index_86746 ? add_89220 : sel_89217;
  assign add_89224 = sel_89221 + 8'h01;
  assign sel_89225 = array_index_89160 == array_index_86752 ? add_89224 : sel_89221;
  assign add_89228 = sel_89225 + 8'h01;
  assign sel_89229 = array_index_89160 == array_index_86758 ? add_89228 : sel_89225;
  assign add_89232 = sel_89229 + 8'h01;
  assign sel_89233 = array_index_89160 == array_index_86764 ? add_89232 : sel_89229;
  assign add_89236 = sel_89233 + 8'h01;
  assign sel_89237 = array_index_89160 == array_index_86770 ? add_89236 : sel_89233;
  assign add_89240 = sel_89237 + 8'h01;
  assign sel_89241 = array_index_89160 == array_index_86776 ? add_89240 : sel_89237;
  assign add_89244 = sel_89241 + 8'h01;
  assign sel_89245 = array_index_89160 == array_index_86782 ? add_89244 : sel_89241;
  assign add_89248 = sel_89245 + 8'h01;
  assign sel_89249 = array_index_89160 == array_index_86788 ? add_89248 : sel_89245;
  assign add_89252 = sel_89249 + 8'h01;
  assign sel_89253 = array_index_89160 == array_index_86794 ? add_89252 : sel_89249;
  assign add_89256 = sel_89253 + 8'h01;
  assign sel_89257 = array_index_89160 == array_index_86800 ? add_89256 : sel_89253;
  assign add_89260 = sel_89257 + 8'h01;
  assign sel_89261 = array_index_89160 == array_index_86806 ? add_89260 : sel_89257;
  assign add_89264 = sel_89261 + 8'h01;
  assign sel_89265 = array_index_89160 == array_index_86812 ? add_89264 : sel_89261;
  assign add_89268 = sel_89265 + 8'h01;
  assign sel_89269 = array_index_89160 == array_index_86818 ? add_89268 : sel_89265;
  assign add_89272 = sel_89269 + 8'h01;
  assign sel_89273 = array_index_89160 == array_index_86824 ? add_89272 : sel_89269;
  assign add_89276 = sel_89273 + 8'h01;
  assign sel_89277 = array_index_89160 == array_index_86830 ? add_89276 : sel_89273;
  assign add_89281 = sel_89277 + 8'h01;
  assign array_index_89282 = set1_unflattened[5'h15];
  assign sel_89283 = array_index_89160 == array_index_86836 ? add_89281 : sel_89277;
  assign add_89286 = sel_89283 + 8'h01;
  assign sel_89287 = array_index_89282 == array_index_86652 ? add_89286 : sel_89283;
  assign add_89290 = sel_89287 + 8'h01;
  assign sel_89291 = array_index_89282 == array_index_86656 ? add_89290 : sel_89287;
  assign add_89294 = sel_89291 + 8'h01;
  assign sel_89295 = array_index_89282 == array_index_86664 ? add_89294 : sel_89291;
  assign add_89298 = sel_89295 + 8'h01;
  assign sel_89299 = array_index_89282 == array_index_86672 ? add_89298 : sel_89295;
  assign add_89302 = sel_89299 + 8'h01;
  assign sel_89303 = array_index_89282 == array_index_86680 ? add_89302 : sel_89299;
  assign add_89306 = sel_89303 + 8'h01;
  assign sel_89307 = array_index_89282 == array_index_86688 ? add_89306 : sel_89303;
  assign add_89310 = sel_89307 + 8'h01;
  assign sel_89311 = array_index_89282 == array_index_86696 ? add_89310 : sel_89307;
  assign add_89314 = sel_89311 + 8'h01;
  assign sel_89315 = array_index_89282 == array_index_86704 ? add_89314 : sel_89311;
  assign add_89318 = sel_89315 + 8'h01;
  assign sel_89319 = array_index_89282 == array_index_86710 ? add_89318 : sel_89315;
  assign add_89322 = sel_89319 + 8'h01;
  assign sel_89323 = array_index_89282 == array_index_86716 ? add_89322 : sel_89319;
  assign add_89326 = sel_89323 + 8'h01;
  assign sel_89327 = array_index_89282 == array_index_86722 ? add_89326 : sel_89323;
  assign add_89330 = sel_89327 + 8'h01;
  assign sel_89331 = array_index_89282 == array_index_86728 ? add_89330 : sel_89327;
  assign add_89334 = sel_89331 + 8'h01;
  assign sel_89335 = array_index_89282 == array_index_86734 ? add_89334 : sel_89331;
  assign add_89338 = sel_89335 + 8'h01;
  assign sel_89339 = array_index_89282 == array_index_86740 ? add_89338 : sel_89335;
  assign add_89342 = sel_89339 + 8'h01;
  assign sel_89343 = array_index_89282 == array_index_86746 ? add_89342 : sel_89339;
  assign add_89346 = sel_89343 + 8'h01;
  assign sel_89347 = array_index_89282 == array_index_86752 ? add_89346 : sel_89343;
  assign add_89350 = sel_89347 + 8'h01;
  assign sel_89351 = array_index_89282 == array_index_86758 ? add_89350 : sel_89347;
  assign add_89354 = sel_89351 + 8'h01;
  assign sel_89355 = array_index_89282 == array_index_86764 ? add_89354 : sel_89351;
  assign add_89358 = sel_89355 + 8'h01;
  assign sel_89359 = array_index_89282 == array_index_86770 ? add_89358 : sel_89355;
  assign add_89362 = sel_89359 + 8'h01;
  assign sel_89363 = array_index_89282 == array_index_86776 ? add_89362 : sel_89359;
  assign add_89366 = sel_89363 + 8'h01;
  assign sel_89367 = array_index_89282 == array_index_86782 ? add_89366 : sel_89363;
  assign add_89370 = sel_89367 + 8'h01;
  assign sel_89371 = array_index_89282 == array_index_86788 ? add_89370 : sel_89367;
  assign add_89374 = sel_89371 + 8'h01;
  assign sel_89375 = array_index_89282 == array_index_86794 ? add_89374 : sel_89371;
  assign add_89378 = sel_89375 + 8'h01;
  assign sel_89379 = array_index_89282 == array_index_86800 ? add_89378 : sel_89375;
  assign add_89382 = sel_89379 + 8'h01;
  assign sel_89383 = array_index_89282 == array_index_86806 ? add_89382 : sel_89379;
  assign add_89386 = sel_89383 + 8'h01;
  assign sel_89387 = array_index_89282 == array_index_86812 ? add_89386 : sel_89383;
  assign add_89390 = sel_89387 + 8'h01;
  assign sel_89391 = array_index_89282 == array_index_86818 ? add_89390 : sel_89387;
  assign add_89394 = sel_89391 + 8'h01;
  assign sel_89395 = array_index_89282 == array_index_86824 ? add_89394 : sel_89391;
  assign add_89398 = sel_89395 + 8'h01;
  assign sel_89399 = array_index_89282 == array_index_86830 ? add_89398 : sel_89395;
  assign add_89403 = sel_89399 + 8'h01;
  assign array_index_89404 = set1_unflattened[5'h16];
  assign sel_89405 = array_index_89282 == array_index_86836 ? add_89403 : sel_89399;
  assign add_89408 = sel_89405 + 8'h01;
  assign sel_89409 = array_index_89404 == array_index_86652 ? add_89408 : sel_89405;
  assign add_89412 = sel_89409 + 8'h01;
  assign sel_89413 = array_index_89404 == array_index_86656 ? add_89412 : sel_89409;
  assign add_89416 = sel_89413 + 8'h01;
  assign sel_89417 = array_index_89404 == array_index_86664 ? add_89416 : sel_89413;
  assign add_89420 = sel_89417 + 8'h01;
  assign sel_89421 = array_index_89404 == array_index_86672 ? add_89420 : sel_89417;
  assign add_89424 = sel_89421 + 8'h01;
  assign sel_89425 = array_index_89404 == array_index_86680 ? add_89424 : sel_89421;
  assign add_89428 = sel_89425 + 8'h01;
  assign sel_89429 = array_index_89404 == array_index_86688 ? add_89428 : sel_89425;
  assign add_89432 = sel_89429 + 8'h01;
  assign sel_89433 = array_index_89404 == array_index_86696 ? add_89432 : sel_89429;
  assign add_89436 = sel_89433 + 8'h01;
  assign sel_89437 = array_index_89404 == array_index_86704 ? add_89436 : sel_89433;
  assign add_89440 = sel_89437 + 8'h01;
  assign sel_89441 = array_index_89404 == array_index_86710 ? add_89440 : sel_89437;
  assign add_89444 = sel_89441 + 8'h01;
  assign sel_89445 = array_index_89404 == array_index_86716 ? add_89444 : sel_89441;
  assign add_89448 = sel_89445 + 8'h01;
  assign sel_89449 = array_index_89404 == array_index_86722 ? add_89448 : sel_89445;
  assign add_89452 = sel_89449 + 8'h01;
  assign sel_89453 = array_index_89404 == array_index_86728 ? add_89452 : sel_89449;
  assign add_89456 = sel_89453 + 8'h01;
  assign sel_89457 = array_index_89404 == array_index_86734 ? add_89456 : sel_89453;
  assign add_89460 = sel_89457 + 8'h01;
  assign sel_89461 = array_index_89404 == array_index_86740 ? add_89460 : sel_89457;
  assign add_89464 = sel_89461 + 8'h01;
  assign sel_89465 = array_index_89404 == array_index_86746 ? add_89464 : sel_89461;
  assign add_89468 = sel_89465 + 8'h01;
  assign sel_89469 = array_index_89404 == array_index_86752 ? add_89468 : sel_89465;
  assign add_89472 = sel_89469 + 8'h01;
  assign sel_89473 = array_index_89404 == array_index_86758 ? add_89472 : sel_89469;
  assign add_89476 = sel_89473 + 8'h01;
  assign sel_89477 = array_index_89404 == array_index_86764 ? add_89476 : sel_89473;
  assign add_89480 = sel_89477 + 8'h01;
  assign sel_89481 = array_index_89404 == array_index_86770 ? add_89480 : sel_89477;
  assign add_89484 = sel_89481 + 8'h01;
  assign sel_89485 = array_index_89404 == array_index_86776 ? add_89484 : sel_89481;
  assign add_89488 = sel_89485 + 8'h01;
  assign sel_89489 = array_index_89404 == array_index_86782 ? add_89488 : sel_89485;
  assign add_89492 = sel_89489 + 8'h01;
  assign sel_89493 = array_index_89404 == array_index_86788 ? add_89492 : sel_89489;
  assign add_89496 = sel_89493 + 8'h01;
  assign sel_89497 = array_index_89404 == array_index_86794 ? add_89496 : sel_89493;
  assign add_89500 = sel_89497 + 8'h01;
  assign sel_89501 = array_index_89404 == array_index_86800 ? add_89500 : sel_89497;
  assign add_89504 = sel_89501 + 8'h01;
  assign sel_89505 = array_index_89404 == array_index_86806 ? add_89504 : sel_89501;
  assign add_89508 = sel_89505 + 8'h01;
  assign sel_89509 = array_index_89404 == array_index_86812 ? add_89508 : sel_89505;
  assign add_89512 = sel_89509 + 8'h01;
  assign sel_89513 = array_index_89404 == array_index_86818 ? add_89512 : sel_89509;
  assign add_89516 = sel_89513 + 8'h01;
  assign sel_89517 = array_index_89404 == array_index_86824 ? add_89516 : sel_89513;
  assign add_89520 = sel_89517 + 8'h01;
  assign sel_89521 = array_index_89404 == array_index_86830 ? add_89520 : sel_89517;
  assign add_89525 = sel_89521 + 8'h01;
  assign array_index_89526 = set1_unflattened[5'h17];
  assign sel_89527 = array_index_89404 == array_index_86836 ? add_89525 : sel_89521;
  assign add_89530 = sel_89527 + 8'h01;
  assign sel_89531 = array_index_89526 == array_index_86652 ? add_89530 : sel_89527;
  assign add_89534 = sel_89531 + 8'h01;
  assign sel_89535 = array_index_89526 == array_index_86656 ? add_89534 : sel_89531;
  assign add_89538 = sel_89535 + 8'h01;
  assign sel_89539 = array_index_89526 == array_index_86664 ? add_89538 : sel_89535;
  assign add_89542 = sel_89539 + 8'h01;
  assign sel_89543 = array_index_89526 == array_index_86672 ? add_89542 : sel_89539;
  assign add_89546 = sel_89543 + 8'h01;
  assign sel_89547 = array_index_89526 == array_index_86680 ? add_89546 : sel_89543;
  assign add_89550 = sel_89547 + 8'h01;
  assign sel_89551 = array_index_89526 == array_index_86688 ? add_89550 : sel_89547;
  assign add_89554 = sel_89551 + 8'h01;
  assign sel_89555 = array_index_89526 == array_index_86696 ? add_89554 : sel_89551;
  assign add_89558 = sel_89555 + 8'h01;
  assign sel_89559 = array_index_89526 == array_index_86704 ? add_89558 : sel_89555;
  assign add_89562 = sel_89559 + 8'h01;
  assign sel_89563 = array_index_89526 == array_index_86710 ? add_89562 : sel_89559;
  assign add_89566 = sel_89563 + 8'h01;
  assign sel_89567 = array_index_89526 == array_index_86716 ? add_89566 : sel_89563;
  assign add_89570 = sel_89567 + 8'h01;
  assign sel_89571 = array_index_89526 == array_index_86722 ? add_89570 : sel_89567;
  assign add_89574 = sel_89571 + 8'h01;
  assign sel_89575 = array_index_89526 == array_index_86728 ? add_89574 : sel_89571;
  assign add_89578 = sel_89575 + 8'h01;
  assign sel_89579 = array_index_89526 == array_index_86734 ? add_89578 : sel_89575;
  assign add_89582 = sel_89579 + 8'h01;
  assign sel_89583 = array_index_89526 == array_index_86740 ? add_89582 : sel_89579;
  assign add_89586 = sel_89583 + 8'h01;
  assign sel_89587 = array_index_89526 == array_index_86746 ? add_89586 : sel_89583;
  assign add_89590 = sel_89587 + 8'h01;
  assign sel_89591 = array_index_89526 == array_index_86752 ? add_89590 : sel_89587;
  assign add_89594 = sel_89591 + 8'h01;
  assign sel_89595 = array_index_89526 == array_index_86758 ? add_89594 : sel_89591;
  assign add_89598 = sel_89595 + 8'h01;
  assign sel_89599 = array_index_89526 == array_index_86764 ? add_89598 : sel_89595;
  assign add_89602 = sel_89599 + 8'h01;
  assign sel_89603 = array_index_89526 == array_index_86770 ? add_89602 : sel_89599;
  assign add_89606 = sel_89603 + 8'h01;
  assign sel_89607 = array_index_89526 == array_index_86776 ? add_89606 : sel_89603;
  assign add_89610 = sel_89607 + 8'h01;
  assign sel_89611 = array_index_89526 == array_index_86782 ? add_89610 : sel_89607;
  assign add_89614 = sel_89611 + 8'h01;
  assign sel_89615 = array_index_89526 == array_index_86788 ? add_89614 : sel_89611;
  assign add_89618 = sel_89615 + 8'h01;
  assign sel_89619 = array_index_89526 == array_index_86794 ? add_89618 : sel_89615;
  assign add_89622 = sel_89619 + 8'h01;
  assign sel_89623 = array_index_89526 == array_index_86800 ? add_89622 : sel_89619;
  assign add_89626 = sel_89623 + 8'h01;
  assign sel_89627 = array_index_89526 == array_index_86806 ? add_89626 : sel_89623;
  assign add_89630 = sel_89627 + 8'h01;
  assign sel_89631 = array_index_89526 == array_index_86812 ? add_89630 : sel_89627;
  assign add_89634 = sel_89631 + 8'h01;
  assign sel_89635 = array_index_89526 == array_index_86818 ? add_89634 : sel_89631;
  assign add_89638 = sel_89635 + 8'h01;
  assign sel_89639 = array_index_89526 == array_index_86824 ? add_89638 : sel_89635;
  assign add_89642 = sel_89639 + 8'h01;
  assign sel_89643 = array_index_89526 == array_index_86830 ? add_89642 : sel_89639;
  assign add_89647 = sel_89643 + 8'h01;
  assign array_index_89648 = set1_unflattened[5'h18];
  assign sel_89649 = array_index_89526 == array_index_86836 ? add_89647 : sel_89643;
  assign add_89652 = sel_89649 + 8'h01;
  assign sel_89653 = array_index_89648 == array_index_86652 ? add_89652 : sel_89649;
  assign add_89656 = sel_89653 + 8'h01;
  assign sel_89657 = array_index_89648 == array_index_86656 ? add_89656 : sel_89653;
  assign add_89660 = sel_89657 + 8'h01;
  assign sel_89661 = array_index_89648 == array_index_86664 ? add_89660 : sel_89657;
  assign add_89664 = sel_89661 + 8'h01;
  assign sel_89665 = array_index_89648 == array_index_86672 ? add_89664 : sel_89661;
  assign add_89668 = sel_89665 + 8'h01;
  assign sel_89669 = array_index_89648 == array_index_86680 ? add_89668 : sel_89665;
  assign add_89672 = sel_89669 + 8'h01;
  assign sel_89673 = array_index_89648 == array_index_86688 ? add_89672 : sel_89669;
  assign add_89676 = sel_89673 + 8'h01;
  assign sel_89677 = array_index_89648 == array_index_86696 ? add_89676 : sel_89673;
  assign add_89680 = sel_89677 + 8'h01;
  assign sel_89681 = array_index_89648 == array_index_86704 ? add_89680 : sel_89677;
  assign add_89684 = sel_89681 + 8'h01;
  assign sel_89685 = array_index_89648 == array_index_86710 ? add_89684 : sel_89681;
  assign add_89688 = sel_89685 + 8'h01;
  assign sel_89689 = array_index_89648 == array_index_86716 ? add_89688 : sel_89685;
  assign add_89692 = sel_89689 + 8'h01;
  assign sel_89693 = array_index_89648 == array_index_86722 ? add_89692 : sel_89689;
  assign add_89696 = sel_89693 + 8'h01;
  assign sel_89697 = array_index_89648 == array_index_86728 ? add_89696 : sel_89693;
  assign add_89700 = sel_89697 + 8'h01;
  assign sel_89701 = array_index_89648 == array_index_86734 ? add_89700 : sel_89697;
  assign add_89704 = sel_89701 + 8'h01;
  assign sel_89705 = array_index_89648 == array_index_86740 ? add_89704 : sel_89701;
  assign add_89708 = sel_89705 + 8'h01;
  assign sel_89709 = array_index_89648 == array_index_86746 ? add_89708 : sel_89705;
  assign add_89712 = sel_89709 + 8'h01;
  assign sel_89713 = array_index_89648 == array_index_86752 ? add_89712 : sel_89709;
  assign add_89716 = sel_89713 + 8'h01;
  assign sel_89717 = array_index_89648 == array_index_86758 ? add_89716 : sel_89713;
  assign add_89720 = sel_89717 + 8'h01;
  assign sel_89721 = array_index_89648 == array_index_86764 ? add_89720 : sel_89717;
  assign add_89724 = sel_89721 + 8'h01;
  assign sel_89725 = array_index_89648 == array_index_86770 ? add_89724 : sel_89721;
  assign add_89728 = sel_89725 + 8'h01;
  assign sel_89729 = array_index_89648 == array_index_86776 ? add_89728 : sel_89725;
  assign add_89732 = sel_89729 + 8'h01;
  assign sel_89733 = array_index_89648 == array_index_86782 ? add_89732 : sel_89729;
  assign add_89736 = sel_89733 + 8'h01;
  assign sel_89737 = array_index_89648 == array_index_86788 ? add_89736 : sel_89733;
  assign add_89740 = sel_89737 + 8'h01;
  assign sel_89741 = array_index_89648 == array_index_86794 ? add_89740 : sel_89737;
  assign add_89744 = sel_89741 + 8'h01;
  assign sel_89745 = array_index_89648 == array_index_86800 ? add_89744 : sel_89741;
  assign add_89748 = sel_89745 + 8'h01;
  assign sel_89749 = array_index_89648 == array_index_86806 ? add_89748 : sel_89745;
  assign add_89752 = sel_89749 + 8'h01;
  assign sel_89753 = array_index_89648 == array_index_86812 ? add_89752 : sel_89749;
  assign add_89756 = sel_89753 + 8'h01;
  assign sel_89757 = array_index_89648 == array_index_86818 ? add_89756 : sel_89753;
  assign add_89760 = sel_89757 + 8'h01;
  assign sel_89761 = array_index_89648 == array_index_86824 ? add_89760 : sel_89757;
  assign add_89764 = sel_89761 + 8'h01;
  assign sel_89765 = array_index_89648 == array_index_86830 ? add_89764 : sel_89761;
  assign add_89769 = sel_89765 + 8'h01;
  assign array_index_89770 = set1_unflattened[5'h19];
  assign sel_89771 = array_index_89648 == array_index_86836 ? add_89769 : sel_89765;
  assign add_89774 = sel_89771 + 8'h01;
  assign sel_89775 = array_index_89770 == array_index_86652 ? add_89774 : sel_89771;
  assign add_89778 = sel_89775 + 8'h01;
  assign sel_89779 = array_index_89770 == array_index_86656 ? add_89778 : sel_89775;
  assign add_89782 = sel_89779 + 8'h01;
  assign sel_89783 = array_index_89770 == array_index_86664 ? add_89782 : sel_89779;
  assign add_89786 = sel_89783 + 8'h01;
  assign sel_89787 = array_index_89770 == array_index_86672 ? add_89786 : sel_89783;
  assign add_89790 = sel_89787 + 8'h01;
  assign sel_89791 = array_index_89770 == array_index_86680 ? add_89790 : sel_89787;
  assign add_89794 = sel_89791 + 8'h01;
  assign sel_89795 = array_index_89770 == array_index_86688 ? add_89794 : sel_89791;
  assign add_89798 = sel_89795 + 8'h01;
  assign sel_89799 = array_index_89770 == array_index_86696 ? add_89798 : sel_89795;
  assign add_89802 = sel_89799 + 8'h01;
  assign sel_89803 = array_index_89770 == array_index_86704 ? add_89802 : sel_89799;
  assign add_89806 = sel_89803 + 8'h01;
  assign sel_89807 = array_index_89770 == array_index_86710 ? add_89806 : sel_89803;
  assign add_89810 = sel_89807 + 8'h01;
  assign sel_89811 = array_index_89770 == array_index_86716 ? add_89810 : sel_89807;
  assign add_89814 = sel_89811 + 8'h01;
  assign sel_89815 = array_index_89770 == array_index_86722 ? add_89814 : sel_89811;
  assign add_89818 = sel_89815 + 8'h01;
  assign sel_89819 = array_index_89770 == array_index_86728 ? add_89818 : sel_89815;
  assign add_89822 = sel_89819 + 8'h01;
  assign sel_89823 = array_index_89770 == array_index_86734 ? add_89822 : sel_89819;
  assign add_89826 = sel_89823 + 8'h01;
  assign sel_89827 = array_index_89770 == array_index_86740 ? add_89826 : sel_89823;
  assign add_89830 = sel_89827 + 8'h01;
  assign sel_89831 = array_index_89770 == array_index_86746 ? add_89830 : sel_89827;
  assign add_89834 = sel_89831 + 8'h01;
  assign sel_89835 = array_index_89770 == array_index_86752 ? add_89834 : sel_89831;
  assign add_89838 = sel_89835 + 8'h01;
  assign sel_89839 = array_index_89770 == array_index_86758 ? add_89838 : sel_89835;
  assign add_89842 = sel_89839 + 8'h01;
  assign sel_89843 = array_index_89770 == array_index_86764 ? add_89842 : sel_89839;
  assign add_89846 = sel_89843 + 8'h01;
  assign sel_89847 = array_index_89770 == array_index_86770 ? add_89846 : sel_89843;
  assign add_89850 = sel_89847 + 8'h01;
  assign sel_89851 = array_index_89770 == array_index_86776 ? add_89850 : sel_89847;
  assign add_89854 = sel_89851 + 8'h01;
  assign sel_89855 = array_index_89770 == array_index_86782 ? add_89854 : sel_89851;
  assign add_89858 = sel_89855 + 8'h01;
  assign sel_89859 = array_index_89770 == array_index_86788 ? add_89858 : sel_89855;
  assign add_89862 = sel_89859 + 8'h01;
  assign sel_89863 = array_index_89770 == array_index_86794 ? add_89862 : sel_89859;
  assign add_89866 = sel_89863 + 8'h01;
  assign sel_89867 = array_index_89770 == array_index_86800 ? add_89866 : sel_89863;
  assign add_89870 = sel_89867 + 8'h01;
  assign sel_89871 = array_index_89770 == array_index_86806 ? add_89870 : sel_89867;
  assign add_89874 = sel_89871 + 8'h01;
  assign sel_89875 = array_index_89770 == array_index_86812 ? add_89874 : sel_89871;
  assign add_89878 = sel_89875 + 8'h01;
  assign sel_89879 = array_index_89770 == array_index_86818 ? add_89878 : sel_89875;
  assign add_89882 = sel_89879 + 8'h01;
  assign sel_89883 = array_index_89770 == array_index_86824 ? add_89882 : sel_89879;
  assign add_89886 = sel_89883 + 8'h01;
  assign sel_89887 = array_index_89770 == array_index_86830 ? add_89886 : sel_89883;
  assign add_89891 = sel_89887 + 8'h01;
  assign array_index_89892 = set1_unflattened[5'h1a];
  assign sel_89893 = array_index_89770 == array_index_86836 ? add_89891 : sel_89887;
  assign add_89896 = sel_89893 + 8'h01;
  assign sel_89897 = array_index_89892 == array_index_86652 ? add_89896 : sel_89893;
  assign add_89900 = sel_89897 + 8'h01;
  assign sel_89901 = array_index_89892 == array_index_86656 ? add_89900 : sel_89897;
  assign add_89904 = sel_89901 + 8'h01;
  assign sel_89905 = array_index_89892 == array_index_86664 ? add_89904 : sel_89901;
  assign add_89908 = sel_89905 + 8'h01;
  assign sel_89909 = array_index_89892 == array_index_86672 ? add_89908 : sel_89905;
  assign add_89912 = sel_89909 + 8'h01;
  assign sel_89913 = array_index_89892 == array_index_86680 ? add_89912 : sel_89909;
  assign add_89916 = sel_89913 + 8'h01;
  assign sel_89917 = array_index_89892 == array_index_86688 ? add_89916 : sel_89913;
  assign add_89920 = sel_89917 + 8'h01;
  assign sel_89921 = array_index_89892 == array_index_86696 ? add_89920 : sel_89917;
  assign add_89924 = sel_89921 + 8'h01;
  assign sel_89925 = array_index_89892 == array_index_86704 ? add_89924 : sel_89921;
  assign add_89928 = sel_89925 + 8'h01;
  assign sel_89929 = array_index_89892 == array_index_86710 ? add_89928 : sel_89925;
  assign add_89932 = sel_89929 + 8'h01;
  assign sel_89933 = array_index_89892 == array_index_86716 ? add_89932 : sel_89929;
  assign add_89936 = sel_89933 + 8'h01;
  assign sel_89937 = array_index_89892 == array_index_86722 ? add_89936 : sel_89933;
  assign add_89940 = sel_89937 + 8'h01;
  assign sel_89941 = array_index_89892 == array_index_86728 ? add_89940 : sel_89937;
  assign add_89944 = sel_89941 + 8'h01;
  assign sel_89945 = array_index_89892 == array_index_86734 ? add_89944 : sel_89941;
  assign add_89948 = sel_89945 + 8'h01;
  assign sel_89949 = array_index_89892 == array_index_86740 ? add_89948 : sel_89945;
  assign add_89952 = sel_89949 + 8'h01;
  assign sel_89953 = array_index_89892 == array_index_86746 ? add_89952 : sel_89949;
  assign add_89956 = sel_89953 + 8'h01;
  assign sel_89957 = array_index_89892 == array_index_86752 ? add_89956 : sel_89953;
  assign add_89960 = sel_89957 + 8'h01;
  assign sel_89961 = array_index_89892 == array_index_86758 ? add_89960 : sel_89957;
  assign add_89964 = sel_89961 + 8'h01;
  assign sel_89965 = array_index_89892 == array_index_86764 ? add_89964 : sel_89961;
  assign add_89968 = sel_89965 + 8'h01;
  assign sel_89969 = array_index_89892 == array_index_86770 ? add_89968 : sel_89965;
  assign add_89972 = sel_89969 + 8'h01;
  assign sel_89973 = array_index_89892 == array_index_86776 ? add_89972 : sel_89969;
  assign add_89976 = sel_89973 + 8'h01;
  assign sel_89977 = array_index_89892 == array_index_86782 ? add_89976 : sel_89973;
  assign add_89980 = sel_89977 + 8'h01;
  assign sel_89981 = array_index_89892 == array_index_86788 ? add_89980 : sel_89977;
  assign add_89984 = sel_89981 + 8'h01;
  assign sel_89985 = array_index_89892 == array_index_86794 ? add_89984 : sel_89981;
  assign add_89988 = sel_89985 + 8'h01;
  assign sel_89989 = array_index_89892 == array_index_86800 ? add_89988 : sel_89985;
  assign add_89992 = sel_89989 + 8'h01;
  assign sel_89993 = array_index_89892 == array_index_86806 ? add_89992 : sel_89989;
  assign add_89996 = sel_89993 + 8'h01;
  assign sel_89997 = array_index_89892 == array_index_86812 ? add_89996 : sel_89993;
  assign add_90000 = sel_89997 + 8'h01;
  assign sel_90001 = array_index_89892 == array_index_86818 ? add_90000 : sel_89997;
  assign add_90004 = sel_90001 + 8'h01;
  assign sel_90005 = array_index_89892 == array_index_86824 ? add_90004 : sel_90001;
  assign add_90008 = sel_90005 + 8'h01;
  assign sel_90009 = array_index_89892 == array_index_86830 ? add_90008 : sel_90005;
  assign add_90013 = sel_90009 + 8'h01;
  assign array_index_90014 = set1_unflattened[5'h1b];
  assign sel_90015 = array_index_89892 == array_index_86836 ? add_90013 : sel_90009;
  assign add_90018 = sel_90015 + 8'h01;
  assign sel_90019 = array_index_90014 == array_index_86652 ? add_90018 : sel_90015;
  assign add_90022 = sel_90019 + 8'h01;
  assign sel_90023 = array_index_90014 == array_index_86656 ? add_90022 : sel_90019;
  assign add_90026 = sel_90023 + 8'h01;
  assign sel_90027 = array_index_90014 == array_index_86664 ? add_90026 : sel_90023;
  assign add_90030 = sel_90027 + 8'h01;
  assign sel_90031 = array_index_90014 == array_index_86672 ? add_90030 : sel_90027;
  assign add_90034 = sel_90031 + 8'h01;
  assign sel_90035 = array_index_90014 == array_index_86680 ? add_90034 : sel_90031;
  assign add_90038 = sel_90035 + 8'h01;
  assign sel_90039 = array_index_90014 == array_index_86688 ? add_90038 : sel_90035;
  assign add_90042 = sel_90039 + 8'h01;
  assign sel_90043 = array_index_90014 == array_index_86696 ? add_90042 : sel_90039;
  assign add_90046 = sel_90043 + 8'h01;
  assign sel_90047 = array_index_90014 == array_index_86704 ? add_90046 : sel_90043;
  assign add_90050 = sel_90047 + 8'h01;
  assign sel_90051 = array_index_90014 == array_index_86710 ? add_90050 : sel_90047;
  assign add_90054 = sel_90051 + 8'h01;
  assign sel_90055 = array_index_90014 == array_index_86716 ? add_90054 : sel_90051;
  assign add_90058 = sel_90055 + 8'h01;
  assign sel_90059 = array_index_90014 == array_index_86722 ? add_90058 : sel_90055;
  assign add_90062 = sel_90059 + 8'h01;
  assign sel_90063 = array_index_90014 == array_index_86728 ? add_90062 : sel_90059;
  assign add_90066 = sel_90063 + 8'h01;
  assign sel_90067 = array_index_90014 == array_index_86734 ? add_90066 : sel_90063;
  assign add_90070 = sel_90067 + 8'h01;
  assign sel_90071 = array_index_90014 == array_index_86740 ? add_90070 : sel_90067;
  assign add_90074 = sel_90071 + 8'h01;
  assign sel_90075 = array_index_90014 == array_index_86746 ? add_90074 : sel_90071;
  assign add_90078 = sel_90075 + 8'h01;
  assign sel_90079 = array_index_90014 == array_index_86752 ? add_90078 : sel_90075;
  assign add_90082 = sel_90079 + 8'h01;
  assign sel_90083 = array_index_90014 == array_index_86758 ? add_90082 : sel_90079;
  assign add_90086 = sel_90083 + 8'h01;
  assign sel_90087 = array_index_90014 == array_index_86764 ? add_90086 : sel_90083;
  assign add_90090 = sel_90087 + 8'h01;
  assign sel_90091 = array_index_90014 == array_index_86770 ? add_90090 : sel_90087;
  assign add_90094 = sel_90091 + 8'h01;
  assign sel_90095 = array_index_90014 == array_index_86776 ? add_90094 : sel_90091;
  assign add_90098 = sel_90095 + 8'h01;
  assign sel_90099 = array_index_90014 == array_index_86782 ? add_90098 : sel_90095;
  assign add_90102 = sel_90099 + 8'h01;
  assign sel_90103 = array_index_90014 == array_index_86788 ? add_90102 : sel_90099;
  assign add_90106 = sel_90103 + 8'h01;
  assign sel_90107 = array_index_90014 == array_index_86794 ? add_90106 : sel_90103;
  assign add_90110 = sel_90107 + 8'h01;
  assign sel_90111 = array_index_90014 == array_index_86800 ? add_90110 : sel_90107;
  assign add_90114 = sel_90111 + 8'h01;
  assign sel_90115 = array_index_90014 == array_index_86806 ? add_90114 : sel_90111;
  assign add_90118 = sel_90115 + 8'h01;
  assign sel_90119 = array_index_90014 == array_index_86812 ? add_90118 : sel_90115;
  assign add_90122 = sel_90119 + 8'h01;
  assign sel_90123 = array_index_90014 == array_index_86818 ? add_90122 : sel_90119;
  assign add_90126 = sel_90123 + 8'h01;
  assign sel_90127 = array_index_90014 == array_index_86824 ? add_90126 : sel_90123;
  assign add_90130 = sel_90127 + 8'h01;
  assign sel_90131 = array_index_90014 == array_index_86830 ? add_90130 : sel_90127;
  assign add_90135 = sel_90131 + 8'h01;
  assign array_index_90136 = set1_unflattened[5'h1c];
  assign sel_90137 = array_index_90014 == array_index_86836 ? add_90135 : sel_90131;
  assign add_90140 = sel_90137 + 8'h01;
  assign sel_90141 = array_index_90136 == array_index_86652 ? add_90140 : sel_90137;
  assign add_90144 = sel_90141 + 8'h01;
  assign sel_90145 = array_index_90136 == array_index_86656 ? add_90144 : sel_90141;
  assign add_90148 = sel_90145 + 8'h01;
  assign sel_90149 = array_index_90136 == array_index_86664 ? add_90148 : sel_90145;
  assign add_90152 = sel_90149 + 8'h01;
  assign sel_90153 = array_index_90136 == array_index_86672 ? add_90152 : sel_90149;
  assign add_90156 = sel_90153 + 8'h01;
  assign sel_90157 = array_index_90136 == array_index_86680 ? add_90156 : sel_90153;
  assign add_90160 = sel_90157 + 8'h01;
  assign sel_90161 = array_index_90136 == array_index_86688 ? add_90160 : sel_90157;
  assign add_90164 = sel_90161 + 8'h01;
  assign sel_90165 = array_index_90136 == array_index_86696 ? add_90164 : sel_90161;
  assign add_90168 = sel_90165 + 8'h01;
  assign sel_90169 = array_index_90136 == array_index_86704 ? add_90168 : sel_90165;
  assign add_90172 = sel_90169 + 8'h01;
  assign sel_90173 = array_index_90136 == array_index_86710 ? add_90172 : sel_90169;
  assign add_90176 = sel_90173 + 8'h01;
  assign sel_90177 = array_index_90136 == array_index_86716 ? add_90176 : sel_90173;
  assign add_90180 = sel_90177 + 8'h01;
  assign sel_90181 = array_index_90136 == array_index_86722 ? add_90180 : sel_90177;
  assign add_90184 = sel_90181 + 8'h01;
  assign sel_90185 = array_index_90136 == array_index_86728 ? add_90184 : sel_90181;
  assign add_90188 = sel_90185 + 8'h01;
  assign sel_90189 = array_index_90136 == array_index_86734 ? add_90188 : sel_90185;
  assign add_90192 = sel_90189 + 8'h01;
  assign sel_90193 = array_index_90136 == array_index_86740 ? add_90192 : sel_90189;
  assign add_90196 = sel_90193 + 8'h01;
  assign sel_90197 = array_index_90136 == array_index_86746 ? add_90196 : sel_90193;
  assign add_90200 = sel_90197 + 8'h01;
  assign sel_90201 = array_index_90136 == array_index_86752 ? add_90200 : sel_90197;
  assign add_90204 = sel_90201 + 8'h01;
  assign sel_90205 = array_index_90136 == array_index_86758 ? add_90204 : sel_90201;
  assign add_90208 = sel_90205 + 8'h01;
  assign sel_90209 = array_index_90136 == array_index_86764 ? add_90208 : sel_90205;
  assign add_90212 = sel_90209 + 8'h01;
  assign sel_90213 = array_index_90136 == array_index_86770 ? add_90212 : sel_90209;
  assign add_90216 = sel_90213 + 8'h01;
  assign sel_90217 = array_index_90136 == array_index_86776 ? add_90216 : sel_90213;
  assign add_90220 = sel_90217 + 8'h01;
  assign sel_90221 = array_index_90136 == array_index_86782 ? add_90220 : sel_90217;
  assign add_90224 = sel_90221 + 8'h01;
  assign sel_90225 = array_index_90136 == array_index_86788 ? add_90224 : sel_90221;
  assign add_90228 = sel_90225 + 8'h01;
  assign sel_90229 = array_index_90136 == array_index_86794 ? add_90228 : sel_90225;
  assign add_90232 = sel_90229 + 8'h01;
  assign sel_90233 = array_index_90136 == array_index_86800 ? add_90232 : sel_90229;
  assign add_90236 = sel_90233 + 8'h01;
  assign sel_90237 = array_index_90136 == array_index_86806 ? add_90236 : sel_90233;
  assign add_90240 = sel_90237 + 8'h01;
  assign sel_90241 = array_index_90136 == array_index_86812 ? add_90240 : sel_90237;
  assign add_90244 = sel_90241 + 8'h01;
  assign sel_90245 = array_index_90136 == array_index_86818 ? add_90244 : sel_90241;
  assign add_90248 = sel_90245 + 8'h01;
  assign sel_90249 = array_index_90136 == array_index_86824 ? add_90248 : sel_90245;
  assign add_90252 = sel_90249 + 8'h01;
  assign sel_90253 = array_index_90136 == array_index_86830 ? add_90252 : sel_90249;
  assign add_90257 = sel_90253 + 8'h01;
  assign array_index_90258 = set1_unflattened[5'h1d];
  assign sel_90259 = array_index_90136 == array_index_86836 ? add_90257 : sel_90253;
  assign add_90262 = sel_90259 + 8'h01;
  assign sel_90263 = array_index_90258 == array_index_86652 ? add_90262 : sel_90259;
  assign add_90266 = sel_90263 + 8'h01;
  assign sel_90267 = array_index_90258 == array_index_86656 ? add_90266 : sel_90263;
  assign add_90270 = sel_90267 + 8'h01;
  assign sel_90271 = array_index_90258 == array_index_86664 ? add_90270 : sel_90267;
  assign add_90274 = sel_90271 + 8'h01;
  assign sel_90275 = array_index_90258 == array_index_86672 ? add_90274 : sel_90271;
  assign add_90278 = sel_90275 + 8'h01;
  assign sel_90279 = array_index_90258 == array_index_86680 ? add_90278 : sel_90275;
  assign add_90282 = sel_90279 + 8'h01;
  assign sel_90283 = array_index_90258 == array_index_86688 ? add_90282 : sel_90279;
  assign add_90286 = sel_90283 + 8'h01;
  assign sel_90287 = array_index_90258 == array_index_86696 ? add_90286 : sel_90283;
  assign add_90290 = sel_90287 + 8'h01;
  assign sel_90291 = array_index_90258 == array_index_86704 ? add_90290 : sel_90287;
  assign add_90294 = sel_90291 + 8'h01;
  assign sel_90295 = array_index_90258 == array_index_86710 ? add_90294 : sel_90291;
  assign add_90298 = sel_90295 + 8'h01;
  assign sel_90299 = array_index_90258 == array_index_86716 ? add_90298 : sel_90295;
  assign add_90302 = sel_90299 + 8'h01;
  assign sel_90303 = array_index_90258 == array_index_86722 ? add_90302 : sel_90299;
  assign add_90306 = sel_90303 + 8'h01;
  assign sel_90307 = array_index_90258 == array_index_86728 ? add_90306 : sel_90303;
  assign add_90310 = sel_90307 + 8'h01;
  assign sel_90311 = array_index_90258 == array_index_86734 ? add_90310 : sel_90307;
  assign add_90314 = sel_90311 + 8'h01;
  assign sel_90315 = array_index_90258 == array_index_86740 ? add_90314 : sel_90311;
  assign add_90318 = sel_90315 + 8'h01;
  assign sel_90319 = array_index_90258 == array_index_86746 ? add_90318 : sel_90315;
  assign add_90322 = sel_90319 + 8'h01;
  assign sel_90323 = array_index_90258 == array_index_86752 ? add_90322 : sel_90319;
  assign add_90326 = sel_90323 + 8'h01;
  assign sel_90327 = array_index_90258 == array_index_86758 ? add_90326 : sel_90323;
  assign add_90330 = sel_90327 + 8'h01;
  assign sel_90331 = array_index_90258 == array_index_86764 ? add_90330 : sel_90327;
  assign add_90334 = sel_90331 + 8'h01;
  assign sel_90335 = array_index_90258 == array_index_86770 ? add_90334 : sel_90331;
  assign add_90338 = sel_90335 + 8'h01;
  assign sel_90339 = array_index_90258 == array_index_86776 ? add_90338 : sel_90335;
  assign add_90342 = sel_90339 + 8'h01;
  assign sel_90343 = array_index_90258 == array_index_86782 ? add_90342 : sel_90339;
  assign add_90346 = sel_90343 + 8'h01;
  assign sel_90347 = array_index_90258 == array_index_86788 ? add_90346 : sel_90343;
  assign add_90350 = sel_90347 + 8'h01;
  assign sel_90351 = array_index_90258 == array_index_86794 ? add_90350 : sel_90347;
  assign add_90354 = sel_90351 + 8'h01;
  assign sel_90355 = array_index_90258 == array_index_86800 ? add_90354 : sel_90351;
  assign add_90358 = sel_90355 + 8'h01;
  assign sel_90359 = array_index_90258 == array_index_86806 ? add_90358 : sel_90355;
  assign add_90362 = sel_90359 + 8'h01;
  assign sel_90363 = array_index_90258 == array_index_86812 ? add_90362 : sel_90359;
  assign add_90366 = sel_90363 + 8'h01;
  assign sel_90367 = array_index_90258 == array_index_86818 ? add_90366 : sel_90363;
  assign add_90370 = sel_90367 + 8'h01;
  assign sel_90371 = array_index_90258 == array_index_86824 ? add_90370 : sel_90367;
  assign add_90374 = sel_90371 + 8'h01;
  assign sel_90375 = array_index_90258 == array_index_86830 ? add_90374 : sel_90371;
  assign add_90378 = sel_90375 + 8'h01;
  assign out = {array_index_90258 == array_index_86836 ? add_90378 : sel_90375, {set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
