module min_hash(
  input wire [159:0] set1,
  input wire [159:0] set2,
  output wire [335:0] out
);
  wire [15:0] set1_unflattened[10];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  wire [15:0] set2_unflattened[10];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  wire [15:0] array_index_18141;
  wire [15:0] array_index_18142;
  wire [11:0] add_18149;
  wire [11:0] add_18152;
  wire [15:0] array_index_18157;
  wire [15:0] array_index_18160;
  wire [10:0] add_18164;
  wire [10:0] add_18167;
  wire [11:0] add_18183;
  wire [11:0] sel_18185;
  wire [11:0] add_18188;
  wire [11:0] sel_18190;
  wire [15:0] array_index_18205;
  wire [15:0] array_index_18208;
  wire [8:0] add_18212;
  wire [8:0] add_18215;
  wire [10:0] add_18218;
  wire [11:0] sel_18221;
  wire [10:0] add_18223;
  wire [11:0] sel_18226;
  wire [11:0] add_18243;
  wire [11:0] sel_18245;
  wire [11:0] add_18248;
  wire [11:0] sel_18250;
  wire [15:0] array_index_18271;
  wire [15:0] array_index_18274;
  wire [10:0] add_18278;
  wire [10:0] add_18280;
  wire [8:0] add_18282;
  wire [11:0] sel_18285;
  wire [8:0] add_18287;
  wire [11:0] sel_18290;
  wire [10:0] add_18292;
  wire [11:0] sel_18295;
  wire [10:0] add_18297;
  wire [11:0] sel_18300;
  wire [11:0] add_18321;
  wire [11:0] sel_18323;
  wire [11:0] add_18326;
  wire [11:0] sel_18328;
  wire [15:0] array_index_18355;
  wire [15:0] array_index_18358;
  wire [10:0] add_18362;
  wire [10:0] add_18364;
  wire [10:0] add_18366;
  wire [11:0] sel_18368;
  wire [10:0] add_18370;
  wire [11:0] sel_18372;
  wire [8:0] add_18374;
  wire [11:0] sel_18377;
  wire [8:0] add_18379;
  wire [11:0] sel_18382;
  wire [10:0] add_18384;
  wire [11:0] sel_18387;
  wire [10:0] add_18389;
  wire [11:0] sel_18392;
  wire [11:0] add_18417;
  wire [11:0] sel_18419;
  wire [11:0] add_18422;
  wire [11:0] sel_18424;
  wire [15:0] array_index_18455;
  wire [15:0] array_index_18458;
  wire [10:0] add_18462;
  wire [11:0] sel_18464;
  wire [10:0] add_18466;
  wire [11:0] sel_18468;
  wire [10:0] add_18470;
  wire [11:0] sel_18472;
  wire [10:0] add_18474;
  wire [11:0] sel_18476;
  wire [8:0] add_18478;
  wire [11:0] sel_18481;
  wire [8:0] add_18483;
  wire [11:0] sel_18486;
  wire [10:0] add_18488;
  wire [11:0] sel_18491;
  wire [10:0] add_18493;
  wire [11:0] sel_18496;
  wire [11:0] add_18521;
  wire [11:0] sel_18523;
  wire [11:0] add_18526;
  wire [11:0] sel_18528;
  wire [15:0] array_index_18557;
  wire [15:0] array_index_18560;
  wire [10:0] add_18564;
  wire [11:0] sel_18566;
  wire [10:0] add_18568;
  wire [11:0] sel_18570;
  wire [10:0] add_18572;
  wire [11:0] sel_18574;
  wire [10:0] add_18576;
  wire [11:0] sel_18578;
  wire [8:0] add_18580;
  wire [11:0] sel_18583;
  wire [8:0] add_18585;
  wire [11:0] sel_18588;
  wire [10:0] add_18590;
  wire [11:0] sel_18593;
  wire [10:0] add_18595;
  wire [11:0] sel_18598;
  wire [11:0] add_18623;
  wire [11:0] sel_18625;
  wire [11:0] add_18628;
  wire [11:0] sel_18630;
  wire [15:0] array_index_18659;
  wire [15:0] array_index_18662;
  wire [10:0] add_18666;
  wire [11:0] sel_18668;
  wire [10:0] add_18670;
  wire [11:0] sel_18672;
  wire [10:0] add_18674;
  wire [11:0] sel_18676;
  wire [10:0] add_18678;
  wire [11:0] sel_18680;
  wire [8:0] add_18682;
  wire [11:0] sel_18685;
  wire [8:0] add_18687;
  wire [11:0] sel_18690;
  wire [10:0] add_18692;
  wire [11:0] sel_18695;
  wire [10:0] add_18697;
  wire [11:0] sel_18700;
  wire [11:0] add_18725;
  wire [11:0] sel_18727;
  wire [11:0] add_18730;
  wire [11:0] sel_18732;
  wire [15:0] array_index_18761;
  wire [15:0] array_index_18764;
  wire [10:0] add_18768;
  wire [11:0] sel_18770;
  wire [10:0] add_18772;
  wire [11:0] sel_18774;
  wire [10:0] add_18776;
  wire [11:0] sel_18778;
  wire [10:0] add_18780;
  wire [11:0] sel_18782;
  wire [8:0] add_18784;
  wire [11:0] sel_18787;
  wire [8:0] add_18789;
  wire [11:0] sel_18792;
  wire [10:0] add_18794;
  wire [11:0] sel_18797;
  wire [10:0] add_18799;
  wire [11:0] sel_18802;
  wire [11:0] add_18827;
  wire [11:0] sel_18829;
  wire [11:0] add_18832;
  wire [11:0] sel_18834;
  wire [15:0] array_index_18863;
  wire [15:0] array_index_18866;
  wire [10:0] add_18870;
  wire [11:0] sel_18872;
  wire [10:0] add_18874;
  wire [11:0] sel_18876;
  wire [10:0] add_18878;
  wire [11:0] sel_18880;
  wire [10:0] add_18882;
  wire [11:0] sel_18884;
  wire [8:0] add_18886;
  wire [11:0] sel_18889;
  wire [8:0] add_18891;
  wire [11:0] sel_18894;
  wire [10:0] add_18896;
  wire [11:0] sel_18899;
  wire [10:0] add_18901;
  wire [11:0] sel_18904;
  wire [11:0] add_18928;
  wire [11:0] sel_18930;
  wire [11:0] add_18932;
  wire [11:0] sel_18934;
  wire [10:0] add_18968;
  wire [11:0] sel_18970;
  wire [10:0] add_18972;
  wire [11:0] sel_18974;
  wire [10:0] add_18976;
  wire [11:0] sel_18978;
  wire [10:0] add_18980;
  wire [11:0] sel_18982;
  wire [8:0] add_18984;
  wire [11:0] sel_18987;
  wire [8:0] add_18989;
  wire [11:0] sel_18992;
  wire [10:0] add_18994;
  wire [11:0] sel_18997;
  wire [10:0] add_18999;
  wire [11:0] sel_19002;
  wire [10:0] add_19050;
  wire [11:0] sel_19052;
  wire [10:0] add_19054;
  wire [11:0] sel_19056;
  wire [10:0] add_19058;
  wire [11:0] sel_19060;
  wire [10:0] add_19062;
  wire [11:0] sel_19064;
  wire [8:0] add_19066;
  wire [11:0] sel_19069;
  wire [8:0] add_19071;
  wire [11:0] sel_19074;
  wire [1:0] concat_19077;
  wire [1:0] add_19092;
  wire [10:0] add_19112;
  wire [11:0] sel_19114;
  wire [10:0] add_19116;
  wire [11:0] sel_19118;
  wire [10:0] add_19120;
  wire [11:0] sel_19122;
  wire [10:0] add_19124;
  wire [11:0] sel_19126;
  wire [2:0] concat_19129;
  wire [2:0] add_19140;
  wire [10:0] add_19154;
  wire [11:0] sel_19156;
  wire [10:0] add_19158;
  wire [11:0] sel_19160;
  wire [3:0] concat_19163;
  wire [3:0] add_19170;
  wire [4:0] concat_19179;
  wire [4:0] add_19182;
  assign array_index_18141 = set1_unflattened[4'h0];
  assign array_index_18142 = set2_unflattened[4'h0];
  assign add_18149 = array_index_18141[11:0] + 12'h247;
  assign add_18152 = array_index_18142[11:0] + 12'h247;
  assign array_index_18157 = set1_unflattened[4'h1];
  assign array_index_18160 = set2_unflattened[4'h1];
  assign add_18164 = array_index_18141[11:1] + 11'h247;
  assign add_18167 = array_index_18142[11:1] + 11'h247;
  assign add_18183 = array_index_18157[11:0] + 12'h247;
  assign sel_18185 = $signed({1'h0, add_18149}) < $signed(13'h0fff) ? add_18149 : 12'hfff;
  assign add_18188 = array_index_18160[11:0] + 12'h247;
  assign sel_18190 = $signed({1'h0, add_18152}) < $signed(13'h0fff) ? add_18152 : 12'hfff;
  assign array_index_18205 = set1_unflattened[4'h2];
  assign array_index_18208 = set2_unflattened[4'h2];
  assign add_18212 = array_index_18141[11:3] + 9'h0bd;
  assign add_18215 = array_index_18142[11:3] + 9'h0bd;
  assign add_18218 = array_index_18157[11:1] + 11'h247;
  assign sel_18221 = $signed({1'h0, add_18164, array_index_18141[0]}) < $signed(13'h0fff) ? {add_18164, array_index_18141[0]} : 12'hfff;
  assign add_18223 = array_index_18160[11:1] + 11'h247;
  assign sel_18226 = $signed({1'h0, add_18167, array_index_18142[0]}) < $signed(13'h0fff) ? {add_18167, array_index_18142[0]} : 12'hfff;
  assign add_18243 = array_index_18205[11:0] + 12'h247;
  assign sel_18245 = $signed({1'h0, add_18183}) < $signed({1'h0, sel_18185}) ? add_18183 : sel_18185;
  assign add_18248 = array_index_18208[11:0] + 12'h247;
  assign sel_18250 = $signed({1'h0, add_18188}) < $signed({1'h0, sel_18190}) ? add_18188 : sel_18190;
  assign array_index_18271 = set1_unflattened[4'h3];
  assign array_index_18274 = set2_unflattened[4'h3];
  assign add_18278 = array_index_18141[11:1] + 11'h347;
  assign add_18280 = array_index_18142[11:1] + 11'h347;
  assign add_18282 = array_index_18157[11:3] + 9'h0bd;
  assign sel_18285 = $signed({1'h0, add_18212, array_index_18141[2:0]}) < $signed(13'h0fff) ? {add_18212, array_index_18141[2:0]} : 12'hfff;
  assign add_18287 = array_index_18160[11:3] + 9'h0bd;
  assign sel_18290 = $signed({1'h0, add_18215, array_index_18142[2:0]}) < $signed(13'h0fff) ? {add_18215, array_index_18142[2:0]} : 12'hfff;
  assign add_18292 = array_index_18205[11:1] + 11'h247;
  assign sel_18295 = $signed({1'h0, add_18218, array_index_18157[0]}) < $signed({1'h0, sel_18221}) ? {add_18218, array_index_18157[0]} : sel_18221;
  assign add_18297 = array_index_18208[11:1] + 11'h247;
  assign sel_18300 = $signed({1'h0, add_18223, array_index_18160[0]}) < $signed({1'h0, sel_18226}) ? {add_18223, array_index_18160[0]} : sel_18226;
  assign add_18321 = array_index_18271[11:0] + 12'h247;
  assign sel_18323 = $signed({1'h0, add_18243}) < $signed({1'h0, sel_18245}) ? add_18243 : sel_18245;
  assign add_18326 = array_index_18274[11:0] + 12'h247;
  assign sel_18328 = $signed({1'h0, add_18248}) < $signed({1'h0, sel_18250}) ? add_18248 : sel_18250;
  assign array_index_18355 = set1_unflattened[4'h4];
  assign array_index_18358 = set2_unflattened[4'h4];
  assign add_18362 = array_index_18141[11:1] + 11'h79d;
  assign add_18364 = array_index_18142[11:1] + 11'h79d;
  assign add_18366 = array_index_18157[11:1] + 11'h347;
  assign sel_18368 = $signed({1'h0, add_18278, array_index_18141[0]}) < $signed(13'h0fff) ? {add_18278, array_index_18141[0]} : 12'hfff;
  assign add_18370 = array_index_18160[11:1] + 11'h347;
  assign sel_18372 = $signed({1'h0, add_18280, array_index_18142[0]}) < $signed(13'h0fff) ? {add_18280, array_index_18142[0]} : 12'hfff;
  assign add_18374 = array_index_18205[11:3] + 9'h0bd;
  assign sel_18377 = $signed({1'h0, add_18282, array_index_18157[2:0]}) < $signed({1'h0, sel_18285}) ? {add_18282, array_index_18157[2:0]} : sel_18285;
  assign add_18379 = array_index_18208[11:3] + 9'h0bd;
  assign sel_18382 = $signed({1'h0, add_18287, array_index_18160[2:0]}) < $signed({1'h0, sel_18290}) ? {add_18287, array_index_18160[2:0]} : sel_18290;
  assign add_18384 = array_index_18271[11:1] + 11'h247;
  assign sel_18387 = $signed({1'h0, add_18292, array_index_18205[0]}) < $signed({1'h0, sel_18295}) ? {add_18292, array_index_18205[0]} : sel_18295;
  assign add_18389 = array_index_18274[11:1] + 11'h247;
  assign sel_18392 = $signed({1'h0, add_18297, array_index_18208[0]}) < $signed({1'h0, sel_18300}) ? {add_18297, array_index_18208[0]} : sel_18300;
  assign add_18417 = array_index_18355[11:0] + 12'h247;
  assign sel_18419 = $signed({1'h0, add_18321}) < $signed({1'h0, sel_18323}) ? add_18321 : sel_18323;
  assign add_18422 = array_index_18358[11:0] + 12'h247;
  assign sel_18424 = $signed({1'h0, add_18326}) < $signed({1'h0, sel_18328}) ? add_18326 : sel_18328;
  assign array_index_18455 = set1_unflattened[4'h5];
  assign array_index_18458 = set2_unflattened[4'h5];
  assign add_18462 = array_index_18157[11:1] + 11'h79d;
  assign sel_18464 = $signed({1'h0, add_18362, array_index_18141[0]}) < $signed(13'h0fff) ? {add_18362, array_index_18141[0]} : 12'hfff;
  assign add_18466 = array_index_18160[11:1] + 11'h79d;
  assign sel_18468 = $signed({1'h0, add_18364, array_index_18142[0]}) < $signed(13'h0fff) ? {add_18364, array_index_18142[0]} : 12'hfff;
  assign add_18470 = array_index_18205[11:1] + 11'h347;
  assign sel_18472 = $signed({1'h0, add_18366, array_index_18157[0]}) < $signed({1'h0, sel_18368}) ? {add_18366, array_index_18157[0]} : sel_18368;
  assign add_18474 = array_index_18208[11:1] + 11'h347;
  assign sel_18476 = $signed({1'h0, add_18370, array_index_18160[0]}) < $signed({1'h0, sel_18372}) ? {add_18370, array_index_18160[0]} : sel_18372;
  assign add_18478 = array_index_18271[11:3] + 9'h0bd;
  assign sel_18481 = $signed({1'h0, add_18374, array_index_18205[2:0]}) < $signed({1'h0, sel_18377}) ? {add_18374, array_index_18205[2:0]} : sel_18377;
  assign add_18483 = array_index_18274[11:3] + 9'h0bd;
  assign sel_18486 = $signed({1'h0, add_18379, array_index_18208[2:0]}) < $signed({1'h0, sel_18382}) ? {add_18379, array_index_18208[2:0]} : sel_18382;
  assign add_18488 = array_index_18355[11:1] + 11'h247;
  assign sel_18491 = $signed({1'h0, add_18384, array_index_18271[0]}) < $signed({1'h0, sel_18387}) ? {add_18384, array_index_18271[0]} : sel_18387;
  assign add_18493 = array_index_18358[11:1] + 11'h247;
  assign sel_18496 = $signed({1'h0, add_18389, array_index_18274[0]}) < $signed({1'h0, sel_18392}) ? {add_18389, array_index_18274[0]} : sel_18392;
  assign add_18521 = array_index_18455[11:0] + 12'h247;
  assign sel_18523 = $signed({1'h0, add_18417}) < $signed({1'h0, sel_18419}) ? add_18417 : sel_18419;
  assign add_18526 = array_index_18458[11:0] + 12'h247;
  assign sel_18528 = $signed({1'h0, add_18422}) < $signed({1'h0, sel_18424}) ? add_18422 : sel_18424;
  assign array_index_18557 = set1_unflattened[4'h6];
  assign array_index_18560 = set2_unflattened[4'h6];
  assign add_18564 = array_index_18205[11:1] + 11'h79d;
  assign sel_18566 = $signed({1'h0, add_18462, array_index_18157[0]}) < $signed({1'h0, sel_18464}) ? {add_18462, array_index_18157[0]} : sel_18464;
  assign add_18568 = array_index_18208[11:1] + 11'h79d;
  assign sel_18570 = $signed({1'h0, add_18466, array_index_18160[0]}) < $signed({1'h0, sel_18468}) ? {add_18466, array_index_18160[0]} : sel_18468;
  assign add_18572 = array_index_18271[11:1] + 11'h347;
  assign sel_18574 = $signed({1'h0, add_18470, array_index_18205[0]}) < $signed({1'h0, sel_18472}) ? {add_18470, array_index_18205[0]} : sel_18472;
  assign add_18576 = array_index_18274[11:1] + 11'h347;
  assign sel_18578 = $signed({1'h0, add_18474, array_index_18208[0]}) < $signed({1'h0, sel_18476}) ? {add_18474, array_index_18208[0]} : sel_18476;
  assign add_18580 = array_index_18355[11:3] + 9'h0bd;
  assign sel_18583 = $signed({1'h0, add_18478, array_index_18271[2:0]}) < $signed({1'h0, sel_18481}) ? {add_18478, array_index_18271[2:0]} : sel_18481;
  assign add_18585 = array_index_18358[11:3] + 9'h0bd;
  assign sel_18588 = $signed({1'h0, add_18483, array_index_18274[2:0]}) < $signed({1'h0, sel_18486}) ? {add_18483, array_index_18274[2:0]} : sel_18486;
  assign add_18590 = array_index_18455[11:1] + 11'h247;
  assign sel_18593 = $signed({1'h0, add_18488, array_index_18355[0]}) < $signed({1'h0, sel_18491}) ? {add_18488, array_index_18355[0]} : sel_18491;
  assign add_18595 = array_index_18458[11:1] + 11'h247;
  assign sel_18598 = $signed({1'h0, add_18493, array_index_18358[0]}) < $signed({1'h0, sel_18496}) ? {add_18493, array_index_18358[0]} : sel_18496;
  assign add_18623 = array_index_18557[11:0] + 12'h247;
  assign sel_18625 = $signed({1'h0, add_18521}) < $signed({1'h0, sel_18523}) ? add_18521 : sel_18523;
  assign add_18628 = array_index_18560[11:0] + 12'h247;
  assign sel_18630 = $signed({1'h0, add_18526}) < $signed({1'h0, sel_18528}) ? add_18526 : sel_18528;
  assign array_index_18659 = set1_unflattened[4'h7];
  assign array_index_18662 = set2_unflattened[4'h7];
  assign add_18666 = array_index_18271[11:1] + 11'h79d;
  assign sel_18668 = $signed({1'h0, add_18564, array_index_18205[0]}) < $signed({1'h0, sel_18566}) ? {add_18564, array_index_18205[0]} : sel_18566;
  assign add_18670 = array_index_18274[11:1] + 11'h79d;
  assign sel_18672 = $signed({1'h0, add_18568, array_index_18208[0]}) < $signed({1'h0, sel_18570}) ? {add_18568, array_index_18208[0]} : sel_18570;
  assign add_18674 = array_index_18355[11:1] + 11'h347;
  assign sel_18676 = $signed({1'h0, add_18572, array_index_18271[0]}) < $signed({1'h0, sel_18574}) ? {add_18572, array_index_18271[0]} : sel_18574;
  assign add_18678 = array_index_18358[11:1] + 11'h347;
  assign sel_18680 = $signed({1'h0, add_18576, array_index_18274[0]}) < $signed({1'h0, sel_18578}) ? {add_18576, array_index_18274[0]} : sel_18578;
  assign add_18682 = array_index_18455[11:3] + 9'h0bd;
  assign sel_18685 = $signed({1'h0, add_18580, array_index_18355[2:0]}) < $signed({1'h0, sel_18583}) ? {add_18580, array_index_18355[2:0]} : sel_18583;
  assign add_18687 = array_index_18458[11:3] + 9'h0bd;
  assign sel_18690 = $signed({1'h0, add_18585, array_index_18358[2:0]}) < $signed({1'h0, sel_18588}) ? {add_18585, array_index_18358[2:0]} : sel_18588;
  assign add_18692 = array_index_18557[11:1] + 11'h247;
  assign sel_18695 = $signed({1'h0, add_18590, array_index_18455[0]}) < $signed({1'h0, sel_18593}) ? {add_18590, array_index_18455[0]} : sel_18593;
  assign add_18697 = array_index_18560[11:1] + 11'h247;
  assign sel_18700 = $signed({1'h0, add_18595, array_index_18458[0]}) < $signed({1'h0, sel_18598}) ? {add_18595, array_index_18458[0]} : sel_18598;
  assign add_18725 = array_index_18659[11:0] + 12'h247;
  assign sel_18727 = $signed({1'h0, add_18623}) < $signed({1'h0, sel_18625}) ? add_18623 : sel_18625;
  assign add_18730 = array_index_18662[11:0] + 12'h247;
  assign sel_18732 = $signed({1'h0, add_18628}) < $signed({1'h0, sel_18630}) ? add_18628 : sel_18630;
  assign array_index_18761 = set1_unflattened[4'h8];
  assign array_index_18764 = set2_unflattened[4'h8];
  assign add_18768 = array_index_18355[11:1] + 11'h79d;
  assign sel_18770 = $signed({1'h0, add_18666, array_index_18271[0]}) < $signed({1'h0, sel_18668}) ? {add_18666, array_index_18271[0]} : sel_18668;
  assign add_18772 = array_index_18358[11:1] + 11'h79d;
  assign sel_18774 = $signed({1'h0, add_18670, array_index_18274[0]}) < $signed({1'h0, sel_18672}) ? {add_18670, array_index_18274[0]} : sel_18672;
  assign add_18776 = array_index_18455[11:1] + 11'h347;
  assign sel_18778 = $signed({1'h0, add_18674, array_index_18355[0]}) < $signed({1'h0, sel_18676}) ? {add_18674, array_index_18355[0]} : sel_18676;
  assign add_18780 = array_index_18458[11:1] + 11'h347;
  assign sel_18782 = $signed({1'h0, add_18678, array_index_18358[0]}) < $signed({1'h0, sel_18680}) ? {add_18678, array_index_18358[0]} : sel_18680;
  assign add_18784 = array_index_18557[11:3] + 9'h0bd;
  assign sel_18787 = $signed({1'h0, add_18682, array_index_18455[2:0]}) < $signed({1'h0, sel_18685}) ? {add_18682, array_index_18455[2:0]} : sel_18685;
  assign add_18789 = array_index_18560[11:3] + 9'h0bd;
  assign sel_18792 = $signed({1'h0, add_18687, array_index_18458[2:0]}) < $signed({1'h0, sel_18690}) ? {add_18687, array_index_18458[2:0]} : sel_18690;
  assign add_18794 = array_index_18659[11:1] + 11'h247;
  assign sel_18797 = $signed({1'h0, add_18692, array_index_18557[0]}) < $signed({1'h0, sel_18695}) ? {add_18692, array_index_18557[0]} : sel_18695;
  assign add_18799 = array_index_18662[11:1] + 11'h247;
  assign sel_18802 = $signed({1'h0, add_18697, array_index_18560[0]}) < $signed({1'h0, sel_18700}) ? {add_18697, array_index_18560[0]} : sel_18700;
  assign add_18827 = array_index_18761[11:0] + 12'h247;
  assign sel_18829 = $signed({1'h0, add_18725}) < $signed({1'h0, sel_18727}) ? add_18725 : sel_18727;
  assign add_18832 = array_index_18764[11:0] + 12'h247;
  assign sel_18834 = $signed({1'h0, add_18730}) < $signed({1'h0, sel_18732}) ? add_18730 : sel_18732;
  assign array_index_18863 = set1_unflattened[4'h9];
  assign array_index_18866 = set2_unflattened[4'h9];
  assign add_18870 = array_index_18455[11:1] + 11'h79d;
  assign sel_18872 = $signed({1'h0, add_18768, array_index_18355[0]}) < $signed({1'h0, sel_18770}) ? {add_18768, array_index_18355[0]} : sel_18770;
  assign add_18874 = array_index_18458[11:1] + 11'h79d;
  assign sel_18876 = $signed({1'h0, add_18772, array_index_18358[0]}) < $signed({1'h0, sel_18774}) ? {add_18772, array_index_18358[0]} : sel_18774;
  assign add_18878 = array_index_18557[11:1] + 11'h347;
  assign sel_18880 = $signed({1'h0, add_18776, array_index_18455[0]}) < $signed({1'h0, sel_18778}) ? {add_18776, array_index_18455[0]} : sel_18778;
  assign add_18882 = array_index_18560[11:1] + 11'h347;
  assign sel_18884 = $signed({1'h0, add_18780, array_index_18458[0]}) < $signed({1'h0, sel_18782}) ? {add_18780, array_index_18458[0]} : sel_18782;
  assign add_18886 = array_index_18659[11:3] + 9'h0bd;
  assign sel_18889 = $signed({1'h0, add_18784, array_index_18557[2:0]}) < $signed({1'h0, sel_18787}) ? {add_18784, array_index_18557[2:0]} : sel_18787;
  assign add_18891 = array_index_18662[11:3] + 9'h0bd;
  assign sel_18894 = $signed({1'h0, add_18789, array_index_18560[2:0]}) < $signed({1'h0, sel_18792}) ? {add_18789, array_index_18560[2:0]} : sel_18792;
  assign add_18896 = array_index_18761[11:1] + 11'h247;
  assign sel_18899 = $signed({1'h0, add_18794, array_index_18659[0]}) < $signed({1'h0, sel_18797}) ? {add_18794, array_index_18659[0]} : sel_18797;
  assign add_18901 = array_index_18764[11:1] + 11'h247;
  assign sel_18904 = $signed({1'h0, add_18799, array_index_18662[0]}) < $signed({1'h0, sel_18802}) ? {add_18799, array_index_18662[0]} : sel_18802;
  assign add_18928 = array_index_18863[11:0] + 12'h247;
  assign sel_18930 = $signed({1'h0, add_18827}) < $signed({1'h0, sel_18829}) ? add_18827 : sel_18829;
  assign add_18932 = array_index_18866[11:0] + 12'h247;
  assign sel_18934 = $signed({1'h0, add_18832}) < $signed({1'h0, sel_18834}) ? add_18832 : sel_18834;
  assign add_18968 = array_index_18557[11:1] + 11'h79d;
  assign sel_18970 = $signed({1'h0, add_18870, array_index_18455[0]}) < $signed({1'h0, sel_18872}) ? {add_18870, array_index_18455[0]} : sel_18872;
  assign add_18972 = array_index_18560[11:1] + 11'h79d;
  assign sel_18974 = $signed({1'h0, add_18874, array_index_18458[0]}) < $signed({1'h0, sel_18876}) ? {add_18874, array_index_18458[0]} : sel_18876;
  assign add_18976 = array_index_18659[11:1] + 11'h347;
  assign sel_18978 = $signed({1'h0, add_18878, array_index_18557[0]}) < $signed({1'h0, sel_18880}) ? {add_18878, array_index_18557[0]} : sel_18880;
  assign add_18980 = array_index_18662[11:1] + 11'h347;
  assign sel_18982 = $signed({1'h0, add_18882, array_index_18560[0]}) < $signed({1'h0, sel_18884}) ? {add_18882, array_index_18560[0]} : sel_18884;
  assign add_18984 = array_index_18761[11:3] + 9'h0bd;
  assign sel_18987 = $signed({1'h0, add_18886, array_index_18659[2:0]}) < $signed({1'h0, sel_18889}) ? {add_18886, array_index_18659[2:0]} : sel_18889;
  assign add_18989 = array_index_18764[11:3] + 9'h0bd;
  assign sel_18992 = $signed({1'h0, add_18891, array_index_18662[2:0]}) < $signed({1'h0, sel_18894}) ? {add_18891, array_index_18662[2:0]} : sel_18894;
  assign add_18994 = array_index_18863[11:1] + 11'h247;
  assign sel_18997 = $signed({1'h0, add_18896, array_index_18761[0]}) < $signed({1'h0, sel_18899}) ? {add_18896, array_index_18761[0]} : sel_18899;
  assign add_18999 = array_index_18866[11:1] + 11'h247;
  assign sel_19002 = $signed({1'h0, add_18901, array_index_18764[0]}) < $signed({1'h0, sel_18904}) ? {add_18901, array_index_18764[0]} : sel_18904;
  assign add_19050 = array_index_18659[11:1] + 11'h79d;
  assign sel_19052 = $signed({1'h0, add_18968, array_index_18557[0]}) < $signed({1'h0, sel_18970}) ? {add_18968, array_index_18557[0]} : sel_18970;
  assign add_19054 = array_index_18662[11:1] + 11'h79d;
  assign sel_19056 = $signed({1'h0, add_18972, array_index_18560[0]}) < $signed({1'h0, sel_18974}) ? {add_18972, array_index_18560[0]} : sel_18974;
  assign add_19058 = array_index_18761[11:1] + 11'h347;
  assign sel_19060 = $signed({1'h0, add_18976, array_index_18659[0]}) < $signed({1'h0, sel_18978}) ? {add_18976, array_index_18659[0]} : sel_18978;
  assign add_19062 = array_index_18764[11:1] + 11'h347;
  assign sel_19064 = $signed({1'h0, add_18980, array_index_18662[0]}) < $signed({1'h0, sel_18982}) ? {add_18980, array_index_18662[0]} : sel_18982;
  assign add_19066 = array_index_18863[11:3] + 9'h0bd;
  assign sel_19069 = $signed({1'h0, add_18984, array_index_18761[2:0]}) < $signed({1'h0, sel_18987}) ? {add_18984, array_index_18761[2:0]} : sel_18987;
  assign add_19071 = array_index_18866[11:3] + 9'h0bd;
  assign sel_19074 = $signed({1'h0, add_18989, array_index_18764[2:0]}) < $signed({1'h0, sel_18992}) ? {add_18989, array_index_18764[2:0]} : sel_18992;
  assign concat_19077 = {1'h0, ($signed({1'h0, add_18928}) < $signed({1'h0, sel_18930}) ? add_18928 : sel_18930) == ($signed({1'h0, add_18932}) < $signed({1'h0, sel_18934}) ? add_18932 : sel_18934)};
  assign add_19092 = concat_19077 + 2'h1;
  assign add_19112 = array_index_18761[11:1] + 11'h79d;
  assign sel_19114 = $signed({1'h0, add_19050, array_index_18659[0]}) < $signed({1'h0, sel_19052}) ? {add_19050, array_index_18659[0]} : sel_19052;
  assign add_19116 = array_index_18764[11:1] + 11'h79d;
  assign sel_19118 = $signed({1'h0, add_19054, array_index_18662[0]}) < $signed({1'h0, sel_19056}) ? {add_19054, array_index_18662[0]} : sel_19056;
  assign add_19120 = array_index_18863[11:1] + 11'h347;
  assign sel_19122 = $signed({1'h0, add_19058, array_index_18761[0]}) < $signed({1'h0, sel_19060}) ? {add_19058, array_index_18761[0]} : sel_19060;
  assign add_19124 = array_index_18866[11:1] + 11'h347;
  assign sel_19126 = $signed({1'h0, add_19062, array_index_18764[0]}) < $signed({1'h0, sel_19064}) ? {add_19062, array_index_18764[0]} : sel_19064;
  assign concat_19129 = {1'h0, ($signed({1'h0, add_18994, array_index_18863[0]}) < $signed({1'h0, sel_18997}) ? {add_18994, array_index_18863[0]} : sel_18997) == ($signed({1'h0, add_18999, array_index_18866[0]}) < $signed({1'h0, sel_19002}) ? {add_18999, array_index_18866[0]} : sel_19002) ? add_19092 : concat_19077};
  assign add_19140 = concat_19129 + 3'h1;
  assign add_19154 = array_index_18863[11:1] + 11'h79d;
  assign sel_19156 = $signed({1'h0, add_19112, array_index_18761[0]}) < $signed({1'h0, sel_19114}) ? {add_19112, array_index_18761[0]} : sel_19114;
  assign add_19158 = array_index_18866[11:1] + 11'h79d;
  assign sel_19160 = $signed({1'h0, add_19116, array_index_18764[0]}) < $signed({1'h0, sel_19118}) ? {add_19116, array_index_18764[0]} : sel_19118;
  assign concat_19163 = {1'h0, ($signed({1'h0, add_19066, array_index_18863[2:0]}) < $signed({1'h0, sel_19069}) ? {add_19066, array_index_18863[2:0]} : sel_19069) == ($signed({1'h0, add_19071, array_index_18866[2:0]}) < $signed({1'h0, sel_19074}) ? {add_19071, array_index_18866[2:0]} : sel_19074) ? add_19140 : concat_19129};
  assign add_19170 = concat_19163 + 4'h1;
  assign concat_19179 = {1'h0, ($signed({1'h0, add_19120, array_index_18863[0]}) < $signed({1'h0, sel_19122}) ? {add_19120, array_index_18863[0]} : sel_19122) == ($signed({1'h0, add_19124, array_index_18866[0]}) < $signed({1'h0, sel_19126}) ? {add_19124, array_index_18866[0]} : sel_19126) ? add_19170 : concat_19163};
  assign add_19182 = concat_19179 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_19154, array_index_18863[0]}) < $signed({1'h0, sel_19156}) ? {add_19154, array_index_18863[0]} : sel_19156) == ($signed({1'h0, add_19158, array_index_18866[0]}) < $signed({1'h0, sel_19160}) ? {add_19158, array_index_18866[0]} : sel_19160) ? add_19182 : concat_19179}, {set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
