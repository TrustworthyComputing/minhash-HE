module min_hash(
  input wire [799:0] set1,
  input wire [799:0] set2,
  output wire [1615:0] out
);
  wire [15:0] set1_unflattened[50];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  wire [15:0] set2_unflattened[50];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  wire [15:0] array_index_87063;
  wire [15:0] array_index_87064;
  wire [11:0] add_87071;
  wire [11:0] add_87074;
  wire [15:0] array_index_87079;
  wire [15:0] array_index_87082;
  wire [10:0] add_87086;
  wire [10:0] add_87089;
  wire [11:0] add_87105;
  wire [11:0] sel_87107;
  wire [11:0] add_87110;
  wire [11:0] sel_87112;
  wire [15:0] array_index_87127;
  wire [15:0] array_index_87130;
  wire [8:0] add_87134;
  wire [8:0] add_87137;
  wire [10:0] add_87140;
  wire [11:0] sel_87143;
  wire [10:0] add_87145;
  wire [11:0] sel_87148;
  wire [11:0] add_87165;
  wire [11:0] sel_87167;
  wire [11:0] add_87170;
  wire [11:0] sel_87172;
  wire [15:0] array_index_87193;
  wire [15:0] array_index_87196;
  wire [10:0] add_87200;
  wire [10:0] add_87202;
  wire [8:0] add_87204;
  wire [11:0] sel_87207;
  wire [8:0] add_87209;
  wire [11:0] sel_87212;
  wire [10:0] add_87214;
  wire [11:0] sel_87217;
  wire [10:0] add_87219;
  wire [11:0] sel_87222;
  wire [11:0] add_87243;
  wire [11:0] sel_87245;
  wire [11:0] add_87248;
  wire [11:0] sel_87250;
  wire [15:0] array_index_87277;
  wire [15:0] array_index_87280;
  wire [10:0] add_87284;
  wire [10:0] add_87286;
  wire [10:0] add_87288;
  wire [11:0] sel_87290;
  wire [10:0] add_87292;
  wire [11:0] sel_87294;
  wire [8:0] add_87296;
  wire [11:0] sel_87299;
  wire [8:0] add_87301;
  wire [11:0] sel_87304;
  wire [10:0] add_87306;
  wire [11:0] sel_87309;
  wire [10:0] add_87311;
  wire [11:0] sel_87314;
  wire [11:0] add_87339;
  wire [11:0] sel_87341;
  wire [11:0] add_87344;
  wire [11:0] sel_87346;
  wire [15:0] array_index_87377;
  wire [15:0] array_index_87380;
  wire [10:0] add_87384;
  wire [11:0] sel_87386;
  wire [10:0] add_87388;
  wire [11:0] sel_87390;
  wire [10:0] add_87392;
  wire [11:0] sel_87394;
  wire [10:0] add_87396;
  wire [11:0] sel_87398;
  wire [8:0] add_87400;
  wire [11:0] sel_87403;
  wire [8:0] add_87405;
  wire [11:0] sel_87408;
  wire [10:0] add_87410;
  wire [11:0] sel_87413;
  wire [10:0] add_87415;
  wire [11:0] sel_87418;
  wire [11:0] add_87443;
  wire [11:0] sel_87445;
  wire [11:0] add_87448;
  wire [11:0] sel_87450;
  wire [15:0] array_index_87479;
  wire [15:0] array_index_87482;
  wire [10:0] add_87486;
  wire [11:0] sel_87488;
  wire [10:0] add_87490;
  wire [11:0] sel_87492;
  wire [10:0] add_87494;
  wire [11:0] sel_87496;
  wire [10:0] add_87498;
  wire [11:0] sel_87500;
  wire [8:0] add_87502;
  wire [11:0] sel_87505;
  wire [8:0] add_87507;
  wire [11:0] sel_87510;
  wire [10:0] add_87512;
  wire [11:0] sel_87515;
  wire [10:0] add_87517;
  wire [11:0] sel_87520;
  wire [11:0] add_87545;
  wire [11:0] sel_87547;
  wire [11:0] add_87550;
  wire [11:0] sel_87552;
  wire [15:0] array_index_87581;
  wire [15:0] array_index_87584;
  wire [10:0] add_87588;
  wire [11:0] sel_87590;
  wire [10:0] add_87592;
  wire [11:0] sel_87594;
  wire [10:0] add_87596;
  wire [11:0] sel_87598;
  wire [10:0] add_87600;
  wire [11:0] sel_87602;
  wire [8:0] add_87604;
  wire [11:0] sel_87607;
  wire [8:0] add_87609;
  wire [11:0] sel_87612;
  wire [10:0] add_87614;
  wire [11:0] sel_87617;
  wire [10:0] add_87619;
  wire [11:0] sel_87622;
  wire [11:0] add_87647;
  wire [11:0] sel_87649;
  wire [11:0] add_87652;
  wire [11:0] sel_87654;
  wire [15:0] array_index_87683;
  wire [15:0] array_index_87686;
  wire [10:0] add_87690;
  wire [11:0] sel_87692;
  wire [10:0] add_87694;
  wire [11:0] sel_87696;
  wire [10:0] add_87698;
  wire [11:0] sel_87700;
  wire [10:0] add_87702;
  wire [11:0] sel_87704;
  wire [8:0] add_87706;
  wire [11:0] sel_87709;
  wire [8:0] add_87711;
  wire [11:0] sel_87714;
  wire [10:0] add_87716;
  wire [11:0] sel_87719;
  wire [10:0] add_87721;
  wire [11:0] sel_87724;
  wire [11:0] add_87749;
  wire [11:0] sel_87751;
  wire [11:0] add_87754;
  wire [11:0] sel_87756;
  wire [15:0] array_index_87785;
  wire [15:0] array_index_87788;
  wire [10:0] add_87792;
  wire [11:0] sel_87794;
  wire [10:0] add_87796;
  wire [11:0] sel_87798;
  wire [10:0] add_87800;
  wire [11:0] sel_87802;
  wire [10:0] add_87804;
  wire [11:0] sel_87806;
  wire [8:0] add_87808;
  wire [11:0] sel_87811;
  wire [8:0] add_87813;
  wire [11:0] sel_87816;
  wire [10:0] add_87818;
  wire [11:0] sel_87821;
  wire [10:0] add_87823;
  wire [11:0] sel_87826;
  wire [11:0] add_87851;
  wire [11:0] sel_87853;
  wire [11:0] add_87856;
  wire [11:0] sel_87858;
  wire [15:0] array_index_87887;
  wire [15:0] array_index_87890;
  wire [10:0] add_87894;
  wire [11:0] sel_87896;
  wire [10:0] add_87898;
  wire [11:0] sel_87900;
  wire [10:0] add_87902;
  wire [11:0] sel_87904;
  wire [10:0] add_87906;
  wire [11:0] sel_87908;
  wire [8:0] add_87910;
  wire [11:0] sel_87913;
  wire [8:0] add_87915;
  wire [11:0] sel_87918;
  wire [10:0] add_87920;
  wire [11:0] sel_87923;
  wire [10:0] add_87925;
  wire [11:0] sel_87928;
  wire [11:0] add_87953;
  wire [11:0] sel_87955;
  wire [11:0] add_87958;
  wire [11:0] sel_87960;
  wire [15:0] array_index_87989;
  wire [15:0] array_index_87992;
  wire [10:0] add_87996;
  wire [11:0] sel_87998;
  wire [10:0] add_88000;
  wire [11:0] sel_88002;
  wire [10:0] add_88004;
  wire [11:0] sel_88006;
  wire [10:0] add_88008;
  wire [11:0] sel_88010;
  wire [8:0] add_88012;
  wire [11:0] sel_88015;
  wire [8:0] add_88017;
  wire [11:0] sel_88020;
  wire [10:0] add_88022;
  wire [11:0] sel_88025;
  wire [10:0] add_88027;
  wire [11:0] sel_88030;
  wire [11:0] add_88055;
  wire [11:0] sel_88057;
  wire [11:0] add_88060;
  wire [11:0] sel_88062;
  wire [15:0] array_index_88091;
  wire [15:0] array_index_88094;
  wire [10:0] add_88098;
  wire [11:0] sel_88100;
  wire [10:0] add_88102;
  wire [11:0] sel_88104;
  wire [10:0] add_88106;
  wire [11:0] sel_88108;
  wire [10:0] add_88110;
  wire [11:0] sel_88112;
  wire [8:0] add_88114;
  wire [11:0] sel_88117;
  wire [8:0] add_88119;
  wire [11:0] sel_88122;
  wire [10:0] add_88124;
  wire [11:0] sel_88127;
  wire [10:0] add_88129;
  wire [11:0] sel_88132;
  wire [11:0] add_88157;
  wire [11:0] sel_88159;
  wire [11:0] add_88162;
  wire [11:0] sel_88164;
  wire [15:0] array_index_88193;
  wire [15:0] array_index_88196;
  wire [10:0] add_88200;
  wire [11:0] sel_88202;
  wire [10:0] add_88204;
  wire [11:0] sel_88206;
  wire [10:0] add_88208;
  wire [11:0] sel_88210;
  wire [10:0] add_88212;
  wire [11:0] sel_88214;
  wire [8:0] add_88216;
  wire [11:0] sel_88219;
  wire [8:0] add_88221;
  wire [11:0] sel_88224;
  wire [10:0] add_88226;
  wire [11:0] sel_88229;
  wire [10:0] add_88231;
  wire [11:0] sel_88234;
  wire [11:0] add_88259;
  wire [11:0] sel_88261;
  wire [11:0] add_88264;
  wire [11:0] sel_88266;
  wire [15:0] array_index_88295;
  wire [15:0] array_index_88298;
  wire [10:0] add_88302;
  wire [11:0] sel_88304;
  wire [10:0] add_88306;
  wire [11:0] sel_88308;
  wire [10:0] add_88310;
  wire [11:0] sel_88312;
  wire [10:0] add_88314;
  wire [11:0] sel_88316;
  wire [8:0] add_88318;
  wire [11:0] sel_88321;
  wire [8:0] add_88323;
  wire [11:0] sel_88326;
  wire [10:0] add_88328;
  wire [11:0] sel_88331;
  wire [10:0] add_88333;
  wire [11:0] sel_88336;
  wire [11:0] add_88361;
  wire [11:0] sel_88363;
  wire [11:0] add_88366;
  wire [11:0] sel_88368;
  wire [15:0] array_index_88397;
  wire [15:0] array_index_88400;
  wire [10:0] add_88404;
  wire [11:0] sel_88406;
  wire [10:0] add_88408;
  wire [11:0] sel_88410;
  wire [10:0] add_88412;
  wire [11:0] sel_88414;
  wire [10:0] add_88416;
  wire [11:0] sel_88418;
  wire [8:0] add_88420;
  wire [11:0] sel_88423;
  wire [8:0] add_88425;
  wire [11:0] sel_88428;
  wire [10:0] add_88430;
  wire [11:0] sel_88433;
  wire [10:0] add_88435;
  wire [11:0] sel_88438;
  wire [11:0] add_88463;
  wire [11:0] sel_88465;
  wire [11:0] add_88468;
  wire [11:0] sel_88470;
  wire [15:0] array_index_88499;
  wire [15:0] array_index_88502;
  wire [10:0] add_88506;
  wire [11:0] sel_88508;
  wire [10:0] add_88510;
  wire [11:0] sel_88512;
  wire [10:0] add_88514;
  wire [11:0] sel_88516;
  wire [10:0] add_88518;
  wire [11:0] sel_88520;
  wire [8:0] add_88522;
  wire [11:0] sel_88525;
  wire [8:0] add_88527;
  wire [11:0] sel_88530;
  wire [10:0] add_88532;
  wire [11:0] sel_88535;
  wire [10:0] add_88537;
  wire [11:0] sel_88540;
  wire [11:0] add_88565;
  wire [11:0] sel_88567;
  wire [11:0] add_88570;
  wire [11:0] sel_88572;
  wire [15:0] array_index_88601;
  wire [15:0] array_index_88604;
  wire [10:0] add_88608;
  wire [11:0] sel_88610;
  wire [10:0] add_88612;
  wire [11:0] sel_88614;
  wire [10:0] add_88616;
  wire [11:0] sel_88618;
  wire [10:0] add_88620;
  wire [11:0] sel_88622;
  wire [8:0] add_88624;
  wire [11:0] sel_88627;
  wire [8:0] add_88629;
  wire [11:0] sel_88632;
  wire [10:0] add_88634;
  wire [11:0] sel_88637;
  wire [10:0] add_88639;
  wire [11:0] sel_88642;
  wire [11:0] add_88667;
  wire [11:0] sel_88669;
  wire [11:0] add_88672;
  wire [11:0] sel_88674;
  wire [15:0] array_index_88703;
  wire [15:0] array_index_88706;
  wire [10:0] add_88710;
  wire [11:0] sel_88712;
  wire [10:0] add_88714;
  wire [11:0] sel_88716;
  wire [10:0] add_88718;
  wire [11:0] sel_88720;
  wire [10:0] add_88722;
  wire [11:0] sel_88724;
  wire [8:0] add_88726;
  wire [11:0] sel_88729;
  wire [8:0] add_88731;
  wire [11:0] sel_88734;
  wire [10:0] add_88736;
  wire [11:0] sel_88739;
  wire [10:0] add_88741;
  wire [11:0] sel_88744;
  wire [11:0] add_88769;
  wire [11:0] sel_88771;
  wire [11:0] add_88774;
  wire [11:0] sel_88776;
  wire [15:0] array_index_88805;
  wire [15:0] array_index_88808;
  wire [10:0] add_88812;
  wire [11:0] sel_88814;
  wire [10:0] add_88816;
  wire [11:0] sel_88818;
  wire [10:0] add_88820;
  wire [11:0] sel_88822;
  wire [10:0] add_88824;
  wire [11:0] sel_88826;
  wire [8:0] add_88828;
  wire [11:0] sel_88831;
  wire [8:0] add_88833;
  wire [11:0] sel_88836;
  wire [10:0] add_88838;
  wire [11:0] sel_88841;
  wire [10:0] add_88843;
  wire [11:0] sel_88846;
  wire [11:0] add_88871;
  wire [11:0] sel_88873;
  wire [11:0] add_88876;
  wire [11:0] sel_88878;
  wire [15:0] array_index_88907;
  wire [15:0] array_index_88910;
  wire [10:0] add_88914;
  wire [11:0] sel_88916;
  wire [10:0] add_88918;
  wire [11:0] sel_88920;
  wire [10:0] add_88922;
  wire [11:0] sel_88924;
  wire [10:0] add_88926;
  wire [11:0] sel_88928;
  wire [8:0] add_88930;
  wire [11:0] sel_88933;
  wire [8:0] add_88935;
  wire [11:0] sel_88938;
  wire [10:0] add_88940;
  wire [11:0] sel_88943;
  wire [10:0] add_88945;
  wire [11:0] sel_88948;
  wire [11:0] add_88973;
  wire [11:0] sel_88975;
  wire [11:0] add_88978;
  wire [11:0] sel_88980;
  wire [15:0] array_index_89009;
  wire [15:0] array_index_89012;
  wire [10:0] add_89016;
  wire [11:0] sel_89018;
  wire [10:0] add_89020;
  wire [11:0] sel_89022;
  wire [10:0] add_89024;
  wire [11:0] sel_89026;
  wire [10:0] add_89028;
  wire [11:0] sel_89030;
  wire [8:0] add_89032;
  wire [11:0] sel_89035;
  wire [8:0] add_89037;
  wire [11:0] sel_89040;
  wire [10:0] add_89042;
  wire [11:0] sel_89045;
  wire [10:0] add_89047;
  wire [11:0] sel_89050;
  wire [11:0] add_89075;
  wire [11:0] sel_89077;
  wire [11:0] add_89080;
  wire [11:0] sel_89082;
  wire [15:0] array_index_89111;
  wire [15:0] array_index_89114;
  wire [10:0] add_89118;
  wire [11:0] sel_89120;
  wire [10:0] add_89122;
  wire [11:0] sel_89124;
  wire [10:0] add_89126;
  wire [11:0] sel_89128;
  wire [10:0] add_89130;
  wire [11:0] sel_89132;
  wire [8:0] add_89134;
  wire [11:0] sel_89137;
  wire [8:0] add_89139;
  wire [11:0] sel_89142;
  wire [10:0] add_89144;
  wire [11:0] sel_89147;
  wire [10:0] add_89149;
  wire [11:0] sel_89152;
  wire [11:0] add_89177;
  wire [11:0] sel_89179;
  wire [11:0] add_89182;
  wire [11:0] sel_89184;
  wire [15:0] array_index_89213;
  wire [15:0] array_index_89216;
  wire [10:0] add_89220;
  wire [11:0] sel_89222;
  wire [10:0] add_89224;
  wire [11:0] sel_89226;
  wire [10:0] add_89228;
  wire [11:0] sel_89230;
  wire [10:0] add_89232;
  wire [11:0] sel_89234;
  wire [8:0] add_89236;
  wire [11:0] sel_89239;
  wire [8:0] add_89241;
  wire [11:0] sel_89244;
  wire [10:0] add_89246;
  wire [11:0] sel_89249;
  wire [10:0] add_89251;
  wire [11:0] sel_89254;
  wire [11:0] add_89279;
  wire [11:0] sel_89281;
  wire [11:0] add_89284;
  wire [11:0] sel_89286;
  wire [15:0] array_index_89315;
  wire [15:0] array_index_89318;
  wire [10:0] add_89322;
  wire [11:0] sel_89324;
  wire [10:0] add_89326;
  wire [11:0] sel_89328;
  wire [10:0] add_89330;
  wire [11:0] sel_89332;
  wire [10:0] add_89334;
  wire [11:0] sel_89336;
  wire [8:0] add_89338;
  wire [11:0] sel_89341;
  wire [8:0] add_89343;
  wire [11:0] sel_89346;
  wire [10:0] add_89348;
  wire [11:0] sel_89351;
  wire [10:0] add_89353;
  wire [11:0] sel_89356;
  wire [11:0] add_89381;
  wire [11:0] sel_89383;
  wire [11:0] add_89386;
  wire [11:0] sel_89388;
  wire [15:0] array_index_89417;
  wire [15:0] array_index_89420;
  wire [10:0] add_89424;
  wire [11:0] sel_89426;
  wire [10:0] add_89428;
  wire [11:0] sel_89430;
  wire [10:0] add_89432;
  wire [11:0] sel_89434;
  wire [10:0] add_89436;
  wire [11:0] sel_89438;
  wire [8:0] add_89440;
  wire [11:0] sel_89443;
  wire [8:0] add_89445;
  wire [11:0] sel_89448;
  wire [10:0] add_89450;
  wire [11:0] sel_89453;
  wire [10:0] add_89455;
  wire [11:0] sel_89458;
  wire [11:0] add_89483;
  wire [11:0] sel_89485;
  wire [11:0] add_89488;
  wire [11:0] sel_89490;
  wire [15:0] array_index_89519;
  wire [15:0] array_index_89522;
  wire [10:0] add_89526;
  wire [11:0] sel_89528;
  wire [10:0] add_89530;
  wire [11:0] sel_89532;
  wire [10:0] add_89534;
  wire [11:0] sel_89536;
  wire [10:0] add_89538;
  wire [11:0] sel_89540;
  wire [8:0] add_89542;
  wire [11:0] sel_89545;
  wire [8:0] add_89547;
  wire [11:0] sel_89550;
  wire [10:0] add_89552;
  wire [11:0] sel_89555;
  wire [10:0] add_89557;
  wire [11:0] sel_89560;
  wire [11:0] add_89585;
  wire [11:0] sel_89587;
  wire [11:0] add_89590;
  wire [11:0] sel_89592;
  wire [15:0] array_index_89621;
  wire [15:0] array_index_89624;
  wire [10:0] add_89628;
  wire [11:0] sel_89630;
  wire [10:0] add_89632;
  wire [11:0] sel_89634;
  wire [10:0] add_89636;
  wire [11:0] sel_89638;
  wire [10:0] add_89640;
  wire [11:0] sel_89642;
  wire [8:0] add_89644;
  wire [11:0] sel_89647;
  wire [8:0] add_89649;
  wire [11:0] sel_89652;
  wire [10:0] add_89654;
  wire [11:0] sel_89657;
  wire [10:0] add_89659;
  wire [11:0] sel_89662;
  wire [11:0] add_89687;
  wire [11:0] sel_89689;
  wire [11:0] add_89692;
  wire [11:0] sel_89694;
  wire [15:0] array_index_89723;
  wire [15:0] array_index_89726;
  wire [10:0] add_89730;
  wire [11:0] sel_89732;
  wire [10:0] add_89734;
  wire [11:0] sel_89736;
  wire [10:0] add_89738;
  wire [11:0] sel_89740;
  wire [10:0] add_89742;
  wire [11:0] sel_89744;
  wire [8:0] add_89746;
  wire [11:0] sel_89749;
  wire [8:0] add_89751;
  wire [11:0] sel_89754;
  wire [10:0] add_89756;
  wire [11:0] sel_89759;
  wire [10:0] add_89761;
  wire [11:0] sel_89764;
  wire [11:0] add_89789;
  wire [11:0] sel_89791;
  wire [11:0] add_89794;
  wire [11:0] sel_89796;
  wire [15:0] array_index_89825;
  wire [15:0] array_index_89828;
  wire [10:0] add_89832;
  wire [11:0] sel_89834;
  wire [10:0] add_89836;
  wire [11:0] sel_89838;
  wire [10:0] add_89840;
  wire [11:0] sel_89842;
  wire [10:0] add_89844;
  wire [11:0] sel_89846;
  wire [8:0] add_89848;
  wire [11:0] sel_89851;
  wire [8:0] add_89853;
  wire [11:0] sel_89856;
  wire [10:0] add_89858;
  wire [11:0] sel_89861;
  wire [10:0] add_89863;
  wire [11:0] sel_89866;
  wire [11:0] add_89891;
  wire [11:0] sel_89893;
  wire [11:0] add_89896;
  wire [11:0] sel_89898;
  wire [15:0] array_index_89927;
  wire [15:0] array_index_89930;
  wire [10:0] add_89934;
  wire [11:0] sel_89936;
  wire [10:0] add_89938;
  wire [11:0] sel_89940;
  wire [10:0] add_89942;
  wire [11:0] sel_89944;
  wire [10:0] add_89946;
  wire [11:0] sel_89948;
  wire [8:0] add_89950;
  wire [11:0] sel_89953;
  wire [8:0] add_89955;
  wire [11:0] sel_89958;
  wire [10:0] add_89960;
  wire [11:0] sel_89963;
  wire [10:0] add_89965;
  wire [11:0] sel_89968;
  wire [11:0] add_89993;
  wire [11:0] sel_89995;
  wire [11:0] add_89998;
  wire [11:0] sel_90000;
  wire [15:0] array_index_90029;
  wire [15:0] array_index_90032;
  wire [10:0] add_90036;
  wire [11:0] sel_90038;
  wire [10:0] add_90040;
  wire [11:0] sel_90042;
  wire [10:0] add_90044;
  wire [11:0] sel_90046;
  wire [10:0] add_90048;
  wire [11:0] sel_90050;
  wire [8:0] add_90052;
  wire [11:0] sel_90055;
  wire [8:0] add_90057;
  wire [11:0] sel_90060;
  wire [10:0] add_90062;
  wire [11:0] sel_90065;
  wire [10:0] add_90067;
  wire [11:0] sel_90070;
  wire [11:0] add_90095;
  wire [11:0] sel_90097;
  wire [11:0] add_90100;
  wire [11:0] sel_90102;
  wire [15:0] array_index_90131;
  wire [15:0] array_index_90134;
  wire [10:0] add_90138;
  wire [11:0] sel_90140;
  wire [10:0] add_90142;
  wire [11:0] sel_90144;
  wire [10:0] add_90146;
  wire [11:0] sel_90148;
  wire [10:0] add_90150;
  wire [11:0] sel_90152;
  wire [8:0] add_90154;
  wire [11:0] sel_90157;
  wire [8:0] add_90159;
  wire [11:0] sel_90162;
  wire [10:0] add_90164;
  wire [11:0] sel_90167;
  wire [10:0] add_90169;
  wire [11:0] sel_90172;
  wire [11:0] add_90197;
  wire [11:0] sel_90199;
  wire [11:0] add_90202;
  wire [11:0] sel_90204;
  wire [15:0] array_index_90233;
  wire [15:0] array_index_90236;
  wire [10:0] add_90240;
  wire [11:0] sel_90242;
  wire [10:0] add_90244;
  wire [11:0] sel_90246;
  wire [10:0] add_90248;
  wire [11:0] sel_90250;
  wire [10:0] add_90252;
  wire [11:0] sel_90254;
  wire [8:0] add_90256;
  wire [11:0] sel_90259;
  wire [8:0] add_90261;
  wire [11:0] sel_90264;
  wire [10:0] add_90266;
  wire [11:0] sel_90269;
  wire [10:0] add_90271;
  wire [11:0] sel_90274;
  wire [11:0] add_90299;
  wire [11:0] sel_90301;
  wire [11:0] add_90304;
  wire [11:0] sel_90306;
  wire [15:0] array_index_90335;
  wire [15:0] array_index_90338;
  wire [10:0] add_90342;
  wire [11:0] sel_90344;
  wire [10:0] add_90346;
  wire [11:0] sel_90348;
  wire [10:0] add_90350;
  wire [11:0] sel_90352;
  wire [10:0] add_90354;
  wire [11:0] sel_90356;
  wire [8:0] add_90358;
  wire [11:0] sel_90361;
  wire [8:0] add_90363;
  wire [11:0] sel_90366;
  wire [10:0] add_90368;
  wire [11:0] sel_90371;
  wire [10:0] add_90373;
  wire [11:0] sel_90376;
  wire [11:0] add_90401;
  wire [11:0] sel_90403;
  wire [11:0] add_90406;
  wire [11:0] sel_90408;
  wire [15:0] array_index_90437;
  wire [15:0] array_index_90440;
  wire [10:0] add_90444;
  wire [11:0] sel_90446;
  wire [10:0] add_90448;
  wire [11:0] sel_90450;
  wire [10:0] add_90452;
  wire [11:0] sel_90454;
  wire [10:0] add_90456;
  wire [11:0] sel_90458;
  wire [8:0] add_90460;
  wire [11:0] sel_90463;
  wire [8:0] add_90465;
  wire [11:0] sel_90468;
  wire [10:0] add_90470;
  wire [11:0] sel_90473;
  wire [10:0] add_90475;
  wire [11:0] sel_90478;
  wire [11:0] add_90503;
  wire [11:0] sel_90505;
  wire [11:0] add_90508;
  wire [11:0] sel_90510;
  wire [15:0] array_index_90539;
  wire [15:0] array_index_90542;
  wire [10:0] add_90546;
  wire [11:0] sel_90548;
  wire [10:0] add_90550;
  wire [11:0] sel_90552;
  wire [10:0] add_90554;
  wire [11:0] sel_90556;
  wire [10:0] add_90558;
  wire [11:0] sel_90560;
  wire [8:0] add_90562;
  wire [11:0] sel_90565;
  wire [8:0] add_90567;
  wire [11:0] sel_90570;
  wire [10:0] add_90572;
  wire [11:0] sel_90575;
  wire [10:0] add_90577;
  wire [11:0] sel_90580;
  wire [11:0] add_90605;
  wire [11:0] sel_90607;
  wire [11:0] add_90610;
  wire [11:0] sel_90612;
  wire [15:0] array_index_90641;
  wire [15:0] array_index_90644;
  wire [10:0] add_90648;
  wire [11:0] sel_90650;
  wire [10:0] add_90652;
  wire [11:0] sel_90654;
  wire [10:0] add_90656;
  wire [11:0] sel_90658;
  wire [10:0] add_90660;
  wire [11:0] sel_90662;
  wire [8:0] add_90664;
  wire [11:0] sel_90667;
  wire [8:0] add_90669;
  wire [11:0] sel_90672;
  wire [10:0] add_90674;
  wire [11:0] sel_90677;
  wire [10:0] add_90679;
  wire [11:0] sel_90682;
  wire [11:0] add_90707;
  wire [11:0] sel_90709;
  wire [11:0] add_90712;
  wire [11:0] sel_90714;
  wire [15:0] array_index_90743;
  wire [15:0] array_index_90746;
  wire [10:0] add_90750;
  wire [11:0] sel_90752;
  wire [10:0] add_90754;
  wire [11:0] sel_90756;
  wire [10:0] add_90758;
  wire [11:0] sel_90760;
  wire [10:0] add_90762;
  wire [11:0] sel_90764;
  wire [8:0] add_90766;
  wire [11:0] sel_90769;
  wire [8:0] add_90771;
  wire [11:0] sel_90774;
  wire [10:0] add_90776;
  wire [11:0] sel_90779;
  wire [10:0] add_90781;
  wire [11:0] sel_90784;
  wire [11:0] add_90809;
  wire [11:0] sel_90811;
  wire [11:0] add_90814;
  wire [11:0] sel_90816;
  wire [15:0] array_index_90845;
  wire [15:0] array_index_90848;
  wire [10:0] add_90852;
  wire [11:0] sel_90854;
  wire [10:0] add_90856;
  wire [11:0] sel_90858;
  wire [10:0] add_90860;
  wire [11:0] sel_90862;
  wire [10:0] add_90864;
  wire [11:0] sel_90866;
  wire [8:0] add_90868;
  wire [11:0] sel_90871;
  wire [8:0] add_90873;
  wire [11:0] sel_90876;
  wire [10:0] add_90878;
  wire [11:0] sel_90881;
  wire [10:0] add_90883;
  wire [11:0] sel_90886;
  wire [11:0] add_90911;
  wire [11:0] sel_90913;
  wire [11:0] add_90916;
  wire [11:0] sel_90918;
  wire [15:0] array_index_90947;
  wire [15:0] array_index_90950;
  wire [10:0] add_90954;
  wire [11:0] sel_90956;
  wire [10:0] add_90958;
  wire [11:0] sel_90960;
  wire [10:0] add_90962;
  wire [11:0] sel_90964;
  wire [10:0] add_90966;
  wire [11:0] sel_90968;
  wire [8:0] add_90970;
  wire [11:0] sel_90973;
  wire [8:0] add_90975;
  wire [11:0] sel_90978;
  wire [10:0] add_90980;
  wire [11:0] sel_90983;
  wire [10:0] add_90985;
  wire [11:0] sel_90988;
  wire [11:0] add_91013;
  wire [11:0] sel_91015;
  wire [11:0] add_91018;
  wire [11:0] sel_91020;
  wire [15:0] array_index_91049;
  wire [15:0] array_index_91052;
  wire [10:0] add_91056;
  wire [11:0] sel_91058;
  wire [10:0] add_91060;
  wire [11:0] sel_91062;
  wire [10:0] add_91064;
  wire [11:0] sel_91066;
  wire [10:0] add_91068;
  wire [11:0] sel_91070;
  wire [8:0] add_91072;
  wire [11:0] sel_91075;
  wire [8:0] add_91077;
  wire [11:0] sel_91080;
  wire [10:0] add_91082;
  wire [11:0] sel_91085;
  wire [10:0] add_91087;
  wire [11:0] sel_91090;
  wire [11:0] add_91115;
  wire [11:0] sel_91117;
  wire [11:0] add_91120;
  wire [11:0] sel_91122;
  wire [15:0] array_index_91151;
  wire [15:0] array_index_91154;
  wire [10:0] add_91158;
  wire [11:0] sel_91160;
  wire [10:0] add_91162;
  wire [11:0] sel_91164;
  wire [10:0] add_91166;
  wire [11:0] sel_91168;
  wire [10:0] add_91170;
  wire [11:0] sel_91172;
  wire [8:0] add_91174;
  wire [11:0] sel_91177;
  wire [8:0] add_91179;
  wire [11:0] sel_91182;
  wire [10:0] add_91184;
  wire [11:0] sel_91187;
  wire [10:0] add_91189;
  wire [11:0] sel_91192;
  wire [11:0] add_91217;
  wire [11:0] sel_91219;
  wire [11:0] add_91222;
  wire [11:0] sel_91224;
  wire [15:0] array_index_91253;
  wire [15:0] array_index_91256;
  wire [10:0] add_91260;
  wire [11:0] sel_91262;
  wire [10:0] add_91264;
  wire [11:0] sel_91266;
  wire [10:0] add_91268;
  wire [11:0] sel_91270;
  wire [10:0] add_91272;
  wire [11:0] sel_91274;
  wire [8:0] add_91276;
  wire [11:0] sel_91279;
  wire [8:0] add_91281;
  wire [11:0] sel_91284;
  wire [10:0] add_91286;
  wire [11:0] sel_91289;
  wire [10:0] add_91291;
  wire [11:0] sel_91294;
  wire [11:0] add_91319;
  wire [11:0] sel_91321;
  wire [11:0] add_91324;
  wire [11:0] sel_91326;
  wire [15:0] array_index_91355;
  wire [15:0] array_index_91358;
  wire [10:0] add_91362;
  wire [11:0] sel_91364;
  wire [10:0] add_91366;
  wire [11:0] sel_91368;
  wire [10:0] add_91370;
  wire [11:0] sel_91372;
  wire [10:0] add_91374;
  wire [11:0] sel_91376;
  wire [8:0] add_91378;
  wire [11:0] sel_91381;
  wire [8:0] add_91383;
  wire [11:0] sel_91386;
  wire [10:0] add_91388;
  wire [11:0] sel_91391;
  wire [10:0] add_91393;
  wire [11:0] sel_91396;
  wire [11:0] add_91421;
  wire [11:0] sel_91423;
  wire [11:0] add_91426;
  wire [11:0] sel_91428;
  wire [15:0] array_index_91457;
  wire [15:0] array_index_91460;
  wire [10:0] add_91464;
  wire [11:0] sel_91466;
  wire [10:0] add_91468;
  wire [11:0] sel_91470;
  wire [10:0] add_91472;
  wire [11:0] sel_91474;
  wire [10:0] add_91476;
  wire [11:0] sel_91478;
  wire [8:0] add_91480;
  wire [11:0] sel_91483;
  wire [8:0] add_91485;
  wire [11:0] sel_91488;
  wire [10:0] add_91490;
  wire [11:0] sel_91493;
  wire [10:0] add_91495;
  wire [11:0] sel_91498;
  wire [11:0] add_91523;
  wire [11:0] sel_91525;
  wire [11:0] add_91528;
  wire [11:0] sel_91530;
  wire [15:0] array_index_91559;
  wire [15:0] array_index_91562;
  wire [10:0] add_91566;
  wire [11:0] sel_91568;
  wire [10:0] add_91570;
  wire [11:0] sel_91572;
  wire [10:0] add_91574;
  wire [11:0] sel_91576;
  wire [10:0] add_91578;
  wire [11:0] sel_91580;
  wire [8:0] add_91582;
  wire [11:0] sel_91585;
  wire [8:0] add_91587;
  wire [11:0] sel_91590;
  wire [10:0] add_91592;
  wire [11:0] sel_91595;
  wire [10:0] add_91597;
  wire [11:0] sel_91600;
  wire [11:0] add_91625;
  wire [11:0] sel_91627;
  wire [11:0] add_91630;
  wire [11:0] sel_91632;
  wire [15:0] array_index_91661;
  wire [15:0] array_index_91664;
  wire [10:0] add_91668;
  wire [11:0] sel_91670;
  wire [10:0] add_91672;
  wire [11:0] sel_91674;
  wire [10:0] add_91676;
  wire [11:0] sel_91678;
  wire [10:0] add_91680;
  wire [11:0] sel_91682;
  wire [8:0] add_91684;
  wire [11:0] sel_91687;
  wire [8:0] add_91689;
  wire [11:0] sel_91692;
  wire [10:0] add_91694;
  wire [11:0] sel_91697;
  wire [10:0] add_91699;
  wire [11:0] sel_91702;
  wire [11:0] add_91727;
  wire [11:0] sel_91729;
  wire [11:0] add_91732;
  wire [11:0] sel_91734;
  wire [15:0] array_index_91763;
  wire [15:0] array_index_91766;
  wire [10:0] add_91770;
  wire [11:0] sel_91772;
  wire [10:0] add_91774;
  wire [11:0] sel_91776;
  wire [10:0] add_91778;
  wire [11:0] sel_91780;
  wire [10:0] add_91782;
  wire [11:0] sel_91784;
  wire [8:0] add_91786;
  wire [11:0] sel_91789;
  wire [8:0] add_91791;
  wire [11:0] sel_91794;
  wire [10:0] add_91796;
  wire [11:0] sel_91799;
  wire [10:0] add_91801;
  wire [11:0] sel_91804;
  wire [11:0] add_91829;
  wire [11:0] sel_91831;
  wire [11:0] add_91834;
  wire [11:0] sel_91836;
  wire [15:0] array_index_91865;
  wire [15:0] array_index_91868;
  wire [10:0] add_91872;
  wire [11:0] sel_91874;
  wire [10:0] add_91876;
  wire [11:0] sel_91878;
  wire [10:0] add_91880;
  wire [11:0] sel_91882;
  wire [10:0] add_91884;
  wire [11:0] sel_91886;
  wire [8:0] add_91888;
  wire [11:0] sel_91891;
  wire [8:0] add_91893;
  wire [11:0] sel_91896;
  wire [10:0] add_91898;
  wire [11:0] sel_91901;
  wire [10:0] add_91903;
  wire [11:0] sel_91906;
  wire [11:0] add_91930;
  wire [11:0] sel_91932;
  wire [11:0] add_91934;
  wire [11:0] sel_91936;
  wire [10:0] add_91970;
  wire [11:0] sel_91972;
  wire [10:0] add_91974;
  wire [11:0] sel_91976;
  wire [10:0] add_91978;
  wire [11:0] sel_91980;
  wire [10:0] add_91982;
  wire [11:0] sel_91984;
  wire [8:0] add_91986;
  wire [11:0] sel_91989;
  wire [8:0] add_91991;
  wire [11:0] sel_91994;
  wire [10:0] add_91996;
  wire [11:0] sel_91999;
  wire [10:0] add_92001;
  wire [11:0] sel_92004;
  wire [10:0] add_92052;
  wire [11:0] sel_92054;
  wire [10:0] add_92056;
  wire [11:0] sel_92058;
  wire [10:0] add_92060;
  wire [11:0] sel_92062;
  wire [10:0] add_92064;
  wire [11:0] sel_92066;
  wire [8:0] add_92068;
  wire [11:0] sel_92071;
  wire [8:0] add_92073;
  wire [11:0] sel_92076;
  wire [1:0] concat_92079;
  wire [1:0] add_92094;
  wire [10:0] add_92114;
  wire [11:0] sel_92116;
  wire [10:0] add_92118;
  wire [11:0] sel_92120;
  wire [10:0] add_92122;
  wire [11:0] sel_92124;
  wire [10:0] add_92126;
  wire [11:0] sel_92128;
  wire [2:0] concat_92131;
  wire [2:0] add_92142;
  wire [10:0] add_92156;
  wire [11:0] sel_92158;
  wire [10:0] add_92160;
  wire [11:0] sel_92162;
  wire [3:0] concat_92165;
  wire [3:0] add_92172;
  wire [4:0] concat_92181;
  wire [4:0] add_92184;
  assign array_index_87063 = set1_unflattened[6'h00];
  assign array_index_87064 = set2_unflattened[6'h00];
  assign add_87071 = array_index_87063[11:0] + 12'h247;
  assign add_87074 = array_index_87064[11:0] + 12'h247;
  assign array_index_87079 = set1_unflattened[6'h01];
  assign array_index_87082 = set2_unflattened[6'h01];
  assign add_87086 = array_index_87063[11:1] + 11'h247;
  assign add_87089 = array_index_87064[11:1] + 11'h247;
  assign add_87105 = array_index_87079[11:0] + 12'h247;
  assign sel_87107 = $signed({1'h0, add_87071}) < $signed(13'h0fff) ? add_87071 : 12'hfff;
  assign add_87110 = array_index_87082[11:0] + 12'h247;
  assign sel_87112 = $signed({1'h0, add_87074}) < $signed(13'h0fff) ? add_87074 : 12'hfff;
  assign array_index_87127 = set1_unflattened[6'h02];
  assign array_index_87130 = set2_unflattened[6'h02];
  assign add_87134 = array_index_87063[11:3] + 9'h0bd;
  assign add_87137 = array_index_87064[11:3] + 9'h0bd;
  assign add_87140 = array_index_87079[11:1] + 11'h247;
  assign sel_87143 = $signed({1'h0, add_87086, array_index_87063[0]}) < $signed(13'h0fff) ? {add_87086, array_index_87063[0]} : 12'hfff;
  assign add_87145 = array_index_87082[11:1] + 11'h247;
  assign sel_87148 = $signed({1'h0, add_87089, array_index_87064[0]}) < $signed(13'h0fff) ? {add_87089, array_index_87064[0]} : 12'hfff;
  assign add_87165 = array_index_87127[11:0] + 12'h247;
  assign sel_87167 = $signed({1'h0, add_87105}) < $signed({1'h0, sel_87107}) ? add_87105 : sel_87107;
  assign add_87170 = array_index_87130[11:0] + 12'h247;
  assign sel_87172 = $signed({1'h0, add_87110}) < $signed({1'h0, sel_87112}) ? add_87110 : sel_87112;
  assign array_index_87193 = set1_unflattened[6'h03];
  assign array_index_87196 = set2_unflattened[6'h03];
  assign add_87200 = array_index_87063[11:1] + 11'h347;
  assign add_87202 = array_index_87064[11:1] + 11'h347;
  assign add_87204 = array_index_87079[11:3] + 9'h0bd;
  assign sel_87207 = $signed({1'h0, add_87134, array_index_87063[2:0]}) < $signed(13'h0fff) ? {add_87134, array_index_87063[2:0]} : 12'hfff;
  assign add_87209 = array_index_87082[11:3] + 9'h0bd;
  assign sel_87212 = $signed({1'h0, add_87137, array_index_87064[2:0]}) < $signed(13'h0fff) ? {add_87137, array_index_87064[2:0]} : 12'hfff;
  assign add_87214 = array_index_87127[11:1] + 11'h247;
  assign sel_87217 = $signed({1'h0, add_87140, array_index_87079[0]}) < $signed({1'h0, sel_87143}) ? {add_87140, array_index_87079[0]} : sel_87143;
  assign add_87219 = array_index_87130[11:1] + 11'h247;
  assign sel_87222 = $signed({1'h0, add_87145, array_index_87082[0]}) < $signed({1'h0, sel_87148}) ? {add_87145, array_index_87082[0]} : sel_87148;
  assign add_87243 = array_index_87193[11:0] + 12'h247;
  assign sel_87245 = $signed({1'h0, add_87165}) < $signed({1'h0, sel_87167}) ? add_87165 : sel_87167;
  assign add_87248 = array_index_87196[11:0] + 12'h247;
  assign sel_87250 = $signed({1'h0, add_87170}) < $signed({1'h0, sel_87172}) ? add_87170 : sel_87172;
  assign array_index_87277 = set1_unflattened[6'h04];
  assign array_index_87280 = set2_unflattened[6'h04];
  assign add_87284 = array_index_87063[11:1] + 11'h79d;
  assign add_87286 = array_index_87064[11:1] + 11'h79d;
  assign add_87288 = array_index_87079[11:1] + 11'h347;
  assign sel_87290 = $signed({1'h0, add_87200, array_index_87063[0]}) < $signed(13'h0fff) ? {add_87200, array_index_87063[0]} : 12'hfff;
  assign add_87292 = array_index_87082[11:1] + 11'h347;
  assign sel_87294 = $signed({1'h0, add_87202, array_index_87064[0]}) < $signed(13'h0fff) ? {add_87202, array_index_87064[0]} : 12'hfff;
  assign add_87296 = array_index_87127[11:3] + 9'h0bd;
  assign sel_87299 = $signed({1'h0, add_87204, array_index_87079[2:0]}) < $signed({1'h0, sel_87207}) ? {add_87204, array_index_87079[2:0]} : sel_87207;
  assign add_87301 = array_index_87130[11:3] + 9'h0bd;
  assign sel_87304 = $signed({1'h0, add_87209, array_index_87082[2:0]}) < $signed({1'h0, sel_87212}) ? {add_87209, array_index_87082[2:0]} : sel_87212;
  assign add_87306 = array_index_87193[11:1] + 11'h247;
  assign sel_87309 = $signed({1'h0, add_87214, array_index_87127[0]}) < $signed({1'h0, sel_87217}) ? {add_87214, array_index_87127[0]} : sel_87217;
  assign add_87311 = array_index_87196[11:1] + 11'h247;
  assign sel_87314 = $signed({1'h0, add_87219, array_index_87130[0]}) < $signed({1'h0, sel_87222}) ? {add_87219, array_index_87130[0]} : sel_87222;
  assign add_87339 = array_index_87277[11:0] + 12'h247;
  assign sel_87341 = $signed({1'h0, add_87243}) < $signed({1'h0, sel_87245}) ? add_87243 : sel_87245;
  assign add_87344 = array_index_87280[11:0] + 12'h247;
  assign sel_87346 = $signed({1'h0, add_87248}) < $signed({1'h0, sel_87250}) ? add_87248 : sel_87250;
  assign array_index_87377 = set1_unflattened[6'h05];
  assign array_index_87380 = set2_unflattened[6'h05];
  assign add_87384 = array_index_87079[11:1] + 11'h79d;
  assign sel_87386 = $signed({1'h0, add_87284, array_index_87063[0]}) < $signed(13'h0fff) ? {add_87284, array_index_87063[0]} : 12'hfff;
  assign add_87388 = array_index_87082[11:1] + 11'h79d;
  assign sel_87390 = $signed({1'h0, add_87286, array_index_87064[0]}) < $signed(13'h0fff) ? {add_87286, array_index_87064[0]} : 12'hfff;
  assign add_87392 = array_index_87127[11:1] + 11'h347;
  assign sel_87394 = $signed({1'h0, add_87288, array_index_87079[0]}) < $signed({1'h0, sel_87290}) ? {add_87288, array_index_87079[0]} : sel_87290;
  assign add_87396 = array_index_87130[11:1] + 11'h347;
  assign sel_87398 = $signed({1'h0, add_87292, array_index_87082[0]}) < $signed({1'h0, sel_87294}) ? {add_87292, array_index_87082[0]} : sel_87294;
  assign add_87400 = array_index_87193[11:3] + 9'h0bd;
  assign sel_87403 = $signed({1'h0, add_87296, array_index_87127[2:0]}) < $signed({1'h0, sel_87299}) ? {add_87296, array_index_87127[2:0]} : sel_87299;
  assign add_87405 = array_index_87196[11:3] + 9'h0bd;
  assign sel_87408 = $signed({1'h0, add_87301, array_index_87130[2:0]}) < $signed({1'h0, sel_87304}) ? {add_87301, array_index_87130[2:0]} : sel_87304;
  assign add_87410 = array_index_87277[11:1] + 11'h247;
  assign sel_87413 = $signed({1'h0, add_87306, array_index_87193[0]}) < $signed({1'h0, sel_87309}) ? {add_87306, array_index_87193[0]} : sel_87309;
  assign add_87415 = array_index_87280[11:1] + 11'h247;
  assign sel_87418 = $signed({1'h0, add_87311, array_index_87196[0]}) < $signed({1'h0, sel_87314}) ? {add_87311, array_index_87196[0]} : sel_87314;
  assign add_87443 = array_index_87377[11:0] + 12'h247;
  assign sel_87445 = $signed({1'h0, add_87339}) < $signed({1'h0, sel_87341}) ? add_87339 : sel_87341;
  assign add_87448 = array_index_87380[11:0] + 12'h247;
  assign sel_87450 = $signed({1'h0, add_87344}) < $signed({1'h0, sel_87346}) ? add_87344 : sel_87346;
  assign array_index_87479 = set1_unflattened[6'h06];
  assign array_index_87482 = set2_unflattened[6'h06];
  assign add_87486 = array_index_87127[11:1] + 11'h79d;
  assign sel_87488 = $signed({1'h0, add_87384, array_index_87079[0]}) < $signed({1'h0, sel_87386}) ? {add_87384, array_index_87079[0]} : sel_87386;
  assign add_87490 = array_index_87130[11:1] + 11'h79d;
  assign sel_87492 = $signed({1'h0, add_87388, array_index_87082[0]}) < $signed({1'h0, sel_87390}) ? {add_87388, array_index_87082[0]} : sel_87390;
  assign add_87494 = array_index_87193[11:1] + 11'h347;
  assign sel_87496 = $signed({1'h0, add_87392, array_index_87127[0]}) < $signed({1'h0, sel_87394}) ? {add_87392, array_index_87127[0]} : sel_87394;
  assign add_87498 = array_index_87196[11:1] + 11'h347;
  assign sel_87500 = $signed({1'h0, add_87396, array_index_87130[0]}) < $signed({1'h0, sel_87398}) ? {add_87396, array_index_87130[0]} : sel_87398;
  assign add_87502 = array_index_87277[11:3] + 9'h0bd;
  assign sel_87505 = $signed({1'h0, add_87400, array_index_87193[2:0]}) < $signed({1'h0, sel_87403}) ? {add_87400, array_index_87193[2:0]} : sel_87403;
  assign add_87507 = array_index_87280[11:3] + 9'h0bd;
  assign sel_87510 = $signed({1'h0, add_87405, array_index_87196[2:0]}) < $signed({1'h0, sel_87408}) ? {add_87405, array_index_87196[2:0]} : sel_87408;
  assign add_87512 = array_index_87377[11:1] + 11'h247;
  assign sel_87515 = $signed({1'h0, add_87410, array_index_87277[0]}) < $signed({1'h0, sel_87413}) ? {add_87410, array_index_87277[0]} : sel_87413;
  assign add_87517 = array_index_87380[11:1] + 11'h247;
  assign sel_87520 = $signed({1'h0, add_87415, array_index_87280[0]}) < $signed({1'h0, sel_87418}) ? {add_87415, array_index_87280[0]} : sel_87418;
  assign add_87545 = array_index_87479[11:0] + 12'h247;
  assign sel_87547 = $signed({1'h0, add_87443}) < $signed({1'h0, sel_87445}) ? add_87443 : sel_87445;
  assign add_87550 = array_index_87482[11:0] + 12'h247;
  assign sel_87552 = $signed({1'h0, add_87448}) < $signed({1'h0, sel_87450}) ? add_87448 : sel_87450;
  assign array_index_87581 = set1_unflattened[6'h07];
  assign array_index_87584 = set2_unflattened[6'h07];
  assign add_87588 = array_index_87193[11:1] + 11'h79d;
  assign sel_87590 = $signed({1'h0, add_87486, array_index_87127[0]}) < $signed({1'h0, sel_87488}) ? {add_87486, array_index_87127[0]} : sel_87488;
  assign add_87592 = array_index_87196[11:1] + 11'h79d;
  assign sel_87594 = $signed({1'h0, add_87490, array_index_87130[0]}) < $signed({1'h0, sel_87492}) ? {add_87490, array_index_87130[0]} : sel_87492;
  assign add_87596 = array_index_87277[11:1] + 11'h347;
  assign sel_87598 = $signed({1'h0, add_87494, array_index_87193[0]}) < $signed({1'h0, sel_87496}) ? {add_87494, array_index_87193[0]} : sel_87496;
  assign add_87600 = array_index_87280[11:1] + 11'h347;
  assign sel_87602 = $signed({1'h0, add_87498, array_index_87196[0]}) < $signed({1'h0, sel_87500}) ? {add_87498, array_index_87196[0]} : sel_87500;
  assign add_87604 = array_index_87377[11:3] + 9'h0bd;
  assign sel_87607 = $signed({1'h0, add_87502, array_index_87277[2:0]}) < $signed({1'h0, sel_87505}) ? {add_87502, array_index_87277[2:0]} : sel_87505;
  assign add_87609 = array_index_87380[11:3] + 9'h0bd;
  assign sel_87612 = $signed({1'h0, add_87507, array_index_87280[2:0]}) < $signed({1'h0, sel_87510}) ? {add_87507, array_index_87280[2:0]} : sel_87510;
  assign add_87614 = array_index_87479[11:1] + 11'h247;
  assign sel_87617 = $signed({1'h0, add_87512, array_index_87377[0]}) < $signed({1'h0, sel_87515}) ? {add_87512, array_index_87377[0]} : sel_87515;
  assign add_87619 = array_index_87482[11:1] + 11'h247;
  assign sel_87622 = $signed({1'h0, add_87517, array_index_87380[0]}) < $signed({1'h0, sel_87520}) ? {add_87517, array_index_87380[0]} : sel_87520;
  assign add_87647 = array_index_87581[11:0] + 12'h247;
  assign sel_87649 = $signed({1'h0, add_87545}) < $signed({1'h0, sel_87547}) ? add_87545 : sel_87547;
  assign add_87652 = array_index_87584[11:0] + 12'h247;
  assign sel_87654 = $signed({1'h0, add_87550}) < $signed({1'h0, sel_87552}) ? add_87550 : sel_87552;
  assign array_index_87683 = set1_unflattened[6'h08];
  assign array_index_87686 = set2_unflattened[6'h08];
  assign add_87690 = array_index_87277[11:1] + 11'h79d;
  assign sel_87692 = $signed({1'h0, add_87588, array_index_87193[0]}) < $signed({1'h0, sel_87590}) ? {add_87588, array_index_87193[0]} : sel_87590;
  assign add_87694 = array_index_87280[11:1] + 11'h79d;
  assign sel_87696 = $signed({1'h0, add_87592, array_index_87196[0]}) < $signed({1'h0, sel_87594}) ? {add_87592, array_index_87196[0]} : sel_87594;
  assign add_87698 = array_index_87377[11:1] + 11'h347;
  assign sel_87700 = $signed({1'h0, add_87596, array_index_87277[0]}) < $signed({1'h0, sel_87598}) ? {add_87596, array_index_87277[0]} : sel_87598;
  assign add_87702 = array_index_87380[11:1] + 11'h347;
  assign sel_87704 = $signed({1'h0, add_87600, array_index_87280[0]}) < $signed({1'h0, sel_87602}) ? {add_87600, array_index_87280[0]} : sel_87602;
  assign add_87706 = array_index_87479[11:3] + 9'h0bd;
  assign sel_87709 = $signed({1'h0, add_87604, array_index_87377[2:0]}) < $signed({1'h0, sel_87607}) ? {add_87604, array_index_87377[2:0]} : sel_87607;
  assign add_87711 = array_index_87482[11:3] + 9'h0bd;
  assign sel_87714 = $signed({1'h0, add_87609, array_index_87380[2:0]}) < $signed({1'h0, sel_87612}) ? {add_87609, array_index_87380[2:0]} : sel_87612;
  assign add_87716 = array_index_87581[11:1] + 11'h247;
  assign sel_87719 = $signed({1'h0, add_87614, array_index_87479[0]}) < $signed({1'h0, sel_87617}) ? {add_87614, array_index_87479[0]} : sel_87617;
  assign add_87721 = array_index_87584[11:1] + 11'h247;
  assign sel_87724 = $signed({1'h0, add_87619, array_index_87482[0]}) < $signed({1'h0, sel_87622}) ? {add_87619, array_index_87482[0]} : sel_87622;
  assign add_87749 = array_index_87683[11:0] + 12'h247;
  assign sel_87751 = $signed({1'h0, add_87647}) < $signed({1'h0, sel_87649}) ? add_87647 : sel_87649;
  assign add_87754 = array_index_87686[11:0] + 12'h247;
  assign sel_87756 = $signed({1'h0, add_87652}) < $signed({1'h0, sel_87654}) ? add_87652 : sel_87654;
  assign array_index_87785 = set1_unflattened[6'h09];
  assign array_index_87788 = set2_unflattened[6'h09];
  assign add_87792 = array_index_87377[11:1] + 11'h79d;
  assign sel_87794 = $signed({1'h0, add_87690, array_index_87277[0]}) < $signed({1'h0, sel_87692}) ? {add_87690, array_index_87277[0]} : sel_87692;
  assign add_87796 = array_index_87380[11:1] + 11'h79d;
  assign sel_87798 = $signed({1'h0, add_87694, array_index_87280[0]}) < $signed({1'h0, sel_87696}) ? {add_87694, array_index_87280[0]} : sel_87696;
  assign add_87800 = array_index_87479[11:1] + 11'h347;
  assign sel_87802 = $signed({1'h0, add_87698, array_index_87377[0]}) < $signed({1'h0, sel_87700}) ? {add_87698, array_index_87377[0]} : sel_87700;
  assign add_87804 = array_index_87482[11:1] + 11'h347;
  assign sel_87806 = $signed({1'h0, add_87702, array_index_87380[0]}) < $signed({1'h0, sel_87704}) ? {add_87702, array_index_87380[0]} : sel_87704;
  assign add_87808 = array_index_87581[11:3] + 9'h0bd;
  assign sel_87811 = $signed({1'h0, add_87706, array_index_87479[2:0]}) < $signed({1'h0, sel_87709}) ? {add_87706, array_index_87479[2:0]} : sel_87709;
  assign add_87813 = array_index_87584[11:3] + 9'h0bd;
  assign sel_87816 = $signed({1'h0, add_87711, array_index_87482[2:0]}) < $signed({1'h0, sel_87714}) ? {add_87711, array_index_87482[2:0]} : sel_87714;
  assign add_87818 = array_index_87683[11:1] + 11'h247;
  assign sel_87821 = $signed({1'h0, add_87716, array_index_87581[0]}) < $signed({1'h0, sel_87719}) ? {add_87716, array_index_87581[0]} : sel_87719;
  assign add_87823 = array_index_87686[11:1] + 11'h247;
  assign sel_87826 = $signed({1'h0, add_87721, array_index_87584[0]}) < $signed({1'h0, sel_87724}) ? {add_87721, array_index_87584[0]} : sel_87724;
  assign add_87851 = array_index_87785[11:0] + 12'h247;
  assign sel_87853 = $signed({1'h0, add_87749}) < $signed({1'h0, sel_87751}) ? add_87749 : sel_87751;
  assign add_87856 = array_index_87788[11:0] + 12'h247;
  assign sel_87858 = $signed({1'h0, add_87754}) < $signed({1'h0, sel_87756}) ? add_87754 : sel_87756;
  assign array_index_87887 = set1_unflattened[6'h0a];
  assign array_index_87890 = set2_unflattened[6'h0a];
  assign add_87894 = array_index_87479[11:1] + 11'h79d;
  assign sel_87896 = $signed({1'h0, add_87792, array_index_87377[0]}) < $signed({1'h0, sel_87794}) ? {add_87792, array_index_87377[0]} : sel_87794;
  assign add_87898 = array_index_87482[11:1] + 11'h79d;
  assign sel_87900 = $signed({1'h0, add_87796, array_index_87380[0]}) < $signed({1'h0, sel_87798}) ? {add_87796, array_index_87380[0]} : sel_87798;
  assign add_87902 = array_index_87581[11:1] + 11'h347;
  assign sel_87904 = $signed({1'h0, add_87800, array_index_87479[0]}) < $signed({1'h0, sel_87802}) ? {add_87800, array_index_87479[0]} : sel_87802;
  assign add_87906 = array_index_87584[11:1] + 11'h347;
  assign sel_87908 = $signed({1'h0, add_87804, array_index_87482[0]}) < $signed({1'h0, sel_87806}) ? {add_87804, array_index_87482[0]} : sel_87806;
  assign add_87910 = array_index_87683[11:3] + 9'h0bd;
  assign sel_87913 = $signed({1'h0, add_87808, array_index_87581[2:0]}) < $signed({1'h0, sel_87811}) ? {add_87808, array_index_87581[2:0]} : sel_87811;
  assign add_87915 = array_index_87686[11:3] + 9'h0bd;
  assign sel_87918 = $signed({1'h0, add_87813, array_index_87584[2:0]}) < $signed({1'h0, sel_87816}) ? {add_87813, array_index_87584[2:0]} : sel_87816;
  assign add_87920 = array_index_87785[11:1] + 11'h247;
  assign sel_87923 = $signed({1'h0, add_87818, array_index_87683[0]}) < $signed({1'h0, sel_87821}) ? {add_87818, array_index_87683[0]} : sel_87821;
  assign add_87925 = array_index_87788[11:1] + 11'h247;
  assign sel_87928 = $signed({1'h0, add_87823, array_index_87686[0]}) < $signed({1'h0, sel_87826}) ? {add_87823, array_index_87686[0]} : sel_87826;
  assign add_87953 = array_index_87887[11:0] + 12'h247;
  assign sel_87955 = $signed({1'h0, add_87851}) < $signed({1'h0, sel_87853}) ? add_87851 : sel_87853;
  assign add_87958 = array_index_87890[11:0] + 12'h247;
  assign sel_87960 = $signed({1'h0, add_87856}) < $signed({1'h0, sel_87858}) ? add_87856 : sel_87858;
  assign array_index_87989 = set1_unflattened[6'h0b];
  assign array_index_87992 = set2_unflattened[6'h0b];
  assign add_87996 = array_index_87581[11:1] + 11'h79d;
  assign sel_87998 = $signed({1'h0, add_87894, array_index_87479[0]}) < $signed({1'h0, sel_87896}) ? {add_87894, array_index_87479[0]} : sel_87896;
  assign add_88000 = array_index_87584[11:1] + 11'h79d;
  assign sel_88002 = $signed({1'h0, add_87898, array_index_87482[0]}) < $signed({1'h0, sel_87900}) ? {add_87898, array_index_87482[0]} : sel_87900;
  assign add_88004 = array_index_87683[11:1] + 11'h347;
  assign sel_88006 = $signed({1'h0, add_87902, array_index_87581[0]}) < $signed({1'h0, sel_87904}) ? {add_87902, array_index_87581[0]} : sel_87904;
  assign add_88008 = array_index_87686[11:1] + 11'h347;
  assign sel_88010 = $signed({1'h0, add_87906, array_index_87584[0]}) < $signed({1'h0, sel_87908}) ? {add_87906, array_index_87584[0]} : sel_87908;
  assign add_88012 = array_index_87785[11:3] + 9'h0bd;
  assign sel_88015 = $signed({1'h0, add_87910, array_index_87683[2:0]}) < $signed({1'h0, sel_87913}) ? {add_87910, array_index_87683[2:0]} : sel_87913;
  assign add_88017 = array_index_87788[11:3] + 9'h0bd;
  assign sel_88020 = $signed({1'h0, add_87915, array_index_87686[2:0]}) < $signed({1'h0, sel_87918}) ? {add_87915, array_index_87686[2:0]} : sel_87918;
  assign add_88022 = array_index_87887[11:1] + 11'h247;
  assign sel_88025 = $signed({1'h0, add_87920, array_index_87785[0]}) < $signed({1'h0, sel_87923}) ? {add_87920, array_index_87785[0]} : sel_87923;
  assign add_88027 = array_index_87890[11:1] + 11'h247;
  assign sel_88030 = $signed({1'h0, add_87925, array_index_87788[0]}) < $signed({1'h0, sel_87928}) ? {add_87925, array_index_87788[0]} : sel_87928;
  assign add_88055 = array_index_87989[11:0] + 12'h247;
  assign sel_88057 = $signed({1'h0, add_87953}) < $signed({1'h0, sel_87955}) ? add_87953 : sel_87955;
  assign add_88060 = array_index_87992[11:0] + 12'h247;
  assign sel_88062 = $signed({1'h0, add_87958}) < $signed({1'h0, sel_87960}) ? add_87958 : sel_87960;
  assign array_index_88091 = set1_unflattened[6'h0c];
  assign array_index_88094 = set2_unflattened[6'h0c];
  assign add_88098 = array_index_87683[11:1] + 11'h79d;
  assign sel_88100 = $signed({1'h0, add_87996, array_index_87581[0]}) < $signed({1'h0, sel_87998}) ? {add_87996, array_index_87581[0]} : sel_87998;
  assign add_88102 = array_index_87686[11:1] + 11'h79d;
  assign sel_88104 = $signed({1'h0, add_88000, array_index_87584[0]}) < $signed({1'h0, sel_88002}) ? {add_88000, array_index_87584[0]} : sel_88002;
  assign add_88106 = array_index_87785[11:1] + 11'h347;
  assign sel_88108 = $signed({1'h0, add_88004, array_index_87683[0]}) < $signed({1'h0, sel_88006}) ? {add_88004, array_index_87683[0]} : sel_88006;
  assign add_88110 = array_index_87788[11:1] + 11'h347;
  assign sel_88112 = $signed({1'h0, add_88008, array_index_87686[0]}) < $signed({1'h0, sel_88010}) ? {add_88008, array_index_87686[0]} : sel_88010;
  assign add_88114 = array_index_87887[11:3] + 9'h0bd;
  assign sel_88117 = $signed({1'h0, add_88012, array_index_87785[2:0]}) < $signed({1'h0, sel_88015}) ? {add_88012, array_index_87785[2:0]} : sel_88015;
  assign add_88119 = array_index_87890[11:3] + 9'h0bd;
  assign sel_88122 = $signed({1'h0, add_88017, array_index_87788[2:0]}) < $signed({1'h0, sel_88020}) ? {add_88017, array_index_87788[2:0]} : sel_88020;
  assign add_88124 = array_index_87989[11:1] + 11'h247;
  assign sel_88127 = $signed({1'h0, add_88022, array_index_87887[0]}) < $signed({1'h0, sel_88025}) ? {add_88022, array_index_87887[0]} : sel_88025;
  assign add_88129 = array_index_87992[11:1] + 11'h247;
  assign sel_88132 = $signed({1'h0, add_88027, array_index_87890[0]}) < $signed({1'h0, sel_88030}) ? {add_88027, array_index_87890[0]} : sel_88030;
  assign add_88157 = array_index_88091[11:0] + 12'h247;
  assign sel_88159 = $signed({1'h0, add_88055}) < $signed({1'h0, sel_88057}) ? add_88055 : sel_88057;
  assign add_88162 = array_index_88094[11:0] + 12'h247;
  assign sel_88164 = $signed({1'h0, add_88060}) < $signed({1'h0, sel_88062}) ? add_88060 : sel_88062;
  assign array_index_88193 = set1_unflattened[6'h0d];
  assign array_index_88196 = set2_unflattened[6'h0d];
  assign add_88200 = array_index_87785[11:1] + 11'h79d;
  assign sel_88202 = $signed({1'h0, add_88098, array_index_87683[0]}) < $signed({1'h0, sel_88100}) ? {add_88098, array_index_87683[0]} : sel_88100;
  assign add_88204 = array_index_87788[11:1] + 11'h79d;
  assign sel_88206 = $signed({1'h0, add_88102, array_index_87686[0]}) < $signed({1'h0, sel_88104}) ? {add_88102, array_index_87686[0]} : sel_88104;
  assign add_88208 = array_index_87887[11:1] + 11'h347;
  assign sel_88210 = $signed({1'h0, add_88106, array_index_87785[0]}) < $signed({1'h0, sel_88108}) ? {add_88106, array_index_87785[0]} : sel_88108;
  assign add_88212 = array_index_87890[11:1] + 11'h347;
  assign sel_88214 = $signed({1'h0, add_88110, array_index_87788[0]}) < $signed({1'h0, sel_88112}) ? {add_88110, array_index_87788[0]} : sel_88112;
  assign add_88216 = array_index_87989[11:3] + 9'h0bd;
  assign sel_88219 = $signed({1'h0, add_88114, array_index_87887[2:0]}) < $signed({1'h0, sel_88117}) ? {add_88114, array_index_87887[2:0]} : sel_88117;
  assign add_88221 = array_index_87992[11:3] + 9'h0bd;
  assign sel_88224 = $signed({1'h0, add_88119, array_index_87890[2:0]}) < $signed({1'h0, sel_88122}) ? {add_88119, array_index_87890[2:0]} : sel_88122;
  assign add_88226 = array_index_88091[11:1] + 11'h247;
  assign sel_88229 = $signed({1'h0, add_88124, array_index_87989[0]}) < $signed({1'h0, sel_88127}) ? {add_88124, array_index_87989[0]} : sel_88127;
  assign add_88231 = array_index_88094[11:1] + 11'h247;
  assign sel_88234 = $signed({1'h0, add_88129, array_index_87992[0]}) < $signed({1'h0, sel_88132}) ? {add_88129, array_index_87992[0]} : sel_88132;
  assign add_88259 = array_index_88193[11:0] + 12'h247;
  assign sel_88261 = $signed({1'h0, add_88157}) < $signed({1'h0, sel_88159}) ? add_88157 : sel_88159;
  assign add_88264 = array_index_88196[11:0] + 12'h247;
  assign sel_88266 = $signed({1'h0, add_88162}) < $signed({1'h0, sel_88164}) ? add_88162 : sel_88164;
  assign array_index_88295 = set1_unflattened[6'h0e];
  assign array_index_88298 = set2_unflattened[6'h0e];
  assign add_88302 = array_index_87887[11:1] + 11'h79d;
  assign sel_88304 = $signed({1'h0, add_88200, array_index_87785[0]}) < $signed({1'h0, sel_88202}) ? {add_88200, array_index_87785[0]} : sel_88202;
  assign add_88306 = array_index_87890[11:1] + 11'h79d;
  assign sel_88308 = $signed({1'h0, add_88204, array_index_87788[0]}) < $signed({1'h0, sel_88206}) ? {add_88204, array_index_87788[0]} : sel_88206;
  assign add_88310 = array_index_87989[11:1] + 11'h347;
  assign sel_88312 = $signed({1'h0, add_88208, array_index_87887[0]}) < $signed({1'h0, sel_88210}) ? {add_88208, array_index_87887[0]} : sel_88210;
  assign add_88314 = array_index_87992[11:1] + 11'h347;
  assign sel_88316 = $signed({1'h0, add_88212, array_index_87890[0]}) < $signed({1'h0, sel_88214}) ? {add_88212, array_index_87890[0]} : sel_88214;
  assign add_88318 = array_index_88091[11:3] + 9'h0bd;
  assign sel_88321 = $signed({1'h0, add_88216, array_index_87989[2:0]}) < $signed({1'h0, sel_88219}) ? {add_88216, array_index_87989[2:0]} : sel_88219;
  assign add_88323 = array_index_88094[11:3] + 9'h0bd;
  assign sel_88326 = $signed({1'h0, add_88221, array_index_87992[2:0]}) < $signed({1'h0, sel_88224}) ? {add_88221, array_index_87992[2:0]} : sel_88224;
  assign add_88328 = array_index_88193[11:1] + 11'h247;
  assign sel_88331 = $signed({1'h0, add_88226, array_index_88091[0]}) < $signed({1'h0, sel_88229}) ? {add_88226, array_index_88091[0]} : sel_88229;
  assign add_88333 = array_index_88196[11:1] + 11'h247;
  assign sel_88336 = $signed({1'h0, add_88231, array_index_88094[0]}) < $signed({1'h0, sel_88234}) ? {add_88231, array_index_88094[0]} : sel_88234;
  assign add_88361 = array_index_88295[11:0] + 12'h247;
  assign sel_88363 = $signed({1'h0, add_88259}) < $signed({1'h0, sel_88261}) ? add_88259 : sel_88261;
  assign add_88366 = array_index_88298[11:0] + 12'h247;
  assign sel_88368 = $signed({1'h0, add_88264}) < $signed({1'h0, sel_88266}) ? add_88264 : sel_88266;
  assign array_index_88397 = set1_unflattened[6'h0f];
  assign array_index_88400 = set2_unflattened[6'h0f];
  assign add_88404 = array_index_87989[11:1] + 11'h79d;
  assign sel_88406 = $signed({1'h0, add_88302, array_index_87887[0]}) < $signed({1'h0, sel_88304}) ? {add_88302, array_index_87887[0]} : sel_88304;
  assign add_88408 = array_index_87992[11:1] + 11'h79d;
  assign sel_88410 = $signed({1'h0, add_88306, array_index_87890[0]}) < $signed({1'h0, sel_88308}) ? {add_88306, array_index_87890[0]} : sel_88308;
  assign add_88412 = array_index_88091[11:1] + 11'h347;
  assign sel_88414 = $signed({1'h0, add_88310, array_index_87989[0]}) < $signed({1'h0, sel_88312}) ? {add_88310, array_index_87989[0]} : sel_88312;
  assign add_88416 = array_index_88094[11:1] + 11'h347;
  assign sel_88418 = $signed({1'h0, add_88314, array_index_87992[0]}) < $signed({1'h0, sel_88316}) ? {add_88314, array_index_87992[0]} : sel_88316;
  assign add_88420 = array_index_88193[11:3] + 9'h0bd;
  assign sel_88423 = $signed({1'h0, add_88318, array_index_88091[2:0]}) < $signed({1'h0, sel_88321}) ? {add_88318, array_index_88091[2:0]} : sel_88321;
  assign add_88425 = array_index_88196[11:3] + 9'h0bd;
  assign sel_88428 = $signed({1'h0, add_88323, array_index_88094[2:0]}) < $signed({1'h0, sel_88326}) ? {add_88323, array_index_88094[2:0]} : sel_88326;
  assign add_88430 = array_index_88295[11:1] + 11'h247;
  assign sel_88433 = $signed({1'h0, add_88328, array_index_88193[0]}) < $signed({1'h0, sel_88331}) ? {add_88328, array_index_88193[0]} : sel_88331;
  assign add_88435 = array_index_88298[11:1] + 11'h247;
  assign sel_88438 = $signed({1'h0, add_88333, array_index_88196[0]}) < $signed({1'h0, sel_88336}) ? {add_88333, array_index_88196[0]} : sel_88336;
  assign add_88463 = array_index_88397[11:0] + 12'h247;
  assign sel_88465 = $signed({1'h0, add_88361}) < $signed({1'h0, sel_88363}) ? add_88361 : sel_88363;
  assign add_88468 = array_index_88400[11:0] + 12'h247;
  assign sel_88470 = $signed({1'h0, add_88366}) < $signed({1'h0, sel_88368}) ? add_88366 : sel_88368;
  assign array_index_88499 = set1_unflattened[6'h10];
  assign array_index_88502 = set2_unflattened[6'h10];
  assign add_88506 = array_index_88091[11:1] + 11'h79d;
  assign sel_88508 = $signed({1'h0, add_88404, array_index_87989[0]}) < $signed({1'h0, sel_88406}) ? {add_88404, array_index_87989[0]} : sel_88406;
  assign add_88510 = array_index_88094[11:1] + 11'h79d;
  assign sel_88512 = $signed({1'h0, add_88408, array_index_87992[0]}) < $signed({1'h0, sel_88410}) ? {add_88408, array_index_87992[0]} : sel_88410;
  assign add_88514 = array_index_88193[11:1] + 11'h347;
  assign sel_88516 = $signed({1'h0, add_88412, array_index_88091[0]}) < $signed({1'h0, sel_88414}) ? {add_88412, array_index_88091[0]} : sel_88414;
  assign add_88518 = array_index_88196[11:1] + 11'h347;
  assign sel_88520 = $signed({1'h0, add_88416, array_index_88094[0]}) < $signed({1'h0, sel_88418}) ? {add_88416, array_index_88094[0]} : sel_88418;
  assign add_88522 = array_index_88295[11:3] + 9'h0bd;
  assign sel_88525 = $signed({1'h0, add_88420, array_index_88193[2:0]}) < $signed({1'h0, sel_88423}) ? {add_88420, array_index_88193[2:0]} : sel_88423;
  assign add_88527 = array_index_88298[11:3] + 9'h0bd;
  assign sel_88530 = $signed({1'h0, add_88425, array_index_88196[2:0]}) < $signed({1'h0, sel_88428}) ? {add_88425, array_index_88196[2:0]} : sel_88428;
  assign add_88532 = array_index_88397[11:1] + 11'h247;
  assign sel_88535 = $signed({1'h0, add_88430, array_index_88295[0]}) < $signed({1'h0, sel_88433}) ? {add_88430, array_index_88295[0]} : sel_88433;
  assign add_88537 = array_index_88400[11:1] + 11'h247;
  assign sel_88540 = $signed({1'h0, add_88435, array_index_88298[0]}) < $signed({1'h0, sel_88438}) ? {add_88435, array_index_88298[0]} : sel_88438;
  assign add_88565 = array_index_88499[11:0] + 12'h247;
  assign sel_88567 = $signed({1'h0, add_88463}) < $signed({1'h0, sel_88465}) ? add_88463 : sel_88465;
  assign add_88570 = array_index_88502[11:0] + 12'h247;
  assign sel_88572 = $signed({1'h0, add_88468}) < $signed({1'h0, sel_88470}) ? add_88468 : sel_88470;
  assign array_index_88601 = set1_unflattened[6'h11];
  assign array_index_88604 = set2_unflattened[6'h11];
  assign add_88608 = array_index_88193[11:1] + 11'h79d;
  assign sel_88610 = $signed({1'h0, add_88506, array_index_88091[0]}) < $signed({1'h0, sel_88508}) ? {add_88506, array_index_88091[0]} : sel_88508;
  assign add_88612 = array_index_88196[11:1] + 11'h79d;
  assign sel_88614 = $signed({1'h0, add_88510, array_index_88094[0]}) < $signed({1'h0, sel_88512}) ? {add_88510, array_index_88094[0]} : sel_88512;
  assign add_88616 = array_index_88295[11:1] + 11'h347;
  assign sel_88618 = $signed({1'h0, add_88514, array_index_88193[0]}) < $signed({1'h0, sel_88516}) ? {add_88514, array_index_88193[0]} : sel_88516;
  assign add_88620 = array_index_88298[11:1] + 11'h347;
  assign sel_88622 = $signed({1'h0, add_88518, array_index_88196[0]}) < $signed({1'h0, sel_88520}) ? {add_88518, array_index_88196[0]} : sel_88520;
  assign add_88624 = array_index_88397[11:3] + 9'h0bd;
  assign sel_88627 = $signed({1'h0, add_88522, array_index_88295[2:0]}) < $signed({1'h0, sel_88525}) ? {add_88522, array_index_88295[2:0]} : sel_88525;
  assign add_88629 = array_index_88400[11:3] + 9'h0bd;
  assign sel_88632 = $signed({1'h0, add_88527, array_index_88298[2:0]}) < $signed({1'h0, sel_88530}) ? {add_88527, array_index_88298[2:0]} : sel_88530;
  assign add_88634 = array_index_88499[11:1] + 11'h247;
  assign sel_88637 = $signed({1'h0, add_88532, array_index_88397[0]}) < $signed({1'h0, sel_88535}) ? {add_88532, array_index_88397[0]} : sel_88535;
  assign add_88639 = array_index_88502[11:1] + 11'h247;
  assign sel_88642 = $signed({1'h0, add_88537, array_index_88400[0]}) < $signed({1'h0, sel_88540}) ? {add_88537, array_index_88400[0]} : sel_88540;
  assign add_88667 = array_index_88601[11:0] + 12'h247;
  assign sel_88669 = $signed({1'h0, add_88565}) < $signed({1'h0, sel_88567}) ? add_88565 : sel_88567;
  assign add_88672 = array_index_88604[11:0] + 12'h247;
  assign sel_88674 = $signed({1'h0, add_88570}) < $signed({1'h0, sel_88572}) ? add_88570 : sel_88572;
  assign array_index_88703 = set1_unflattened[6'h12];
  assign array_index_88706 = set2_unflattened[6'h12];
  assign add_88710 = array_index_88295[11:1] + 11'h79d;
  assign sel_88712 = $signed({1'h0, add_88608, array_index_88193[0]}) < $signed({1'h0, sel_88610}) ? {add_88608, array_index_88193[0]} : sel_88610;
  assign add_88714 = array_index_88298[11:1] + 11'h79d;
  assign sel_88716 = $signed({1'h0, add_88612, array_index_88196[0]}) < $signed({1'h0, sel_88614}) ? {add_88612, array_index_88196[0]} : sel_88614;
  assign add_88718 = array_index_88397[11:1] + 11'h347;
  assign sel_88720 = $signed({1'h0, add_88616, array_index_88295[0]}) < $signed({1'h0, sel_88618}) ? {add_88616, array_index_88295[0]} : sel_88618;
  assign add_88722 = array_index_88400[11:1] + 11'h347;
  assign sel_88724 = $signed({1'h0, add_88620, array_index_88298[0]}) < $signed({1'h0, sel_88622}) ? {add_88620, array_index_88298[0]} : sel_88622;
  assign add_88726 = array_index_88499[11:3] + 9'h0bd;
  assign sel_88729 = $signed({1'h0, add_88624, array_index_88397[2:0]}) < $signed({1'h0, sel_88627}) ? {add_88624, array_index_88397[2:0]} : sel_88627;
  assign add_88731 = array_index_88502[11:3] + 9'h0bd;
  assign sel_88734 = $signed({1'h0, add_88629, array_index_88400[2:0]}) < $signed({1'h0, sel_88632}) ? {add_88629, array_index_88400[2:0]} : sel_88632;
  assign add_88736 = array_index_88601[11:1] + 11'h247;
  assign sel_88739 = $signed({1'h0, add_88634, array_index_88499[0]}) < $signed({1'h0, sel_88637}) ? {add_88634, array_index_88499[0]} : sel_88637;
  assign add_88741 = array_index_88604[11:1] + 11'h247;
  assign sel_88744 = $signed({1'h0, add_88639, array_index_88502[0]}) < $signed({1'h0, sel_88642}) ? {add_88639, array_index_88502[0]} : sel_88642;
  assign add_88769 = array_index_88703[11:0] + 12'h247;
  assign sel_88771 = $signed({1'h0, add_88667}) < $signed({1'h0, sel_88669}) ? add_88667 : sel_88669;
  assign add_88774 = array_index_88706[11:0] + 12'h247;
  assign sel_88776 = $signed({1'h0, add_88672}) < $signed({1'h0, sel_88674}) ? add_88672 : sel_88674;
  assign array_index_88805 = set1_unflattened[6'h13];
  assign array_index_88808 = set2_unflattened[6'h13];
  assign add_88812 = array_index_88397[11:1] + 11'h79d;
  assign sel_88814 = $signed({1'h0, add_88710, array_index_88295[0]}) < $signed({1'h0, sel_88712}) ? {add_88710, array_index_88295[0]} : sel_88712;
  assign add_88816 = array_index_88400[11:1] + 11'h79d;
  assign sel_88818 = $signed({1'h0, add_88714, array_index_88298[0]}) < $signed({1'h0, sel_88716}) ? {add_88714, array_index_88298[0]} : sel_88716;
  assign add_88820 = array_index_88499[11:1] + 11'h347;
  assign sel_88822 = $signed({1'h0, add_88718, array_index_88397[0]}) < $signed({1'h0, sel_88720}) ? {add_88718, array_index_88397[0]} : sel_88720;
  assign add_88824 = array_index_88502[11:1] + 11'h347;
  assign sel_88826 = $signed({1'h0, add_88722, array_index_88400[0]}) < $signed({1'h0, sel_88724}) ? {add_88722, array_index_88400[0]} : sel_88724;
  assign add_88828 = array_index_88601[11:3] + 9'h0bd;
  assign sel_88831 = $signed({1'h0, add_88726, array_index_88499[2:0]}) < $signed({1'h0, sel_88729}) ? {add_88726, array_index_88499[2:0]} : sel_88729;
  assign add_88833 = array_index_88604[11:3] + 9'h0bd;
  assign sel_88836 = $signed({1'h0, add_88731, array_index_88502[2:0]}) < $signed({1'h0, sel_88734}) ? {add_88731, array_index_88502[2:0]} : sel_88734;
  assign add_88838 = array_index_88703[11:1] + 11'h247;
  assign sel_88841 = $signed({1'h0, add_88736, array_index_88601[0]}) < $signed({1'h0, sel_88739}) ? {add_88736, array_index_88601[0]} : sel_88739;
  assign add_88843 = array_index_88706[11:1] + 11'h247;
  assign sel_88846 = $signed({1'h0, add_88741, array_index_88604[0]}) < $signed({1'h0, sel_88744}) ? {add_88741, array_index_88604[0]} : sel_88744;
  assign add_88871 = array_index_88805[11:0] + 12'h247;
  assign sel_88873 = $signed({1'h0, add_88769}) < $signed({1'h0, sel_88771}) ? add_88769 : sel_88771;
  assign add_88876 = array_index_88808[11:0] + 12'h247;
  assign sel_88878 = $signed({1'h0, add_88774}) < $signed({1'h0, sel_88776}) ? add_88774 : sel_88776;
  assign array_index_88907 = set1_unflattened[6'h14];
  assign array_index_88910 = set2_unflattened[6'h14];
  assign add_88914 = array_index_88499[11:1] + 11'h79d;
  assign sel_88916 = $signed({1'h0, add_88812, array_index_88397[0]}) < $signed({1'h0, sel_88814}) ? {add_88812, array_index_88397[0]} : sel_88814;
  assign add_88918 = array_index_88502[11:1] + 11'h79d;
  assign sel_88920 = $signed({1'h0, add_88816, array_index_88400[0]}) < $signed({1'h0, sel_88818}) ? {add_88816, array_index_88400[0]} : sel_88818;
  assign add_88922 = array_index_88601[11:1] + 11'h347;
  assign sel_88924 = $signed({1'h0, add_88820, array_index_88499[0]}) < $signed({1'h0, sel_88822}) ? {add_88820, array_index_88499[0]} : sel_88822;
  assign add_88926 = array_index_88604[11:1] + 11'h347;
  assign sel_88928 = $signed({1'h0, add_88824, array_index_88502[0]}) < $signed({1'h0, sel_88826}) ? {add_88824, array_index_88502[0]} : sel_88826;
  assign add_88930 = array_index_88703[11:3] + 9'h0bd;
  assign sel_88933 = $signed({1'h0, add_88828, array_index_88601[2:0]}) < $signed({1'h0, sel_88831}) ? {add_88828, array_index_88601[2:0]} : sel_88831;
  assign add_88935 = array_index_88706[11:3] + 9'h0bd;
  assign sel_88938 = $signed({1'h0, add_88833, array_index_88604[2:0]}) < $signed({1'h0, sel_88836}) ? {add_88833, array_index_88604[2:0]} : sel_88836;
  assign add_88940 = array_index_88805[11:1] + 11'h247;
  assign sel_88943 = $signed({1'h0, add_88838, array_index_88703[0]}) < $signed({1'h0, sel_88841}) ? {add_88838, array_index_88703[0]} : sel_88841;
  assign add_88945 = array_index_88808[11:1] + 11'h247;
  assign sel_88948 = $signed({1'h0, add_88843, array_index_88706[0]}) < $signed({1'h0, sel_88846}) ? {add_88843, array_index_88706[0]} : sel_88846;
  assign add_88973 = array_index_88907[11:0] + 12'h247;
  assign sel_88975 = $signed({1'h0, add_88871}) < $signed({1'h0, sel_88873}) ? add_88871 : sel_88873;
  assign add_88978 = array_index_88910[11:0] + 12'h247;
  assign sel_88980 = $signed({1'h0, add_88876}) < $signed({1'h0, sel_88878}) ? add_88876 : sel_88878;
  assign array_index_89009 = set1_unflattened[6'h15];
  assign array_index_89012 = set2_unflattened[6'h15];
  assign add_89016 = array_index_88601[11:1] + 11'h79d;
  assign sel_89018 = $signed({1'h0, add_88914, array_index_88499[0]}) < $signed({1'h0, sel_88916}) ? {add_88914, array_index_88499[0]} : sel_88916;
  assign add_89020 = array_index_88604[11:1] + 11'h79d;
  assign sel_89022 = $signed({1'h0, add_88918, array_index_88502[0]}) < $signed({1'h0, sel_88920}) ? {add_88918, array_index_88502[0]} : sel_88920;
  assign add_89024 = array_index_88703[11:1] + 11'h347;
  assign sel_89026 = $signed({1'h0, add_88922, array_index_88601[0]}) < $signed({1'h0, sel_88924}) ? {add_88922, array_index_88601[0]} : sel_88924;
  assign add_89028 = array_index_88706[11:1] + 11'h347;
  assign sel_89030 = $signed({1'h0, add_88926, array_index_88604[0]}) < $signed({1'h0, sel_88928}) ? {add_88926, array_index_88604[0]} : sel_88928;
  assign add_89032 = array_index_88805[11:3] + 9'h0bd;
  assign sel_89035 = $signed({1'h0, add_88930, array_index_88703[2:0]}) < $signed({1'h0, sel_88933}) ? {add_88930, array_index_88703[2:0]} : sel_88933;
  assign add_89037 = array_index_88808[11:3] + 9'h0bd;
  assign sel_89040 = $signed({1'h0, add_88935, array_index_88706[2:0]}) < $signed({1'h0, sel_88938}) ? {add_88935, array_index_88706[2:0]} : sel_88938;
  assign add_89042 = array_index_88907[11:1] + 11'h247;
  assign sel_89045 = $signed({1'h0, add_88940, array_index_88805[0]}) < $signed({1'h0, sel_88943}) ? {add_88940, array_index_88805[0]} : sel_88943;
  assign add_89047 = array_index_88910[11:1] + 11'h247;
  assign sel_89050 = $signed({1'h0, add_88945, array_index_88808[0]}) < $signed({1'h0, sel_88948}) ? {add_88945, array_index_88808[0]} : sel_88948;
  assign add_89075 = array_index_89009[11:0] + 12'h247;
  assign sel_89077 = $signed({1'h0, add_88973}) < $signed({1'h0, sel_88975}) ? add_88973 : sel_88975;
  assign add_89080 = array_index_89012[11:0] + 12'h247;
  assign sel_89082 = $signed({1'h0, add_88978}) < $signed({1'h0, sel_88980}) ? add_88978 : sel_88980;
  assign array_index_89111 = set1_unflattened[6'h16];
  assign array_index_89114 = set2_unflattened[6'h16];
  assign add_89118 = array_index_88703[11:1] + 11'h79d;
  assign sel_89120 = $signed({1'h0, add_89016, array_index_88601[0]}) < $signed({1'h0, sel_89018}) ? {add_89016, array_index_88601[0]} : sel_89018;
  assign add_89122 = array_index_88706[11:1] + 11'h79d;
  assign sel_89124 = $signed({1'h0, add_89020, array_index_88604[0]}) < $signed({1'h0, sel_89022}) ? {add_89020, array_index_88604[0]} : sel_89022;
  assign add_89126 = array_index_88805[11:1] + 11'h347;
  assign sel_89128 = $signed({1'h0, add_89024, array_index_88703[0]}) < $signed({1'h0, sel_89026}) ? {add_89024, array_index_88703[0]} : sel_89026;
  assign add_89130 = array_index_88808[11:1] + 11'h347;
  assign sel_89132 = $signed({1'h0, add_89028, array_index_88706[0]}) < $signed({1'h0, sel_89030}) ? {add_89028, array_index_88706[0]} : sel_89030;
  assign add_89134 = array_index_88907[11:3] + 9'h0bd;
  assign sel_89137 = $signed({1'h0, add_89032, array_index_88805[2:0]}) < $signed({1'h0, sel_89035}) ? {add_89032, array_index_88805[2:0]} : sel_89035;
  assign add_89139 = array_index_88910[11:3] + 9'h0bd;
  assign sel_89142 = $signed({1'h0, add_89037, array_index_88808[2:0]}) < $signed({1'h0, sel_89040}) ? {add_89037, array_index_88808[2:0]} : sel_89040;
  assign add_89144 = array_index_89009[11:1] + 11'h247;
  assign sel_89147 = $signed({1'h0, add_89042, array_index_88907[0]}) < $signed({1'h0, sel_89045}) ? {add_89042, array_index_88907[0]} : sel_89045;
  assign add_89149 = array_index_89012[11:1] + 11'h247;
  assign sel_89152 = $signed({1'h0, add_89047, array_index_88910[0]}) < $signed({1'h0, sel_89050}) ? {add_89047, array_index_88910[0]} : sel_89050;
  assign add_89177 = array_index_89111[11:0] + 12'h247;
  assign sel_89179 = $signed({1'h0, add_89075}) < $signed({1'h0, sel_89077}) ? add_89075 : sel_89077;
  assign add_89182 = array_index_89114[11:0] + 12'h247;
  assign sel_89184 = $signed({1'h0, add_89080}) < $signed({1'h0, sel_89082}) ? add_89080 : sel_89082;
  assign array_index_89213 = set1_unflattened[6'h17];
  assign array_index_89216 = set2_unflattened[6'h17];
  assign add_89220 = array_index_88805[11:1] + 11'h79d;
  assign sel_89222 = $signed({1'h0, add_89118, array_index_88703[0]}) < $signed({1'h0, sel_89120}) ? {add_89118, array_index_88703[0]} : sel_89120;
  assign add_89224 = array_index_88808[11:1] + 11'h79d;
  assign sel_89226 = $signed({1'h0, add_89122, array_index_88706[0]}) < $signed({1'h0, sel_89124}) ? {add_89122, array_index_88706[0]} : sel_89124;
  assign add_89228 = array_index_88907[11:1] + 11'h347;
  assign sel_89230 = $signed({1'h0, add_89126, array_index_88805[0]}) < $signed({1'h0, sel_89128}) ? {add_89126, array_index_88805[0]} : sel_89128;
  assign add_89232 = array_index_88910[11:1] + 11'h347;
  assign sel_89234 = $signed({1'h0, add_89130, array_index_88808[0]}) < $signed({1'h0, sel_89132}) ? {add_89130, array_index_88808[0]} : sel_89132;
  assign add_89236 = array_index_89009[11:3] + 9'h0bd;
  assign sel_89239 = $signed({1'h0, add_89134, array_index_88907[2:0]}) < $signed({1'h0, sel_89137}) ? {add_89134, array_index_88907[2:0]} : sel_89137;
  assign add_89241 = array_index_89012[11:3] + 9'h0bd;
  assign sel_89244 = $signed({1'h0, add_89139, array_index_88910[2:0]}) < $signed({1'h0, sel_89142}) ? {add_89139, array_index_88910[2:0]} : sel_89142;
  assign add_89246 = array_index_89111[11:1] + 11'h247;
  assign sel_89249 = $signed({1'h0, add_89144, array_index_89009[0]}) < $signed({1'h0, sel_89147}) ? {add_89144, array_index_89009[0]} : sel_89147;
  assign add_89251 = array_index_89114[11:1] + 11'h247;
  assign sel_89254 = $signed({1'h0, add_89149, array_index_89012[0]}) < $signed({1'h0, sel_89152}) ? {add_89149, array_index_89012[0]} : sel_89152;
  assign add_89279 = array_index_89213[11:0] + 12'h247;
  assign sel_89281 = $signed({1'h0, add_89177}) < $signed({1'h0, sel_89179}) ? add_89177 : sel_89179;
  assign add_89284 = array_index_89216[11:0] + 12'h247;
  assign sel_89286 = $signed({1'h0, add_89182}) < $signed({1'h0, sel_89184}) ? add_89182 : sel_89184;
  assign array_index_89315 = set1_unflattened[6'h18];
  assign array_index_89318 = set2_unflattened[6'h18];
  assign add_89322 = array_index_88907[11:1] + 11'h79d;
  assign sel_89324 = $signed({1'h0, add_89220, array_index_88805[0]}) < $signed({1'h0, sel_89222}) ? {add_89220, array_index_88805[0]} : sel_89222;
  assign add_89326 = array_index_88910[11:1] + 11'h79d;
  assign sel_89328 = $signed({1'h0, add_89224, array_index_88808[0]}) < $signed({1'h0, sel_89226}) ? {add_89224, array_index_88808[0]} : sel_89226;
  assign add_89330 = array_index_89009[11:1] + 11'h347;
  assign sel_89332 = $signed({1'h0, add_89228, array_index_88907[0]}) < $signed({1'h0, sel_89230}) ? {add_89228, array_index_88907[0]} : sel_89230;
  assign add_89334 = array_index_89012[11:1] + 11'h347;
  assign sel_89336 = $signed({1'h0, add_89232, array_index_88910[0]}) < $signed({1'h0, sel_89234}) ? {add_89232, array_index_88910[0]} : sel_89234;
  assign add_89338 = array_index_89111[11:3] + 9'h0bd;
  assign sel_89341 = $signed({1'h0, add_89236, array_index_89009[2:0]}) < $signed({1'h0, sel_89239}) ? {add_89236, array_index_89009[2:0]} : sel_89239;
  assign add_89343 = array_index_89114[11:3] + 9'h0bd;
  assign sel_89346 = $signed({1'h0, add_89241, array_index_89012[2:0]}) < $signed({1'h0, sel_89244}) ? {add_89241, array_index_89012[2:0]} : sel_89244;
  assign add_89348 = array_index_89213[11:1] + 11'h247;
  assign sel_89351 = $signed({1'h0, add_89246, array_index_89111[0]}) < $signed({1'h0, sel_89249}) ? {add_89246, array_index_89111[0]} : sel_89249;
  assign add_89353 = array_index_89216[11:1] + 11'h247;
  assign sel_89356 = $signed({1'h0, add_89251, array_index_89114[0]}) < $signed({1'h0, sel_89254}) ? {add_89251, array_index_89114[0]} : sel_89254;
  assign add_89381 = array_index_89315[11:0] + 12'h247;
  assign sel_89383 = $signed({1'h0, add_89279}) < $signed({1'h0, sel_89281}) ? add_89279 : sel_89281;
  assign add_89386 = array_index_89318[11:0] + 12'h247;
  assign sel_89388 = $signed({1'h0, add_89284}) < $signed({1'h0, sel_89286}) ? add_89284 : sel_89286;
  assign array_index_89417 = set1_unflattened[6'h19];
  assign array_index_89420 = set2_unflattened[6'h19];
  assign add_89424 = array_index_89009[11:1] + 11'h79d;
  assign sel_89426 = $signed({1'h0, add_89322, array_index_88907[0]}) < $signed({1'h0, sel_89324}) ? {add_89322, array_index_88907[0]} : sel_89324;
  assign add_89428 = array_index_89012[11:1] + 11'h79d;
  assign sel_89430 = $signed({1'h0, add_89326, array_index_88910[0]}) < $signed({1'h0, sel_89328}) ? {add_89326, array_index_88910[0]} : sel_89328;
  assign add_89432 = array_index_89111[11:1] + 11'h347;
  assign sel_89434 = $signed({1'h0, add_89330, array_index_89009[0]}) < $signed({1'h0, sel_89332}) ? {add_89330, array_index_89009[0]} : sel_89332;
  assign add_89436 = array_index_89114[11:1] + 11'h347;
  assign sel_89438 = $signed({1'h0, add_89334, array_index_89012[0]}) < $signed({1'h0, sel_89336}) ? {add_89334, array_index_89012[0]} : sel_89336;
  assign add_89440 = array_index_89213[11:3] + 9'h0bd;
  assign sel_89443 = $signed({1'h0, add_89338, array_index_89111[2:0]}) < $signed({1'h0, sel_89341}) ? {add_89338, array_index_89111[2:0]} : sel_89341;
  assign add_89445 = array_index_89216[11:3] + 9'h0bd;
  assign sel_89448 = $signed({1'h0, add_89343, array_index_89114[2:0]}) < $signed({1'h0, sel_89346}) ? {add_89343, array_index_89114[2:0]} : sel_89346;
  assign add_89450 = array_index_89315[11:1] + 11'h247;
  assign sel_89453 = $signed({1'h0, add_89348, array_index_89213[0]}) < $signed({1'h0, sel_89351}) ? {add_89348, array_index_89213[0]} : sel_89351;
  assign add_89455 = array_index_89318[11:1] + 11'h247;
  assign sel_89458 = $signed({1'h0, add_89353, array_index_89216[0]}) < $signed({1'h0, sel_89356}) ? {add_89353, array_index_89216[0]} : sel_89356;
  assign add_89483 = array_index_89417[11:0] + 12'h247;
  assign sel_89485 = $signed({1'h0, add_89381}) < $signed({1'h0, sel_89383}) ? add_89381 : sel_89383;
  assign add_89488 = array_index_89420[11:0] + 12'h247;
  assign sel_89490 = $signed({1'h0, add_89386}) < $signed({1'h0, sel_89388}) ? add_89386 : sel_89388;
  assign array_index_89519 = set1_unflattened[6'h1a];
  assign array_index_89522 = set2_unflattened[6'h1a];
  assign add_89526 = array_index_89111[11:1] + 11'h79d;
  assign sel_89528 = $signed({1'h0, add_89424, array_index_89009[0]}) < $signed({1'h0, sel_89426}) ? {add_89424, array_index_89009[0]} : sel_89426;
  assign add_89530 = array_index_89114[11:1] + 11'h79d;
  assign sel_89532 = $signed({1'h0, add_89428, array_index_89012[0]}) < $signed({1'h0, sel_89430}) ? {add_89428, array_index_89012[0]} : sel_89430;
  assign add_89534 = array_index_89213[11:1] + 11'h347;
  assign sel_89536 = $signed({1'h0, add_89432, array_index_89111[0]}) < $signed({1'h0, sel_89434}) ? {add_89432, array_index_89111[0]} : sel_89434;
  assign add_89538 = array_index_89216[11:1] + 11'h347;
  assign sel_89540 = $signed({1'h0, add_89436, array_index_89114[0]}) < $signed({1'h0, sel_89438}) ? {add_89436, array_index_89114[0]} : sel_89438;
  assign add_89542 = array_index_89315[11:3] + 9'h0bd;
  assign sel_89545 = $signed({1'h0, add_89440, array_index_89213[2:0]}) < $signed({1'h0, sel_89443}) ? {add_89440, array_index_89213[2:0]} : sel_89443;
  assign add_89547 = array_index_89318[11:3] + 9'h0bd;
  assign sel_89550 = $signed({1'h0, add_89445, array_index_89216[2:0]}) < $signed({1'h0, sel_89448}) ? {add_89445, array_index_89216[2:0]} : sel_89448;
  assign add_89552 = array_index_89417[11:1] + 11'h247;
  assign sel_89555 = $signed({1'h0, add_89450, array_index_89315[0]}) < $signed({1'h0, sel_89453}) ? {add_89450, array_index_89315[0]} : sel_89453;
  assign add_89557 = array_index_89420[11:1] + 11'h247;
  assign sel_89560 = $signed({1'h0, add_89455, array_index_89318[0]}) < $signed({1'h0, sel_89458}) ? {add_89455, array_index_89318[0]} : sel_89458;
  assign add_89585 = array_index_89519[11:0] + 12'h247;
  assign sel_89587 = $signed({1'h0, add_89483}) < $signed({1'h0, sel_89485}) ? add_89483 : sel_89485;
  assign add_89590 = array_index_89522[11:0] + 12'h247;
  assign sel_89592 = $signed({1'h0, add_89488}) < $signed({1'h0, sel_89490}) ? add_89488 : sel_89490;
  assign array_index_89621 = set1_unflattened[6'h1b];
  assign array_index_89624 = set2_unflattened[6'h1b];
  assign add_89628 = array_index_89213[11:1] + 11'h79d;
  assign sel_89630 = $signed({1'h0, add_89526, array_index_89111[0]}) < $signed({1'h0, sel_89528}) ? {add_89526, array_index_89111[0]} : sel_89528;
  assign add_89632 = array_index_89216[11:1] + 11'h79d;
  assign sel_89634 = $signed({1'h0, add_89530, array_index_89114[0]}) < $signed({1'h0, sel_89532}) ? {add_89530, array_index_89114[0]} : sel_89532;
  assign add_89636 = array_index_89315[11:1] + 11'h347;
  assign sel_89638 = $signed({1'h0, add_89534, array_index_89213[0]}) < $signed({1'h0, sel_89536}) ? {add_89534, array_index_89213[0]} : sel_89536;
  assign add_89640 = array_index_89318[11:1] + 11'h347;
  assign sel_89642 = $signed({1'h0, add_89538, array_index_89216[0]}) < $signed({1'h0, sel_89540}) ? {add_89538, array_index_89216[0]} : sel_89540;
  assign add_89644 = array_index_89417[11:3] + 9'h0bd;
  assign sel_89647 = $signed({1'h0, add_89542, array_index_89315[2:0]}) < $signed({1'h0, sel_89545}) ? {add_89542, array_index_89315[2:0]} : sel_89545;
  assign add_89649 = array_index_89420[11:3] + 9'h0bd;
  assign sel_89652 = $signed({1'h0, add_89547, array_index_89318[2:0]}) < $signed({1'h0, sel_89550}) ? {add_89547, array_index_89318[2:0]} : sel_89550;
  assign add_89654 = array_index_89519[11:1] + 11'h247;
  assign sel_89657 = $signed({1'h0, add_89552, array_index_89417[0]}) < $signed({1'h0, sel_89555}) ? {add_89552, array_index_89417[0]} : sel_89555;
  assign add_89659 = array_index_89522[11:1] + 11'h247;
  assign sel_89662 = $signed({1'h0, add_89557, array_index_89420[0]}) < $signed({1'h0, sel_89560}) ? {add_89557, array_index_89420[0]} : sel_89560;
  assign add_89687 = array_index_89621[11:0] + 12'h247;
  assign sel_89689 = $signed({1'h0, add_89585}) < $signed({1'h0, sel_89587}) ? add_89585 : sel_89587;
  assign add_89692 = array_index_89624[11:0] + 12'h247;
  assign sel_89694 = $signed({1'h0, add_89590}) < $signed({1'h0, sel_89592}) ? add_89590 : sel_89592;
  assign array_index_89723 = set1_unflattened[6'h1c];
  assign array_index_89726 = set2_unflattened[6'h1c];
  assign add_89730 = array_index_89315[11:1] + 11'h79d;
  assign sel_89732 = $signed({1'h0, add_89628, array_index_89213[0]}) < $signed({1'h0, sel_89630}) ? {add_89628, array_index_89213[0]} : sel_89630;
  assign add_89734 = array_index_89318[11:1] + 11'h79d;
  assign sel_89736 = $signed({1'h0, add_89632, array_index_89216[0]}) < $signed({1'h0, sel_89634}) ? {add_89632, array_index_89216[0]} : sel_89634;
  assign add_89738 = array_index_89417[11:1] + 11'h347;
  assign sel_89740 = $signed({1'h0, add_89636, array_index_89315[0]}) < $signed({1'h0, sel_89638}) ? {add_89636, array_index_89315[0]} : sel_89638;
  assign add_89742 = array_index_89420[11:1] + 11'h347;
  assign sel_89744 = $signed({1'h0, add_89640, array_index_89318[0]}) < $signed({1'h0, sel_89642}) ? {add_89640, array_index_89318[0]} : sel_89642;
  assign add_89746 = array_index_89519[11:3] + 9'h0bd;
  assign sel_89749 = $signed({1'h0, add_89644, array_index_89417[2:0]}) < $signed({1'h0, sel_89647}) ? {add_89644, array_index_89417[2:0]} : sel_89647;
  assign add_89751 = array_index_89522[11:3] + 9'h0bd;
  assign sel_89754 = $signed({1'h0, add_89649, array_index_89420[2:0]}) < $signed({1'h0, sel_89652}) ? {add_89649, array_index_89420[2:0]} : sel_89652;
  assign add_89756 = array_index_89621[11:1] + 11'h247;
  assign sel_89759 = $signed({1'h0, add_89654, array_index_89519[0]}) < $signed({1'h0, sel_89657}) ? {add_89654, array_index_89519[0]} : sel_89657;
  assign add_89761 = array_index_89624[11:1] + 11'h247;
  assign sel_89764 = $signed({1'h0, add_89659, array_index_89522[0]}) < $signed({1'h0, sel_89662}) ? {add_89659, array_index_89522[0]} : sel_89662;
  assign add_89789 = array_index_89723[11:0] + 12'h247;
  assign sel_89791 = $signed({1'h0, add_89687}) < $signed({1'h0, sel_89689}) ? add_89687 : sel_89689;
  assign add_89794 = array_index_89726[11:0] + 12'h247;
  assign sel_89796 = $signed({1'h0, add_89692}) < $signed({1'h0, sel_89694}) ? add_89692 : sel_89694;
  assign array_index_89825 = set1_unflattened[6'h1d];
  assign array_index_89828 = set2_unflattened[6'h1d];
  assign add_89832 = array_index_89417[11:1] + 11'h79d;
  assign sel_89834 = $signed({1'h0, add_89730, array_index_89315[0]}) < $signed({1'h0, sel_89732}) ? {add_89730, array_index_89315[0]} : sel_89732;
  assign add_89836 = array_index_89420[11:1] + 11'h79d;
  assign sel_89838 = $signed({1'h0, add_89734, array_index_89318[0]}) < $signed({1'h0, sel_89736}) ? {add_89734, array_index_89318[0]} : sel_89736;
  assign add_89840 = array_index_89519[11:1] + 11'h347;
  assign sel_89842 = $signed({1'h0, add_89738, array_index_89417[0]}) < $signed({1'h0, sel_89740}) ? {add_89738, array_index_89417[0]} : sel_89740;
  assign add_89844 = array_index_89522[11:1] + 11'h347;
  assign sel_89846 = $signed({1'h0, add_89742, array_index_89420[0]}) < $signed({1'h0, sel_89744}) ? {add_89742, array_index_89420[0]} : sel_89744;
  assign add_89848 = array_index_89621[11:3] + 9'h0bd;
  assign sel_89851 = $signed({1'h0, add_89746, array_index_89519[2:0]}) < $signed({1'h0, sel_89749}) ? {add_89746, array_index_89519[2:0]} : sel_89749;
  assign add_89853 = array_index_89624[11:3] + 9'h0bd;
  assign sel_89856 = $signed({1'h0, add_89751, array_index_89522[2:0]}) < $signed({1'h0, sel_89754}) ? {add_89751, array_index_89522[2:0]} : sel_89754;
  assign add_89858 = array_index_89723[11:1] + 11'h247;
  assign sel_89861 = $signed({1'h0, add_89756, array_index_89621[0]}) < $signed({1'h0, sel_89759}) ? {add_89756, array_index_89621[0]} : sel_89759;
  assign add_89863 = array_index_89726[11:1] + 11'h247;
  assign sel_89866 = $signed({1'h0, add_89761, array_index_89624[0]}) < $signed({1'h0, sel_89764}) ? {add_89761, array_index_89624[0]} : sel_89764;
  assign add_89891 = array_index_89825[11:0] + 12'h247;
  assign sel_89893 = $signed({1'h0, add_89789}) < $signed({1'h0, sel_89791}) ? add_89789 : sel_89791;
  assign add_89896 = array_index_89828[11:0] + 12'h247;
  assign sel_89898 = $signed({1'h0, add_89794}) < $signed({1'h0, sel_89796}) ? add_89794 : sel_89796;
  assign array_index_89927 = set1_unflattened[6'h1e];
  assign array_index_89930 = set2_unflattened[6'h1e];
  assign add_89934 = array_index_89519[11:1] + 11'h79d;
  assign sel_89936 = $signed({1'h0, add_89832, array_index_89417[0]}) < $signed({1'h0, sel_89834}) ? {add_89832, array_index_89417[0]} : sel_89834;
  assign add_89938 = array_index_89522[11:1] + 11'h79d;
  assign sel_89940 = $signed({1'h0, add_89836, array_index_89420[0]}) < $signed({1'h0, sel_89838}) ? {add_89836, array_index_89420[0]} : sel_89838;
  assign add_89942 = array_index_89621[11:1] + 11'h347;
  assign sel_89944 = $signed({1'h0, add_89840, array_index_89519[0]}) < $signed({1'h0, sel_89842}) ? {add_89840, array_index_89519[0]} : sel_89842;
  assign add_89946 = array_index_89624[11:1] + 11'h347;
  assign sel_89948 = $signed({1'h0, add_89844, array_index_89522[0]}) < $signed({1'h0, sel_89846}) ? {add_89844, array_index_89522[0]} : sel_89846;
  assign add_89950 = array_index_89723[11:3] + 9'h0bd;
  assign sel_89953 = $signed({1'h0, add_89848, array_index_89621[2:0]}) < $signed({1'h0, sel_89851}) ? {add_89848, array_index_89621[2:0]} : sel_89851;
  assign add_89955 = array_index_89726[11:3] + 9'h0bd;
  assign sel_89958 = $signed({1'h0, add_89853, array_index_89624[2:0]}) < $signed({1'h0, sel_89856}) ? {add_89853, array_index_89624[2:0]} : sel_89856;
  assign add_89960 = array_index_89825[11:1] + 11'h247;
  assign sel_89963 = $signed({1'h0, add_89858, array_index_89723[0]}) < $signed({1'h0, sel_89861}) ? {add_89858, array_index_89723[0]} : sel_89861;
  assign add_89965 = array_index_89828[11:1] + 11'h247;
  assign sel_89968 = $signed({1'h0, add_89863, array_index_89726[0]}) < $signed({1'h0, sel_89866}) ? {add_89863, array_index_89726[0]} : sel_89866;
  assign add_89993 = array_index_89927[11:0] + 12'h247;
  assign sel_89995 = $signed({1'h0, add_89891}) < $signed({1'h0, sel_89893}) ? add_89891 : sel_89893;
  assign add_89998 = array_index_89930[11:0] + 12'h247;
  assign sel_90000 = $signed({1'h0, add_89896}) < $signed({1'h0, sel_89898}) ? add_89896 : sel_89898;
  assign array_index_90029 = set1_unflattened[6'h1f];
  assign array_index_90032 = set2_unflattened[6'h1f];
  assign add_90036 = array_index_89621[11:1] + 11'h79d;
  assign sel_90038 = $signed({1'h0, add_89934, array_index_89519[0]}) < $signed({1'h0, sel_89936}) ? {add_89934, array_index_89519[0]} : sel_89936;
  assign add_90040 = array_index_89624[11:1] + 11'h79d;
  assign sel_90042 = $signed({1'h0, add_89938, array_index_89522[0]}) < $signed({1'h0, sel_89940}) ? {add_89938, array_index_89522[0]} : sel_89940;
  assign add_90044 = array_index_89723[11:1] + 11'h347;
  assign sel_90046 = $signed({1'h0, add_89942, array_index_89621[0]}) < $signed({1'h0, sel_89944}) ? {add_89942, array_index_89621[0]} : sel_89944;
  assign add_90048 = array_index_89726[11:1] + 11'h347;
  assign sel_90050 = $signed({1'h0, add_89946, array_index_89624[0]}) < $signed({1'h0, sel_89948}) ? {add_89946, array_index_89624[0]} : sel_89948;
  assign add_90052 = array_index_89825[11:3] + 9'h0bd;
  assign sel_90055 = $signed({1'h0, add_89950, array_index_89723[2:0]}) < $signed({1'h0, sel_89953}) ? {add_89950, array_index_89723[2:0]} : sel_89953;
  assign add_90057 = array_index_89828[11:3] + 9'h0bd;
  assign sel_90060 = $signed({1'h0, add_89955, array_index_89726[2:0]}) < $signed({1'h0, sel_89958}) ? {add_89955, array_index_89726[2:0]} : sel_89958;
  assign add_90062 = array_index_89927[11:1] + 11'h247;
  assign sel_90065 = $signed({1'h0, add_89960, array_index_89825[0]}) < $signed({1'h0, sel_89963}) ? {add_89960, array_index_89825[0]} : sel_89963;
  assign add_90067 = array_index_89930[11:1] + 11'h247;
  assign sel_90070 = $signed({1'h0, add_89965, array_index_89828[0]}) < $signed({1'h0, sel_89968}) ? {add_89965, array_index_89828[0]} : sel_89968;
  assign add_90095 = array_index_90029[11:0] + 12'h247;
  assign sel_90097 = $signed({1'h0, add_89993}) < $signed({1'h0, sel_89995}) ? add_89993 : sel_89995;
  assign add_90100 = array_index_90032[11:0] + 12'h247;
  assign sel_90102 = $signed({1'h0, add_89998}) < $signed({1'h0, sel_90000}) ? add_89998 : sel_90000;
  assign array_index_90131 = set1_unflattened[6'h20];
  assign array_index_90134 = set2_unflattened[6'h20];
  assign add_90138 = array_index_89723[11:1] + 11'h79d;
  assign sel_90140 = $signed({1'h0, add_90036, array_index_89621[0]}) < $signed({1'h0, sel_90038}) ? {add_90036, array_index_89621[0]} : sel_90038;
  assign add_90142 = array_index_89726[11:1] + 11'h79d;
  assign sel_90144 = $signed({1'h0, add_90040, array_index_89624[0]}) < $signed({1'h0, sel_90042}) ? {add_90040, array_index_89624[0]} : sel_90042;
  assign add_90146 = array_index_89825[11:1] + 11'h347;
  assign sel_90148 = $signed({1'h0, add_90044, array_index_89723[0]}) < $signed({1'h0, sel_90046}) ? {add_90044, array_index_89723[0]} : sel_90046;
  assign add_90150 = array_index_89828[11:1] + 11'h347;
  assign sel_90152 = $signed({1'h0, add_90048, array_index_89726[0]}) < $signed({1'h0, sel_90050}) ? {add_90048, array_index_89726[0]} : sel_90050;
  assign add_90154 = array_index_89927[11:3] + 9'h0bd;
  assign sel_90157 = $signed({1'h0, add_90052, array_index_89825[2:0]}) < $signed({1'h0, sel_90055}) ? {add_90052, array_index_89825[2:0]} : sel_90055;
  assign add_90159 = array_index_89930[11:3] + 9'h0bd;
  assign sel_90162 = $signed({1'h0, add_90057, array_index_89828[2:0]}) < $signed({1'h0, sel_90060}) ? {add_90057, array_index_89828[2:0]} : sel_90060;
  assign add_90164 = array_index_90029[11:1] + 11'h247;
  assign sel_90167 = $signed({1'h0, add_90062, array_index_89927[0]}) < $signed({1'h0, sel_90065}) ? {add_90062, array_index_89927[0]} : sel_90065;
  assign add_90169 = array_index_90032[11:1] + 11'h247;
  assign sel_90172 = $signed({1'h0, add_90067, array_index_89930[0]}) < $signed({1'h0, sel_90070}) ? {add_90067, array_index_89930[0]} : sel_90070;
  assign add_90197 = array_index_90131[11:0] + 12'h247;
  assign sel_90199 = $signed({1'h0, add_90095}) < $signed({1'h0, sel_90097}) ? add_90095 : sel_90097;
  assign add_90202 = array_index_90134[11:0] + 12'h247;
  assign sel_90204 = $signed({1'h0, add_90100}) < $signed({1'h0, sel_90102}) ? add_90100 : sel_90102;
  assign array_index_90233 = set1_unflattened[6'h21];
  assign array_index_90236 = set2_unflattened[6'h21];
  assign add_90240 = array_index_89825[11:1] + 11'h79d;
  assign sel_90242 = $signed({1'h0, add_90138, array_index_89723[0]}) < $signed({1'h0, sel_90140}) ? {add_90138, array_index_89723[0]} : sel_90140;
  assign add_90244 = array_index_89828[11:1] + 11'h79d;
  assign sel_90246 = $signed({1'h0, add_90142, array_index_89726[0]}) < $signed({1'h0, sel_90144}) ? {add_90142, array_index_89726[0]} : sel_90144;
  assign add_90248 = array_index_89927[11:1] + 11'h347;
  assign sel_90250 = $signed({1'h0, add_90146, array_index_89825[0]}) < $signed({1'h0, sel_90148}) ? {add_90146, array_index_89825[0]} : sel_90148;
  assign add_90252 = array_index_89930[11:1] + 11'h347;
  assign sel_90254 = $signed({1'h0, add_90150, array_index_89828[0]}) < $signed({1'h0, sel_90152}) ? {add_90150, array_index_89828[0]} : sel_90152;
  assign add_90256 = array_index_90029[11:3] + 9'h0bd;
  assign sel_90259 = $signed({1'h0, add_90154, array_index_89927[2:0]}) < $signed({1'h0, sel_90157}) ? {add_90154, array_index_89927[2:0]} : sel_90157;
  assign add_90261 = array_index_90032[11:3] + 9'h0bd;
  assign sel_90264 = $signed({1'h0, add_90159, array_index_89930[2:0]}) < $signed({1'h0, sel_90162}) ? {add_90159, array_index_89930[2:0]} : sel_90162;
  assign add_90266 = array_index_90131[11:1] + 11'h247;
  assign sel_90269 = $signed({1'h0, add_90164, array_index_90029[0]}) < $signed({1'h0, sel_90167}) ? {add_90164, array_index_90029[0]} : sel_90167;
  assign add_90271 = array_index_90134[11:1] + 11'h247;
  assign sel_90274 = $signed({1'h0, add_90169, array_index_90032[0]}) < $signed({1'h0, sel_90172}) ? {add_90169, array_index_90032[0]} : sel_90172;
  assign add_90299 = array_index_90233[11:0] + 12'h247;
  assign sel_90301 = $signed({1'h0, add_90197}) < $signed({1'h0, sel_90199}) ? add_90197 : sel_90199;
  assign add_90304 = array_index_90236[11:0] + 12'h247;
  assign sel_90306 = $signed({1'h0, add_90202}) < $signed({1'h0, sel_90204}) ? add_90202 : sel_90204;
  assign array_index_90335 = set1_unflattened[6'h22];
  assign array_index_90338 = set2_unflattened[6'h22];
  assign add_90342 = array_index_89927[11:1] + 11'h79d;
  assign sel_90344 = $signed({1'h0, add_90240, array_index_89825[0]}) < $signed({1'h0, sel_90242}) ? {add_90240, array_index_89825[0]} : sel_90242;
  assign add_90346 = array_index_89930[11:1] + 11'h79d;
  assign sel_90348 = $signed({1'h0, add_90244, array_index_89828[0]}) < $signed({1'h0, sel_90246}) ? {add_90244, array_index_89828[0]} : sel_90246;
  assign add_90350 = array_index_90029[11:1] + 11'h347;
  assign sel_90352 = $signed({1'h0, add_90248, array_index_89927[0]}) < $signed({1'h0, sel_90250}) ? {add_90248, array_index_89927[0]} : sel_90250;
  assign add_90354 = array_index_90032[11:1] + 11'h347;
  assign sel_90356 = $signed({1'h0, add_90252, array_index_89930[0]}) < $signed({1'h0, sel_90254}) ? {add_90252, array_index_89930[0]} : sel_90254;
  assign add_90358 = array_index_90131[11:3] + 9'h0bd;
  assign sel_90361 = $signed({1'h0, add_90256, array_index_90029[2:0]}) < $signed({1'h0, sel_90259}) ? {add_90256, array_index_90029[2:0]} : sel_90259;
  assign add_90363 = array_index_90134[11:3] + 9'h0bd;
  assign sel_90366 = $signed({1'h0, add_90261, array_index_90032[2:0]}) < $signed({1'h0, sel_90264}) ? {add_90261, array_index_90032[2:0]} : sel_90264;
  assign add_90368 = array_index_90233[11:1] + 11'h247;
  assign sel_90371 = $signed({1'h0, add_90266, array_index_90131[0]}) < $signed({1'h0, sel_90269}) ? {add_90266, array_index_90131[0]} : sel_90269;
  assign add_90373 = array_index_90236[11:1] + 11'h247;
  assign sel_90376 = $signed({1'h0, add_90271, array_index_90134[0]}) < $signed({1'h0, sel_90274}) ? {add_90271, array_index_90134[0]} : sel_90274;
  assign add_90401 = array_index_90335[11:0] + 12'h247;
  assign sel_90403 = $signed({1'h0, add_90299}) < $signed({1'h0, sel_90301}) ? add_90299 : sel_90301;
  assign add_90406 = array_index_90338[11:0] + 12'h247;
  assign sel_90408 = $signed({1'h0, add_90304}) < $signed({1'h0, sel_90306}) ? add_90304 : sel_90306;
  assign array_index_90437 = set1_unflattened[6'h23];
  assign array_index_90440 = set2_unflattened[6'h23];
  assign add_90444 = array_index_90029[11:1] + 11'h79d;
  assign sel_90446 = $signed({1'h0, add_90342, array_index_89927[0]}) < $signed({1'h0, sel_90344}) ? {add_90342, array_index_89927[0]} : sel_90344;
  assign add_90448 = array_index_90032[11:1] + 11'h79d;
  assign sel_90450 = $signed({1'h0, add_90346, array_index_89930[0]}) < $signed({1'h0, sel_90348}) ? {add_90346, array_index_89930[0]} : sel_90348;
  assign add_90452 = array_index_90131[11:1] + 11'h347;
  assign sel_90454 = $signed({1'h0, add_90350, array_index_90029[0]}) < $signed({1'h0, sel_90352}) ? {add_90350, array_index_90029[0]} : sel_90352;
  assign add_90456 = array_index_90134[11:1] + 11'h347;
  assign sel_90458 = $signed({1'h0, add_90354, array_index_90032[0]}) < $signed({1'h0, sel_90356}) ? {add_90354, array_index_90032[0]} : sel_90356;
  assign add_90460 = array_index_90233[11:3] + 9'h0bd;
  assign sel_90463 = $signed({1'h0, add_90358, array_index_90131[2:0]}) < $signed({1'h0, sel_90361}) ? {add_90358, array_index_90131[2:0]} : sel_90361;
  assign add_90465 = array_index_90236[11:3] + 9'h0bd;
  assign sel_90468 = $signed({1'h0, add_90363, array_index_90134[2:0]}) < $signed({1'h0, sel_90366}) ? {add_90363, array_index_90134[2:0]} : sel_90366;
  assign add_90470 = array_index_90335[11:1] + 11'h247;
  assign sel_90473 = $signed({1'h0, add_90368, array_index_90233[0]}) < $signed({1'h0, sel_90371}) ? {add_90368, array_index_90233[0]} : sel_90371;
  assign add_90475 = array_index_90338[11:1] + 11'h247;
  assign sel_90478 = $signed({1'h0, add_90373, array_index_90236[0]}) < $signed({1'h0, sel_90376}) ? {add_90373, array_index_90236[0]} : sel_90376;
  assign add_90503 = array_index_90437[11:0] + 12'h247;
  assign sel_90505 = $signed({1'h0, add_90401}) < $signed({1'h0, sel_90403}) ? add_90401 : sel_90403;
  assign add_90508 = array_index_90440[11:0] + 12'h247;
  assign sel_90510 = $signed({1'h0, add_90406}) < $signed({1'h0, sel_90408}) ? add_90406 : sel_90408;
  assign array_index_90539 = set1_unflattened[6'h24];
  assign array_index_90542 = set2_unflattened[6'h24];
  assign add_90546 = array_index_90131[11:1] + 11'h79d;
  assign sel_90548 = $signed({1'h0, add_90444, array_index_90029[0]}) < $signed({1'h0, sel_90446}) ? {add_90444, array_index_90029[0]} : sel_90446;
  assign add_90550 = array_index_90134[11:1] + 11'h79d;
  assign sel_90552 = $signed({1'h0, add_90448, array_index_90032[0]}) < $signed({1'h0, sel_90450}) ? {add_90448, array_index_90032[0]} : sel_90450;
  assign add_90554 = array_index_90233[11:1] + 11'h347;
  assign sel_90556 = $signed({1'h0, add_90452, array_index_90131[0]}) < $signed({1'h0, sel_90454}) ? {add_90452, array_index_90131[0]} : sel_90454;
  assign add_90558 = array_index_90236[11:1] + 11'h347;
  assign sel_90560 = $signed({1'h0, add_90456, array_index_90134[0]}) < $signed({1'h0, sel_90458}) ? {add_90456, array_index_90134[0]} : sel_90458;
  assign add_90562 = array_index_90335[11:3] + 9'h0bd;
  assign sel_90565 = $signed({1'h0, add_90460, array_index_90233[2:0]}) < $signed({1'h0, sel_90463}) ? {add_90460, array_index_90233[2:0]} : sel_90463;
  assign add_90567 = array_index_90338[11:3] + 9'h0bd;
  assign sel_90570 = $signed({1'h0, add_90465, array_index_90236[2:0]}) < $signed({1'h0, sel_90468}) ? {add_90465, array_index_90236[2:0]} : sel_90468;
  assign add_90572 = array_index_90437[11:1] + 11'h247;
  assign sel_90575 = $signed({1'h0, add_90470, array_index_90335[0]}) < $signed({1'h0, sel_90473}) ? {add_90470, array_index_90335[0]} : sel_90473;
  assign add_90577 = array_index_90440[11:1] + 11'h247;
  assign sel_90580 = $signed({1'h0, add_90475, array_index_90338[0]}) < $signed({1'h0, sel_90478}) ? {add_90475, array_index_90338[0]} : sel_90478;
  assign add_90605 = array_index_90539[11:0] + 12'h247;
  assign sel_90607 = $signed({1'h0, add_90503}) < $signed({1'h0, sel_90505}) ? add_90503 : sel_90505;
  assign add_90610 = array_index_90542[11:0] + 12'h247;
  assign sel_90612 = $signed({1'h0, add_90508}) < $signed({1'h0, sel_90510}) ? add_90508 : sel_90510;
  assign array_index_90641 = set1_unflattened[6'h25];
  assign array_index_90644 = set2_unflattened[6'h25];
  assign add_90648 = array_index_90233[11:1] + 11'h79d;
  assign sel_90650 = $signed({1'h0, add_90546, array_index_90131[0]}) < $signed({1'h0, sel_90548}) ? {add_90546, array_index_90131[0]} : sel_90548;
  assign add_90652 = array_index_90236[11:1] + 11'h79d;
  assign sel_90654 = $signed({1'h0, add_90550, array_index_90134[0]}) < $signed({1'h0, sel_90552}) ? {add_90550, array_index_90134[0]} : sel_90552;
  assign add_90656 = array_index_90335[11:1] + 11'h347;
  assign sel_90658 = $signed({1'h0, add_90554, array_index_90233[0]}) < $signed({1'h0, sel_90556}) ? {add_90554, array_index_90233[0]} : sel_90556;
  assign add_90660 = array_index_90338[11:1] + 11'h347;
  assign sel_90662 = $signed({1'h0, add_90558, array_index_90236[0]}) < $signed({1'h0, sel_90560}) ? {add_90558, array_index_90236[0]} : sel_90560;
  assign add_90664 = array_index_90437[11:3] + 9'h0bd;
  assign sel_90667 = $signed({1'h0, add_90562, array_index_90335[2:0]}) < $signed({1'h0, sel_90565}) ? {add_90562, array_index_90335[2:0]} : sel_90565;
  assign add_90669 = array_index_90440[11:3] + 9'h0bd;
  assign sel_90672 = $signed({1'h0, add_90567, array_index_90338[2:0]}) < $signed({1'h0, sel_90570}) ? {add_90567, array_index_90338[2:0]} : sel_90570;
  assign add_90674 = array_index_90539[11:1] + 11'h247;
  assign sel_90677 = $signed({1'h0, add_90572, array_index_90437[0]}) < $signed({1'h0, sel_90575}) ? {add_90572, array_index_90437[0]} : sel_90575;
  assign add_90679 = array_index_90542[11:1] + 11'h247;
  assign sel_90682 = $signed({1'h0, add_90577, array_index_90440[0]}) < $signed({1'h0, sel_90580}) ? {add_90577, array_index_90440[0]} : sel_90580;
  assign add_90707 = array_index_90641[11:0] + 12'h247;
  assign sel_90709 = $signed({1'h0, add_90605}) < $signed({1'h0, sel_90607}) ? add_90605 : sel_90607;
  assign add_90712 = array_index_90644[11:0] + 12'h247;
  assign sel_90714 = $signed({1'h0, add_90610}) < $signed({1'h0, sel_90612}) ? add_90610 : sel_90612;
  assign array_index_90743 = set1_unflattened[6'h26];
  assign array_index_90746 = set2_unflattened[6'h26];
  assign add_90750 = array_index_90335[11:1] + 11'h79d;
  assign sel_90752 = $signed({1'h0, add_90648, array_index_90233[0]}) < $signed({1'h0, sel_90650}) ? {add_90648, array_index_90233[0]} : sel_90650;
  assign add_90754 = array_index_90338[11:1] + 11'h79d;
  assign sel_90756 = $signed({1'h0, add_90652, array_index_90236[0]}) < $signed({1'h0, sel_90654}) ? {add_90652, array_index_90236[0]} : sel_90654;
  assign add_90758 = array_index_90437[11:1] + 11'h347;
  assign sel_90760 = $signed({1'h0, add_90656, array_index_90335[0]}) < $signed({1'h0, sel_90658}) ? {add_90656, array_index_90335[0]} : sel_90658;
  assign add_90762 = array_index_90440[11:1] + 11'h347;
  assign sel_90764 = $signed({1'h0, add_90660, array_index_90338[0]}) < $signed({1'h0, sel_90662}) ? {add_90660, array_index_90338[0]} : sel_90662;
  assign add_90766 = array_index_90539[11:3] + 9'h0bd;
  assign sel_90769 = $signed({1'h0, add_90664, array_index_90437[2:0]}) < $signed({1'h0, sel_90667}) ? {add_90664, array_index_90437[2:0]} : sel_90667;
  assign add_90771 = array_index_90542[11:3] + 9'h0bd;
  assign sel_90774 = $signed({1'h0, add_90669, array_index_90440[2:0]}) < $signed({1'h0, sel_90672}) ? {add_90669, array_index_90440[2:0]} : sel_90672;
  assign add_90776 = array_index_90641[11:1] + 11'h247;
  assign sel_90779 = $signed({1'h0, add_90674, array_index_90539[0]}) < $signed({1'h0, sel_90677}) ? {add_90674, array_index_90539[0]} : sel_90677;
  assign add_90781 = array_index_90644[11:1] + 11'h247;
  assign sel_90784 = $signed({1'h0, add_90679, array_index_90542[0]}) < $signed({1'h0, sel_90682}) ? {add_90679, array_index_90542[0]} : sel_90682;
  assign add_90809 = array_index_90743[11:0] + 12'h247;
  assign sel_90811 = $signed({1'h0, add_90707}) < $signed({1'h0, sel_90709}) ? add_90707 : sel_90709;
  assign add_90814 = array_index_90746[11:0] + 12'h247;
  assign sel_90816 = $signed({1'h0, add_90712}) < $signed({1'h0, sel_90714}) ? add_90712 : sel_90714;
  assign array_index_90845 = set1_unflattened[6'h27];
  assign array_index_90848 = set2_unflattened[6'h27];
  assign add_90852 = array_index_90437[11:1] + 11'h79d;
  assign sel_90854 = $signed({1'h0, add_90750, array_index_90335[0]}) < $signed({1'h0, sel_90752}) ? {add_90750, array_index_90335[0]} : sel_90752;
  assign add_90856 = array_index_90440[11:1] + 11'h79d;
  assign sel_90858 = $signed({1'h0, add_90754, array_index_90338[0]}) < $signed({1'h0, sel_90756}) ? {add_90754, array_index_90338[0]} : sel_90756;
  assign add_90860 = array_index_90539[11:1] + 11'h347;
  assign sel_90862 = $signed({1'h0, add_90758, array_index_90437[0]}) < $signed({1'h0, sel_90760}) ? {add_90758, array_index_90437[0]} : sel_90760;
  assign add_90864 = array_index_90542[11:1] + 11'h347;
  assign sel_90866 = $signed({1'h0, add_90762, array_index_90440[0]}) < $signed({1'h0, sel_90764}) ? {add_90762, array_index_90440[0]} : sel_90764;
  assign add_90868 = array_index_90641[11:3] + 9'h0bd;
  assign sel_90871 = $signed({1'h0, add_90766, array_index_90539[2:0]}) < $signed({1'h0, sel_90769}) ? {add_90766, array_index_90539[2:0]} : sel_90769;
  assign add_90873 = array_index_90644[11:3] + 9'h0bd;
  assign sel_90876 = $signed({1'h0, add_90771, array_index_90542[2:0]}) < $signed({1'h0, sel_90774}) ? {add_90771, array_index_90542[2:0]} : sel_90774;
  assign add_90878 = array_index_90743[11:1] + 11'h247;
  assign sel_90881 = $signed({1'h0, add_90776, array_index_90641[0]}) < $signed({1'h0, sel_90779}) ? {add_90776, array_index_90641[0]} : sel_90779;
  assign add_90883 = array_index_90746[11:1] + 11'h247;
  assign sel_90886 = $signed({1'h0, add_90781, array_index_90644[0]}) < $signed({1'h0, sel_90784}) ? {add_90781, array_index_90644[0]} : sel_90784;
  assign add_90911 = array_index_90845[11:0] + 12'h247;
  assign sel_90913 = $signed({1'h0, add_90809}) < $signed({1'h0, sel_90811}) ? add_90809 : sel_90811;
  assign add_90916 = array_index_90848[11:0] + 12'h247;
  assign sel_90918 = $signed({1'h0, add_90814}) < $signed({1'h0, sel_90816}) ? add_90814 : sel_90816;
  assign array_index_90947 = set1_unflattened[6'h28];
  assign array_index_90950 = set2_unflattened[6'h28];
  assign add_90954 = array_index_90539[11:1] + 11'h79d;
  assign sel_90956 = $signed({1'h0, add_90852, array_index_90437[0]}) < $signed({1'h0, sel_90854}) ? {add_90852, array_index_90437[0]} : sel_90854;
  assign add_90958 = array_index_90542[11:1] + 11'h79d;
  assign sel_90960 = $signed({1'h0, add_90856, array_index_90440[0]}) < $signed({1'h0, sel_90858}) ? {add_90856, array_index_90440[0]} : sel_90858;
  assign add_90962 = array_index_90641[11:1] + 11'h347;
  assign sel_90964 = $signed({1'h0, add_90860, array_index_90539[0]}) < $signed({1'h0, sel_90862}) ? {add_90860, array_index_90539[0]} : sel_90862;
  assign add_90966 = array_index_90644[11:1] + 11'h347;
  assign sel_90968 = $signed({1'h0, add_90864, array_index_90542[0]}) < $signed({1'h0, sel_90866}) ? {add_90864, array_index_90542[0]} : sel_90866;
  assign add_90970 = array_index_90743[11:3] + 9'h0bd;
  assign sel_90973 = $signed({1'h0, add_90868, array_index_90641[2:0]}) < $signed({1'h0, sel_90871}) ? {add_90868, array_index_90641[2:0]} : sel_90871;
  assign add_90975 = array_index_90746[11:3] + 9'h0bd;
  assign sel_90978 = $signed({1'h0, add_90873, array_index_90644[2:0]}) < $signed({1'h0, sel_90876}) ? {add_90873, array_index_90644[2:0]} : sel_90876;
  assign add_90980 = array_index_90845[11:1] + 11'h247;
  assign sel_90983 = $signed({1'h0, add_90878, array_index_90743[0]}) < $signed({1'h0, sel_90881}) ? {add_90878, array_index_90743[0]} : sel_90881;
  assign add_90985 = array_index_90848[11:1] + 11'h247;
  assign sel_90988 = $signed({1'h0, add_90883, array_index_90746[0]}) < $signed({1'h0, sel_90886}) ? {add_90883, array_index_90746[0]} : sel_90886;
  assign add_91013 = array_index_90947[11:0] + 12'h247;
  assign sel_91015 = $signed({1'h0, add_90911}) < $signed({1'h0, sel_90913}) ? add_90911 : sel_90913;
  assign add_91018 = array_index_90950[11:0] + 12'h247;
  assign sel_91020 = $signed({1'h0, add_90916}) < $signed({1'h0, sel_90918}) ? add_90916 : sel_90918;
  assign array_index_91049 = set1_unflattened[6'h29];
  assign array_index_91052 = set2_unflattened[6'h29];
  assign add_91056 = array_index_90641[11:1] + 11'h79d;
  assign sel_91058 = $signed({1'h0, add_90954, array_index_90539[0]}) < $signed({1'h0, sel_90956}) ? {add_90954, array_index_90539[0]} : sel_90956;
  assign add_91060 = array_index_90644[11:1] + 11'h79d;
  assign sel_91062 = $signed({1'h0, add_90958, array_index_90542[0]}) < $signed({1'h0, sel_90960}) ? {add_90958, array_index_90542[0]} : sel_90960;
  assign add_91064 = array_index_90743[11:1] + 11'h347;
  assign sel_91066 = $signed({1'h0, add_90962, array_index_90641[0]}) < $signed({1'h0, sel_90964}) ? {add_90962, array_index_90641[0]} : sel_90964;
  assign add_91068 = array_index_90746[11:1] + 11'h347;
  assign sel_91070 = $signed({1'h0, add_90966, array_index_90644[0]}) < $signed({1'h0, sel_90968}) ? {add_90966, array_index_90644[0]} : sel_90968;
  assign add_91072 = array_index_90845[11:3] + 9'h0bd;
  assign sel_91075 = $signed({1'h0, add_90970, array_index_90743[2:0]}) < $signed({1'h0, sel_90973}) ? {add_90970, array_index_90743[2:0]} : sel_90973;
  assign add_91077 = array_index_90848[11:3] + 9'h0bd;
  assign sel_91080 = $signed({1'h0, add_90975, array_index_90746[2:0]}) < $signed({1'h0, sel_90978}) ? {add_90975, array_index_90746[2:0]} : sel_90978;
  assign add_91082 = array_index_90947[11:1] + 11'h247;
  assign sel_91085 = $signed({1'h0, add_90980, array_index_90845[0]}) < $signed({1'h0, sel_90983}) ? {add_90980, array_index_90845[0]} : sel_90983;
  assign add_91087 = array_index_90950[11:1] + 11'h247;
  assign sel_91090 = $signed({1'h0, add_90985, array_index_90848[0]}) < $signed({1'h0, sel_90988}) ? {add_90985, array_index_90848[0]} : sel_90988;
  assign add_91115 = array_index_91049[11:0] + 12'h247;
  assign sel_91117 = $signed({1'h0, add_91013}) < $signed({1'h0, sel_91015}) ? add_91013 : sel_91015;
  assign add_91120 = array_index_91052[11:0] + 12'h247;
  assign sel_91122 = $signed({1'h0, add_91018}) < $signed({1'h0, sel_91020}) ? add_91018 : sel_91020;
  assign array_index_91151 = set1_unflattened[6'h2a];
  assign array_index_91154 = set2_unflattened[6'h2a];
  assign add_91158 = array_index_90743[11:1] + 11'h79d;
  assign sel_91160 = $signed({1'h0, add_91056, array_index_90641[0]}) < $signed({1'h0, sel_91058}) ? {add_91056, array_index_90641[0]} : sel_91058;
  assign add_91162 = array_index_90746[11:1] + 11'h79d;
  assign sel_91164 = $signed({1'h0, add_91060, array_index_90644[0]}) < $signed({1'h0, sel_91062}) ? {add_91060, array_index_90644[0]} : sel_91062;
  assign add_91166 = array_index_90845[11:1] + 11'h347;
  assign sel_91168 = $signed({1'h0, add_91064, array_index_90743[0]}) < $signed({1'h0, sel_91066}) ? {add_91064, array_index_90743[0]} : sel_91066;
  assign add_91170 = array_index_90848[11:1] + 11'h347;
  assign sel_91172 = $signed({1'h0, add_91068, array_index_90746[0]}) < $signed({1'h0, sel_91070}) ? {add_91068, array_index_90746[0]} : sel_91070;
  assign add_91174 = array_index_90947[11:3] + 9'h0bd;
  assign sel_91177 = $signed({1'h0, add_91072, array_index_90845[2:0]}) < $signed({1'h0, sel_91075}) ? {add_91072, array_index_90845[2:0]} : sel_91075;
  assign add_91179 = array_index_90950[11:3] + 9'h0bd;
  assign sel_91182 = $signed({1'h0, add_91077, array_index_90848[2:0]}) < $signed({1'h0, sel_91080}) ? {add_91077, array_index_90848[2:0]} : sel_91080;
  assign add_91184 = array_index_91049[11:1] + 11'h247;
  assign sel_91187 = $signed({1'h0, add_91082, array_index_90947[0]}) < $signed({1'h0, sel_91085}) ? {add_91082, array_index_90947[0]} : sel_91085;
  assign add_91189 = array_index_91052[11:1] + 11'h247;
  assign sel_91192 = $signed({1'h0, add_91087, array_index_90950[0]}) < $signed({1'h0, sel_91090}) ? {add_91087, array_index_90950[0]} : sel_91090;
  assign add_91217 = array_index_91151[11:0] + 12'h247;
  assign sel_91219 = $signed({1'h0, add_91115}) < $signed({1'h0, sel_91117}) ? add_91115 : sel_91117;
  assign add_91222 = array_index_91154[11:0] + 12'h247;
  assign sel_91224 = $signed({1'h0, add_91120}) < $signed({1'h0, sel_91122}) ? add_91120 : sel_91122;
  assign array_index_91253 = set1_unflattened[6'h2b];
  assign array_index_91256 = set2_unflattened[6'h2b];
  assign add_91260 = array_index_90845[11:1] + 11'h79d;
  assign sel_91262 = $signed({1'h0, add_91158, array_index_90743[0]}) < $signed({1'h0, sel_91160}) ? {add_91158, array_index_90743[0]} : sel_91160;
  assign add_91264 = array_index_90848[11:1] + 11'h79d;
  assign sel_91266 = $signed({1'h0, add_91162, array_index_90746[0]}) < $signed({1'h0, sel_91164}) ? {add_91162, array_index_90746[0]} : sel_91164;
  assign add_91268 = array_index_90947[11:1] + 11'h347;
  assign sel_91270 = $signed({1'h0, add_91166, array_index_90845[0]}) < $signed({1'h0, sel_91168}) ? {add_91166, array_index_90845[0]} : sel_91168;
  assign add_91272 = array_index_90950[11:1] + 11'h347;
  assign sel_91274 = $signed({1'h0, add_91170, array_index_90848[0]}) < $signed({1'h0, sel_91172}) ? {add_91170, array_index_90848[0]} : sel_91172;
  assign add_91276 = array_index_91049[11:3] + 9'h0bd;
  assign sel_91279 = $signed({1'h0, add_91174, array_index_90947[2:0]}) < $signed({1'h0, sel_91177}) ? {add_91174, array_index_90947[2:0]} : sel_91177;
  assign add_91281 = array_index_91052[11:3] + 9'h0bd;
  assign sel_91284 = $signed({1'h0, add_91179, array_index_90950[2:0]}) < $signed({1'h0, sel_91182}) ? {add_91179, array_index_90950[2:0]} : sel_91182;
  assign add_91286 = array_index_91151[11:1] + 11'h247;
  assign sel_91289 = $signed({1'h0, add_91184, array_index_91049[0]}) < $signed({1'h0, sel_91187}) ? {add_91184, array_index_91049[0]} : sel_91187;
  assign add_91291 = array_index_91154[11:1] + 11'h247;
  assign sel_91294 = $signed({1'h0, add_91189, array_index_91052[0]}) < $signed({1'h0, sel_91192}) ? {add_91189, array_index_91052[0]} : sel_91192;
  assign add_91319 = array_index_91253[11:0] + 12'h247;
  assign sel_91321 = $signed({1'h0, add_91217}) < $signed({1'h0, sel_91219}) ? add_91217 : sel_91219;
  assign add_91324 = array_index_91256[11:0] + 12'h247;
  assign sel_91326 = $signed({1'h0, add_91222}) < $signed({1'h0, sel_91224}) ? add_91222 : sel_91224;
  assign array_index_91355 = set1_unflattened[6'h2c];
  assign array_index_91358 = set2_unflattened[6'h2c];
  assign add_91362 = array_index_90947[11:1] + 11'h79d;
  assign sel_91364 = $signed({1'h0, add_91260, array_index_90845[0]}) < $signed({1'h0, sel_91262}) ? {add_91260, array_index_90845[0]} : sel_91262;
  assign add_91366 = array_index_90950[11:1] + 11'h79d;
  assign sel_91368 = $signed({1'h0, add_91264, array_index_90848[0]}) < $signed({1'h0, sel_91266}) ? {add_91264, array_index_90848[0]} : sel_91266;
  assign add_91370 = array_index_91049[11:1] + 11'h347;
  assign sel_91372 = $signed({1'h0, add_91268, array_index_90947[0]}) < $signed({1'h0, sel_91270}) ? {add_91268, array_index_90947[0]} : sel_91270;
  assign add_91374 = array_index_91052[11:1] + 11'h347;
  assign sel_91376 = $signed({1'h0, add_91272, array_index_90950[0]}) < $signed({1'h0, sel_91274}) ? {add_91272, array_index_90950[0]} : sel_91274;
  assign add_91378 = array_index_91151[11:3] + 9'h0bd;
  assign sel_91381 = $signed({1'h0, add_91276, array_index_91049[2:0]}) < $signed({1'h0, sel_91279}) ? {add_91276, array_index_91049[2:0]} : sel_91279;
  assign add_91383 = array_index_91154[11:3] + 9'h0bd;
  assign sel_91386 = $signed({1'h0, add_91281, array_index_91052[2:0]}) < $signed({1'h0, sel_91284}) ? {add_91281, array_index_91052[2:0]} : sel_91284;
  assign add_91388 = array_index_91253[11:1] + 11'h247;
  assign sel_91391 = $signed({1'h0, add_91286, array_index_91151[0]}) < $signed({1'h0, sel_91289}) ? {add_91286, array_index_91151[0]} : sel_91289;
  assign add_91393 = array_index_91256[11:1] + 11'h247;
  assign sel_91396 = $signed({1'h0, add_91291, array_index_91154[0]}) < $signed({1'h0, sel_91294}) ? {add_91291, array_index_91154[0]} : sel_91294;
  assign add_91421 = array_index_91355[11:0] + 12'h247;
  assign sel_91423 = $signed({1'h0, add_91319}) < $signed({1'h0, sel_91321}) ? add_91319 : sel_91321;
  assign add_91426 = array_index_91358[11:0] + 12'h247;
  assign sel_91428 = $signed({1'h0, add_91324}) < $signed({1'h0, sel_91326}) ? add_91324 : sel_91326;
  assign array_index_91457 = set1_unflattened[6'h2d];
  assign array_index_91460 = set2_unflattened[6'h2d];
  assign add_91464 = array_index_91049[11:1] + 11'h79d;
  assign sel_91466 = $signed({1'h0, add_91362, array_index_90947[0]}) < $signed({1'h0, sel_91364}) ? {add_91362, array_index_90947[0]} : sel_91364;
  assign add_91468 = array_index_91052[11:1] + 11'h79d;
  assign sel_91470 = $signed({1'h0, add_91366, array_index_90950[0]}) < $signed({1'h0, sel_91368}) ? {add_91366, array_index_90950[0]} : sel_91368;
  assign add_91472 = array_index_91151[11:1] + 11'h347;
  assign sel_91474 = $signed({1'h0, add_91370, array_index_91049[0]}) < $signed({1'h0, sel_91372}) ? {add_91370, array_index_91049[0]} : sel_91372;
  assign add_91476 = array_index_91154[11:1] + 11'h347;
  assign sel_91478 = $signed({1'h0, add_91374, array_index_91052[0]}) < $signed({1'h0, sel_91376}) ? {add_91374, array_index_91052[0]} : sel_91376;
  assign add_91480 = array_index_91253[11:3] + 9'h0bd;
  assign sel_91483 = $signed({1'h0, add_91378, array_index_91151[2:0]}) < $signed({1'h0, sel_91381}) ? {add_91378, array_index_91151[2:0]} : sel_91381;
  assign add_91485 = array_index_91256[11:3] + 9'h0bd;
  assign sel_91488 = $signed({1'h0, add_91383, array_index_91154[2:0]}) < $signed({1'h0, sel_91386}) ? {add_91383, array_index_91154[2:0]} : sel_91386;
  assign add_91490 = array_index_91355[11:1] + 11'h247;
  assign sel_91493 = $signed({1'h0, add_91388, array_index_91253[0]}) < $signed({1'h0, sel_91391}) ? {add_91388, array_index_91253[0]} : sel_91391;
  assign add_91495 = array_index_91358[11:1] + 11'h247;
  assign sel_91498 = $signed({1'h0, add_91393, array_index_91256[0]}) < $signed({1'h0, sel_91396}) ? {add_91393, array_index_91256[0]} : sel_91396;
  assign add_91523 = array_index_91457[11:0] + 12'h247;
  assign sel_91525 = $signed({1'h0, add_91421}) < $signed({1'h0, sel_91423}) ? add_91421 : sel_91423;
  assign add_91528 = array_index_91460[11:0] + 12'h247;
  assign sel_91530 = $signed({1'h0, add_91426}) < $signed({1'h0, sel_91428}) ? add_91426 : sel_91428;
  assign array_index_91559 = set1_unflattened[6'h2e];
  assign array_index_91562 = set2_unflattened[6'h2e];
  assign add_91566 = array_index_91151[11:1] + 11'h79d;
  assign sel_91568 = $signed({1'h0, add_91464, array_index_91049[0]}) < $signed({1'h0, sel_91466}) ? {add_91464, array_index_91049[0]} : sel_91466;
  assign add_91570 = array_index_91154[11:1] + 11'h79d;
  assign sel_91572 = $signed({1'h0, add_91468, array_index_91052[0]}) < $signed({1'h0, sel_91470}) ? {add_91468, array_index_91052[0]} : sel_91470;
  assign add_91574 = array_index_91253[11:1] + 11'h347;
  assign sel_91576 = $signed({1'h0, add_91472, array_index_91151[0]}) < $signed({1'h0, sel_91474}) ? {add_91472, array_index_91151[0]} : sel_91474;
  assign add_91578 = array_index_91256[11:1] + 11'h347;
  assign sel_91580 = $signed({1'h0, add_91476, array_index_91154[0]}) < $signed({1'h0, sel_91478}) ? {add_91476, array_index_91154[0]} : sel_91478;
  assign add_91582 = array_index_91355[11:3] + 9'h0bd;
  assign sel_91585 = $signed({1'h0, add_91480, array_index_91253[2:0]}) < $signed({1'h0, sel_91483}) ? {add_91480, array_index_91253[2:0]} : sel_91483;
  assign add_91587 = array_index_91358[11:3] + 9'h0bd;
  assign sel_91590 = $signed({1'h0, add_91485, array_index_91256[2:0]}) < $signed({1'h0, sel_91488}) ? {add_91485, array_index_91256[2:0]} : sel_91488;
  assign add_91592 = array_index_91457[11:1] + 11'h247;
  assign sel_91595 = $signed({1'h0, add_91490, array_index_91355[0]}) < $signed({1'h0, sel_91493}) ? {add_91490, array_index_91355[0]} : sel_91493;
  assign add_91597 = array_index_91460[11:1] + 11'h247;
  assign sel_91600 = $signed({1'h0, add_91495, array_index_91358[0]}) < $signed({1'h0, sel_91498}) ? {add_91495, array_index_91358[0]} : sel_91498;
  assign add_91625 = array_index_91559[11:0] + 12'h247;
  assign sel_91627 = $signed({1'h0, add_91523}) < $signed({1'h0, sel_91525}) ? add_91523 : sel_91525;
  assign add_91630 = array_index_91562[11:0] + 12'h247;
  assign sel_91632 = $signed({1'h0, add_91528}) < $signed({1'h0, sel_91530}) ? add_91528 : sel_91530;
  assign array_index_91661 = set1_unflattened[6'h2f];
  assign array_index_91664 = set2_unflattened[6'h2f];
  assign add_91668 = array_index_91253[11:1] + 11'h79d;
  assign sel_91670 = $signed({1'h0, add_91566, array_index_91151[0]}) < $signed({1'h0, sel_91568}) ? {add_91566, array_index_91151[0]} : sel_91568;
  assign add_91672 = array_index_91256[11:1] + 11'h79d;
  assign sel_91674 = $signed({1'h0, add_91570, array_index_91154[0]}) < $signed({1'h0, sel_91572}) ? {add_91570, array_index_91154[0]} : sel_91572;
  assign add_91676 = array_index_91355[11:1] + 11'h347;
  assign sel_91678 = $signed({1'h0, add_91574, array_index_91253[0]}) < $signed({1'h0, sel_91576}) ? {add_91574, array_index_91253[0]} : sel_91576;
  assign add_91680 = array_index_91358[11:1] + 11'h347;
  assign sel_91682 = $signed({1'h0, add_91578, array_index_91256[0]}) < $signed({1'h0, sel_91580}) ? {add_91578, array_index_91256[0]} : sel_91580;
  assign add_91684 = array_index_91457[11:3] + 9'h0bd;
  assign sel_91687 = $signed({1'h0, add_91582, array_index_91355[2:0]}) < $signed({1'h0, sel_91585}) ? {add_91582, array_index_91355[2:0]} : sel_91585;
  assign add_91689 = array_index_91460[11:3] + 9'h0bd;
  assign sel_91692 = $signed({1'h0, add_91587, array_index_91358[2:0]}) < $signed({1'h0, sel_91590}) ? {add_91587, array_index_91358[2:0]} : sel_91590;
  assign add_91694 = array_index_91559[11:1] + 11'h247;
  assign sel_91697 = $signed({1'h0, add_91592, array_index_91457[0]}) < $signed({1'h0, sel_91595}) ? {add_91592, array_index_91457[0]} : sel_91595;
  assign add_91699 = array_index_91562[11:1] + 11'h247;
  assign sel_91702 = $signed({1'h0, add_91597, array_index_91460[0]}) < $signed({1'h0, sel_91600}) ? {add_91597, array_index_91460[0]} : sel_91600;
  assign add_91727 = array_index_91661[11:0] + 12'h247;
  assign sel_91729 = $signed({1'h0, add_91625}) < $signed({1'h0, sel_91627}) ? add_91625 : sel_91627;
  assign add_91732 = array_index_91664[11:0] + 12'h247;
  assign sel_91734 = $signed({1'h0, add_91630}) < $signed({1'h0, sel_91632}) ? add_91630 : sel_91632;
  assign array_index_91763 = set1_unflattened[6'h30];
  assign array_index_91766 = set2_unflattened[6'h30];
  assign add_91770 = array_index_91355[11:1] + 11'h79d;
  assign sel_91772 = $signed({1'h0, add_91668, array_index_91253[0]}) < $signed({1'h0, sel_91670}) ? {add_91668, array_index_91253[0]} : sel_91670;
  assign add_91774 = array_index_91358[11:1] + 11'h79d;
  assign sel_91776 = $signed({1'h0, add_91672, array_index_91256[0]}) < $signed({1'h0, sel_91674}) ? {add_91672, array_index_91256[0]} : sel_91674;
  assign add_91778 = array_index_91457[11:1] + 11'h347;
  assign sel_91780 = $signed({1'h0, add_91676, array_index_91355[0]}) < $signed({1'h0, sel_91678}) ? {add_91676, array_index_91355[0]} : sel_91678;
  assign add_91782 = array_index_91460[11:1] + 11'h347;
  assign sel_91784 = $signed({1'h0, add_91680, array_index_91358[0]}) < $signed({1'h0, sel_91682}) ? {add_91680, array_index_91358[0]} : sel_91682;
  assign add_91786 = array_index_91559[11:3] + 9'h0bd;
  assign sel_91789 = $signed({1'h0, add_91684, array_index_91457[2:0]}) < $signed({1'h0, sel_91687}) ? {add_91684, array_index_91457[2:0]} : sel_91687;
  assign add_91791 = array_index_91562[11:3] + 9'h0bd;
  assign sel_91794 = $signed({1'h0, add_91689, array_index_91460[2:0]}) < $signed({1'h0, sel_91692}) ? {add_91689, array_index_91460[2:0]} : sel_91692;
  assign add_91796 = array_index_91661[11:1] + 11'h247;
  assign sel_91799 = $signed({1'h0, add_91694, array_index_91559[0]}) < $signed({1'h0, sel_91697}) ? {add_91694, array_index_91559[0]} : sel_91697;
  assign add_91801 = array_index_91664[11:1] + 11'h247;
  assign sel_91804 = $signed({1'h0, add_91699, array_index_91562[0]}) < $signed({1'h0, sel_91702}) ? {add_91699, array_index_91562[0]} : sel_91702;
  assign add_91829 = array_index_91763[11:0] + 12'h247;
  assign sel_91831 = $signed({1'h0, add_91727}) < $signed({1'h0, sel_91729}) ? add_91727 : sel_91729;
  assign add_91834 = array_index_91766[11:0] + 12'h247;
  assign sel_91836 = $signed({1'h0, add_91732}) < $signed({1'h0, sel_91734}) ? add_91732 : sel_91734;
  assign array_index_91865 = set1_unflattened[6'h31];
  assign array_index_91868 = set2_unflattened[6'h31];
  assign add_91872 = array_index_91457[11:1] + 11'h79d;
  assign sel_91874 = $signed({1'h0, add_91770, array_index_91355[0]}) < $signed({1'h0, sel_91772}) ? {add_91770, array_index_91355[0]} : sel_91772;
  assign add_91876 = array_index_91460[11:1] + 11'h79d;
  assign sel_91878 = $signed({1'h0, add_91774, array_index_91358[0]}) < $signed({1'h0, sel_91776}) ? {add_91774, array_index_91358[0]} : sel_91776;
  assign add_91880 = array_index_91559[11:1] + 11'h347;
  assign sel_91882 = $signed({1'h0, add_91778, array_index_91457[0]}) < $signed({1'h0, sel_91780}) ? {add_91778, array_index_91457[0]} : sel_91780;
  assign add_91884 = array_index_91562[11:1] + 11'h347;
  assign sel_91886 = $signed({1'h0, add_91782, array_index_91460[0]}) < $signed({1'h0, sel_91784}) ? {add_91782, array_index_91460[0]} : sel_91784;
  assign add_91888 = array_index_91661[11:3] + 9'h0bd;
  assign sel_91891 = $signed({1'h0, add_91786, array_index_91559[2:0]}) < $signed({1'h0, sel_91789}) ? {add_91786, array_index_91559[2:0]} : sel_91789;
  assign add_91893 = array_index_91664[11:3] + 9'h0bd;
  assign sel_91896 = $signed({1'h0, add_91791, array_index_91562[2:0]}) < $signed({1'h0, sel_91794}) ? {add_91791, array_index_91562[2:0]} : sel_91794;
  assign add_91898 = array_index_91763[11:1] + 11'h247;
  assign sel_91901 = $signed({1'h0, add_91796, array_index_91661[0]}) < $signed({1'h0, sel_91799}) ? {add_91796, array_index_91661[0]} : sel_91799;
  assign add_91903 = array_index_91766[11:1] + 11'h247;
  assign sel_91906 = $signed({1'h0, add_91801, array_index_91664[0]}) < $signed({1'h0, sel_91804}) ? {add_91801, array_index_91664[0]} : sel_91804;
  assign add_91930 = array_index_91865[11:0] + 12'h247;
  assign sel_91932 = $signed({1'h0, add_91829}) < $signed({1'h0, sel_91831}) ? add_91829 : sel_91831;
  assign add_91934 = array_index_91868[11:0] + 12'h247;
  assign sel_91936 = $signed({1'h0, add_91834}) < $signed({1'h0, sel_91836}) ? add_91834 : sel_91836;
  assign add_91970 = array_index_91559[11:1] + 11'h79d;
  assign sel_91972 = $signed({1'h0, add_91872, array_index_91457[0]}) < $signed({1'h0, sel_91874}) ? {add_91872, array_index_91457[0]} : sel_91874;
  assign add_91974 = array_index_91562[11:1] + 11'h79d;
  assign sel_91976 = $signed({1'h0, add_91876, array_index_91460[0]}) < $signed({1'h0, sel_91878}) ? {add_91876, array_index_91460[0]} : sel_91878;
  assign add_91978 = array_index_91661[11:1] + 11'h347;
  assign sel_91980 = $signed({1'h0, add_91880, array_index_91559[0]}) < $signed({1'h0, sel_91882}) ? {add_91880, array_index_91559[0]} : sel_91882;
  assign add_91982 = array_index_91664[11:1] + 11'h347;
  assign sel_91984 = $signed({1'h0, add_91884, array_index_91562[0]}) < $signed({1'h0, sel_91886}) ? {add_91884, array_index_91562[0]} : sel_91886;
  assign add_91986 = array_index_91763[11:3] + 9'h0bd;
  assign sel_91989 = $signed({1'h0, add_91888, array_index_91661[2:0]}) < $signed({1'h0, sel_91891}) ? {add_91888, array_index_91661[2:0]} : sel_91891;
  assign add_91991 = array_index_91766[11:3] + 9'h0bd;
  assign sel_91994 = $signed({1'h0, add_91893, array_index_91664[2:0]}) < $signed({1'h0, sel_91896}) ? {add_91893, array_index_91664[2:0]} : sel_91896;
  assign add_91996 = array_index_91865[11:1] + 11'h247;
  assign sel_91999 = $signed({1'h0, add_91898, array_index_91763[0]}) < $signed({1'h0, sel_91901}) ? {add_91898, array_index_91763[0]} : sel_91901;
  assign add_92001 = array_index_91868[11:1] + 11'h247;
  assign sel_92004 = $signed({1'h0, add_91903, array_index_91766[0]}) < $signed({1'h0, sel_91906}) ? {add_91903, array_index_91766[0]} : sel_91906;
  assign add_92052 = array_index_91661[11:1] + 11'h79d;
  assign sel_92054 = $signed({1'h0, add_91970, array_index_91559[0]}) < $signed({1'h0, sel_91972}) ? {add_91970, array_index_91559[0]} : sel_91972;
  assign add_92056 = array_index_91664[11:1] + 11'h79d;
  assign sel_92058 = $signed({1'h0, add_91974, array_index_91562[0]}) < $signed({1'h0, sel_91976}) ? {add_91974, array_index_91562[0]} : sel_91976;
  assign add_92060 = array_index_91763[11:1] + 11'h347;
  assign sel_92062 = $signed({1'h0, add_91978, array_index_91661[0]}) < $signed({1'h0, sel_91980}) ? {add_91978, array_index_91661[0]} : sel_91980;
  assign add_92064 = array_index_91766[11:1] + 11'h347;
  assign sel_92066 = $signed({1'h0, add_91982, array_index_91664[0]}) < $signed({1'h0, sel_91984}) ? {add_91982, array_index_91664[0]} : sel_91984;
  assign add_92068 = array_index_91865[11:3] + 9'h0bd;
  assign sel_92071 = $signed({1'h0, add_91986, array_index_91763[2:0]}) < $signed({1'h0, sel_91989}) ? {add_91986, array_index_91763[2:0]} : sel_91989;
  assign add_92073 = array_index_91868[11:3] + 9'h0bd;
  assign sel_92076 = $signed({1'h0, add_91991, array_index_91766[2:0]}) < $signed({1'h0, sel_91994}) ? {add_91991, array_index_91766[2:0]} : sel_91994;
  assign concat_92079 = {1'h0, ($signed({1'h0, add_91930}) < $signed({1'h0, sel_91932}) ? add_91930 : sel_91932) == ($signed({1'h0, add_91934}) < $signed({1'h0, sel_91936}) ? add_91934 : sel_91936)};
  assign add_92094 = concat_92079 + 2'h1;
  assign add_92114 = array_index_91763[11:1] + 11'h79d;
  assign sel_92116 = $signed({1'h0, add_92052, array_index_91661[0]}) < $signed({1'h0, sel_92054}) ? {add_92052, array_index_91661[0]} : sel_92054;
  assign add_92118 = array_index_91766[11:1] + 11'h79d;
  assign sel_92120 = $signed({1'h0, add_92056, array_index_91664[0]}) < $signed({1'h0, sel_92058}) ? {add_92056, array_index_91664[0]} : sel_92058;
  assign add_92122 = array_index_91865[11:1] + 11'h347;
  assign sel_92124 = $signed({1'h0, add_92060, array_index_91763[0]}) < $signed({1'h0, sel_92062}) ? {add_92060, array_index_91763[0]} : sel_92062;
  assign add_92126 = array_index_91868[11:1] + 11'h347;
  assign sel_92128 = $signed({1'h0, add_92064, array_index_91766[0]}) < $signed({1'h0, sel_92066}) ? {add_92064, array_index_91766[0]} : sel_92066;
  assign concat_92131 = {1'h0, ($signed({1'h0, add_91996, array_index_91865[0]}) < $signed({1'h0, sel_91999}) ? {add_91996, array_index_91865[0]} : sel_91999) == ($signed({1'h0, add_92001, array_index_91868[0]}) < $signed({1'h0, sel_92004}) ? {add_92001, array_index_91868[0]} : sel_92004) ? add_92094 : concat_92079};
  assign add_92142 = concat_92131 + 3'h1;
  assign add_92156 = array_index_91865[11:1] + 11'h79d;
  assign sel_92158 = $signed({1'h0, add_92114, array_index_91763[0]}) < $signed({1'h0, sel_92116}) ? {add_92114, array_index_91763[0]} : sel_92116;
  assign add_92160 = array_index_91868[11:1] + 11'h79d;
  assign sel_92162 = $signed({1'h0, add_92118, array_index_91766[0]}) < $signed({1'h0, sel_92120}) ? {add_92118, array_index_91766[0]} : sel_92120;
  assign concat_92165 = {1'h0, ($signed({1'h0, add_92068, array_index_91865[2:0]}) < $signed({1'h0, sel_92071}) ? {add_92068, array_index_91865[2:0]} : sel_92071) == ($signed({1'h0, add_92073, array_index_91868[2:0]}) < $signed({1'h0, sel_92076}) ? {add_92073, array_index_91868[2:0]} : sel_92076) ? add_92142 : concat_92131};
  assign add_92172 = concat_92165 + 4'h1;
  assign concat_92181 = {1'h0, ($signed({1'h0, add_92122, array_index_91865[0]}) < $signed({1'h0, sel_92124}) ? {add_92122, array_index_91865[0]} : sel_92124) == ($signed({1'h0, add_92126, array_index_91868[0]}) < $signed({1'h0, sel_92128}) ? {add_92126, array_index_91868[0]} : sel_92128) ? add_92172 : concat_92165};
  assign add_92184 = concat_92181 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_92156, array_index_91865[0]}) < $signed({1'h0, sel_92158}) ? {add_92156, array_index_91865[0]} : sel_92158) == ($signed({1'h0, add_92160, array_index_91868[0]}) < $signed({1'h0, sel_92162}) ? {add_92160, array_index_91868[0]} : sel_92162) ? add_92184 : concat_92181}, {set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
