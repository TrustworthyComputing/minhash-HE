module min_hash(set1, set2, out);
  wire _000000_, _000001_, _000002_, _000003_, _000004_, _000005_, _000006_, _000007_, _000008_, _000009_, _000010_, _000011_, _000012_, _000013_, _000014_, _000015_, _000016_, _000017_, _000018_, _000019_, _000020_, _000021_, _000022_, _000023_, _000024_, _000025_, _000026_, _000027_, _000028_, _000029_, _000030_, _000031_, _000032_, _000033_, _000034_, _000035_, _000036_, _000037_, _000038_, _000039_, _000040_, _000041_, _000042_, _000043_, _000044_, _000045_, _000046_, _000047_, _000048_, _000049_, _000050_, _000051_, _000052_, _000053_, _000054_, _000055_, _000056_, _000057_, _000058_, _000059_, _000060_, _000061_, _000062_, _000063_, _000064_, _000065_, _000066_, _000067_, _000068_, _000069_, _000070_, _000071_, _000072_, _000073_, _000074_, _000075_, _000076_, _000077_, _000078_, _000079_, _000080_, _000081_, _000082_, _000083_, _000084_, _000085_, _000086_, _000087_, _000088_, _000089_, _000090_, _000091_, _000092_, _000093_, _000094_, _000095_, _000096_, _000097_, _000098_, _000099_, _000100_, _000101_, _000102_, _000103_, _000104_, _000105_, _000106_, _000107_, _000108_, _000109_, _000110_, _000111_, _000112_, _000113_, _000114_, _000115_, _000116_, _000117_, _000118_, _000119_, _000120_, _000121_, _000122_, _000123_, _000124_, _000125_, _000126_, _000127_, _000128_, _000129_, _000130_, _000131_, _000132_, _000133_, _000134_, _000135_, _000136_, _000137_, _000138_, _000139_, _000140_, _000141_, _000142_, _000143_, _000144_, _000145_, _000146_, _000147_, _000148_, _000149_, _000150_, _000151_, _000152_, _000153_, _000154_, _000155_, _000156_, _000157_, _000158_, _000159_, _000160_, _000161_, _000162_, _000163_, _000164_, _000165_, _000166_, _000167_, _000168_, _000169_, _000170_, _000171_, _000172_, _000173_, _000174_, _000175_, _000176_, _000177_, _000178_, _000179_, _000180_, _000181_, _000182_, _000183_, _000184_, _000185_, _000186_, _000187_, _000188_, _000189_, _000190_, _000191_, _000192_, _000193_, _000194_, _000195_, _000196_, _000197_, _000198_, _000199_, _000200_, _000201_, _000202_, _000203_, _000204_, _000205_, _000206_, _000207_, _000208_, _000209_, _000210_, _000211_, _000212_, _000213_, _000214_, _000215_, _000216_, _000217_, _000218_, _000219_, _000220_, _000221_, _000222_, _000223_, _000224_, _000225_, _000226_, _000227_, _000228_, _000229_, _000230_, _000231_, _000232_, _000233_, _000234_, _000235_, _000236_, _000237_, _000238_, _000239_, _000240_, _000241_, _000242_, _000243_, _000244_, _000245_, _000246_, _000247_, _000248_, _000249_, _000250_, _000251_, _000252_, _000253_, _000254_, _000255_, _000256_, _000257_, _000258_, _000259_, _000260_, _000261_, _000262_, _000263_, _000264_, _000265_, _000266_, _000267_, _000268_, _000269_, _000270_, _000271_, _000272_, _000273_, _000274_, _000275_, _000276_, _000277_, _000278_, _000279_, _000280_, _000281_, _000282_, _000283_, _000284_, _000285_, _000286_, _000287_, _000288_, _000289_, _000290_, _000291_, _000292_, _000293_, _000294_, _000295_, _000296_, _000297_, _000298_, _000299_, _000300_, _000301_, _000302_, _000303_, _000304_, _000305_, _000306_, _000307_, _000308_, _000309_, _000310_, _000311_, _000312_, _000313_, _000314_, _000315_, _000316_, _000317_, _000318_, _000319_, _000320_, _000321_, _000322_, _000323_, _000324_, _000325_, _000326_, _000327_, _000328_, _000329_, _000330_, _000331_, _000332_, _000333_, _000334_, _000335_, _000336_, _000337_, _000338_, _000339_, _000340_, _000341_, _000342_, _000343_, _000344_, _000345_, _000346_, _000347_, _000348_, _000349_, _000350_, _000351_, _000352_, _000353_, _000354_, _000355_, _000356_, _000357_, _000358_, _000359_, _000360_, _000361_, _000362_, _000363_, _000364_, _000365_, _000366_, _000367_, _000368_, _000369_, _000370_, _000371_, _000372_, _000373_, _000374_, _000375_, _000376_, _000377_, _000378_, _000379_, _000380_, _000381_, _000382_, _000383_, _000384_, _000385_, _000386_, _000387_, _000388_, _000389_, _000390_, _000391_, _000392_, _000393_, _000394_, _000395_, _000396_, _000397_, _000398_, _000399_, _000400_, _000401_, _000402_, _000403_, _000404_, _000405_, _000406_, _000407_, _000408_, _000409_, _000410_, _000411_, _000412_, _000413_, _000414_, _000415_, _000416_, _000417_, _000418_, _000419_, _000420_, _000421_, _000422_, _000423_, _000424_, _000425_, _000426_, _000427_, _000428_, _000429_, _000430_, _000431_, _000432_, _000433_, _000434_, _000435_, _000436_, _000437_, _000438_, _000439_, _000440_, _000441_, _000442_, _000443_, _000444_, _000445_, _000446_, _000447_, _000448_, _000449_, _000450_, _000451_, _000452_, _000453_, _000454_, _000455_, _000456_, _000457_, _000458_, _000459_, _000460_, _000461_, _000462_, _000463_, _000464_, _000465_, _000466_, _000467_, _000468_, _000469_, _000470_, _000471_, _000472_, _000473_, _000474_, _000475_, _000476_, _000477_, _000478_, _000479_, _000480_, _000481_, _000482_, _000483_, _000484_, _000485_, _000486_, _000487_, _000488_, _000489_, _000490_, _000491_, _000492_, _000493_, _000494_, _000495_, _000496_, _000497_, _000498_, _000499_, _000500_, _000501_, _000502_, _000503_, _000504_, _000505_, _000506_, _000507_, _000508_, _000509_, _000510_, _000511_, _000512_, _000513_, _000514_, _000515_, _000516_, _000517_, _000518_, _000519_, _000520_, _000521_, _000522_, _000523_, _000524_, _000525_, _000526_, _000527_, _000528_, _000529_, _000530_, _000531_, _000532_, _000533_, _000534_, _000535_, _000536_, _000537_, _000538_, _000539_, _000540_, _000541_, _000542_, _000543_, _000544_, _000545_, _000546_, _000547_, _000548_, _000549_, _000550_, _000551_, _000552_, _000553_, _000554_, _000555_, _000556_, _000557_, _000558_, _000559_, _000560_, _000561_, _000562_, _000563_, _000564_, _000565_, _000566_, _000567_, _000568_, _000569_, _000570_, _000571_, _000572_, _000573_, _000574_, _000575_, _000576_, _000577_, _000578_, _000579_, _000580_, _000581_, _000582_, _000583_, _000584_, _000585_, _000586_, _000587_, _000588_, _000589_, _000590_, _000591_, _000592_, _000593_, _000594_, _000595_, _000596_, _000597_, _000598_, _000599_, _000600_, _000601_, _000602_, _000603_, _000604_, _000605_, _000606_, _000607_, _000608_, _000609_, _000610_, _000611_, _000612_, _000613_, _000614_, _000615_, _000616_, _000617_, _000618_, _000619_, _000620_, _000621_, _000622_, _000623_, _000624_, _000625_, _000626_, _000627_, _000628_, _000629_, _000630_, _000631_, _000632_, _000633_, _000634_, _000635_, _000636_, _000637_, _000638_, _000639_, _000640_, _000641_, _000642_, _000643_, _000644_, _000645_, _000646_, _000647_, _000648_, _000649_, _000650_, _000651_, _000652_, _000653_, _000654_, _000655_, _000656_, _000657_, _000658_, _000659_, _000660_, _000661_, _000662_, _000663_, _000664_, _000665_, _000666_, _000667_, _000668_, _000669_, _000670_, _000671_, _000672_, _000673_, _000674_, _000675_, _000676_, _000677_, _000678_, _000679_, _000680_, _000681_, _000682_, _000683_, _000684_, _000685_, _000686_, _000687_, _000688_, _000689_, _000690_, _000691_, _000692_, _000693_, _000694_, _000695_, _000696_, _000697_, _000698_, _000699_, _000700_, _000701_, _000702_, _000703_, _000704_, _000705_, _000706_, _000707_, _000708_, _000709_, _000710_, _000711_, _000712_, _000713_, _000714_, _000715_, _000716_, _000717_, _000718_, _000719_, _000720_, _000721_, _000722_, _000723_, _000724_, _000725_, _000726_, _000727_, _000728_, _000729_, _000730_, _000731_, _000732_, _000733_, _000734_, _000735_, _000736_, _000737_, _000738_, _000739_, _000740_, _000741_, _000742_, _000743_, _000744_, _000745_, _000746_, _000747_, _000748_, _000749_, _000750_, _000751_, _000752_, _000753_, _000754_, _000755_, _000756_, _000757_, _000758_, _000759_, _000760_, _000761_, _000762_, _000763_, _000764_, _000765_, _000766_, _000767_, _000768_, _000769_, _000770_, _000771_, _000772_, _000773_, _000774_, _000775_, _000776_, _000777_, _000778_, _000779_, _000780_, _000781_, _000782_, _000783_, _000784_, _000785_, _000786_, _000787_, _000788_, _000789_, _000790_, _000791_, _000792_, _000793_, _000794_, _000795_, _000796_, _000797_, _000798_, _000799_, _000800_, _000801_, _000802_, _000803_, _000804_, _000805_, _000806_, _000807_, _000808_, _000809_, _000810_, _000811_, _000812_, _000813_, _000814_, _000815_, _000816_, _000817_, _000818_, _000819_, _000820_, _000821_, _000822_, _000823_, _000824_, _000825_, _000826_, _000827_, _000828_, _000829_, _000830_, _000831_, _000832_, _000833_, _000834_, _000835_, _000836_, _000837_, _000838_, _000839_, _000840_, _000841_, _000842_, _000843_, _000844_, _000845_, _000846_, _000847_, _000848_, _000849_, _000850_, _000851_, _000852_, _000853_, _000854_, _000855_, _000856_, _000857_, _000858_, _000859_, _000860_, _000861_, _000862_, _000863_, _000864_, _000865_, _000866_, _000867_, _000868_, _000869_, _000870_, _000871_, _000872_, _000873_, _000874_, _000875_, _000876_, _000877_, _000878_, _000879_, _000880_, _000881_, _000882_, _000883_, _000884_, _000885_, _000886_, _000887_, _000888_, _000889_, _000890_, _000891_, _000892_, _000893_, _000894_, _000895_, _000896_, _000897_, _000898_, _000899_, _000900_, _000901_, _000902_, _000903_, _000904_, _000905_, _000906_, _000907_, _000908_, _000909_, _000910_, _000911_, _000912_, _000913_, _000914_, _000915_, _000916_, _000917_, _000918_, _000919_, _000920_, _000921_, _000922_, _000923_, _000924_, _000925_, _000926_, _000927_, _000928_, _000929_, _000930_, _000931_, _000932_, _000933_, _000934_, _000935_, _000936_, _000937_, _000938_, _000939_, _000940_, _000941_, _000942_, _000943_, _000944_, _000945_, _000946_, _000947_, _000948_, _000949_, _000950_, _000951_, _000952_, _000953_, _000954_, _000955_, _000956_, _000957_, _000958_, _000959_, _000960_, _000961_, _000962_, _000963_, _000964_, _000965_, _000966_, _000967_, _000968_, _000969_, _000970_, _000971_, _000972_, _000973_, _000974_, _000975_, _000976_, _000977_, _000978_, _000979_, _000980_, _000981_, _000982_, _000983_, _000984_, _000985_, _000986_, _000987_, _000988_, _000989_, _000990_, _000991_, _000992_, _000993_, _000994_, _000995_, _000996_, _000997_, _000998_, _000999_, _001000_, _001001_, _001002_, _001003_, _001004_, _001005_, _001006_, _001007_, _001008_, _001009_, _001010_, _001011_, _001012_, _001013_, _001014_, _001015_, _001016_, _001017_, _001018_, _001019_, _001020_, _001021_, _001022_, _001023_, _001024_, _001025_, _001026_, _001027_, _001028_, _001029_, _001030_, _001031_, _001032_, _001033_, _001034_, _001035_, _001036_, _001037_, _001038_, _001039_, _001040_, _001041_, _001042_, _001043_, _001044_, _001045_, _001046_, _001047_, _001048_, _001049_, _001050_, _001051_, _001052_, _001053_, _001054_, _001055_, _001056_, _001057_, _001058_, _001059_, _001060_, _001061_, _001062_, _001063_, _001064_, _001065_, _001066_, _001067_, _001068_, _001069_, _001070_, _001071_, _001072_, _001073_, _001074_, _001075_, _001076_, _001077_, _001078_, _001079_, _001080_, _001081_, _001082_, _001083_, _001084_, _001085_, _001086_, _001087_, _001088_, _001089_, _001090_, _001091_, _001092_, _001093_, _001094_, _001095_, _001096_, _001097_, _001098_, _001099_, _001100_, _001101_, _001102_, _001103_, _001104_, _001105_, _001106_, _001107_, _001108_, _001109_, _001110_, _001111_, _001112_, _001113_, _001114_, _001115_, _001116_, _001117_, _001118_, _001119_, _001120_, _001121_, _001122_, _001123_, _001124_, _001125_, _001126_, _001127_, _001128_, _001129_, _001130_, _001131_, _001132_, _001133_, _001134_, _001135_, _001136_, _001137_, _001138_, _001139_, _001140_, _001141_, _001142_, _001143_, _001144_, _001145_, _001146_, _001147_, _001148_, _001149_, _001150_, _001151_, _001152_, _001153_, _001154_, _001155_, _001156_, _001157_, _001158_, _001159_, _001160_, _001161_, _001162_, _001163_, _001164_, _001165_, _001166_, _001167_, _001168_, _001169_, _001170_, _001171_, _001172_, _001173_, _001174_, _001175_, _001176_, _001177_, _001178_, _001179_, _001180_, _001181_, _001182_, _001183_, _001184_, _001185_, _001186_, _001187_, _001188_, _001189_, _001190_, _001191_, _001192_, _001193_, _001194_, _001195_, _001196_, _001197_, _001198_, _001199_, _001200_, _001201_, _001202_, _001203_, _001204_, _001205_, _001206_, _001207_, _001208_, _001209_, _001210_, _001211_, _001212_, _001213_, _001214_, _001215_, _001216_, _001217_, _001218_, _001219_, _001220_, _001221_, _001222_, _001223_, _001224_, _001225_, _001226_, _001227_, _001228_, _001229_, _001230_, _001231_, _001232_, _001233_, _001234_, _001235_, _001236_, _001237_, _001238_, _001239_, _001240_, _001241_, _001242_, _001243_, _001244_, _001245_, _001246_, _001247_, _001248_, _001249_, _001250_, _001251_, _001252_, _001253_, _001254_, _001255_, _001256_, _001257_, _001258_, _001259_, _001260_, _001261_, _001262_, _001263_, _001264_, _001265_, _001266_, _001267_, _001268_, _001269_, _001270_, _001271_, _001272_, _001273_, _001274_, _001275_, _001276_, _001277_, _001278_, _001279_, _001280_, _001281_, _001282_, _001283_, _001284_, _001285_, _001286_, _001287_, _001288_, _001289_, _001290_, _001291_, _001292_, _001293_, _001294_, _001295_, _001296_, _001297_, _001298_, _001299_, _001300_, _001301_, _001302_, _001303_, _001304_, _001305_, _001306_, _001307_, _001308_, _001309_, _001310_, _001311_, _001312_, _001313_, _001314_, _001315_, _001316_, _001317_, _001318_, _001319_, _001320_, _001321_, _001322_, _001323_, _001324_, _001325_, _001326_, _001327_, _001328_, _001329_, _001330_, _001331_, _001332_, _001333_, _001334_, _001335_, _001336_, _001337_, _001338_, _001339_, _001340_, _001341_, _001342_, _001343_, _001344_, _001345_, _001346_, _001347_, _001348_, _001349_, _001350_, _001351_, _001352_, _001353_, _001354_, _001355_, _001356_, _001357_, _001358_, _001359_, _001360_, _001361_, _001362_, _001363_, _001364_, _001365_, _001366_, _001367_, _001368_, _001369_, _001370_, _001371_, _001372_, _001373_, _001374_, _001375_, _001376_, _001377_, _001378_, _001379_, _001380_, _001381_, _001382_, _001383_, _001384_, _001385_, _001386_, _001387_, _001388_, _001389_, _001390_, _001391_, _001392_, _001393_, _001394_, _001395_, _001396_, _001397_, _001398_, _001399_, _001400_, _001401_, _001402_, _001403_, _001404_, _001405_, _001406_, _001407_, _001408_, _001409_, _001410_, _001411_, _001412_, _001413_, _001414_, _001415_, _001416_, _001417_, _001418_, _001419_, _001420_, _001421_, _001422_, _001423_, _001424_, _001425_, _001426_, _001427_, _001428_, _001429_, _001430_, _001431_, _001432_, _001433_, _001434_, _001435_, _001436_, _001437_, _001438_, _001439_, _001440_, _001441_, _001442_, _001443_, _001444_, _001445_, _001446_, _001447_, _001448_, _001449_, _001450_, _001451_, _001452_, _001453_, _001454_, _001455_, _001456_, _001457_, _001458_, _001459_, _001460_, _001461_, _001462_, _001463_, _001464_, _001465_, _001466_, _001467_, _001468_, _001469_, _001470_, _001471_, _001472_, _001473_, _001474_, _001475_, _001476_, _001477_, _001478_, _001479_, _001480_, _001481_, _001482_, _001483_, _001484_, _001485_, _001486_, _001487_, _001488_, _001489_, _001490_, _001491_, _001492_, _001493_, _001494_, _001495_, _001496_, _001497_, _001498_, _001499_, _001500_, _001501_, _001502_, _001503_, _001504_, _001505_, _001506_, _001507_, _001508_, _001509_, _001510_, _001511_, _001512_, _001513_, _001514_, _001515_, _001516_, _001517_, _001518_, _001519_, _001520_, _001521_, _001522_, _001523_, _001524_, _001525_, _001526_, _001527_, _001528_, _001529_, _001530_, _001531_, _001532_, _001533_, _001534_, _001535_, _001536_, _001537_, _001538_, _001539_, _001540_, _001541_, _001542_, _001543_, _001544_, _001545_, _001546_, _001547_, _001548_, _001549_, _001550_, _001551_, _001552_, _001553_, _001554_, _001555_, _001556_, _001557_, _001558_, _001559_, _001560_, _001561_, _001562_, _001563_, _001564_, _001565_, _001566_, _001567_, _001568_, _001569_, _001570_, _001571_, _001572_, _001573_, _001574_, _001575_, _001576_, _001577_, _001578_, _001579_, _001580_, _001581_, _001582_, _001583_, _001584_, _001585_, _001586_, _001587_, _001588_, _001589_, _001590_, _001591_, _001592_, _001593_, _001594_, _001595_, _001596_, _001597_, _001598_, _001599_, _001600_, _001601_, _001602_, _001603_, _001604_, _001605_, _001606_, _001607_, _001608_, _001609_, _001610_, _001611_, _001612_, _001613_, _001614_, _001615_, _001616_, _001617_, _001618_, _001619_, _001620_, _001621_, _001622_, _001623_, _001624_, _001625_, _001626_, _001627_, _001628_, _001629_, _001630_, _001631_, _001632_, _001633_, _001634_, _001635_, _001636_, _001637_, _001638_, _001639_, _001640_, _001641_, _001642_, _001643_, _001644_, _001645_, _001646_, _001647_, _001648_, _001649_, _001650_, _001651_, _001652_, _001653_, _001654_, _001655_, _001656_, _001657_, _001658_, _001659_, _001660_, _001661_, _001662_, _001663_, _001664_, _001665_, _001666_, _001667_, _001668_, _001669_, _001670_, _001671_, _001672_, _001673_, _001674_, _001675_, _001676_, _001677_, _001678_, _001679_, _001680_, _001681_, _001682_, _001683_, _001684_, _001685_, _001686_, _001687_, _001688_, _001689_, _001690_, _001691_, _001692_, _001693_, _001694_, _001695_, _001696_, _001697_, _001698_, _001699_, _001700_, _001701_, _001702_, _001703_, _001704_, _001705_, _001706_, _001707_, _001708_, _001709_, _001710_, _001711_, _001712_, _001713_, _001714_, _001715_, _001716_, _001717_, _001718_, _001719_, _001720_, _001721_, _001722_, _001723_, _001724_, _001725_, _001726_, _001727_, _001728_, _001729_, _001730_, _001731_, _001732_, _001733_, _001734_, _001735_, _001736_, _001737_, _001738_, _001739_, _001740_, _001741_, _001742_, _001743_, _001744_, _001745_, _001746_, _001747_, _001748_, _001749_, _001750_, _001751_, _001752_, _001753_, _001754_, _001755_, _001756_, _001757_, _001758_, _001759_, _001760_, _001761_, _001762_, _001763_, _001764_, _001765_, _001766_, _001767_, _001768_, _001769_, _001770_, _001771_, _001772_, _001773_, _001774_, _001775_, _001776_, _001777_, _001778_, _001779_, _001780_, _001781_, _001782_, _001783_, _001784_, _001785_, _001786_, _001787_, _001788_, _001789_, _001790_, _001791_, _001792_, _001793_, _001794_, _001795_, _001796_, _001797_, _001798_, _001799_, _001800_, _001801_, _001802_, _001803_, _001804_, _001805_, _001806_, _001807_, _001808_, _001809_, _001810_, _001811_, _001812_, _001813_, _001814_, _001815_, _001816_, _001817_, _001818_, _001819_, _001820_, _001821_, _001822_, _001823_, _001824_, _001825_, _001826_, _001827_, _001828_, _001829_, _001830_, _001831_, _001832_, _001833_, _001834_, _001835_, _001836_, _001837_, _001838_, _001839_, _001840_, _001841_, _001842_, _001843_, _001844_, _001845_, _001846_, _001847_, _001848_, _001849_, _001850_, _001851_, _001852_, _001853_, _001854_, _001855_, _001856_, _001857_, _001858_, _001859_, _001860_, _001861_, _001862_, _001863_, _001864_, _001865_, _001866_, _001867_, _001868_, _001869_, _001870_, _001871_, _001872_, _001873_, _001874_, _001875_, _001876_, _001877_, _001878_, _001879_, _001880_, _001881_, _001882_, _001883_, _001884_, _001885_, _001886_, _001887_, _001888_, _001889_, _001890_, _001891_, _001892_, _001893_, _001894_, _001895_, _001896_, _001897_, _001898_, _001899_, _001900_, _001901_, _001902_, _001903_, _001904_, _001905_, _001906_, _001907_, _001908_, _001909_, _001910_, _001911_, _001912_, _001913_, _001914_, _001915_, _001916_, _001917_, _001918_, _001919_, _001920_, _001921_, _001922_, _001923_, _001924_, _001925_, _001926_, _001927_, _001928_, _001929_, _001930_, _001931_, _001932_, _001933_, _001934_, _001935_, _001936_, _001937_, _001938_, _001939_, _001940_, _001941_, _001942_, _001943_, _001944_, _001945_, _001946_, _001947_, _001948_, _001949_, _001950_, _001951_, _001952_, _001953_, _001954_, _001955_, _001956_, _001957_, _001958_, _001959_, _001960_, _001961_, _001962_, _001963_, _001964_, _001965_, _001966_, _001967_, _001968_, _001969_, _001970_, _001971_, _001972_, _001973_, _001974_, _001975_, _001976_, _001977_, _001978_, _001979_, _001980_, _001981_, _001982_, _001983_, _001984_, _001985_, _001986_, _001987_, _001988_, _001989_, _001990_, _001991_, _001992_, _001993_, _001994_, _001995_, _001996_, _001997_, _001998_, _001999_, _002000_, _002001_, _002002_, _002003_, _002004_, _002005_, _002006_, _002007_, _002008_, _002009_, _002010_, _002011_, _002012_, _002013_, _002014_, _002015_, _002016_, _002017_, _002018_, _002019_, _002020_, _002021_, _002022_, _002023_, _002024_, _002025_, _002026_, _002027_, _002028_, _002029_, _002030_, _002031_, _002032_, _002033_, _002034_, _002035_, _002036_, _002037_, _002038_, _002039_, _002040_, _002041_, _002042_, _002043_, _002044_, _002045_, _002046_, _002047_, _002048_, _002049_, _002050_, _002051_, _002052_, _002053_, _002054_, _002055_, _002056_, _002057_, _002058_, _002059_, _002060_, _002061_, _002062_, _002063_, _002064_, _002065_, _002066_, _002067_, _002068_, _002069_, _002070_, _002071_, _002072_, _002073_, _002074_, _002075_, _002076_, _002077_, _002078_, _002079_, _002080_, _002081_, _002082_, _002083_, _002084_, _002085_, _002086_, _002087_, _002088_, _002089_, _002090_, _002091_, _002092_, _002093_, _002094_, _002095_, _002096_, _002097_, _002098_, _002099_, _002100_, _002101_, _002102_, _002103_, _002104_, _002105_, _002106_, _002107_, _002108_, _002109_, _002110_, _002111_, _002112_, _002113_, _002114_, _002115_, _002116_, _002117_, _002118_, _002119_, _002120_, _002121_, _002122_, _002123_, _002124_, _002125_, _002126_, _002127_, _002128_, _002129_, _002130_, _002131_, _002132_, _002133_, _002134_, _002135_, _002136_, _002137_, _002138_, _002139_, _002140_, _002141_, _002142_, _002143_, _002144_, _002145_, _002146_, _002147_, _002148_, _002149_, _002150_, _002151_, _002152_, _002153_, _002154_, _002155_, _002156_, _002157_, _002158_, _002159_, _002160_, _002161_, _002162_, _002163_, _002164_, _002165_, _002166_, _002167_, _002168_, _002169_, _002170_, _002171_, _002172_, _002173_, _002174_, _002175_, _002176_, _002177_, _002178_, _002179_, _002180_, _002181_, _002182_, _002183_, _002184_, _002185_, _002186_, _002187_, _002188_, _002189_, _002190_, _002191_, _002192_, _002193_, _002194_, _002195_, _002196_, _002197_, _002198_, _002199_, _002200_, _002201_, _002202_, _002203_, _002204_, _002205_, _002206_, _002207_, _002208_, _002209_, _002210_, _002211_, _002212_, _002213_, _002214_, _002215_, _002216_, _002217_, _002218_, _002219_, _002220_, _002221_, _002222_, _002223_, _002224_, _002225_, _002226_, _002227_, _002228_, _002229_, _002230_, _002231_, _002232_, _002233_, _002234_, _002235_, _002236_, _002237_, _002238_, _002239_, _002240_, _002241_, _002242_, _002243_, _002244_, _002245_, _002246_, _002247_, _002248_, _002249_, _002250_, _002251_, _002252_, _002253_, _002254_, _002255_, _002256_, _002257_, _002258_, _002259_, _002260_, _002261_, _002262_, _002263_, _002264_, _002265_, _002266_, _002267_, _002268_, _002269_, _002270_, _002271_, _002272_, _002273_, _002274_, _002275_, _002276_, _002277_, _002278_, _002279_, _002280_, _002281_, _002282_, _002283_, _002284_, _002285_, _002286_, _002287_, _002288_, _002289_, _002290_, _002291_, _002292_, _002293_, _002294_, _002295_, _002296_, _002297_, _002298_, _002299_, _002300_, _002301_, _002302_, _002303_, _002304_, _002305_, _002306_, _002307_, _002308_, _002309_, _002310_, _002311_, _002312_, _002313_, _002314_, _002315_, _002316_, _002317_, _002318_, _002319_, _002320_, _002321_, _002322_, _002323_, _002324_, _002325_, _002326_, _002327_, _002328_, _002329_, _002330_, _002331_, _002332_, _002333_, _002334_, _002335_, _002336_, _002337_, _002338_, _002339_, _002340_, _002341_, _002342_, _002343_, _002344_, _002345_, _002346_, _002347_, _002348_, _002349_, _002350_, _002351_, _002352_, _002353_, _002354_, _002355_, _002356_, _002357_, _002358_, _002359_, _002360_, _002361_, _002362_, _002363_, _002364_, _002365_, _002366_, _002367_, _002368_, _002369_, _002370_, _002371_, _002372_, _002373_, _002374_, _002375_, _002376_, _002377_, _002378_, _002379_, _002380_, _002381_, _002382_, _002383_, _002384_, _002385_, _002386_, _002387_, _002388_, _002389_, _002390_, _002391_, _002392_, _002393_, _002394_, _002395_, _002396_, _002397_, _002398_, _002399_, _002400_, _002401_, _002402_, _002403_, _002404_, _002405_, _002406_, _002407_, _002408_, _002409_, _002410_, _002411_, _002412_, _002413_, _002414_, _002415_, _002416_, _002417_, _002418_, _002419_, _002420_, _002421_, _002422_, _002423_, _002424_, _002425_, _002426_, _002427_, _002428_, _002429_, _002430_, _002431_, _002432_, _002433_, _002434_, _002435_, _002436_, _002437_, _002438_, _002439_, _002440_, _002441_, _002442_, _002443_, _002444_, _002445_, _002446_, _002447_, _002448_, _002449_, _002450_, _002451_, _002452_, _002453_, _002454_, _002455_, _002456_, _002457_, _002458_, _002459_, _002460_, _002461_, _002462_, _002463_, _002464_, _002465_, _002466_, _002467_, _002468_, _002469_, _002470_, _002471_, _002472_, _002473_, _002474_, _002475_, _002476_, _002477_, _002478_, _002479_, _002480_, _002481_, _002482_, _002483_, _002484_, _002485_, _002486_, _002487_, _002488_, _002489_, _002490_, _002491_, _002492_, _002493_, _002494_, _002495_, _002496_, _002497_, _002498_, _002499_, _002500_, _002501_, _002502_, _002503_, _002504_, _002505_, _002506_, _002507_, _002508_, _002509_, _002510_, _002511_, _002512_, _002513_, _002514_, _002515_, _002516_, _002517_, _002518_, _002519_, _002520_, _002521_, _002522_, _002523_, _002524_, _002525_, _002526_, _002527_, _002528_, _002529_, _002530_, _002531_, _002532_, _002533_, _002534_, _002535_, _002536_, _002537_, _002538_, _002539_, _002540_, _002541_, _002542_, _002543_, _002544_, _002545_, _002546_, _002547_, _002548_, _002549_, _002550_, _002551_, _002552_, _002553_, _002554_, _002555_, _002556_, _002557_, _002558_, _002559_, _002560_, _002561_, _002562_, _002563_, _002564_, _002565_, _002566_, _002567_, _002568_, _002569_, _002570_, _002571_, _002572_, _002573_, _002574_, _002575_, _002576_, _002577_, _002578_, _002579_, _002580_, _002581_, _002582_, _002583_, _002584_, _002585_, _002586_, _002587_, _002588_, _002589_, _002590_, _002591_, _002592_, _002593_, _002594_, _002595_, _002596_, _002597_, _002598_, _002599_, _002600_, _002601_, _002602_, _002603_, _002604_, _002605_, _002606_, _002607_, _002608_, _002609_, _002610_, _002611_, _002612_, _002613_, _002614_, _002615_, _002616_, _002617_, _002618_, _002619_, _002620_, _002621_, _002622_, _002623_, _002624_, _002625_, _002626_, _002627_, _002628_, _002629_, _002630_, _002631_, _002632_, _002633_, _002634_, _002635_, _002636_, _002637_, _002638_, _002639_, _002640_, _002641_, _002642_, _002643_, _002644_, _002645_, _002646_, _002647_, _002648_, _002649_, _002650_, _002651_, _002652_, _002653_, _002654_, _002655_, _002656_, _002657_, _002658_, _002659_, _002660_, _002661_, _002662_, _002663_, _002664_, _002665_, _002666_, _002667_, _002668_, _002669_, _002670_, _002671_, _002672_, _002673_, _002674_, _002675_, _002676_, _002677_, _002678_, _002679_, _002680_, _002681_, _002682_, _002683_, _002684_, _002685_, _002686_, _002687_, _002688_, _002689_, _002690_, _002691_, _002692_, _002693_, _002694_, _002695_, _002696_, _002697_, _002698_, _002699_, _002700_, _002701_, _002702_, _002703_, _002704_, _002705_, _002706_, _002707_, _002708_, _002709_, _002710_, _002711_, _002712_, _002713_, _002714_, _002715_, _002716_, _002717_, _002718_, _002719_, _002720_, _002721_, _002722_, _002723_, _002724_, _002725_, _002726_, _002727_, _002728_, _002729_, _002730_, _002731_, _002732_, _002733_, _002734_, _002735_, _002736_, _002737_, _002738_, _002739_, _002740_, _002741_, _002742_, _002743_, _002744_, _002745_, _002746_, _002747_, _002748_, _002749_, _002750_, _002751_, _002752_, _002753_, _002754_, _002755_, _002756_, _002757_, _002758_, _002759_, _002760_, _002761_, _002762_, _002763_, _002764_, _002765_, _002766_, _002767_, _002768_, _002769_, _002770_, _002771_, _002772_, _002773_, _002774_, _002775_, _002776_, _002777_, _002778_, _002779_, _002780_, _002781_, _002782_, _002783_, _002784_, _002785_, _002786_, _002787_, _002788_, _002789_, _002790_, _002791_, _002792_, _002793_, _002794_, _002795_, _002796_, _002797_, _002798_, _002799_, _002800_, _002801_, _002802_, _002803_, _002804_, _002805_, _002806_, _002807_, _002808_, _002809_, _002810_, _002811_, _002812_, _002813_, _002814_, _002815_, _002816_, _002817_, _002818_, _002819_, _002820_, _002821_, _002822_, _002823_, _002824_, _002825_, _002826_, _002827_, _002828_, _002829_, _002830_, _002831_, _002832_, _002833_, _002834_, _002835_, _002836_, _002837_, _002838_, _002839_, _002840_, _002841_, _002842_, _002843_, _002844_, _002845_, _002846_, _002847_, _002848_, _002849_, _002850_, _002851_, _002852_, _002853_, _002854_, _002855_, _002856_, _002857_, _002858_, _002859_, _002860_, _002861_, _002862_, _002863_, _002864_, _002865_, _002866_, _002867_, _002868_, _002869_, _002870_, _002871_, _002872_, _002873_, _002874_, _002875_, _002876_, _002877_, _002878_, _002879_, _002880_, _002881_, _002882_, _002883_, _002884_, _002885_, _002886_, _002887_, _002888_, _002889_, _002890_, _002891_, _002892_, _002893_, _002894_, _002895_, _002896_, _002897_, _002898_, _002899_, _002900_, _002901_, _002902_, _002903_, _002904_, _002905_, _002906_, _002907_, _002908_, _002909_, _002910_, _002911_, _002912_, _002913_, _002914_, _002915_, _002916_, _002917_, _002918_, _002919_, _002920_, _002921_, _002922_, _002923_, _002924_, _002925_, _002926_, _002927_, _002928_, _002929_, _002930_, _002931_, _002932_, _002933_, _002934_, _002935_, _002936_, _002937_, _002938_, _002939_, _002940_, _002941_, _002942_, _002943_, _002944_, _002945_, _002946_, _002947_, _002948_, _002949_, _002950_, _002951_, _002952_, _002953_, _002954_, _002955_, _002956_, _002957_, _002958_, _002959_, _002960_, _002961_, _002962_, _002963_, _002964_, _002965_, _002966_, _002967_, _002968_, _002969_, _002970_, _002971_, _002972_, _002973_, _002974_, _002975_, _002976_, _002977_, _002978_, _002979_, _002980_, _002981_, _002982_, _002983_, _002984_, _002985_, _002986_, _002987_, _002988_, _002989_, _002990_, _002991_, _002992_, _002993_, _002994_, _002995_, _002996_, _002997_, _002998_, _002999_, _003000_, _003001_, _003002_, _003003_, _003004_, _003005_, _003006_, _003007_, _003008_, _003009_, _003010_, _003011_, _003012_, _003013_, _003014_, _003015_, _003016_, _003017_, _003018_, _003019_, _003020_, _003021_, _003022_, _003023_, _003024_, _003025_, _003026_, _003027_, _003028_, _003029_, _003030_, _003031_, _003032_, _003033_, _003034_, _003035_, _003036_, _003037_, _003038_, _003039_, _003040_, _003041_, _003042_, _003043_, _003044_, _003045_, _003046_, _003047_, _003048_, _003049_, _003050_, _003051_, _003052_, _003053_, _003054_, _003055_, _003056_, _003057_, _003058_, _003059_, _003060_, _003061_, _003062_, _003063_, _003064_, _003065_, _003066_, _003067_, _003068_, _003069_, _003070_, _003071_, _003072_, _003073_, _003074_, _003075_, _003076_, _003077_, _003078_, _003079_, _003080_, _003081_, _003082_, _003083_, _003084_, _003085_, _003086_, _003087_, _003088_, _003089_, _003090_, _003091_, _003092_, _003093_, _003094_, _003095_, _003096_, _003097_, _003098_, _003099_, _003100_, _003101_, _003102_, _003103_, _003104_, _003105_, _003106_, _003107_, _003108_, _003109_, _003110_, _003111_, _003112_, _003113_, _003114_, _003115_, _003116_, _003117_, _003118_, _003119_, _003120_, _003121_, _003122_, _003123_, _003124_, _003125_, _003126_, _003127_, _003128_, _003129_, _003130_, _003131_, _003132_, _003133_, _003134_, _003135_, _003136_, _003137_, _003138_, _003139_, _003140_, _003141_, _003142_, _003143_, _003144_, _003145_, _003146_, _003147_, _003148_, _003149_, _003150_, _003151_, _003152_, _003153_, _003154_, _003155_, _003156_, _003157_, _003158_, _003159_, _003160_, _003161_, _003162_, _003163_, _003164_, _003165_, _003166_, _003167_, _003168_, _003169_, _003170_, _003171_, _003172_, _003173_, _003174_, _003175_, _003176_, _003177_, _003178_, _003179_, _003180_, _003181_, _003182_, _003183_, _003184_, _003185_, _003186_, _003187_, _003188_, _003189_, _003190_, _003191_, _003192_, _003193_, _003194_, _003195_, _003196_, _003197_, _003198_, _003199_, _003200_, _003201_, _003202_, _003203_, _003204_, _003205_, _003206_, _003207_, _003208_, _003209_, _003210_, _003211_, _003212_, _003213_, _003214_, _003215_, _003216_, _003217_, _003218_, _003219_, _003220_, _003221_, _003222_, _003223_, _003224_, _003225_, _003226_, _003227_, _003228_, _003229_, _003230_, _003231_, _003232_, _003233_, _003234_, _003235_, _003236_, _003237_, _003238_, _003239_, _003240_, _003241_, _003242_, _003243_, _003244_, _003245_, _003246_, _003247_, _003248_, _003249_, _003250_, _003251_, _003252_, _003253_, _003254_, _003255_, _003256_, _003257_, _003258_, _003259_, _003260_, _003261_, _003262_, _003263_, _003264_, _003265_, _003266_, _003267_, _003268_, _003269_, _003270_, _003271_, _003272_, _003273_, _003274_, _003275_, _003276_, _003277_, _003278_, _003279_, _003280_, _003281_, _003282_, _003283_, _003284_, _003285_, _003286_, _003287_, _003288_, _003289_, _003290_, _003291_, _003292_, _003293_, _003294_, _003295_, _003296_, _003297_, _003298_, _003299_, _003300_, _003301_, _003302_, _003303_, _003304_, _003305_, _003306_, _003307_, _003308_, _003309_, _003310_, _003311_, _003312_, _003313_, _003314_, _003315_, _003316_, _003317_, _003318_, _003319_, _003320_, _003321_, _003322_, _003323_, _003324_, _003325_, _003326_, _003327_, _003328_, _003329_, _003330_, _003331_, _003332_, _003333_, _003334_, _003335_, _003336_, _003337_, _003338_, _003339_, _003340_, _003341_, _003342_, _003343_, _003344_, _003345_, _003346_, _003347_, _003348_, _003349_, _003350_, _003351_, _003352_, _003353_, _003354_, _003355_, _003356_, _003357_, _003358_, _003359_, _003360_, _003361_, _003362_, _003363_, _003364_, _003365_, _003366_, _003367_, _003368_, _003369_, _003370_, _003371_, _003372_, _003373_, _003374_, _003375_, _003376_, _003377_, _003378_, _003379_, _003380_, _003381_, _003382_, _003383_, _003384_, _003385_, _003386_, _003387_, _003388_, _003389_, _003390_, _003391_, _003392_, _003393_, _003394_, _003395_, _003396_, _003397_, _003398_, _003399_, _003400_, _003401_, _003402_, _003403_, _003404_, _003405_, _003406_, _003407_, _003408_, _003409_, _003410_, _003411_, _003412_, _003413_, _003414_, _003415_, _003416_, _003417_, _003418_, _003419_, _003420_, _003421_, _003422_, _003423_, _003424_, _003425_, _003426_, _003427_, _003428_, _003429_, _003430_, _003431_, _003432_, _003433_, _003434_, _003435_, _003436_, _003437_, _003438_, _003439_, _003440_, _003441_, _003442_, _003443_, _003444_, _003445_, _003446_, _003447_, _003448_, _003449_, _003450_, _003451_, _003452_, _003453_, _003454_, _003455_, _003456_, _003457_, _003458_, _003459_, _003460_, _003461_, _003462_, _003463_, _003464_, _003465_, _003466_, _003467_, _003468_, _003469_, _003470_, _003471_, _003472_, _003473_, _003474_, _003475_, _003476_, _003477_, _003478_, _003479_, _003480_, _003481_, _003482_, _003483_, _003484_, _003485_, _003486_, _003487_, _003488_, _003489_, _003490_, _003491_, _003492_, _003493_, _003494_, _003495_, _003496_, _003497_, _003498_, _003499_, _003500_, _003501_, _003502_, _003503_, _003504_, _003505_, _003506_, _003507_, _003508_, _003509_, _003510_, _003511_, _003512_, _003513_, _003514_, _003515_, _003516_, _003517_, _003518_, _003519_, _003520_, _003521_, _003522_, _003523_, _003524_, _003525_, _003526_, _003527_, _003528_, _003529_, _003530_, _003531_, _003532_, _003533_, _003534_, _003535_, _003536_, _003537_, _003538_, _003539_, _003540_, _003541_, _003542_, _003543_, _003544_, _003545_, _003546_, _003547_, _003548_, _003549_, _003550_, _003551_, _003552_, _003553_, _003554_, _003555_, _003556_, _003557_, _003558_, _003559_, _003560_, _003561_, _003562_, _003563_, _003564_, _003565_, _003566_, _003567_, _003568_, _003569_, _003570_, _003571_, _003572_, _003573_, _003574_, _003575_, _003576_, _003577_, _003578_, _003579_, _003580_, _003581_, _003582_, _003583_, _003584_, _003585_, _003586_, _003587_, _003588_, _003589_, _003590_, _003591_, _003592_, _003593_, _003594_, _003595_, _003596_, _003597_, _003598_, _003599_, _003600_, _003601_, _003602_, _003603_, _003604_, _003605_, _003606_, _003607_, _003608_, _003609_, _003610_, _003611_, _003612_, _003613_, _003614_, _003615_, _003616_, _003617_, _003618_, _003619_, _003620_, _003621_, _003622_, _003623_, _003624_, _003625_, _003626_, _003627_, _003628_, _003629_, _003630_, _003631_, _003632_, _003633_, _003634_, _003635_, _003636_, _003637_, _003638_, _003639_, _003640_, _003641_, _003642_, _003643_, _003644_, _003645_, _003646_, _003647_, _003648_, _003649_, _003650_, _003651_, _003652_, _003653_, _003654_, _003655_, _003656_, _003657_, _003658_, _003659_, _003660_, _003661_, _003662_, _003663_, _003664_, _003665_, _003666_, _003667_, _003668_, _003669_, _003670_, _003671_, _003672_, _003673_, _003674_, _003675_, _003676_, _003677_, _003678_, _003679_, _003680_, _003681_, _003682_, _003683_, _003684_, _003685_, _003686_, _003687_, _003688_, _003689_, _003690_, _003691_, _003692_, _003693_, _003694_, _003695_, _003696_, _003697_, _003698_, _003699_, _003700_, _003701_, _003702_, _003703_, _003704_, _003705_, _003706_, _003707_, _003708_, _003709_, _003710_, _003711_, _003712_, _003713_, _003714_, _003715_, _003716_, _003717_, _003718_, _003719_, _003720_, _003721_, _003722_, _003723_, _003724_, _003725_, _003726_, _003727_, _003728_, _003729_, _003730_, _003731_, _003732_, _003733_, _003734_, _003735_, _003736_, _003737_, _003738_, _003739_, _003740_, _003741_, _003742_, _003743_, _003744_, _003745_, _003746_, _003747_, _003748_, _003749_, _003750_, _003751_, _003752_, _003753_, _003754_, _003755_, _003756_, _003757_, _003758_, _003759_, _003760_, _003761_, _003762_, _003763_, _003764_, _003765_, _003766_, _003767_, _003768_, _003769_, _003770_, _003771_, _003772_, _003773_, _003774_, _003775_, _003776_, _003777_, _003778_, _003779_, _003780_, _003781_, _003782_, _003783_, _003784_, _003785_, _003786_, _003787_, _003788_, _003789_, _003790_, _003791_, _003792_, _003793_, _003794_, _003795_, _003796_, _003797_, _003798_, _003799_, _003800_, _003801_, _003802_, _003803_, _003804_, _003805_, _003806_, _003807_, _003808_, _003809_, _003810_, _003811_, _003812_, _003813_, _003814_, _003815_, _003816_, _003817_, _003818_, _003819_, _003820_, _003821_, _003822_, _003823_, _003824_, _003825_, _003826_, _003827_, _003828_, _003829_, _003830_, _003831_, _003832_, _003833_, _003834_, _003835_, _003836_, _003837_, _003838_, _003839_, _003840_, _003841_, _003842_, _003843_, _003844_, _003845_, _003846_, _003847_, _003848_, _003849_, _003850_, _003851_, _003852_, _003853_, _003854_, _003855_, _003856_, _003857_, _003858_, _003859_, _003860_, _003861_, _003862_, _003863_, _003864_, _003865_, _003866_, _003867_, _003868_, _003869_, _003870_, _003871_, _003872_, _003873_, _003874_, _003875_, _003876_, _003877_, _003878_, _003879_, _003880_, _003881_, _003882_, _003883_, _003884_, _003885_, _003886_, _003887_, _003888_, _003889_, _003890_, _003891_, _003892_, _003893_, _003894_, _003895_, _003896_, _003897_, _003898_, _003899_, _003900_, _003901_, _003902_, _003903_, _003904_, _003905_, _003906_, _003907_, _003908_, _003909_, _003910_, _003911_, _003912_, _003913_, _003914_, _003915_, _003916_, _003917_, _003918_, _003919_, _003920_, _003921_, _003922_, _003923_, _003924_, _003925_, _003926_, _003927_, _003928_, _003929_, _003930_, _003931_, _003932_, _003933_, _003934_, _003935_, _003936_, _003937_, _003938_, _003939_, _003940_, _003941_, _003942_, _003943_, _003944_, _003945_, _003946_, _003947_, _003948_, _003949_, _003950_, _003951_, _003952_, _003953_, _003954_, _003955_, _003956_, _003957_, _003958_, _003959_, _003960_, _003961_, _003962_, _003963_, _003964_, _003965_, _003966_, _003967_, _003968_, _003969_, _003970_, _003971_, _003972_, _003973_, _003974_, _003975_, _003976_, _003977_, _003978_, _003979_, _003980_, _003981_, _003982_, _003983_, _003984_, _003985_, _003986_, _003987_, _003988_, _003989_, _003990_, _003991_, _003992_, _003993_, _003994_, _003995_, _003996_, _003997_, _003998_, _003999_, _004000_, _004001_, _004002_, _004003_, _004004_, _004005_, _004006_, _004007_, _004008_, _004009_, _004010_, _004011_, _004012_, _004013_, _004014_, _004015_, _004016_, _004017_, _004018_, _004019_, _004020_, _004021_, _004022_, _004023_, _004024_, _004025_, _004026_, _004027_, _004028_, _004029_, _004030_, _004031_, _004032_, _004033_, _004034_, _004035_, _004036_, _004037_, _004038_, _004039_, _004040_, _004041_, _004042_, _004043_, _004044_, _004045_, _004046_, _004047_, _004048_, _004049_, _004050_, _004051_, _004052_, _004053_, _004054_, _004055_, _004056_, _004057_, _004058_, _004059_, _004060_, _004061_, _004062_, _004063_, _004064_, _004065_, _004066_, _004067_, _004068_, _004069_, _004070_, _004071_, _004072_, _004073_, _004074_, _004075_, _004076_, _004077_, _004078_, _004079_, _004080_, _004081_, _004082_, _004083_, _004084_, _004085_, _004086_, _004087_, _004088_, _004089_, _004090_, _004091_, _004092_, _004093_, _004094_, _004095_, _004096_, _004097_, _004098_, _004099_, _004100_, _004101_, _004102_, _004103_, _004104_, _004105_, _004106_, _004107_, _004108_, _004109_, _004110_, _004111_, _004112_, _004113_, _004114_, _004115_, _004116_, _004117_, _004118_, _004119_, _004120_, _004121_, _004122_, _004123_, _004124_, _004125_, _004126_, _004127_, _004128_, _004129_, _004130_, _004131_, _004132_, _004133_, _004134_, _004135_, _004136_, _004137_, _004138_, _004139_, _004140_, _004141_, _004142_, _004143_, _004144_, _004145_, _004146_, _004147_, _004148_, _004149_, _004150_, _004151_, _004152_, _004153_, _004154_, _004155_, _004156_, _004157_, _004158_, _004159_, _004160_, _004161_, _004162_, _004163_, _004164_, _004165_, _004166_, _004167_, _004168_, _004169_, _004170_, _004171_, _004172_, _004173_, _004174_, _004175_, _004176_, _004177_, _004178_, _004179_, _004180_, _004181_, _004182_, _004183_, _004184_, _004185_, _004186_, _004187_, _004188_, _004189_, _004190_, _004191_, _004192_, _004193_, _004194_, _004195_, _004196_, _004197_, _004198_, _004199_, _004200_, _004201_, _004202_, _004203_, _004204_, _004205_, _004206_, _004207_, _004208_, _004209_, _004210_, _004211_, _004212_, _004213_, _004214_, _004215_, _004216_, _004217_, _004218_, _004219_, _004220_, _004221_, _004222_, _004223_, _004224_, _004225_, _004226_, _004227_, _004228_, _004229_, _004230_, _004231_, _004232_, _004233_, _004234_, _004235_, _004236_, _004237_, _004238_, _004239_, _004240_, _004241_, _004242_, _004243_, _004244_, _004245_, _004246_, _004247_, _004248_, _004249_, _004250_, _004251_, _004252_, _004253_, _004254_, _004255_, _004256_, _004257_, _004258_, _004259_, _004260_, _004261_, _004262_, _004263_, _004264_, _004265_, _004266_, _004267_, _004268_, _004269_, _004270_, _004271_, _004272_, _004273_, _004274_, _004275_, _004276_, _004277_, _004278_, _004279_, _004280_, _004281_, _004282_, _004283_, _004284_, _004285_, _004286_, _004287_, _004288_, _004289_, _004290_, _004291_, _004292_, _004293_, _004294_, _004295_, _004296_, _004297_, _004298_, _004299_, _004300_, _004301_, _004302_, _004303_, _004304_, _004305_, _004306_, _004307_, _004308_, _004309_, _004310_, _004311_, _004312_, _004313_, _004314_, _004315_, _004316_, _004317_, _004318_, _004319_, _004320_, _004321_, _004322_, _004323_, _004324_, _004325_, _004326_, _004327_, _004328_, _004329_, _004330_, _004331_, _004332_, _004333_, _004334_, _004335_, _004336_, _004337_, _004338_, _004339_, _004340_, _004341_, _004342_, _004343_, _004344_, _004345_, _004346_, _004347_, _004348_, _004349_, _004350_, _004351_, _004352_, _004353_, _004354_, _004355_, _004356_, _004357_, _004358_, _004359_, _004360_, _004361_, _004362_, _004363_, _004364_, _004365_, _004366_, _004367_, _004368_, _004369_, _004370_, _004371_, _004372_, _004373_, _004374_, _004375_, _004376_, _004377_, _004378_, _004379_, _004380_, _004381_, _004382_, _004383_, _004384_, _004385_, _004386_, _004387_, _004388_, _004389_, _004390_, _004391_, _004392_, _004393_, _004394_, _004395_, _004396_, _004397_, _004398_, _004399_, _004400_, _004401_, _004402_, _004403_, _004404_, _004405_, _004406_, _004407_, _004408_, _004409_, _004410_, _004411_, _004412_, _004413_, _004414_, _004415_, _004416_, _004417_, _004418_, _004419_, _004420_, _004421_, _004422_, _004423_, _004424_, _004425_, _004426_, _004427_, _004428_, _004429_, _004430_, _004431_, _004432_, _004433_, _004434_, _004435_, _004436_, _004437_, _004438_, _004439_, _004440_, _004441_, _004442_, _004443_, _004444_, _004445_, _004446_, _004447_, _004448_, _004449_, _004450_, _004451_, _004452_, _004453_, _004454_, _004455_, _004456_, _004457_, _004458_, _004459_, _004460_, _004461_, _004462_, _004463_, _004464_, _004465_, _004466_, _004467_, _004468_, _004469_, _004470_, _004471_, _004472_, _004473_, _004474_, _004475_, _004476_, _004477_, _004478_, _004479_, _004480_, _004481_, _004482_, _004483_, _004484_, _004485_, _004486_, _004487_, _004488_, _004489_, _004490_, _004491_, _004492_, _004493_, _004494_, _004495_, _004496_, _004497_, _004498_, _004499_, _004500_, _004501_, _004502_, _004503_, _004504_, _004505_, _004506_, _004507_, _004508_, _004509_, _004510_, _004511_, _004512_, _004513_, _004514_, _004515_, _004516_, _004517_, _004518_, _004519_, _004520_, _004521_, _004522_, _004523_, _004524_, _004525_, _004526_, _004527_, _004528_, _004529_, _004530_, _004531_, _004532_, _004533_, _004534_, _004535_, _004536_, _004537_, _004538_, _004539_, _004540_, _004541_, _004542_, _004543_, _004544_, _004545_, _004546_, _004547_, _004548_, _004549_, _004550_, _004551_, _004552_, _004553_, _004554_, _004555_, _004556_, _004557_, _004558_, _004559_, _004560_, _004561_, _004562_, _004563_, _004564_, _004565_, _004566_, _004567_, _004568_, _004569_, _004570_, _004571_, _004572_, _004573_, _004574_, _004575_, _004576_, _004577_, _004578_, _004579_, _004580_, _004581_, _004582_, _004583_, _004584_, _004585_, _004586_, _004587_, _004588_, _004589_, _004590_, _004591_, _004592_, _004593_, _004594_, _004595_, _004596_, _004597_, _004598_, _004599_, _004600_, _004601_, _004602_, _004603_, _004604_, _004605_, _004606_, _004607_, _004608_, _004609_, _004610_, _004611_, _004612_, _004613_, _004614_, _004615_, _004616_, _004617_, _004618_, _004619_, _004620_, _004621_, _004622_, _004623_, _004624_, _004625_, _004626_, _004627_, _004628_, _004629_, _004630_, _004631_, _004632_, _004633_, _004634_, _004635_, _004636_, _004637_, _004638_, _004639_, _004640_, _004641_, _004642_, _004643_, _004644_, _004645_, _004646_, _004647_, _004648_, _004649_, _004650_, _004651_, _004652_, _004653_, _004654_, _004655_, _004656_, _004657_, _004658_, _004659_, _004660_, _004661_, _004662_, _004663_, _004664_, _004665_, _004666_, _004667_, _004668_, _004669_, _004670_, _004671_, _004672_, _004673_, _004674_, _004675_, _004676_, _004677_, _004678_, _004679_, _004680_, _004681_, _004682_, _004683_, _004684_, _004685_, _004686_, _004687_, _004688_, _004689_, _004690_, _004691_, _004692_, _004693_, _004694_, _004695_, _004696_, _004697_, _004698_, _004699_, _004700_, _004701_, _004702_, _004703_, _004704_, _004705_, _004706_, _004707_, _004708_, _004709_, _004710_, _004711_, _004712_, _004713_, _004714_, _004715_, _004716_, _004717_, _004718_, _004719_, _004720_, _004721_, _004722_, _004723_, _004724_, _004725_, _004726_, _004727_, _004728_, _004729_, _004730_, _004731_, _004732_, _004733_, _004734_, _004735_, _004736_, _004737_, _004738_, _004739_, _004740_, _004741_, _004742_, _004743_, _004744_, _004745_, _004746_, _004747_, _004748_, _004749_, _004750_, _004751_, _004752_, _004753_, _004754_, _004755_, _004756_, _004757_, _004758_, _004759_, _004760_, _004761_, _004762_, _004763_, _004764_, _004765_, _004766_, _004767_, _004768_, _004769_, _004770_, _004771_, _004772_, _004773_, _004774_, _004775_, _004776_, _004777_, _004778_, _004779_, _004780_, _004781_, _004782_, _004783_, _004784_, _004785_, _004786_, _004787_, _004788_, _004789_, _004790_, _004791_, _004792_, _004793_, _004794_, _004795_, _004796_, _004797_, _004798_, _004799_, _004800_, _004801_, _004802_, _004803_, _004804_, _004805_, _004806_, _004807_, _004808_, _004809_, _004810_, _004811_, _004812_, _004813_, _004814_, _004815_, _004816_, _004817_, _004818_, _004819_, _004820_, _004821_, _004822_, _004823_, _004824_, _004825_, _004826_, _004827_, _004828_, _004829_, _004830_, _004831_, _004832_, _004833_, _004834_, _004835_, _004836_, _004837_, _004838_, _004839_, _004840_, _004841_, _004842_, _004843_, _004844_, _004845_, _004846_, _004847_, _004848_, _004849_, _004850_, _004851_, _004852_, _004853_, _004854_, _004855_, _004856_, _004857_, _004858_, _004859_, _004860_, _004861_, _004862_, _004863_, _004864_, _004865_, _004866_, _004867_, _004868_, _004869_, _004870_, _004871_, _004872_, _004873_, _004874_, _004875_, _004876_, _004877_, _004878_, _004879_, _004880_, _004881_, _004882_, _004883_, _004884_, _004885_, _004886_, _004887_, _004888_, _004889_, _004890_, _004891_, _004892_, _004893_, _004894_, _004895_, _004896_, _004897_, _004898_, _004899_, _004900_, _004901_, _004902_, _004903_, _004904_, _004905_, _004906_, _004907_, _004908_, _004909_, _004910_, _004911_, _004912_, _004913_, _004914_, _004915_, _004916_, _004917_, _004918_, _004919_, _004920_, _004921_, _004922_, _004923_, _004924_, _004925_, _004926_, _004927_, _004928_, _004929_, _004930_, _004931_, _004932_, _004933_, _004934_, _004935_, _004936_, _004937_, _004938_, _004939_, _004940_, _004941_, _004942_, _004943_, _004944_, _004945_, _004946_, _004947_, _004948_, _004949_, _004950_, _004951_, _004952_, _004953_, _004954_, _004955_, _004956_, _004957_, _004958_, _004959_, _004960_, _004961_, _004962_, _004963_, _004964_, _004965_, _004966_, _004967_, _004968_, _004969_, _004970_, _004971_, _004972_, _004973_, _004974_, _004975_, _004976_, _004977_, _004978_, _004979_, _004980_, _004981_, _004982_, _004983_, _004984_, _004985_, _004986_, _004987_, _004988_, _004989_, _004990_, _004991_, _004992_, _004993_, _004994_, _004995_, _004996_, _004997_, _004998_, _004999_, _005000_, _005001_, _005002_, _005003_, _005004_, _005005_, _005006_, _005007_, _005008_, _005009_, _005010_, _005011_, _005012_, _005013_, _005014_, _005015_, _005016_, _005017_, _005018_, _005019_, _005020_, _005021_, _005022_, _005023_, _005024_, _005025_, _005026_, _005027_, _005028_, _005029_, _005030_, _005031_, _005032_, _005033_, _005034_, _005035_, _005036_, _005037_, _005038_, _005039_, _005040_, _005041_, _005042_, _005043_, _005044_, _005045_, _005046_, _005047_, _005048_, _005049_, _005050_, _005051_, _005052_, _005053_, _005054_, _005055_, _005056_, _005057_, _005058_, _005059_, _005060_, _005061_, _005062_, _005063_, _005064_, _005065_, _005066_, _005067_, _005068_, _005069_, _005070_, _005071_, _005072_, _005073_, _005074_, _005075_, _005076_, _005077_, _005078_, _005079_, _005080_, _005081_, _005082_, _005083_, _005084_, _005085_, _005086_, _005087_, _005088_, _005089_, _005090_, _005091_, _005092_, _005093_, _005094_, _005095_, _005096_, _005097_, _005098_, _005099_, _005100_, _005101_, _005102_, _005103_, _005104_, _005105_, _005106_, _005107_, _005108_, _005109_, _005110_, _005111_, _005112_, _005113_, _005114_, _005115_, _005116_, _005117_, _005118_, _005119_, _005120_, _005121_, _005122_, _005123_, _005124_, _005125_, _005126_, _005127_, _005128_, _005129_, _005130_, _005131_, _005132_, _005133_, _005134_, _005135_, _005136_, _005137_, _005138_, _005139_, _005140_, _005141_, _005142_, _005143_, _005144_, _005145_, _005146_, _005147_, _005148_, _005149_, _005150_, _005151_, _005152_, _005153_, _005154_, _005155_, _005156_, _005157_, _005158_, _005159_, _005160_, _005161_, _005162_, _005163_, _005164_, _005165_, _005166_, _005167_, _005168_, _005169_, _005170_, _005171_, _005172_, _005173_, _005174_, _005175_, _005176_, _005177_, _005178_, _005179_, _005180_, _005181_, _005182_, _005183_, _005184_, _005185_, _005186_, _005187_, _005188_, _005189_, _005190_, _005191_, _005192_, _005193_, _005194_, _005195_, _005196_, _005197_, _005198_, _005199_, _005200_, _005201_, _005202_, _005203_, _005204_, _005205_, _005206_, _005207_, _005208_, _005209_, _005210_, _005211_, _005212_, _005213_, _005214_, _005215_, _005216_, _005217_, _005218_, _005219_, _005220_, _005221_, _005222_, _005223_, _005224_, _005225_, _005226_, _005227_, _005228_, _005229_, _005230_, _005231_, _005232_, _005233_, _005234_, _005235_, _005236_, _005237_, _005238_, _005239_, _005240_, _005241_, _005242_, _005243_, _005244_, _005245_, _005246_, _005247_, _005248_, _005249_, _005250_, _005251_, _005252_, _005253_, _005254_, _005255_, _005256_, _005257_, _005258_, _005259_, _005260_, _005261_, _005262_, _005263_, _005264_, _005265_, _005266_, _005267_, _005268_, _005269_, _005270_, _005271_, _005272_, _005273_, _005274_, _005275_, _005276_, _005277_, _005278_, _005279_, _005280_, _005281_, _005282_, _005283_, _005284_, _005285_, _005286_, _005287_, _005288_, _005289_, _005290_, _005291_, _005292_, _005293_, _005294_, _005295_, _005296_, _005297_, _005298_, _005299_, _005300_, _005301_, _005302_, _005303_, _005304_, _005305_, _005306_, _005307_, _005308_, _005309_, _005310_, _005311_, _005312_, _005313_, _005314_, _005315_, _005316_, _005317_, _005318_, _005319_, _005320_, _005321_, _005322_, _005323_, _005324_, _005325_, _005326_, _005327_, _005328_, _005329_, _005330_, _005331_, _005332_, _005333_, _005334_, _005335_, _005336_, _005337_, _005338_, _005339_, _005340_, _005341_, _005342_, _005343_, _005344_, _005345_, _005346_, _005347_, _005348_, _005349_, _005350_, _005351_, _005352_, _005353_, _005354_, _005355_, _005356_, _005357_, _005358_, _005359_, _005360_, _005361_, _005362_, _005363_, _005364_, _005365_, _005366_, _005367_, _005368_, _005369_, _005370_, _005371_, _005372_, _005373_, _005374_, _005375_, _005376_, _005377_, _005378_, _005379_, _005380_, _005381_, _005382_, _005383_, _005384_, _005385_, _005386_, _005387_, _005388_, _005389_, _005390_, _005391_, _005392_, _005393_, _005394_, _005395_, _005396_, _005397_, _005398_, _005399_, _005400_, _005401_, _005402_, _005403_, _005404_, _005405_, _005406_, _005407_, _005408_, _005409_, _005410_, _005411_, _005412_, _005413_, _005414_, _005415_, _005416_, _005417_, _005418_, _005419_, _005420_, _005421_, _005422_, _005423_, _005424_, _005425_, _005426_, _005427_, _005428_, _005429_, _005430_, _005431_, _005432_, _005433_, _005434_, _005435_, _005436_, _005437_, _005438_, _005439_, _005440_, _005441_, _005442_, _005443_, _005444_, _005445_, _005446_, _005447_, _005448_, _005449_, _005450_, _005451_, _005452_, _005453_, _005454_, _005455_, _005456_, _005457_, _005458_, _005459_, _005460_, _005461_, _005462_, _005463_, _005464_, _005465_, _005466_, _005467_, _005468_, _005469_, _005470_, _005471_, _005472_, _005473_, _005474_, _005475_, _005476_, _005477_, _005478_, _005479_, _005480_, _005481_, _005482_, _005483_, _005484_, _005485_, _005486_, _005487_, _005488_, _005489_, _005490_, _005491_, _005492_, _005493_, _005494_, _005495_, _005496_, _005497_, _005498_, _005499_, _005500_, _005501_, _005502_, _005503_, _005504_, _005505_, _005506_, _005507_, _005508_, _005509_, _005510_, _005511_, _005512_, _005513_, _005514_, _005515_, _005516_, _005517_, _005518_, _005519_, _005520_, _005521_, _005522_, _005523_, _005524_, _005525_, _005526_, _005527_, _005528_, _005529_, _005530_, _005531_, _005532_, _005533_, _005534_, _005535_, _005536_, _005537_, _005538_, _005539_, _005540_, _005541_, _005542_, _005543_, _005544_, _005545_, _005546_, _005547_, _005548_, _005549_, _005550_, _005551_, _005552_, _005553_, _005554_, _005555_, _005556_, _005557_, _005558_, _005559_, _005560_, _005561_, _005562_, _005563_, _005564_, _005565_, _005566_, _005567_, _005568_, _005569_, _005570_, _005571_, _005572_, _005573_, _005574_, _005575_, _005576_, _005577_, _005578_, _005579_, _005580_, _005581_, _005582_, _005583_, _005584_, _005585_, _005586_, _005587_, _005588_, _005589_, _005590_, _005591_, _005592_, _005593_, _005594_, _005595_, _005596_, _005597_, _005598_, _005599_, _005600_, _005601_, _005602_, _005603_, _005604_, _005605_, _005606_, _005607_, _005608_, _005609_, _005610_, _005611_, _005612_, _005613_, _005614_, _005615_, _005616_, _005617_, _005618_, _005619_, _005620_, _005621_, _005622_, _005623_, _005624_, _005625_, _005626_, _005627_, _005628_, _005629_, _005630_, _005631_, _005632_, _005633_, _005634_, _005635_, _005636_, _005637_, _005638_, _005639_, _005640_, _005641_, _005642_, _005643_, _005644_, _005645_, _005646_, _005647_, _005648_, _005649_, _005650_, _005651_, _005652_, _005653_, _005654_, _005655_, _005656_, _005657_, _005658_, _005659_, _005660_, _005661_, _005662_, _005663_, _005664_, _005665_, _005666_, _005667_, _005668_, _005669_, _005670_, _005671_, _005672_, _005673_, _005674_, _005675_, _005676_, _005677_, _005678_, _005679_, _005680_, _005681_, _005682_, _005683_, _005684_, _005685_, _005686_, _005687_, _005688_, _005689_, _005690_, _005691_, _005692_, _005693_, _005694_, _005695_, _005696_, _005697_, _005698_, _005699_, _005700_, _005701_, _005702_, _005703_, _005704_, _005705_, _005706_, _005707_, _005708_, _005709_, _005710_, _005711_, _005712_, _005713_, _005714_, _005715_, _005716_, _005717_, _005718_, _005719_, _005720_, _005721_, _005722_, _005723_, _005724_, _005725_, _005726_, _005727_, _005728_, _005729_, _005730_, _005731_, _005732_, _005733_, _005734_, _005735_, _005736_, _005737_, _005738_, _005739_, _005740_, _005741_, _005742_, _005743_, _005744_, _005745_, _005746_, _005747_, _005748_, _005749_, _005750_, _005751_, _005752_, _005753_, _005754_, _005755_, _005756_, _005757_, _005758_, _005759_, _005760_, _005761_, _005762_, _005763_, _005764_, _005765_, _005766_, _005767_, _005768_, _005769_, _005770_, _005771_, _005772_, _005773_, _005774_, _005775_, _005776_, _005777_, _005778_, _005779_, _005780_, _005781_, _005782_, _005783_, _005784_, _005785_, _005786_, _005787_, _005788_, _005789_, _005790_, _005791_, _005792_, _005793_, _005794_, _005795_, _005796_, _005797_, _005798_, _005799_, _005800_, _005801_, _005802_, _005803_, _005804_, _005805_, _005806_, _005807_, _005808_, _005809_, _005810_, _005811_, _005812_, _005813_, _005814_, _005815_, _005816_, _005817_, _005818_, _005819_, _005820_, _005821_, _005822_, _005823_, _005824_, _005825_, _005826_, _005827_, _005828_, _005829_, _005830_, _005831_, _005832_, _005833_, _005834_, _005835_, _005836_, _005837_, _005838_, _005839_, _005840_, _005841_, _005842_, _005843_, _005844_, _005845_, _005846_, _005847_, _005848_, _005849_, _005850_, _005851_, _005852_, _005853_, _005854_, _005855_, _005856_, _005857_, _005858_, _005859_, _005860_, _005861_, _005862_, _005863_, _005864_, _005865_, _005866_, _005867_, _005868_, _005869_, _005870_, _005871_, _005872_, _005873_, _005874_, _005875_, _005876_, _005877_, _005878_, _005879_, _005880_, _005881_, _005882_, _005883_, _005884_, _005885_, _005886_, _005887_, _005888_, _005889_, _005890_, _005891_, _005892_, _005893_, _005894_, _005895_, _005896_, _005897_, _005898_, _005899_, _005900_, _005901_, _005902_, _005903_, _005904_, _005905_, _005906_, _005907_, _005908_, _005909_, _005910_, _005911_, _005912_, _005913_, _005914_, _005915_, _005916_, _005917_, _005918_, _005919_, _005920_, _005921_, _005922_, _005923_, _005924_, _005925_, _005926_, _005927_, _005928_, _005929_, _005930_, _005931_, _005932_, _005933_, _005934_, _005935_, _005936_, _005937_, _005938_, _005939_, _005940_, _005941_, _005942_, _005943_, _005944_, _005945_, _005946_, _005947_, _005948_, _005949_, _005950_, _005951_, _005952_, _005953_, _005954_, _005955_, _005956_, _005957_, _005958_, _005959_, _005960_, _005961_, _005962_, _005963_, _005964_, _005965_, _005966_, _005967_, _005968_, _005969_, _005970_, _005971_, _005972_, _005973_, _005974_, _005975_, _005976_, _005977_, _005978_, _005979_, _005980_, _005981_, _005982_, _005983_, _005984_, _005985_, _005986_, _005987_, _005988_, _005989_, _005990_, _005991_, _005992_, _005993_, _005994_, _005995_, _005996_, _005997_, _005998_, _005999_, _006000_, _006001_, _006002_, _006003_, _006004_, _006005_, _006006_, _006007_, _006008_, _006009_, _006010_, _006011_, _006012_, _006013_, _006014_, _006015_, _006016_, _006017_, _006018_, _006019_, _006020_, _006021_, _006022_, _006023_, _006024_, _006025_, _006026_, _006027_, _006028_, _006029_, _006030_, _006031_, _006032_, _006033_, _006034_, _006035_, _006036_, _006037_, _006038_, _006039_, _006040_, _006041_, _006042_, _006043_, _006044_, _006045_, _006046_, _006047_, _006048_, _006049_, _006050_, _006051_, _006052_, _006053_, _006054_, _006055_, _006056_, _006057_, _006058_, _006059_, _006060_, _006061_, _006062_, _006063_, _006064_, _006065_, _006066_, _006067_, _006068_, _006069_, _006070_, _006071_, _006072_, _006073_, _006074_, _006075_, _006076_, _006077_, _006078_, _006079_, _006080_, _006081_, _006082_, _006083_, _006084_, _006085_, _006086_, _006087_, _006088_, _006089_, _006090_, _006091_, _006092_, _006093_, _006094_, _006095_, _006096_, _006097_, _006098_, _006099_, _006100_, _006101_, _006102_, _006103_, _006104_, _006105_, _006106_, _006107_, _006108_, _006109_, _006110_, _006111_, _006112_, _006113_, _006114_, _006115_, _006116_, _006117_, _006118_, _006119_, _006120_, _006121_, _006122_, _006123_, _006124_, _006125_, _006126_, _006127_, _006128_, _006129_, _006130_, _006131_, _006132_, _006133_, _006134_, _006135_, _006136_, _006137_, _006138_, _006139_, _006140_, _006141_, _006142_, _006143_, _006144_, _006145_, _006146_, _006147_, _006148_, _006149_, _006150_, _006151_, _006152_, _006153_, _006154_, _006155_, _006156_, _006157_, _006158_, _006159_, _006160_, _006161_, _006162_, _006163_, _006164_, _006165_, _006166_, _006167_, _006168_, _006169_, _006170_, _006171_, _006172_, _006173_, _006174_, _006175_, _006176_, _006177_, _006178_, _006179_, _006180_, _006181_, _006182_, _006183_, _006184_, _006185_, _006186_, _006187_, _006188_, _006189_, _006190_, _006191_, _006192_, _006193_, _006194_, _006195_, _006196_, _006197_, _006198_, _006199_, _006200_, _006201_, _006202_, _006203_, _006204_, _006205_, _006206_, _006207_, _006208_, _006209_, _006210_, _006211_, _006212_, _006213_, _006214_, _006215_, _006216_, _006217_, _006218_, _006219_, _006220_, _006221_, _006222_, _006223_, _006224_, _006225_, _006226_, _006227_, _006228_, _006229_, _006230_, _006231_, _006232_, _006233_, _006234_, _006235_, _006236_, _006237_, _006238_, _006239_, _006240_, _006241_, _006242_, _006243_, _006244_, _006245_, _006246_, _006247_, _006248_, _006249_, _006250_, _006251_, _006252_, _006253_, _006254_, _006255_, _006256_, _006257_, _006258_, _006259_, _006260_, _006261_, _006262_, _006263_, _006264_, _006265_, _006266_, _006267_, _006268_, _006269_, _006270_, _006271_, _006272_, _006273_, _006274_, _006275_, _006276_, _006277_, _006278_, _006279_, _006280_, _006281_, _006282_, _006283_, _006284_, _006285_, _006286_, _006287_, _006288_, _006289_, _006290_, _006291_, _006292_, _006293_, _006294_, _006295_, _006296_, _006297_, _006298_, _006299_, _006300_, _006301_, _006302_, _006303_, _006304_, _006305_, _006306_, _006307_, _006308_, _006309_, _006310_, _006311_, _006312_, _006313_, _006314_, _006315_, _006316_, _006317_, _006318_, _006319_, _006320_, _006321_, _006322_, _006323_, _006324_, _006325_, _006326_, _006327_, _006328_, _006329_, _006330_, _006331_, _006332_, _006333_, _006334_, _006335_, _006336_, _006337_, _006338_, _006339_, _006340_, _006341_, _006342_, _006343_, _006344_, _006345_, _006346_, _006347_, _006348_, _006349_, _006350_, _006351_, _006352_, _006353_, _006354_, _006355_, _006356_, _006357_, _006358_, _006359_, _006360_, _006361_, _006362_, _006363_, _006364_, _006365_, _006366_, _006367_, _006368_, _006369_, _006370_, _006371_, _006372_, _006373_, _006374_, _006375_, _006376_, _006377_, _006378_, _006379_, _006380_, _006381_, _006382_, _006383_, _006384_, _006385_, _006386_, _006387_, _006388_, _006389_, _006390_, _006391_, _006392_, _006393_, _006394_, _006395_, _006396_, _006397_, _006398_, _006399_, _006400_, _006401_, _006402_, _006403_, _006404_, _006405_, _006406_, _006407_, _006408_, _006409_, _006410_, _006411_, _006412_, _006413_, _006414_, _006415_, _006416_, _006417_, _006418_, _006419_, _006420_, _006421_, _006422_, _006423_, _006424_, _006425_, _006426_, _006427_, _006428_, _006429_, _006430_, _006431_, _006432_, _006433_, _006434_, _006435_, _006436_, _006437_, _006438_, _006439_, _006440_, _006441_, _006442_, _006443_, _006444_, _006445_, _006446_, _006447_, _006448_, _006449_, _006450_, _006451_, _006452_, _006453_, _006454_, _006455_, _006456_, _006457_, _006458_, _006459_, _006460_, _006461_, _006462_, _006463_, _006464_, _006465_, _006466_, _006467_, _006468_, _006469_, _006470_, _006471_, _006472_, _006473_, _006474_, _006475_, _006476_, _006477_, _006478_, _006479_, _006480_, _006481_, _006482_, _006483_, _006484_, _006485_, _006486_, _006487_, _006488_, _006489_, _006490_, _006491_, _006492_, _006493_, _006494_, _006495_, _006496_, _006497_, _006498_, _006499_, _006500_, _006501_, _006502_, _006503_, _006504_, _006505_, _006506_, _006507_, _006508_, _006509_, _006510_, _006511_, _006512_, _006513_, _006514_, _006515_, _006516_, _006517_, _006518_, _006519_, _006520_, _006521_, _006522_, _006523_, _006524_, _006525_, _006526_, _006527_, _006528_, _006529_, _006530_, _006531_, _006532_, _006533_, _006534_, _006535_, _006536_, _006537_, _006538_, _006539_, _006540_, _006541_, _006542_, _006543_, _006544_, _006545_, _006546_, _006547_, _006548_, _006549_, _006550_, _006551_, _006552_, _006553_, _006554_, _006555_, _006556_, _006557_, _006558_, _006559_, _006560_, _006561_, _006562_, _006563_, _006564_, _006565_, _006566_, _006567_, _006568_, _006569_, _006570_, _006571_, _006572_, _006573_, _006574_, _006575_, _006576_, _006577_, _006578_, _006579_, _006580_, _006581_, _006582_, _006583_, _006584_, _006585_, _006586_, _006587_, _006588_, _006589_, _006590_, _006591_, _006592_, _006593_, _006594_, _006595_, _006596_, _006597_, _006598_, _006599_, _006600_, _006601_, _006602_, _006603_, _006604_, _006605_, _006606_, _006607_, _006608_, _006609_, _006610_, _006611_, _006612_, _006613_, _006614_, _006615_, _006616_, _006617_, _006618_, _006619_, _006620_, _006621_, _006622_, _006623_, _006624_, _006625_, _006626_, _006627_, _006628_, _006629_, _006630_, _006631_, _006632_, _006633_, _006634_, _006635_, _006636_, _006637_, _006638_, _006639_, _006640_, _006641_, _006642_, _006643_, _006644_, _006645_, _006646_, _006647_, _006648_, _006649_, _006650_, _006651_, _006652_, _006653_, _006654_, _006655_, _006656_, _006657_, _006658_, _006659_, _006660_, _006661_, _006662_, _006663_, _006664_, _006665_, _006666_, _006667_, _006668_, _006669_, _006670_, _006671_, _006672_, _006673_, _006674_, _006675_, _006676_, _006677_, _006678_, _006679_, _006680_, _006681_, _006682_, _006683_, _006684_, _006685_, _006686_, _006687_, _006688_, _006689_, _006690_, _006691_, _006692_, _006693_, _006694_, _006695_, _006696_, _006697_, _006698_, _006699_, _006700_, _006701_, _006702_, _006703_, _006704_, _006705_, _006706_, _006707_, _006708_, _006709_, _006710_, _006711_, _006712_, _006713_, _006714_, _006715_, _006716_, _006717_, _006718_, _006719_, _006720_, _006721_, _006722_, _006723_, _006724_, _006725_, _006726_, _006727_, _006728_, _006729_, _006730_, _006731_, _006732_, _006733_, _006734_, _006735_, _006736_, _006737_, _006738_, _006739_, _006740_, _006741_, _006742_, _006743_, _006744_, _006745_, _006746_, _006747_, _006748_, _006749_, _006750_, _006751_, _006752_, _006753_, _006754_, _006755_, _006756_, _006757_, _006758_, _006759_, _006760_, _006761_, _006762_, _006763_, _006764_, _006765_, _006766_, _006767_, _006768_, _006769_, _006770_, _006771_, _006772_, _006773_, _006774_, _006775_, _006776_, _006777_, _006778_, _006779_, _006780_, _006781_, _006782_, _006783_, _006784_, _006785_, _006786_, _006787_, _006788_, _006789_, _006790_, _006791_, _006792_, _006793_, _006794_, _006795_, _006796_, _006797_, _006798_, _006799_, _006800_, _006801_, _006802_, _006803_, _006804_, _006805_, _006806_, _006807_, _006808_, _006809_, _006810_, _006811_, _006812_, _006813_, _006814_, _006815_, _006816_, _006817_, _006818_, _006819_, _006820_, _006821_, _006822_, _006823_, _006824_, _006825_, _006826_, _006827_, _006828_, _006829_, _006830_, _006831_, _006832_, _006833_, _006834_, _006835_, _006836_, _006837_, _006838_, _006839_, _006840_, _006841_, _006842_, _006843_, _006844_, _006845_, _006846_, _006847_, _006848_, _006849_, _006850_, _006851_, _006852_, _006853_, _006854_, _006855_, _006856_, _006857_, _006858_, _006859_, _006860_, _006861_, _006862_, _006863_, _006864_, _006865_, _006866_, _006867_, _006868_, _006869_, _006870_, _006871_, _006872_, _006873_, _006874_, _006875_, _006876_, _006877_, _006878_, _006879_, _006880_, _006881_, _006882_, _006883_, _006884_, _006885_, _006886_, _006887_, _006888_, _006889_, _006890_, _006891_, _006892_, _006893_, _006894_, _006895_, _006896_, _006897_, _006898_, _006899_, _006900_, _006901_, _006902_, _006903_, _006904_, _006905_, _006906_, _006907_, _006908_, _006909_, _006910_, _006911_, _006912_, _006913_, _006914_, _006915_, _006916_, _006917_, _006918_, _006919_, _006920_, _006921_, _006922_, _006923_, _006924_, _006925_, _006926_, _006927_, _006928_, _006929_, _006930_, _006931_, _006932_, _006933_, _006934_, _006935_, _006936_, _006937_, _006938_, _006939_, _006940_, _006941_, _006942_, _006943_, _006944_, _006945_, _006946_, _006947_, _006948_, _006949_, _006950_, _006951_, _006952_, _006953_, _006954_, _006955_, _006956_, _006957_, _006958_, _006959_, _006960_, _006961_, _006962_, _006963_, _006964_, _006965_, _006966_, _006967_, _006968_, _006969_, _006970_, _006971_, _006972_, _006973_, _006974_, _006975_, _006976_, _006977_, _006978_, _006979_, _006980_, _006981_, _006982_, _006983_, _006984_, _006985_, _006986_, _006987_, _006988_, _006989_, _006990_, _006991_, _006992_, _006993_, _006994_, _006995_, _006996_, _006997_, _006998_, _006999_, _007000_, _007001_, _007002_, _007003_, _007004_, _007005_, _007006_, _007007_, _007008_, _007009_, _007010_, _007011_, _007012_, _007013_, _007014_, _007015_, _007016_, _007017_, _007018_, _007019_, _007020_, _007021_, _007022_, _007023_, _007024_, _007025_, _007026_, _007027_, _007028_, _007029_, _007030_, _007031_, _007032_, _007033_, _007034_, _007035_, _007036_, _007037_, _007038_, _007039_, _007040_, _007041_, _007042_, _007043_, _007044_, _007045_, _007046_, _007047_, _007048_, _007049_, _007050_, _007051_, _007052_, _007053_, _007054_, _007055_, _007056_, _007057_, _007058_, _007059_, _007060_, _007061_, _007062_, _007063_, _007064_, _007065_, _007066_, _007067_, _007068_, _007069_, _007070_, _007071_, _007072_, _007073_, _007074_, _007075_, _007076_, _007077_, _007078_, _007079_, _007080_, _007081_, _007082_, _007083_, _007084_, _007085_, _007086_, _007087_, _007088_, _007089_, _007090_, _007091_, _007092_, _007093_, _007094_, _007095_, _007096_, _007097_, _007098_, _007099_, _007100_, _007101_, _007102_, _007103_, _007104_, _007105_, _007106_, _007107_, _007108_, _007109_, _007110_, _007111_, _007112_, _007113_, _007114_, _007115_, _007116_, _007117_, _007118_, _007119_, _007120_, _007121_, _007122_, _007123_, _007124_, _007125_, _007126_, _007127_, _007128_, _007129_, _007130_, _007131_, _007132_, _007133_, _007134_, _007135_, _007136_, _007137_, _007138_, _007139_, _007140_, _007141_, _007142_, _007143_, _007144_, _007145_, _007146_, _007147_, _007148_, _007149_, _007150_, _007151_, _007152_, _007153_, _007154_, _007155_, _007156_, _007157_, _007158_, _007159_, _007160_, _007161_, _007162_, _007163_, _007164_, _007165_, _007166_, _007167_, _007168_, _007169_, _007170_, _007171_, _007172_, _007173_, _007174_, _007175_, _007176_, _007177_, _007178_, _007179_, _007180_, _007181_, _007182_, _007183_, _007184_, _007185_, _007186_, _007187_, _007188_, _007189_, _007190_, _007191_, _007192_, _007193_, _007194_, _007195_, _007196_, _007197_, _007198_, _007199_, _007200_, _007201_, _007202_, _007203_, _007204_, _007205_, _007206_, _007207_, _007208_, _007209_, _007210_, _007211_, _007212_, _007213_, _007214_, _007215_, _007216_, _007217_, _007218_, _007219_, _007220_, _007221_, _007222_, _007223_, _007224_, _007225_, _007226_, _007227_, _007228_, _007229_, _007230_, _007231_, _007232_, _007233_, _007234_, _007235_, _007236_, _007237_, _007238_, _007239_, _007240_, _007241_, _007242_, _007243_, _007244_, _007245_, _007246_, _007247_, _007248_, _007249_, _007250_, _007251_, _007252_, _007253_, _007254_, _007255_, _007256_, _007257_, _007258_, _007259_, _007260_, _007261_, _007262_, _007263_, _007264_, _007265_, _007266_, _007267_, _007268_, _007269_, _007270_, _007271_, _007272_, _007273_, _007274_, _007275_, _007276_, _007277_, _007278_, _007279_, _007280_, _007281_, _007282_, _007283_, _007284_, _007285_, _007286_, _007287_, _007288_, _007289_, _007290_, _007291_, _007292_, _007293_, _007294_, _007295_, _007296_, _007297_, _007298_, _007299_, _007300_, _007301_, _007302_, _007303_, _007304_, _007305_, _007306_, _007307_, _007308_, _007309_, _007310_, _007311_, _007312_, _007313_, _007314_, _007315_, _007316_, _007317_, _007318_, _007319_, _007320_, _007321_, _007322_, _007323_, _007324_, _007325_, _007326_, _007327_, _007328_, _007329_, _007330_, _007331_, _007332_, _007333_, _007334_, _007335_, _007336_, _007337_, _007338_, _007339_, _007340_, _007341_, _007342_, _007343_, _007344_, _007345_, _007346_, _007347_, _007348_, _007349_, _007350_, _007351_, _007352_, _007353_, _007354_, _007355_, _007356_, _007357_, _007358_, _007359_, _007360_, _007361_, _007362_, _007363_, _007364_, _007365_, _007366_, _007367_, _007368_, _007369_, _007370_, _007371_, _007372_, _007373_, _007374_, _007375_, _007376_, _007377_, _007378_, _007379_, _007380_, _007381_, _007382_, _007383_, _007384_, _007385_, _007386_, _007387_, _007388_, _007389_, _007390_, _007391_, _007392_, _007393_, _007394_, _007395_, _007396_, _007397_, _007398_, _007399_, _007400_, _007401_, _007402_, _007403_, _007404_, _007405_, _007406_, _007407_, _007408_, _007409_, _007410_, _007411_, _007412_, _007413_, _007414_, _007415_, _007416_, _007417_, _007418_, _007419_, _007420_, _007421_, _007422_, _007423_, _007424_, _007425_, _007426_, _007427_, _007428_, _007429_, _007430_, _007431_, _007432_, _007433_, _007434_, _007435_, _007436_, _007437_, _007438_, _007439_, _007440_, _007441_, _007442_, _007443_, _007444_, _007445_, _007446_, _007447_, _007448_, _007449_, _007450_, _007451_, _007452_, _007453_, _007454_, _007455_, _007456_, _007457_, _007458_, _007459_, _007460_, _007461_, _007462_, _007463_, _007464_, _007465_, _007466_, _007467_, _007468_, _007469_, _007470_, _007471_, _007472_, _007473_, _007474_, _007475_, _007476_, _007477_, _007478_, _007479_, _007480_, _007481_, _007482_, _007483_, _007484_, _007485_, _007486_, _007487_, _007488_, _007489_, _007490_, _007491_, _007492_, _007493_, _007494_, _007495_, _007496_, _007497_, _007498_, _007499_, _007500_, _007501_, _007502_, _007503_, _007504_, _007505_, _007506_, _007507_, _007508_, _007509_, _007510_, _007511_, _007512_, _007513_, _007514_, _007515_, _007516_, _007517_, _007518_, _007519_, _007520_, _007521_, _007522_, _007523_, _007524_, _007525_, _007526_, _007527_, _007528_, _007529_, _007530_, _007531_, _007532_, _007533_, _007534_, _007535_, _007536_, _007537_, _007538_, _007539_, _007540_, _007541_, _007542_, _007543_, _007544_, _007545_, _007546_, _007547_, _007548_, _007549_, _007550_, _007551_, _007552_, _007553_, _007554_, _007555_, _007556_, _007557_, _007558_, _007559_, _007560_, _007561_, _007562_, _007563_, _007564_, _007565_, _007566_, _007567_, _007568_, _007569_, _007570_, _007571_, _007572_, _007573_, _007574_, _007575_, _007576_, _007577_, _007578_, _007579_, _007580_, _007581_, _007582_, _007583_, _007584_, _007585_, _007586_, _007587_, _007588_, _007589_, _007590_, _007591_, _007592_, _007593_, _007594_, _007595_, _007596_, _007597_, _007598_, _007599_, _007600_, _007601_, _007602_, _007603_, _007604_, _007605_, _007606_, _007607_, _007608_, _007609_, _007610_, _007611_, _007612_, _007613_, _007614_, _007615_, _007616_, _007617_, _007618_, _007619_, _007620_, _007621_, _007622_, _007623_, _007624_, _007625_, _007626_, _007627_, _007628_, _007629_, _007630_, _007631_, _007632_, _007633_, _007634_, _007635_, _007636_, _007637_, _007638_, _007639_, _007640_, _007641_, _007642_, _007643_, _007644_, _007645_, _007646_, _007647_, _007648_, _007649_, _007650_, _007651_, _007652_, _007653_, _007654_, _007655_, _007656_, _007657_, _007658_, _007659_, _007660_, _007661_, _007662_, _007663_, _007664_, _007665_, _007666_, _007667_, _007668_, _007669_, _007670_, _007671_, _007672_, _007673_, _007674_, _007675_, _007676_, _007677_, _007678_, _007679_, _007680_, _007681_, _007682_, _007683_, _007684_, _007685_, _007686_, _007687_, _007688_, _007689_, _007690_, _007691_, _007692_, _007693_, _007694_, _007695_, _007696_, _007697_, _007698_, _007699_, _007700_, _007701_, _007702_, _007703_, _007704_, _007705_, _007706_, _007707_, _007708_, _007709_, _007710_, _007711_, _007712_, _007713_, _007714_, _007715_, _007716_, _007717_, _007718_, _007719_, _007720_, _007721_, _007722_, _007723_, _007724_, _007725_, _007726_, _007727_, _007728_, _007729_, _007730_, _007731_, _007732_, _007733_, _007734_, _007735_, _007736_, _007737_, _007738_, _007739_, _007740_, _007741_, _007742_, _007743_, _007744_, _007745_, _007746_, _007747_, _007748_, _007749_, _007750_, _007751_, _007752_, _007753_, _007754_, _007755_, _007756_, _007757_, _007758_, _007759_, _007760_, _007761_, _007762_, _007763_, _007764_, _007765_, _007766_, _007767_, _007768_, _007769_, _007770_, _007771_, _007772_, _007773_, _007774_, _007775_, _007776_, _007777_, _007778_, _007779_, _007780_, _007781_, _007782_, _007783_, _007784_, _007785_, _007786_, _007787_, _007788_, _007789_, _007790_, _007791_, _007792_, _007793_, _007794_, _007795_, _007796_, _007797_, _007798_, _007799_, _007800_, _007801_, _007802_, _007803_, _007804_, _007805_, _007806_, _007807_, _007808_, _007809_, _007810_, _007811_, _007812_, _007813_, _007814_, _007815_, _007816_, _007817_, _007818_, _007819_, _007820_, _007821_, _007822_, _007823_, _007824_, _007825_, _007826_, _007827_, _007828_, _007829_, _007830_, _007831_, _007832_, _007833_, _007834_, _007835_, _007836_, _007837_, _007838_, _007839_, _007840_, _007841_, _007842_, _007843_, _007844_, _007845_, _007846_, _007847_, _007848_, _007849_, _007850_, _007851_, _007852_, _007853_, _007854_, _007855_, _007856_, _007857_, _007858_, _007859_, _007860_, _007861_, _007862_, _007863_, _007864_, _007865_, _007866_, _007867_, _007868_, _007869_, _007870_, _007871_, _007872_, _007873_, _007874_, _007875_, _007876_, _007877_, _007878_, _007879_, _007880_, _007881_, _007882_, _007883_, _007884_, _007885_, _007886_, _007887_, _007888_, _007889_, _007890_, _007891_, _007892_, _007893_, _007894_, _007895_, _007896_, _007897_, _007898_, _007899_, _007900_, _007901_, _007902_, _007903_, _007904_, _007905_, _007906_, _007907_, _007908_, _007909_, _007910_, _007911_, _007912_, _007913_, _007914_, _007915_, _007916_, _007917_, _007918_, _007919_, _007920_, _007921_, _007922_, _007923_, _007924_, _007925_, _007926_, _007927_, _007928_, _007929_, _007930_, _007931_, _007932_, _007933_, _007934_, _007935_, _007936_, _007937_, _007938_, _007939_, _007940_, _007941_, _007942_, _007943_, _007944_, _007945_, _007946_, _007947_, _007948_, _007949_, _007950_, _007951_, _007952_, _007953_, _007954_, _007955_, _007956_, _007957_, _007958_, _007959_, _007960_, _007961_, _007962_, _007963_, _007964_, _007965_, _007966_, _007967_, _007968_, _007969_, _007970_, _007971_, _007972_, _007973_, _007974_, _007975_, _007976_, _007977_, _007978_, _007979_, _007980_, _007981_, _007982_, _007983_, _007984_, _007985_, _007986_, _007987_, _007988_, _007989_, _007990_, _007991_, _007992_, _007993_, _007994_, _007995_, _007996_, _007997_, _007998_, _007999_, _008000_, _008001_, _008002_, _008003_, _008004_, _008005_, _008006_, _008007_, _008008_, _008009_, _008010_, _008011_, _008012_, _008013_, _008014_, _008015_, _008016_, _008017_, _008018_, _008019_, _008020_, _008021_, _008022_, _008023_, _008024_, _008025_, _008026_, _008027_, _008028_, _008029_, _008030_, _008031_, _008032_, _008033_, _008034_, _008035_, _008036_, _008037_, _008038_, _008039_, _008040_, _008041_, _008042_, _008043_, _008044_, _008045_, _008046_, _008047_, _008048_, _008049_, _008050_, _008051_, _008052_, _008053_, _008054_, _008055_, _008056_, _008057_, _008058_, _008059_, _008060_, _008061_, _008062_, _008063_, _008064_, _008065_, _008066_, _008067_, _008068_, _008069_, _008070_, _008071_, _008072_, _008073_, _008074_, _008075_, _008076_, _008077_, _008078_, _008079_, _008080_, _008081_, _008082_, _008083_, _008084_, _008085_, _008086_, _008087_, _008088_, _008089_, _008090_, _008091_, _008092_, _008093_, _008094_, _008095_, _008096_, _008097_, _008098_, _008099_, _008100_, _008101_, _008102_, _008103_, _008104_, _008105_, _008106_, _008107_, _008108_, _008109_, _008110_, _008111_, _008112_, _008113_, _008114_, _008115_, _008116_, _008117_, _008118_, _008119_, _008120_, _008121_, _008122_, _008123_, _008124_, _008125_, _008126_, _008127_, _008128_, _008129_, _008130_, _008131_, _008132_, _008133_, _008134_, _008135_, _008136_, _008137_, _008138_, _008139_, _008140_, _008141_, _008142_, _008143_, _008144_, _008145_, _008146_, _008147_, _008148_, _008149_, _008150_, _008151_, _008152_, _008153_, _008154_, _008155_, _008156_, _008157_, _008158_, _008159_, _008160_, _008161_, _008162_, _008163_, _008164_, _008165_, _008166_, _008167_, _008168_, _008169_, _008170_, _008171_, _008172_, _008173_, _008174_, _008175_, _008176_, _008177_, _008178_, _008179_, _008180_, _008181_, _008182_, _008183_, _008184_, _008185_, _008186_, _008187_, _008188_, _008189_, _008190_, _008191_, _008192_, _008193_, _008194_, _008195_, _008196_, _008197_, _008198_, _008199_, _008200_, _008201_, _008202_, _008203_, _008204_, _008205_, _008206_, _008207_, _008208_, _008209_, _008210_, _008211_, _008212_, _008213_, _008214_, _008215_, _008216_, _008217_, _008218_, _008219_, _008220_, _008221_, _008222_, _008223_, _008224_, _008225_, _008226_, _008227_, _008228_, _008229_, _008230_, _008231_, _008232_, _008233_, _008234_, _008235_, _008236_, _008237_, _008238_, _008239_, _008240_, _008241_, _008242_, _008243_, _008244_, _008245_, _008246_, _008247_, _008248_, _008249_, _008250_, _008251_, _008252_, _008253_, _008254_, _008255_, _008256_, _008257_, _008258_, _008259_, _008260_, _008261_, _008262_, _008263_, _008264_, _008265_, _008266_, _008267_, _008268_, _008269_, _008270_, _008271_, _008272_, _008273_, _008274_, _008275_, _008276_, _008277_, _008278_, _008279_, _008280_, _008281_, _008282_, _008283_, _008284_, _008285_, _008286_, _008287_, _008288_, _008289_, _008290_, _008291_, _008292_, _008293_, _008294_, _008295_, _008296_, _008297_, _008298_, _008299_, _008300_, _008301_, _008302_, _008303_, _008304_, _008305_, _008306_, _008307_, _008308_, _008309_, _008310_, _008311_, _008312_, _008313_, _008314_, _008315_, _008316_, _008317_, _008318_, _008319_, _008320_, _008321_, _008322_, _008323_, _008324_, _008325_, _008326_, _008327_, _008328_, _008329_, _008330_, _008331_, _008332_, _008333_, _008334_, _008335_, _008336_, _008337_, _008338_, _008339_, _008340_, _008341_, _008342_, _008343_, _008344_, _008345_, _008346_, _008347_, _008348_, _008349_, _008350_, _008351_, _008352_, _008353_, _008354_, _008355_, _008356_, _008357_, _008358_, _008359_, _008360_, _008361_, _008362_, _008363_, _008364_, _008365_, _008366_, _008367_, _008368_, _008369_, _008370_, _008371_, _008372_, _008373_, _008374_, _008375_, _008376_, _008377_, _008378_, _008379_, _008380_, _008381_, _008382_, _008383_, _008384_, _008385_, _008386_, _008387_, _008388_, _008389_, _008390_, _008391_, _008392_, _008393_, _008394_, _008395_, _008396_, _008397_, _008398_, _008399_, _008400_, _008401_, _008402_, _008403_, _008404_, _008405_, _008406_, _008407_, _008408_, _008409_, _008410_, _008411_, _008412_, _008413_, _008414_, _008415_, _008416_, _008417_, _008418_, _008419_, _008420_, _008421_, _008422_, _008423_, _008424_, _008425_, _008426_, _008427_, _008428_, _008429_, _008430_, _008431_, _008432_, _008433_, _008434_, _008435_, _008436_, _008437_, _008438_, _008439_, _008440_, _008441_, _008442_, _008443_, _008444_, _008445_, _008446_, _008447_, _008448_, _008449_, _008450_, _008451_, _008452_, _008453_, _008454_, _008455_, _008456_, _008457_, _008458_, _008459_, _008460_, _008461_, _008462_, _008463_, _008464_, _008465_, _008466_, _008467_, _008468_, _008469_, _008470_, _008471_, _008472_, _008473_, _008474_, _008475_, _008476_, _008477_, _008478_, _008479_, _008480_, _008481_, _008482_, _008483_, _008484_, _008485_, _008486_, _008487_, _008488_, _008489_, _008490_, _008491_, _008492_, _008493_, _008494_, _008495_, _008496_, _008497_, _008498_, _008499_, _008500_, _008501_, _008502_, _008503_, _008504_, _008505_, _008506_, _008507_, _008508_, _008509_, _008510_, _008511_, _008512_, _008513_, _008514_, _008515_, _008516_, _008517_, _008518_, _008519_, _008520_, _008521_, _008522_, _008523_, _008524_, _008525_, _008526_, _008527_, _008528_, _008529_, _008530_, _008531_, _008532_, _008533_, _008534_, _008535_, _008536_, _008537_, _008538_, _008539_, _008540_, _008541_, _008542_, _008543_, _008544_, _008545_, _008546_, _008547_, _008548_, _008549_, _008550_, _008551_, _008552_, _008553_, _008554_, _008555_, _008556_, _008557_, _008558_, _008559_, _008560_, _008561_, _008562_, _008563_, _008564_, _008565_, _008566_, _008567_, _008568_, _008569_, _008570_, _008571_, _008572_, _008573_, _008574_, _008575_, _008576_, _008577_, _008578_, _008579_, _008580_, _008581_, _008582_, _008583_, _008584_, _008585_, _008586_, _008587_, _008588_, _008589_, _008590_, _008591_, _008592_, _008593_, _008594_, _008595_, _008596_, _008597_, _008598_, _008599_, _008600_, _008601_, _008602_, _008603_, _008604_, _008605_, _008606_, _008607_, _008608_, _008609_, _008610_, _008611_, _008612_, _008613_, _008614_, _008615_, _008616_, _008617_, _008618_, _008619_, _008620_, _008621_, _008622_, _008623_, _008624_, _008625_, _008626_, _008627_, _008628_, _008629_, _008630_, _008631_, _008632_, _008633_, _008634_, _008635_, _008636_, _008637_, _008638_, _008639_, _008640_, _008641_, _008642_, _008643_, _008644_, _008645_, _008646_, _008647_, _008648_, _008649_, _008650_, _008651_, _008652_, _008653_, _008654_, _008655_, _008656_, _008657_, _008658_, _008659_, _008660_, _008661_, _008662_, _008663_, _008664_, _008665_, _008666_, _008667_, _008668_, _008669_, _008670_, _008671_, _008672_, _008673_, _008674_, _008675_, _008676_, _008677_, _008678_, _008679_, _008680_, _008681_, _008682_, _008683_, _008684_, _008685_, _008686_, _008687_, _008688_, _008689_, _008690_, _008691_, _008692_, _008693_, _008694_, _008695_, _008696_, _008697_, _008698_, _008699_, _008700_, _008701_, _008702_, _008703_, _008704_, _008705_, _008706_, _008707_, _008708_, _008709_, _008710_, _008711_, _008712_, _008713_, _008714_, _008715_, _008716_, _008717_, _008718_, _008719_, _008720_, _008721_, _008722_, _008723_, _008724_, _008725_, _008726_, _008727_, _008728_, _008729_, _008730_, _008731_, _008732_, _008733_, _008734_, _008735_, _008736_, _008737_, _008738_, _008739_, _008740_, _008741_, _008742_, _008743_, _008744_, _008745_, _008746_, _008747_, _008748_, _008749_, _008750_, _008751_, _008752_, _008753_, _008754_, _008755_, _008756_, _008757_, _008758_, _008759_, _008760_, _008761_, _008762_, _008763_, _008764_, _008765_, _008766_, _008767_, _008768_, _008769_, _008770_, _008771_, _008772_, _008773_, _008774_, _008775_, _008776_, _008777_, _008778_, _008779_, _008780_, _008781_, _008782_, _008783_, _008784_, _008785_, _008786_, _008787_, _008788_, _008789_, _008790_, _008791_, _008792_, _008793_, _008794_, _008795_, _008796_, _008797_, _008798_, _008799_, _008800_, _008801_, _008802_, _008803_, _008804_, _008805_, _008806_, _008807_, _008808_, _008809_, _008810_, _008811_, _008812_, _008813_, _008814_, _008815_, _008816_, _008817_, _008818_, _008819_, _008820_, _008821_, _008822_, _008823_, _008824_, _008825_, _008826_, _008827_, _008828_, _008829_, _008830_, _008831_, _008832_, _008833_, _008834_, _008835_, _008836_, _008837_, _008838_, _008839_, _008840_, _008841_, _008842_, _008843_, _008844_, _008845_, _008846_, _008847_, _008848_, _008849_, _008850_, _008851_, _008852_, _008853_, _008854_, _008855_, _008856_, _008857_, _008858_, _008859_, _008860_, _008861_, _008862_, _008863_, _008864_, _008865_, _008866_, _008867_, _008868_, _008869_, _008870_, _008871_, _008872_, _008873_, _008874_, _008875_, _008876_, _008877_, _008878_, _008879_, _008880_, _008881_, _008882_, _008883_, _008884_, _008885_, _008886_, _008887_, _008888_, _008889_, _008890_, _008891_, _008892_, _008893_, _008894_, _008895_, _008896_, _008897_, _008898_, _008899_, _008900_, _008901_, _008902_, _008903_, _008904_, _008905_, _008906_, _008907_, _008908_, _008909_, _008910_, _008911_, _008912_, _008913_, _008914_, _008915_, _008916_, _008917_, _008918_, _008919_, _008920_, _008921_, _008922_, _008923_, _008924_, _008925_, _008926_, _008927_, _008928_, _008929_, _008930_, _008931_, _008932_, _008933_, _008934_, _008935_, _008936_, _008937_, _008938_, _008939_, _008940_, _008941_, _008942_, _008943_, _008944_, _008945_, _008946_, _008947_, _008948_, _008949_, _008950_, _008951_, _008952_, _008953_, _008954_, _008955_, _008956_, _008957_, _008958_, _008959_, _008960_, _008961_, _008962_, _008963_, _008964_, _008965_, _008966_, _008967_, _008968_, _008969_, _008970_, _008971_, _008972_, _008973_, _008974_, _008975_, _008976_, _008977_, _008978_, _008979_, _008980_, _008981_, _008982_, _008983_, _008984_, _008985_, _008986_, _008987_, _008988_, _008989_, _008990_, _008991_, _008992_, _008993_, _008994_, _008995_, _008996_, _008997_, _008998_, _008999_, _009000_, _009001_, _009002_, _009003_, _009004_, _009005_, _009006_, _009007_, _009008_, _009009_, _009010_, _009011_, _009012_, _009013_, _009014_, _009015_, _009016_, _009017_, _009018_, _009019_, _009020_, _009021_, _009022_, _009023_, _009024_, _009025_, _009026_, _009027_, _009028_, _009029_, _009030_, _009031_, _009032_, _009033_, _009034_, _009035_, _009036_, _009037_, _009038_, _009039_, _009040_, _009041_, _009042_, _009043_, _009044_, _009045_, _009046_, _009047_, _009048_, _009049_, _009050_, _009051_, _009052_, _009053_, _009054_, _009055_, _009056_, _009057_, _009058_, _009059_, _009060_, _009061_, _009062_, _009063_, _009064_, _009065_, _009066_, _009067_, _009068_, _009069_, _009070_, _009071_, _009072_, _009073_, _009074_, _009075_, _009076_, _009077_, _009078_, _009079_, _009080_, _009081_, _009082_, _009083_, _009084_, _009085_, _009086_, _009087_, _009088_, _009089_, _009090_, _009091_, _009092_, _009093_, _009094_, _009095_, _009096_, _009097_, _009098_, _009099_, _009100_, _009101_, _009102_, _009103_, _009104_, _009105_, _009106_, _009107_, _009108_, _009109_, _009110_, _009111_, _009112_, _009113_, _009114_, _009115_, _009116_, _009117_, _009118_, _009119_, _009120_, _009121_, _009122_, _009123_, _009124_, _009125_, _009126_, _009127_, _009128_, _009129_, _009130_, _009131_, _009132_, _009133_, _009134_, _009135_, _009136_, _009137_, _009138_, _009139_, _009140_, _009141_, _009142_, _009143_, _009144_, _009145_, _009146_, _009147_, _009148_, _009149_, _009150_, _009151_, _009152_, _009153_, _009154_, _009155_, _009156_, _009157_, _009158_, _009159_, _009160_, _009161_, _009162_, _009163_, _009164_, _009165_, _009166_, _009167_, _009168_, _009169_, _009170_, _009171_, _009172_, _009173_, _009174_, _009175_, _009176_, _009177_, _009178_, _009179_, _009180_, _009181_, _009182_, _009183_, _009184_, _009185_, _009186_, _009187_, _009188_, _009189_, _009190_, _009191_, _009192_, _009193_, _009194_, _009195_, _009196_, _009197_, _009198_, _009199_, _009200_, _009201_, _009202_, _009203_, _009204_, _009205_, _009206_, _009207_, _009208_, _009209_, _009210_, _009211_, _009212_, _009213_, _009214_, _009215_, _009216_, _009217_, _009218_, _009219_, _009220_, _009221_, _009222_, _009223_, _009224_, _009225_, _009226_, _009227_, _009228_, _009229_, _009230_, _009231_, _009232_, _009233_, _009234_, _009235_, _009236_, _009237_, _009238_, _009239_, _009240_, _009241_, _009242_, _009243_, _009244_, _009245_, _009246_, _009247_, _009248_, _009249_, _009250_, _009251_, _009252_, _009253_, _009254_, _009255_, _009256_, _009257_, _009258_, _009259_, _009260_, _009261_, _009262_, _009263_, _009264_, _009265_, _009266_, _009267_, _009268_, _009269_, _009270_, _009271_, _009272_, _009273_, _009274_, _009275_, _009276_, _009277_, _009278_, _009279_, _009280_, _009281_, _009282_, _009283_, _009284_, _009285_, _009286_, _009287_, _009288_, _009289_, _009290_, _009291_, _009292_, _009293_, _009294_, _009295_, _009296_, _009297_, _009298_, _009299_, _009300_, _009301_, _009302_, _009303_, _009304_, _009305_, _009306_, _009307_, _009308_, _009309_, _009310_, _009311_, _009312_, _009313_, _009314_, _009315_, _009316_, _009317_, _009318_, _009319_, _009320_, _009321_, _009322_, _009323_, _009324_, _009325_, _009326_, _009327_, _009328_, _009329_, _009330_, _009331_, _009332_, _009333_, _009334_, _009335_, _009336_, _009337_, _009338_, _009339_, _009340_, _009341_, _009342_, _009343_, _009344_, _009345_, _009346_, _009347_, _009348_, _009349_, _009350_, _009351_, _009352_, _009353_, _009354_, _009355_, _009356_, _009357_, _009358_, _009359_, _009360_, _009361_, _009362_, _009363_, _009364_, _009365_, _009366_, _009367_, _009368_, _009369_, _009370_, _009371_, _009372_, _009373_, _009374_, _009375_, _009376_, _009377_, _009378_, _009379_, _009380_, _009381_, _009382_, _009383_, _009384_, _009385_, _009386_, _009387_, _009388_, _009389_, _009390_, _009391_, _009392_, _009393_, _009394_, _009395_, _009396_, _009397_, _009398_, _009399_, _009400_, _009401_, _009402_, _009403_, _009404_, _009405_, _009406_, _009407_, _009408_, _009409_, _009410_, _009411_, _009412_, _009413_, _009414_, _009415_, _009416_, _009417_, _009418_, _009419_, _009420_, _009421_, _009422_, _009423_, _009424_, _009425_, _009426_, _009427_, _009428_, _009429_, _009430_, _009431_, _009432_, _009433_, _009434_, _009435_, _009436_, _009437_, _009438_, _009439_, _009440_, _009441_, _009442_, _009443_, _009444_, _009445_, _009446_, _009447_, _009448_, _009449_, _009450_, _009451_, _009452_, _009453_, _009454_, _009455_, _009456_, _009457_, _009458_, _009459_, _009460_, _009461_, _009462_, _009463_, _009464_, _009465_, _009466_, _009467_, _009468_, _009469_, _009470_, _009471_, _009472_, _009473_, _009474_, _009475_, _009476_, _009477_, _009478_, _009479_, _009480_, _009481_, _009482_, _009483_, _009484_, _009485_, _009486_, _009487_, _009488_, _009489_, _009490_, _009491_, _009492_, _009493_, _009494_, _009495_, _009496_, _009497_, _009498_, _009499_, _009500_, _009501_, _009502_, _009503_, _009504_, _009505_, _009506_, _009507_, _009508_, _009509_, _009510_, _009511_, _009512_, _009513_, _009514_, _009515_, _009516_, _009517_, _009518_, _009519_, _009520_, _009521_, _009522_, _009523_, _009524_, _009525_, _009526_, _009527_, _009528_, _009529_, _009530_, _009531_, _009532_, _009533_, _009534_, _009535_, _009536_, _009537_, _009538_, _009539_, _009540_, _009541_, _009542_, _009543_, _009544_, _009545_, _009546_, _009547_, _009548_, _009549_, _009550_, _009551_, _009552_, _009553_, _009554_, _009555_, _009556_, _009557_, _009558_, _009559_, _009560_, _009561_, _009562_, _009563_, _009564_, _009565_, _009566_, _009567_, _009568_, _009569_, _009570_, _009571_, _009572_, _009573_, _009574_, _009575_, _009576_, _009577_, _009578_, _009579_, _009580_, _009581_, _009582_, _009583_, _009584_, _009585_, _009586_, _009587_, _009588_, _009589_, _009590_, _009591_, _009592_, _009593_, _009594_, _009595_, _009596_, _009597_, _009598_, _009599_, _009600_, _009601_, _009602_, _009603_, _009604_, _009605_, _009606_, _009607_, _009608_, _009609_, _009610_, _009611_, _009612_, _009613_, _009614_, _009615_, _009616_, _009617_, _009618_, _009619_, _009620_, _009621_, _009622_, _009623_, _009624_, _009625_, _009626_, _009627_, _009628_, _009629_, _009630_, _009631_, _009632_, _009633_, _009634_, _009635_, _009636_, _009637_, _009638_, _009639_, _009640_, _009641_, _009642_, _009643_, _009644_, _009645_, _009646_, _009647_, _009648_, _009649_, _009650_, _009651_, _009652_, _009653_, _009654_, _009655_, _009656_, _009657_, _009658_, _009659_, _009660_, _009661_, _009662_, _009663_, _009664_, _009665_, _009666_, _009667_, _009668_, _009669_, _009670_, _009671_, _009672_, _009673_, _009674_, _009675_, _009676_, _009677_, _009678_, _009679_, _009680_, _009681_, _009682_, _009683_, _009684_, _009685_, _009686_, _009687_, _009688_, _009689_, _009690_, _009691_, _009692_, _009693_, _009694_, _009695_, _009696_, _009697_, _009698_, _009699_, _009700_, _009701_, _009702_, _009703_, _009704_, _009705_, _009706_, _009707_, _009708_, _009709_, _009710_, _009711_, _009712_, _009713_, _009714_, _009715_, _009716_, _009717_, _009718_, _009719_, _009720_, _009721_, _009722_, _009723_, _009724_, _009725_, _009726_, _009727_, _009728_, _009729_, _009730_, _009731_, _009732_, _009733_, _009734_, _009735_, _009736_, _009737_, _009738_, _009739_, _009740_, _009741_, _009742_, _009743_, _009744_, _009745_, _009746_, _009747_, _009748_, _009749_, _009750_, _009751_, _009752_, _009753_, _009754_, _009755_, _009756_, _009757_, _009758_, _009759_, _009760_, _009761_, _009762_, _009763_, _009764_, _009765_, _009766_, _009767_, _009768_, _009769_, _009770_, _009771_, _009772_, _009773_, _009774_, _009775_, _009776_, _009777_, _009778_, _009779_, _009780_, _009781_, _009782_, _009783_, _009784_, _009785_, _009786_, _009787_, _009788_, _009789_, _009790_, _009791_, _009792_, _009793_, _009794_, _009795_, _009796_, _009797_, _009798_, _009799_, _009800_, _009801_, _009802_, _009803_, _009804_, _009805_, _009806_, _009807_, _009808_, _009809_, _009810_, _009811_, _009812_, _009813_, _009814_, _009815_, _009816_, _009817_, _009818_, _009819_, _009820_, _009821_, _009822_, _009823_, _009824_, _009825_, _009826_, _009827_, _009828_, _009829_, _009830_, _009831_, _009832_, _009833_, _009834_, _009835_, _009836_, _009837_, _009838_, _009839_, _009840_, _009841_, _009842_, _009843_, _009844_, _009845_, _009846_, _009847_, _009848_, _009849_, _009850_, _009851_, _009852_, _009853_, _009854_, _009855_, _009856_, _009857_, _009858_, _009859_, _009860_, _009861_, _009862_, _009863_, _009864_, _009865_, _009866_, _009867_, _009868_, _009869_, _009870_, _009871_, _009872_, _009873_, _009874_, _009875_, _009876_, _009877_, _009878_, _009879_, _009880_, _009881_, _009882_, _009883_, _009884_, _009885_, _009886_, _009887_, _009888_, _009889_, _009890_, _009891_, _009892_, _009893_, _009894_, _009895_, _009896_, _009897_, _009898_, _009899_, _009900_, _009901_, _009902_, _009903_, _009904_, _009905_, _009906_, _009907_, _009908_, _009909_, _009910_, _009911_, _009912_, _009913_, _009914_, _009915_, _009916_, _009917_, _009918_, _009919_, _009920_, _009921_, _009922_, _009923_, _009924_, _009925_, _009926_, _009927_, _009928_, _009929_, _009930_, _009931_, _009932_, _009933_, _009934_, _009935_, _009936_, _009937_, _009938_, _009939_, _009940_, _009941_, _009942_, _009943_, _009944_, _009945_, _009946_, _009947_, _009948_, _009949_, _009950_, _009951_, _009952_, _009953_, _009954_, _009955_, _009956_, _009957_, _009958_, _009959_, _009960_, _009961_, _009962_, _009963_, _009964_, _009965_, _009966_, _009967_, _009968_, _009969_, _009970_, _009971_, _009972_, _009973_, _009974_, _009975_, _009976_, _009977_, _009978_, _009979_, _009980_, _009981_, _009982_, _009983_, _009984_, _009985_, _009986_, _009987_, _009988_, _009989_, _009990_, _009991_, _009992_, _009993_, _009994_, _009995_, _009996_, _009997_, _009998_, _009999_, _010000_, _010001_, _010002_, _010003_, _010004_, _010005_, _010006_, _010007_, _010008_, _010009_, _010010_, _010011_, _010012_, _010013_, _010014_, _010015_, _010016_, _010017_, _010018_, _010019_, _010020_, _010021_, _010022_, _010023_, _010024_, _010025_, _010026_, _010027_, _010028_, _010029_, _010030_, _010031_, _010032_, _010033_, _010034_, _010035_, _010036_, _010037_, _010038_, _010039_, _010040_, _010041_, _010042_, _010043_, _010044_, _010045_, _010046_, _010047_, _010048_, _010049_, _010050_, _010051_, _010052_, _010053_, _010054_, _010055_, _010056_, _010057_, _010058_, _010059_, _010060_, _010061_, _010062_, _010063_, _010064_, _010065_, _010066_, _010067_, _010068_, _010069_, _010070_, _010071_, _010072_, _010073_, _010074_, _010075_, _010076_, _010077_, _010078_, _010079_, _010080_, _010081_, _010082_, _010083_, _010084_, _010085_, _010086_, _010087_, _010088_, _010089_, _010090_, _010091_, _010092_, _010093_, _010094_, _010095_, _010096_, _010097_, _010098_, _010099_, _010100_, _010101_, _010102_, _010103_, _010104_, _010105_, _010106_, _010107_, _010108_, _010109_, _010110_, _010111_, _010112_, _010113_, _010114_, _010115_, _010116_, _010117_, _010118_, _010119_, _010120_, _010121_, _010122_, _010123_, _010124_, _010125_, _010126_, _010127_, _010128_, _010129_, _010130_, _010131_, _010132_, _010133_, _010134_, _010135_, _010136_, _010137_, _010138_, _010139_, _010140_, _010141_, _010142_, _010143_, _010144_, _010145_, _010146_, _010147_, _010148_, _010149_, _010150_, _010151_, _010152_, _010153_, _010154_, _010155_, _010156_, _010157_, _010158_, _010159_, _010160_, _010161_, _010162_, _010163_, _010164_, _010165_, _010166_, _010167_, _010168_, _010169_, _010170_, _010171_, _010172_, _010173_, _010174_, _010175_, _010176_, _010177_, _010178_, _010179_, _010180_, _010181_, _010182_, _010183_, _010184_, _010185_, _010186_, _010187_, _010188_, _010189_, _010190_, _010191_, _010192_, _010193_, _010194_, _010195_, _010196_, _010197_, _010198_, _010199_, _010200_, _010201_, _010202_, _010203_, _010204_, _010205_, _010206_, _010207_, _010208_, _010209_, _010210_, _010211_, _010212_, _010213_, _010214_, _010215_, _010216_, _010217_, _010218_, _010219_, _010220_, _010221_, _010222_, _010223_, _010224_, _010225_, _010226_, _010227_, _010228_, _010229_, _010230_, _010231_, _010232_, _010233_, _010234_, _010235_, _010236_, _010237_, _010238_, _010239_, _010240_, _010241_, _010242_, _010243_, _010244_, _010245_, _010246_, _010247_, _010248_, _010249_, _010250_, _010251_, _010252_, _010253_, _010254_, _010255_, _010256_, _010257_, _010258_, _010259_, _010260_, _010261_, _010262_, _010263_, _010264_, _010265_, _010266_, _010267_, _010268_, _010269_, _010270_, _010271_, _010272_, _010273_, _010274_, _010275_, _010276_, _010277_, _010278_, _010279_, _010280_, _010281_, _010282_, _010283_, _010284_, _010285_, _010286_, _010287_, _010288_, _010289_, _010290_, _010291_, _010292_, _010293_, _010294_, _010295_, _010296_, _010297_, _010298_, _010299_, _010300_, _010301_, _010302_, _010303_, _010304_, _010305_, _010306_, _010307_, _010308_, _010309_, _010310_, _010311_, _010312_, _010313_, _010314_, _010315_, _010316_, _010317_, _010318_, _010319_, _010320_, _010321_, _010322_, _010323_, _010324_, _010325_, _010326_, _010327_, _010328_, _010329_, _010330_, _010331_, _010332_, _010333_, _010334_, _010335_, _010336_, _010337_, _010338_, _010339_, _010340_, _010341_, _010342_, _010343_, _010344_, _010345_, _010346_, _010347_, _010348_, _010349_, _010350_, _010351_, _010352_, _010353_, _010354_, _010355_, _010356_, _010357_, _010358_, _010359_, _010360_, _010361_, _010362_, _010363_, _010364_, _010365_, _010366_, _010367_, _010368_, _010369_, _010370_, _010371_, _010372_, _010373_, _010374_, _010375_, _010376_, _010377_, _010378_, _010379_, _010380_, _010381_, _010382_, _010383_, _010384_, _010385_, _010386_, _010387_, _010388_, _010389_, _010390_, _010391_, _010392_, _010393_, _010394_, _010395_, _010396_, _010397_, _010398_, _010399_, _010400_, _010401_, _010402_, _010403_, _010404_, _010405_, _010406_, _010407_, _010408_, _010409_, _010410_, _010411_, _010412_, _010413_, _010414_, _010415_, _010416_, _010417_, _010418_, _010419_, _010420_, _010421_, _010422_, _010423_, _010424_, _010425_, _010426_, _010427_, _010428_, _010429_, _010430_, _010431_, _010432_, _010433_, _010434_, _010435_, _010436_, _010437_, _010438_, _010439_, _010440_, _010441_, _010442_, _010443_, _010444_, _010445_, _010446_, _010447_, _010448_, _010449_, _010450_, _010451_, _010452_, _010453_, _010454_, _010455_, _010456_, _010457_, _010458_, _010459_, _010460_, _010461_, _010462_, _010463_, _010464_, _010465_, _010466_, _010467_, _010468_, _010469_, _010470_, _010471_, _010472_, _010473_, _010474_, _010475_, _010476_, _010477_, _010478_, _010479_, _010480_, _010481_, _010482_, _010483_, _010484_, _010485_, _010486_, _010487_, _010488_, _010489_, _010490_, _010491_, _010492_, _010493_, _010494_, _010495_, _010496_, _010497_, _010498_, _010499_, _010500_, _010501_, _010502_, _010503_, _010504_, _010505_, _010506_, _010507_, _010508_, _010509_, _010510_, _010511_, _010512_, _010513_, _010514_, _010515_, _010516_, _010517_, _010518_, _010519_, _010520_, _010521_, _010522_, _010523_, _010524_, _010525_, _010526_, _010527_, _010528_, _010529_, _010530_, _010531_, _010532_, _010533_, _010534_, _010535_, _010536_, _010537_, _010538_, _010539_, _010540_, _010541_, _010542_, _010543_, _010544_, _010545_, _010546_, _010547_, _010548_, _010549_, _010550_, _010551_, _010552_, _010553_, _010554_, _010555_, _010556_, _010557_, _010558_, _010559_, _010560_, _010561_, _010562_, _010563_, _010564_, _010565_, _010566_, _010567_, _010568_, _010569_, _010570_, _010571_, _010572_, _010573_, _010574_, _010575_, _010576_, _010577_, _010578_, _010579_, _010580_, _010581_, _010582_, _010583_, _010584_, _010585_, _010586_, _010587_, _010588_, _010589_, _010590_, _010591_, _010592_, _010593_, _010594_, _010595_, _010596_, _010597_, _010598_, _010599_, _010600_, _010601_, _010602_, _010603_, _010604_, _010605_, _010606_, _010607_, _010608_, _010609_, _010610_, _010611_, _010612_, _010613_, _010614_, _010615_, _010616_, _010617_, _010618_, _010619_, _010620_, _010621_, _010622_, _010623_, _010624_, _010625_, _010626_, _010627_, _010628_, _010629_, _010630_, _010631_, _010632_, _010633_, _010634_, _010635_, _010636_, _010637_, _010638_, _010639_, _010640_, _010641_, _010642_, _010643_, _010644_, _010645_, _010646_, _010647_, _010648_, _010649_, _010650_, _010651_, _010652_, _010653_, _010654_, _010655_, _010656_, _010657_, _010658_, _010659_, _010660_, _010661_, _010662_, _010663_, _010664_, _010665_, _010666_, _010667_, _010668_, _010669_, _010670_, _010671_, _010672_, _010673_, _010674_, _010675_, _010676_, _010677_, _010678_, _010679_, _010680_, _010681_, _010682_, _010683_, _010684_, _010685_, _010686_, _010687_, _010688_, _010689_, _010690_, _010691_, _010692_, _010693_, _010694_, _010695_, _010696_, _010697_, _010698_, _010699_, _010700_, _010701_, _010702_, _010703_, _010704_, _010705_, _010706_, _010707_, _010708_, _010709_, _010710_, _010711_, _010712_, _010713_, _010714_, _010715_, _010716_, _010717_, _010718_, _010719_, _010720_, _010721_, _010722_, _010723_, _010724_, _010725_, _010726_, _010727_, _010728_, _010729_, _010730_, _010731_, _010732_, _010733_, _010734_, _010735_, _010736_, _010737_, _010738_, _010739_, _010740_, _010741_, _010742_, _010743_, _010744_, _010745_, _010746_, _010747_, _010748_, _010749_, _010750_, _010751_, _010752_, _010753_, _010754_, _010755_, _010756_, _010757_, _010758_, _010759_, _010760_, _010761_, _010762_, _010763_, _010764_, _010765_, _010766_, _010767_, _010768_, _010769_, _010770_, _010771_, _010772_, _010773_, _010774_, _010775_, _010776_, _010777_, _010778_, _010779_, _010780_, _010781_, _010782_, _010783_, _010784_, _010785_, _010786_, _010787_, _010788_, _010789_, _010790_, _010791_, _010792_, _010793_, _010794_, _010795_, _010796_, _010797_, _010798_, _010799_, _010800_, _010801_, _010802_, _010803_, _010804_, _010805_, _010806_, _010807_, _010808_, _010809_, _010810_, _010811_, _010812_, _010813_, _010814_, _010815_, _010816_, _010817_, _010818_, _010819_, _010820_, _010821_, _010822_, _010823_, _010824_, _010825_, _010826_, _010827_, _010828_, _010829_, _010830_, _010831_, _010832_, _010833_, _010834_, _010835_, _010836_, _010837_, _010838_, _010839_, _010840_, _010841_, _010842_, _010843_, _010844_, _010845_, _010846_, _010847_, _010848_, _010849_, _010850_, _010851_, _010852_, _010853_, _010854_, _010855_, _010856_, _010857_, _010858_, _010859_, _010860_, _010861_, _010862_, _010863_, _010864_, _010865_, _010866_, _010867_, _010868_, _010869_, _010870_, _010871_, _010872_, _010873_, _010874_, _010875_, _010876_, _010877_, _010878_, _010879_, _010880_, _010881_, _010882_, _010883_, _010884_, _010885_, _010886_, _010887_, _010888_, _010889_, _010890_, _010891_, _010892_, _010893_, _010894_, _010895_, _010896_, _010897_, _010898_, _010899_, _010900_, _010901_, _010902_, _010903_, _010904_, _010905_, _010906_, _010907_, _010908_, _010909_, _010910_, _010911_, _010912_, _010913_, _010914_, _010915_, _010916_, _010917_, _010918_, _010919_, _010920_, _010921_, _010922_, _010923_, _010924_, _010925_, _010926_, _010927_, _010928_, _010929_, _010930_, _010931_, _010932_, _010933_, _010934_, _010935_, _010936_, _010937_, _010938_, _010939_, _010940_, _010941_, _010942_, _010943_, _010944_, _010945_, _010946_, _010947_, _010948_, _010949_, _010950_, _010951_, _010952_, _010953_, _010954_, _010955_, _010956_, _010957_, _010958_, _010959_, _010960_, _010961_, _010962_, _010963_, _010964_, _010965_, _010966_, _010967_, _010968_, _010969_, _010970_, _010971_, _010972_, _010973_, _010974_, _010975_, _010976_, _010977_, _010978_, _010979_, _010980_, _010981_, _010982_, _010983_, _010984_, _010985_, _010986_, _010987_, _010988_, _010989_, _010990_, _010991_, _010992_, _010993_, _010994_, _010995_, _010996_, _010997_, _010998_, _010999_, _011000_, _011001_, _011002_, _011003_, _011004_, _011005_, _011006_, _011007_, _011008_, _011009_, _011010_, _011011_, _011012_, _011013_, _011014_, _011015_, _011016_, _011017_, _011018_, _011019_, _011020_, _011021_, _011022_, _011023_, _011024_, _011025_, _011026_, _011027_, _011028_, _011029_, _011030_, _011031_, _011032_, _011033_, _011034_, _011035_, _011036_, _011037_, _011038_, _011039_, _011040_, _011041_, _011042_, _011043_, _011044_, _011045_, _011046_, _011047_, _011048_, _011049_, _011050_, _011051_, _011052_, _011053_, _011054_, _011055_, _011056_, _011057_, _011058_, _011059_, _011060_, _011061_, _011062_, _011063_, _011064_, _011065_, _011066_, _011067_, _011068_, _011069_, _011070_, _011071_, _011072_, _011073_, _011074_, _011075_, _011076_, _011077_, _011078_, _011079_, _011080_, _011081_, _011082_, _011083_, _011084_, _011085_, _011086_, _011087_, _011088_, _011089_, _011090_, _011091_, _011092_, _011093_, _011094_, _011095_, _011096_, _011097_, _011098_, _011099_, _011100_, _011101_, _011102_, _011103_, _011104_, _011105_, _011106_, _011107_, _011108_, _011109_, _011110_, _011111_, _011112_, _011113_, _011114_, _011115_, _011116_, _011117_, _011118_, _011119_, _011120_, _011121_, _011122_, _011123_, _011124_, _011125_, _011126_, _011127_, _011128_, _011129_, _011130_, _011131_, _011132_, _011133_, _011134_, _011135_, _011136_, _011137_, _011138_, _011139_, _011140_, _011141_, _011142_, _011143_, _011144_, _011145_, _011146_, _011147_, _011148_, _011149_, _011150_, _011151_, _011152_, _011153_, _011154_, _011155_, _011156_, _011157_, _011158_, _011159_, _011160_, _011161_, _011162_, _011163_, _011164_, _011165_, _011166_, _011167_, _011168_, _011169_, _011170_, _011171_, _011172_, _011173_, _011174_, _011175_, _011176_, _011177_, _011178_, _011179_, _011180_, _011181_, _011182_, _011183_, _011184_, _011185_, _011186_, _011187_, _011188_, _011189_, _011190_, _011191_, _011192_, _011193_, _011194_, _011195_, _011196_, _011197_, _011198_, _011199_, _011200_, _011201_, _011202_, _011203_, _011204_, _011205_, _011206_, _011207_, _011208_, _011209_, _011210_, _011211_, _011212_, _011213_, _011214_, _011215_, _011216_, _011217_, _011218_, _011219_, _011220_, _011221_, _011222_, _011223_, _011224_, _011225_, _011226_, _011227_, _011228_, _011229_, _011230_, _011231_, _011232_, _011233_, _011234_, _011235_, _011236_, _011237_, _011238_, _011239_, _011240_, _011241_, _011242_, _011243_, _011244_, _011245_, _011246_, _011247_, _011248_, _011249_, _011250_, _011251_, _011252_, _011253_, _011254_, _011255_, _011256_, _011257_, _011258_, _011259_, _011260_, _011261_, _011262_, _011263_, _011264_, _011265_, _011266_, _011267_, _011268_, _011269_, _011270_, _011271_, _011272_, _011273_, _011274_, _011275_, _011276_, _011277_, _011278_, _011279_, _011280_, _011281_, _011282_, _011283_, _011284_, _011285_, _011286_, _011287_, _011288_, _011289_, _011290_, _011291_, _011292_, _011293_, _011294_, _011295_, _011296_, _011297_, _011298_, _011299_, _011300_, _011301_, _011302_, _011303_, _011304_, _011305_, _011306_, _011307_, _011308_, _011309_, _011310_, _011311_, _011312_, _011313_, _011314_, _011315_, _011316_, _011317_, _011318_, _011319_, _011320_, _011321_, _011322_, _011323_, _011324_, _011325_, _011326_, _011327_, _011328_, _011329_, _011330_, _011331_, _011332_, _011333_, _011334_, _011335_, _011336_, _011337_, _011338_, _011339_, _011340_, _011341_, _011342_, _011343_, _011344_, _011345_, _011346_, _011347_, _011348_, _011349_, _011350_, _011351_, _011352_, _011353_, _011354_, _011355_, _011356_, _011357_, _011358_, _011359_, _011360_, _011361_, _011362_, _011363_, _011364_, _011365_, _011366_, _011367_, _011368_, _011369_, _011370_, _011371_, _011372_, _011373_, _011374_, _011375_, _011376_, _011377_, _011378_, _011379_, _011380_, _011381_, _011382_, _011383_, _011384_, _011385_, _011386_, _011387_, _011388_, _011389_, _011390_, _011391_, _011392_, _011393_, _011394_, _011395_, _011396_, _011397_, _011398_, _011399_, _011400_, _011401_, _011402_, _011403_, _011404_, _011405_, _011406_, _011407_, _011408_, _011409_, _011410_, _011411_, _011412_, _011413_, _011414_, _011415_, _011416_, _011417_, _011418_, _011419_, _011420_, _011421_, _011422_, _011423_, _011424_, _011425_, _011426_, _011427_, _011428_, _011429_, _011430_, _011431_, _011432_, _011433_, _011434_, _011435_, _011436_, _011437_, _011438_, _011439_, _011440_, _011441_, _011442_, _011443_, _011444_, _011445_, _011446_, _011447_, _011448_, _011449_, _011450_, _011451_, _011452_, _011453_, _011454_, _011455_, _011456_, _011457_, _011458_, _011459_, _011460_, _011461_, _011462_, _011463_, _011464_, _011465_, _011466_, _011467_, _011468_, _011469_, _011470_, _011471_, _011472_, _011473_, _011474_, _011475_, _011476_, _011477_, _011478_, _011479_, _011480_, _011481_, _011482_, _011483_, _011484_, _011485_, _011486_, _011487_, _011488_, _011489_, _011490_, _011491_, _011492_, _011493_, _011494_, _011495_, _011496_, _011497_, _011498_, _011499_, _011500_, _011501_, _011502_, _011503_, _011504_, _011505_, _011506_, _011507_, _011508_, _011509_, _011510_, _011511_, _011512_, _011513_, _011514_, _011515_, _011516_, _011517_, _011518_, _011519_, _011520_, _011521_, _011522_, _011523_, _011524_, _011525_, _011526_, _011527_, _011528_, _011529_, _011530_, _011531_, _011532_, _011533_, _011534_, _011535_, _011536_, _011537_, _011538_, _011539_, _011540_, _011541_, _011542_, _011543_, _011544_, _011545_, _011546_, _011547_, _011548_, _011549_, _011550_, _011551_, _011552_, _011553_, _011554_, _011555_, _011556_, _011557_, _011558_, _011559_, _011560_, _011561_, _011562_, _011563_, _011564_, _011565_, _011566_, _011567_, _011568_, _011569_, _011570_, _011571_, _011572_, _011573_, _011574_, _011575_, _011576_, _011577_, _011578_, _011579_, _011580_, _011581_, _011582_, _011583_, _011584_, _011585_, _011586_, _011587_, _011588_, _011589_, _011590_, _011591_, _011592_, _011593_, _011594_, _011595_, _011596_, _011597_, _011598_, _011599_, _011600_, _011601_, _011602_, _011603_, _011604_, _011605_, _011606_, _011607_, _011608_, _011609_, _011610_, _011611_, _011612_, _011613_, _011614_, _011615_, _011616_, _011617_, _011618_, _011619_, _011620_, _011621_, _011622_, _011623_, _011624_, _011625_, _011626_, _011627_, _011628_, _011629_, _011630_, _011631_, _011632_, _011633_, _011634_, _011635_, _011636_, _011637_, _011638_, _011639_, _011640_, _011641_, _011642_, _011643_, _011644_, _011645_, _011646_, _011647_, _011648_, _011649_, _011650_, _011651_, _011652_, _011653_, _011654_, _011655_, _011656_, _011657_, _011658_, _011659_, _011660_, _011661_, _011662_, _011663_, _011664_, _011665_, _011666_, _011667_, _011668_, _011669_, _011670_, _011671_, _011672_, _011673_, _011674_, _011675_, _011676_, _011677_, _011678_, _011679_, _011680_, _011681_, _011682_, _011683_, _011684_, _011685_, _011686_, _011687_, _011688_, _011689_, _011690_, _011691_, _011692_, _011693_, _011694_, _011695_, _011696_, _011697_, _011698_, _011699_, _011700_, _011701_, _011702_, _011703_, _011704_, _011705_, _011706_, _011707_, _011708_, _011709_, _011710_, _011711_, _011712_, _011713_, _011714_, _011715_, _011716_, _011717_, _011718_, _011719_, _011720_, _011721_, _011722_, _011723_, _011724_, _011725_, _011726_, _011727_, _011728_, _011729_, _011730_, _011731_, _011732_, _011733_, _011734_, _011735_, _011736_, _011737_, _011738_, _011739_, _011740_, _011741_, _011742_, _011743_, _011744_, _011745_, _011746_, _011747_, _011748_, _011749_, _011750_, _011751_, _011752_, _011753_, _011754_, _011755_, _011756_, _011757_, _011758_, _011759_, _011760_, _011761_, _011762_, _011763_, _011764_, _011765_, _011766_, _011767_, _011768_, _011769_, _011770_, _011771_, _011772_, _011773_, _011774_, _011775_, _011776_, _011777_, _011778_, _011779_, _011780_, _011781_, _011782_, _011783_, _011784_, _011785_, _011786_, _011787_, _011788_, _011789_, _011790_, _011791_, _011792_, _011793_, _011794_, _011795_, _011796_, _011797_, _011798_, _011799_, _011800_, _011801_, _011802_, _011803_, _011804_, _011805_, _011806_, _011807_, _011808_, _011809_, _011810_, _011811_, _011812_, _011813_, _011814_, _011815_, _011816_, _011817_, _011818_, _011819_, _011820_, _011821_, _011822_, _011823_, _011824_, _011825_, _011826_, _011827_, _011828_, _011829_, _011830_, _011831_, _011832_, _011833_, _011834_, _011835_, _011836_, _011837_, _011838_, _011839_, _011840_, _011841_, _011842_, _011843_, _011844_, _011845_, _011846_, _011847_, _011848_, _011849_, _011850_, _011851_, _011852_, _011853_, _011854_, _011855_, _011856_, _011857_, _011858_, _011859_, _011860_, _011861_, _011862_, _011863_, _011864_, _011865_, _011866_, _011867_, _011868_, _011869_, _011870_, _011871_, _011872_, _011873_, _011874_, _011875_, _011876_, _011877_, _011878_, _011879_, _011880_, _011881_, _011882_, _011883_, _011884_, _011885_, _011886_, _011887_, _011888_, _011889_, _011890_, _011891_, _011892_, _011893_, _011894_, _011895_, _011896_, _011897_, _011898_, _011899_, _011900_, _011901_, _011902_, _011903_, _011904_, _011905_, _011906_, _011907_, _011908_, _011909_, _011910_, _011911_, _011912_, _011913_, _011914_, _011915_, _011916_, _011917_, _011918_, _011919_, _011920_, _011921_, _011922_, _011923_, _011924_, _011925_, _011926_, _011927_, _011928_, _011929_, _011930_, _011931_, _011932_, _011933_, _011934_, _011935_, _011936_, _011937_, _011938_, _011939_, _011940_, _011941_, _011942_, _011943_, _011944_, _011945_, _011946_, _011947_, _011948_, _011949_, _011950_, _011951_, _011952_, _011953_, _011954_, _011955_, _011956_, _011957_, _011958_, _011959_, _011960_, _011961_, _011962_, _011963_, _011964_, _011965_, _011966_, _011967_, _011968_, _011969_, _011970_, _011971_, _011972_, _011973_, _011974_, _011975_, _011976_, _011977_, _011978_, _011979_, _011980_, _011981_, _011982_, _011983_, _011984_, _011985_, _011986_, _011987_, _011988_, _011989_, _011990_, _011991_, _011992_, _011993_, _011994_, _011995_, _011996_, _011997_, _011998_, _011999_, _012000_, _012001_, _012002_, _012003_, _012004_, _012005_, _012006_, _012007_, _012008_, _012009_, _012010_, _012011_, _012012_, _012013_, _012014_, _012015_, _012016_, _012017_, _012018_, _012019_, _012020_, _012021_, _012022_, _012023_, _012024_, _012025_, _012026_, _012027_, _012028_, _012029_, _012030_, _012031_, _012032_, _012033_, _012034_, _012035_, _012036_, _012037_, _012038_, _012039_, _012040_, _012041_, _012042_, _012043_, _012044_, _012045_, _012046_, _012047_, _012048_, _012049_, _012050_, _012051_, _012052_, _012053_, _012054_, _012055_, _012056_, _012057_, _012058_, _012059_, _012060_, _012061_, _012062_, _012063_, _012064_, _012065_, _012066_, _012067_, _012068_, _012069_, _012070_, _012071_, _012072_, _012073_, _012074_, _012075_, _012076_, _012077_, _012078_, _012079_, _012080_, _012081_, _012082_, _012083_, _012084_, _012085_, _012086_, _012087_, _012088_, _012089_, _012090_, _012091_, _012092_, _012093_, _012094_, _012095_, _012096_, _012097_, _012098_, _012099_, _012100_, _012101_, _012102_, _012103_, _012104_, _012105_, _012106_, _012107_, _012108_, _012109_, _012110_, _012111_, _012112_, _012113_, _012114_, _012115_, _012116_, _012117_, _012118_, _012119_, _012120_, _012121_, _012122_, _012123_, _012124_, _012125_, _012126_, _012127_, _012128_, _012129_, _012130_, _012131_, _012132_, _012133_, _012134_, _012135_, _012136_, _012137_, _012138_, _012139_, _012140_, _012141_, _012142_, _012143_, _012144_, _012145_, _012146_, _012147_, _012148_, _012149_, _012150_, _012151_, _012152_, _012153_, _012154_, _012155_, _012156_, _012157_, _012158_, _012159_, _012160_, _012161_, _012162_, _012163_, _012164_, _012165_, _012166_, _012167_, _012168_, _012169_, _012170_, _012171_, _012172_, _012173_, _012174_, _012175_, _012176_, _012177_, _012178_, _012179_, _012180_, _012181_, _012182_, _012183_, _012184_, _012185_, _012186_, _012187_, _012188_, _012189_, _012190_, _012191_, _012192_, _012193_, _012194_, _012195_, _012196_, _012197_, _012198_, _012199_, _012200_, _012201_, _012202_, _012203_, _012204_, _012205_, _012206_, _012207_, _012208_, _012209_, _012210_, _012211_, _012212_, _012213_, _012214_, _012215_, _012216_, _012217_, _012218_, _012219_, _012220_, _012221_, _012222_, _012223_, _012224_, _012225_, _012226_, _012227_, _012228_, _012229_, _012230_, _012231_, _012232_, _012233_, _012234_, _012235_, _012236_, _012237_, _012238_, _012239_, _012240_, _012241_, _012242_, _012243_, _012244_, _012245_, _012246_, _012247_, _012248_, _012249_, _012250_, _012251_, _012252_, _012253_, _012254_, _012255_, _012256_, _012257_, _012258_, _012259_, _012260_, _012261_, _012262_, _012263_, _012264_, _012265_, _012266_, _012267_, _012268_, _012269_, _012270_, _012271_, _012272_, _012273_, _012274_, _012275_, _012276_, _012277_, _012278_, _012279_, _012280_, _012281_, _012282_, _012283_, _012284_, _012285_, _012286_, _012287_, _012288_, _012289_, _012290_, _012291_, _012292_, _012293_, _012294_, _012295_, _012296_, _012297_, _012298_, _012299_, _012300_, _012301_, _012302_, _012303_, _012304_, _012305_, _012306_, _012307_, _012308_, _012309_, _012310_, _012311_, _012312_, _012313_, _012314_, _012315_, _012316_, _012317_, _012318_, _012319_, _012320_, _012321_, _012322_, _012323_, _012324_, _012325_, _012326_, _012327_, _012328_, _012329_, _012330_, _012331_, _012332_, _012333_, _012334_, _012335_, _012336_, _012337_, _012338_, _012339_, _012340_, _012341_, _012342_, _012343_, _012344_, _012345_, _012346_, _012347_, _012348_, _012349_, _012350_, _012351_, _012352_, _012353_, _012354_, _012355_, _012356_, _012357_, _012358_, _012359_, _012360_, _012361_, _012362_, _012363_, _012364_, _012365_, _012366_, _012367_, _012368_, _012369_, _012370_, _012371_, _012372_, _012373_, _012374_, _012375_, _012376_, _012377_, _012378_, _012379_, _012380_, _012381_, _012382_, _012383_, _012384_, _012385_, _012386_, _012387_, _012388_, _012389_, _012390_, _012391_, _012392_, _012393_, _012394_, _012395_, _012396_, _012397_, _012398_, _012399_, _012400_, _012401_, _012402_, _012403_, _012404_, _012405_, _012406_, _012407_, _012408_, _012409_, _012410_, _012411_, _012412_, _012413_, _012414_, _012415_, _012416_, _012417_, _012418_, _012419_, _012420_, _012421_, _012422_, _012423_, _012424_, _012425_, _012426_, _012427_, _012428_, _012429_, _012430_, _012431_, _012432_, _012433_, _012434_, _012435_, _012436_, _012437_, _012438_, _012439_, _012440_, _012441_, _012442_, _012443_, _012444_, _012445_, _012446_, _012447_, _012448_, _012449_, _012450_, _012451_, _012452_, _012453_, _012454_, _012455_, _012456_, _012457_, _012458_, _012459_, _012460_, _012461_, _012462_, _012463_, _012464_, _012465_, _012466_, _012467_, _012468_, _012469_, _012470_, _012471_, _012472_, _012473_, _012474_, _012475_, _012476_, _012477_, _012478_, _012479_, _012480_, _012481_, _012482_, _012483_, _012484_, _012485_, _012486_, _012487_, _012488_, _012489_, _012490_, _012491_, _012492_, _012493_, _012494_, _012495_, _012496_, _012497_, _012498_, _012499_, _012500_, _012501_, _012502_, _012503_, _012504_, _012505_, _012506_, _012507_, _012508_, _012509_, _012510_, _012511_, _012512_, _012513_, _012514_, _012515_, _012516_, _012517_, _012518_, _012519_, _012520_, _012521_, _012522_, _012523_, _012524_, _012525_, _012526_, _012527_, _012528_, _012529_, _012530_, _012531_, _012532_, _012533_, _012534_, _012535_, _012536_, _012537_, _012538_, _012539_, _012540_, _012541_, _012542_, _012543_, _012544_, _012545_, _012546_, _012547_, _012548_, _012549_, _012550_, _012551_, _012552_, _012553_, _012554_, _012555_, _012556_, _012557_, _012558_, _012559_, _012560_, _012561_, _012562_, _012563_, _012564_, _012565_, _012566_, _012567_, _012568_, _012569_, _012570_, _012571_, _012572_, _012573_, _012574_, _012575_, _012576_, _012577_, _012578_, _012579_, _012580_, _012581_, _012582_, _012583_, _012584_, _012585_, _012586_, _012587_, _012588_, _012589_, _012590_, _012591_, _012592_, _012593_, _012594_, _012595_, _012596_, _012597_, _012598_, _012599_, _012600_, _012601_, _012602_, _012603_, _012604_, _012605_, _012606_, _012607_, _012608_, _012609_, _012610_, _012611_, _012612_, _012613_, _012614_, _012615_, _012616_, _012617_, _012618_, _012619_, _012620_, _012621_, _012622_, _012623_, _012624_, _012625_, _012626_, _012627_, _012628_, _012629_, _012630_, _012631_, _012632_, _012633_, _012634_, _012635_, _012636_, _012637_, _012638_, _012639_, _012640_, _012641_, _012642_, _012643_, _012644_, _012645_, _012646_, _012647_, _012648_, _012649_, _012650_, _012651_, _012652_, _012653_, _012654_, _012655_, _012656_, _012657_, _012658_, _012659_, _012660_, _012661_, _012662_, _012663_, _012664_, _012665_, _012666_, _012667_, _012668_, _012669_, _012670_, _012671_, _012672_, _012673_, _012674_, _012675_, _012676_, _012677_, _012678_, _012679_, _012680_, _012681_, _012682_, _012683_, _012684_, _012685_, _012686_, _012687_, _012688_, _012689_, _012690_, _012691_, _012692_, _012693_, _012694_, _012695_, _012696_, _012697_, _012698_, _012699_, _012700_, _012701_, _012702_, _012703_, _012704_, _012705_, _012706_, _012707_, _012708_, _012709_, _012710_, _012711_, _012712_, _012713_, _012714_, _012715_, _012716_, _012717_, _012718_, _012719_, _012720_, _012721_, _012722_, _012723_, _012724_, _012725_, _012726_, _012727_, _012728_, _012729_, _012730_, _012731_, _012732_, _012733_, _012734_, _012735_, _012736_, _012737_, _012738_, _012739_, _012740_, _012741_, _012742_, _012743_, _012744_, _012745_, _012746_, _012747_, _012748_, _012749_, _012750_, _012751_, _012752_, _012753_, _012754_, _012755_, _012756_, _012757_, _012758_, _012759_, _012760_, _012761_, _012762_, _012763_, _012764_, _012765_, _012766_, _012767_, _012768_, _012769_, _012770_, _012771_, _012772_, _012773_, _012774_, _012775_, _012776_, _012777_, _012778_, _012779_, _012780_, _012781_, _012782_, _012783_, _012784_, _012785_, _012786_, _012787_, _012788_, _012789_, _012790_, _012791_, _012792_, _012793_, _012794_, _012795_, _012796_, _012797_, _012798_, _012799_, _012800_, _012801_, _012802_, _012803_, _012804_, _012805_, _012806_, _012807_, _012808_, _012809_, _012810_, _012811_, _012812_, _012813_, _012814_, _012815_, _012816_, _012817_, _012818_, _012819_, _012820_, _012821_, _012822_, _012823_, _012824_, _012825_, _012826_, _012827_, _012828_, _012829_, _012830_, _012831_, _012832_, _012833_, _012834_, _012835_, _012836_, _012837_, _012838_, _012839_, _012840_, _012841_, _012842_, _012843_, _012844_, _012845_, _012846_, _012847_, _012848_, _012849_, _012850_, _012851_, _012852_, _012853_, _012854_, _012855_, _012856_, _012857_, _012858_, _012859_, _012860_, _012861_, _012862_, _012863_, _012864_, _012865_, _012866_, _012867_, _012868_, _012869_, _012870_, _012871_, _012872_, _012873_, _012874_, _012875_, _012876_, _012877_, _012878_, _012879_, _012880_, _012881_, _012882_, _012883_, _012884_, _012885_, _012886_, _012887_, _012888_, _012889_, _012890_, _012891_, _012892_, _012893_, _012894_, _012895_, _012896_, _012897_, _012898_, _012899_, _012900_, _012901_, _012902_, _012903_, _012904_, _012905_, _012906_, _012907_, _012908_, _012909_, _012910_, _012911_, _012912_, _012913_, _012914_, _012915_, _012916_, _012917_, _012918_, _012919_, _012920_, _012921_, _012922_, _012923_, _012924_, _012925_, _012926_, _012927_, _012928_, _012929_, _012930_, _012931_, _012932_, _012933_, _012934_, _012935_, _012936_, _012937_, _012938_, _012939_, _012940_, _012941_, _012942_, _012943_, _012944_, _012945_, _012946_, _012947_, _012948_, _012949_, _012950_, _012951_, _012952_, _012953_, _012954_, _012955_, _012956_, _012957_, _012958_, _012959_, _012960_, _012961_, _012962_, _012963_, _012964_, _012965_, _012966_, _012967_, _012968_, _012969_, _012970_, _012971_, _012972_, _012973_, _012974_, _012975_, _012976_, _012977_, _012978_, _012979_, _012980_, _012981_, _012982_, _012983_, _012984_, _012985_, _012986_, _012987_, _012988_, _012989_, _012990_, _012991_, _012992_, _012993_, _012994_, _012995_, _012996_, _012997_, _012998_, _012999_, _013000_, _013001_, _013002_, _013003_, _013004_, _013005_, _013006_, _013007_, _013008_, _013009_, _013010_, _013011_, _013012_, _013013_, _013014_, _013015_, _013016_, _013017_, _013018_, _013019_, _013020_, _013021_, _013022_, _013023_, _013024_, _013025_, _013026_, _013027_, _013028_, _013029_, _013030_, _013031_, _013032_, _013033_, _013034_, _013035_, _013036_, _013037_, _013038_, _013039_, _013040_, _013041_, _013042_, _013043_, _013044_, _013045_, _013046_, _013047_, _013048_, _013049_, _013050_, _013051_, _013052_, _013053_, _013054_, _013055_, _013056_, _013057_, _013058_, _013059_, _013060_, _013061_, _013062_, _013063_, _013064_, _013065_, _013066_, _013067_, _013068_, _013069_, _013070_, _013071_, _013072_, _013073_, _013074_, _013075_, _013076_, _013077_, _013078_, _013079_, _013080_, _013081_, _013082_, _013083_, _013084_, _013085_, _013086_, _013087_, _013088_, _013089_, _013090_, _013091_, _013092_, _013093_, _013094_, _013095_, _013096_, _013097_, _013098_, _013099_, _013100_, _013101_, _013102_, _013103_, _013104_, _013105_, _013106_, _013107_, _013108_, _013109_, _013110_, _013111_, _013112_, _013113_, _013114_, _013115_, _013116_, _013117_, _013118_, _013119_, _013120_, _013121_, _013122_, _013123_, _013124_, _013125_, _013126_, _013127_, _013128_, _013129_, _013130_, _013131_, _013132_, _013133_, _013134_, _013135_, _013136_, _013137_, _013138_, _013139_, _013140_, _013141_, _013142_, _013143_, _013144_, _013145_, _013146_, _013147_, _013148_, _013149_, _013150_, _013151_, _013152_, _013153_, _013154_, _013155_, _013156_, _013157_, _013158_, _013159_, _013160_, _013161_, _013162_, _013163_, _013164_, _013165_, _013166_, _013167_, _013168_, _013169_, _013170_, _013171_, _013172_, _013173_, _013174_, _013175_, _013176_, _013177_, _013178_, _013179_, _013180_, _013181_, _013182_, _013183_, _013184_, _013185_, _013186_, _013187_, _013188_, _013189_, _013190_, _013191_, _013192_, _013193_, _013194_, _013195_, _013196_, _013197_, _013198_, _013199_, _013200_, _013201_, _013202_, _013203_, _013204_, _013205_, _013206_, _013207_, _013208_, _013209_, _013210_, _013211_, _013212_, _013213_, _013214_, _013215_, _013216_, _013217_, _013218_, _013219_, _013220_, _013221_, _013222_, _013223_, _013224_, _013225_, _013226_, _013227_, _013228_, _013229_, _013230_, _013231_, _013232_, _013233_, _013234_, _013235_, _013236_, _013237_, _013238_, _013239_, _013240_, _013241_, _013242_, _013243_, _013244_, _013245_, _013246_, _013247_, _013248_, _013249_, _013250_, _013251_, _013252_, _013253_, _013254_, _013255_, _013256_, _013257_, _013258_, _013259_, _013260_, _013261_, _013262_, _013263_, _013264_, _013265_, _013266_, _013267_, _013268_, _013269_, _013270_, _013271_, _013272_, _013273_, _013274_, _013275_, _013276_, _013277_, _013278_, _013279_, _013280_, _013281_, _013282_, _013283_, _013284_, _013285_, _013286_, _013287_, _013288_, _013289_, _013290_, _013291_, _013292_, _013293_, _013294_, _013295_, _013296_, _013297_, _013298_, _013299_, _013300_, _013301_, _013302_, _013303_, _013304_, _013305_, _013306_, _013307_, _013308_, _013309_, _013310_, _013311_, _013312_, _013313_, _013314_, _013315_, _013316_, _013317_, _013318_, _013319_, _013320_, _013321_, _013322_, _013323_, _013324_, _013325_, _013326_, _013327_, _013328_, _013329_, _013330_, _013331_, _013332_, _013333_, _013334_, _013335_, _013336_, _013337_, _013338_, _013339_, _013340_, _013341_, _013342_, _013343_, _013344_, _013345_, _013346_, _013347_, _013348_, _013349_, _013350_, _013351_, _013352_, _013353_, _013354_, _013355_, _013356_, _013357_, _013358_, _013359_, _013360_, _013361_, _013362_, _013363_, _013364_, _013365_, _013366_, _013367_, _013368_, _013369_, _013370_, _013371_, _013372_, _013373_, _013374_, _013375_, _013376_, _013377_, _013378_, _013379_, _013380_, _013381_, _013382_, _013383_, _013384_, _013385_, _013386_, _013387_, _013388_, _013389_, _013390_, _013391_, _013392_, _013393_, _013394_, _013395_, _013396_, _013397_, _013398_, _013399_, _013400_, _013401_, _013402_, _013403_, _013404_, _013405_, _013406_, _013407_, _013408_, _013409_, _013410_, _013411_, _013412_, _013413_, _013414_, _013415_, _013416_, _013417_, _013418_, _013419_, _013420_, _013421_, _013422_, _013423_, _013424_, _013425_, _013426_, _013427_, _013428_, _013429_, _013430_, _013431_, _013432_, _013433_, _013434_, _013435_, _013436_, _013437_, _013438_, _013439_, _013440_, _013441_, _013442_, _013443_, _013444_, _013445_, _013446_, _013447_, _013448_, _013449_, _013450_, _013451_, _013452_, _013453_, _013454_, _013455_, _013456_, _013457_, _013458_, _013459_, _013460_, _013461_, _013462_, _013463_, _013464_, _013465_, _013466_, _013467_, _013468_, _013469_, _013470_, _013471_, _013472_, _013473_, _013474_, _013475_, _013476_, _013477_, _013478_, _013479_, _013480_, _013481_, _013482_, _013483_, _013484_, _013485_, _013486_, _013487_, _013488_, _013489_, _013490_, _013491_, _013492_, _013493_, _013494_, _013495_, _013496_, _013497_, _013498_, _013499_, _013500_, _013501_, _013502_, _013503_, _013504_, _013505_, _013506_, _013507_, _013508_, _013509_, _013510_, _013511_, _013512_, _013513_, _013514_, _013515_, _013516_, _013517_, _013518_, _013519_, _013520_, _013521_, _013522_, _013523_, _013524_, _013525_, _013526_, _013527_, _013528_, _013529_, _013530_, _013531_, _013532_, _013533_, _013534_, _013535_, _013536_, _013537_, _013538_, _013539_, _013540_, _013541_, _013542_, _013543_, _013544_, _013545_, _013546_, _013547_, _013548_, _013549_, _013550_, _013551_, _013552_, _013553_, _013554_, _013555_, _013556_, _013557_, _013558_, _013559_, _013560_, _013561_, _013562_, _013563_, _013564_, _013565_, _013566_, _013567_, _013568_, _013569_, _013570_, _013571_, _013572_, _013573_, _013574_, _013575_, _013576_, _013577_, _013578_, _013579_, _013580_, _013581_, _013582_, _013583_, _013584_, _013585_, _013586_, _013587_, _013588_, _013589_, _013590_, _013591_, _013592_, _013593_, _013594_, _013595_, _013596_, _013597_, _013598_, _013599_, _013600_, _013601_, _013602_, _013603_, _013604_, _013605_, _013606_, _013607_, _013608_, _013609_, _013610_, _013611_, _013612_, _013613_, _013614_, _013615_, _013616_, _013617_, _013618_, _013619_, _013620_, _013621_, _013622_, _013623_, _013624_, _013625_, _013626_, _013627_, _013628_, _013629_, _013630_, _013631_, _013632_, _013633_, _013634_, _013635_, _013636_, _013637_, _013638_, _013639_, _013640_, _013641_, _013642_, _013643_, _013644_, _013645_, _013646_, _013647_, _013648_, _013649_, _013650_, _013651_, _013652_, _013653_, _013654_, _013655_, _013656_, _013657_, _013658_, _013659_, _013660_, _013661_, _013662_, _013663_, _013664_, _013665_, _013666_, _013667_, _013668_, _013669_, _013670_, _013671_, _013672_, _013673_, _013674_, _013675_, _013676_, _013677_, _013678_, _013679_, _013680_, _013681_, _013682_, _013683_, _013684_, _013685_, _013686_, _013687_, _013688_, _013689_, _013690_, _013691_, _013692_, _013693_, _013694_, _013695_, _013696_, _013697_, _013698_, _013699_, _013700_, _013701_, _013702_, _013703_, _013704_, _013705_, _013706_, _013707_, _013708_, _013709_, _013710_, _013711_, _013712_, _013713_, _013714_, _013715_, _013716_, _013717_, _013718_, _013719_, _013720_, _013721_, _013722_, _013723_, _013724_, _013725_, _013726_, _013727_, _013728_, _013729_, _013730_, _013731_, _013732_, _013733_, _013734_, _013735_, _013736_, _013737_, _013738_, _013739_, _013740_, _013741_, _013742_, _013743_, _013744_, _013745_, _013746_, _013747_, _013748_, _013749_, _013750_, _013751_, _013752_, _013753_, _013754_, _013755_, _013756_, _013757_, _013758_, _013759_, _013760_, _013761_, _013762_, _013763_, _013764_, _013765_, _013766_, _013767_, _013768_, _013769_, _013770_, _013771_, _013772_, _013773_, _013774_, _013775_, _013776_, _013777_, _013778_, _013779_, _013780_, _013781_, _013782_, _013783_, _013784_, _013785_, _013786_, _013787_, _013788_, _013789_, _013790_, _013791_, _013792_, _013793_, _013794_, _013795_, _013796_, _013797_, _013798_, _013799_, _013800_, _013801_, _013802_, _013803_, _013804_, _013805_, _013806_, _013807_, _013808_, _013809_, _013810_, _013811_, _013812_, _013813_, _013814_, _013815_, _013816_, _013817_, _013818_, _013819_, _013820_, _013821_, _013822_, _013823_, _013824_, _013825_, _013826_, _013827_, _013828_, _013829_, _013830_, _013831_, _013832_, _013833_, _013834_, _013835_, _013836_, _013837_, _013838_, _013839_, _013840_, _013841_, _013842_, _013843_, _013844_, _013845_, _013846_, _013847_, _013848_, _013849_, _013850_, _013851_, _013852_, _013853_, _013854_, _013855_, _013856_, _013857_, _013858_, _013859_, _013860_, _013861_, _013862_, _013863_, _013864_, _013865_, _013866_, _013867_, _013868_, _013869_, _013870_, _013871_, _013872_, _013873_, _013874_, _013875_, _013876_, _013877_, _013878_, _013879_, _013880_, _013881_, _013882_, _013883_, _013884_, _013885_, _013886_, _013887_, _013888_, _013889_, _013890_, _013891_, _013892_, _013893_, _013894_, _013895_, _013896_, _013897_, _013898_, _013899_, _013900_, _013901_, _013902_, _013903_, _013904_, _013905_, _013906_, _013907_, _013908_, _013909_, _013910_, _013911_, _013912_, _013913_, _013914_, _013915_, _013916_, _013917_, _013918_, _013919_, _013920_, _013921_, _013922_, _013923_, _013924_, _013925_, _013926_, _013927_, _013928_, _013929_, _013930_, _013931_, _013932_, _013933_, _013934_, _013935_, _013936_, _013937_, _013938_, _013939_, _013940_, _013941_, _013942_, _013943_, _013944_, _013945_, _013946_, _013947_, _013948_, _013949_, _013950_, _013951_, _013952_, _013953_, _013954_, _013955_, _013956_, _013957_, _013958_, _013959_, _013960_, _013961_, _013962_, _013963_, _013964_, _013965_, _013966_, _013967_, _013968_, _013969_, _013970_, _013971_, _013972_, _013973_, _013974_, _013975_, _013976_, _013977_, _013978_, _013979_, _013980_, _013981_, _013982_, _013983_, _013984_, _013985_, _013986_, _013987_, _013988_, _013989_, _013990_, _013991_, _013992_, _013993_, _013994_, _013995_, _013996_, _013997_, _013998_, _013999_, _014000_, _014001_, _014002_, _014003_, _014004_, _014005_, _014006_, _014007_, _014008_, _014009_, _014010_, _014011_, _014012_, _014013_, _014014_, _014015_, _014016_, _014017_, _014018_, _014019_, _014020_, _014021_, _014022_, _014023_, _014024_, _014025_, _014026_, _014027_, _014028_, _014029_, _014030_, _014031_, _014032_, _014033_, _014034_, _014035_, _014036_, _014037_, _014038_, _014039_, _014040_, _014041_, _014042_, _014043_, _014044_, _014045_, _014046_, _014047_, _014048_, _014049_, _014050_, _014051_, _014052_, _014053_, _014054_, _014055_, _014056_, _014057_, _014058_, _014059_, _014060_, _014061_, _014062_, _014063_, _014064_, _014065_, _014066_, _014067_, _014068_, _014069_, _014070_, _014071_, _014072_, _014073_, _014074_, _014075_, _014076_, _014077_, _014078_, _014079_, _014080_, _014081_, _014082_, _014083_, _014084_, _014085_, _014086_, _014087_, _014088_, _014089_, _014090_, _014091_, _014092_, _014093_, _014094_, _014095_, _014096_, _014097_, _014098_, _014099_, _014100_, _014101_, _014102_, _014103_, _014104_, _014105_, _014106_, _014107_, _014108_, _014109_, _014110_, _014111_, _014112_, _014113_, _014114_, _014115_, _014116_, _014117_, _014118_, _014119_, _014120_, _014121_, _014122_, _014123_, _014124_, _014125_, _014126_, _014127_, _014128_, _014129_, _014130_, _014131_, _014132_, _014133_, _014134_, _014135_, _014136_, _014137_, _014138_, _014139_, _014140_, _014141_, _014142_, _014143_, _014144_, _014145_, _014146_, _014147_, _014148_, _014149_, _014150_, _014151_, _014152_, _014153_, _014154_, _014155_, _014156_, _014157_, _014158_, _014159_, _014160_, _014161_, _014162_, _014163_, _014164_, _014165_, _014166_, _014167_, _014168_, _014169_, _014170_, _014171_, _014172_, _014173_, _014174_, _014175_, _014176_, _014177_, _014178_, _014179_, _014180_, _014181_, _014182_, _014183_, _014184_, _014185_, _014186_, _014187_, _014188_, _014189_, _014190_, _014191_, _014192_, _014193_, _014194_, _014195_, _014196_, _014197_, _014198_, _014199_, _014200_, _014201_, _014202_, _014203_, _014204_, _014205_, _014206_, _014207_, _014208_, _014209_, _014210_, _014211_, _014212_, _014213_, _014214_, _014215_, _014216_, _014217_, _014218_, _014219_, _014220_, _014221_, _014222_, _014223_, _014224_, _014225_, _014226_, _014227_, _014228_, _014229_, _014230_, _014231_, _014232_, _014233_, _014234_, _014235_, _014236_, _014237_, _014238_, _014239_, _014240_, _014241_, _014242_, _014243_, _014244_, _014245_, _014246_, _014247_, _014248_, _014249_, _014250_, _014251_, _014252_, _014253_, _014254_, _014255_, _014256_, _014257_, _014258_, _014259_, _014260_, _014261_, _014262_, _014263_, _014264_, _014265_, _014266_, _014267_, _014268_, _014269_, _014270_, _014271_, _014272_, _014273_, _014274_, _014275_, _014276_, _014277_, _014278_, _014279_, _014280_, _014281_, _014282_, _014283_, _014284_, _014285_, _014286_, _014287_, _014288_, _014289_, _014290_, _014291_, _014292_, _014293_, _014294_, _014295_, _014296_, _014297_, _014298_, _014299_, _014300_, _014301_, _014302_, _014303_, _014304_, _014305_, _014306_, _014307_, _014308_, _014309_, _014310_, _014311_, _014312_, _014313_, _014314_, _014315_, _014316_, _014317_, _014318_, _014319_, _014320_, _014321_, _014322_, _014323_, _014324_, _014325_, _014326_, _014327_, _014328_, _014329_, _014330_, _014331_, _014332_, _014333_, _014334_, _014335_, _014336_, _014337_, _014338_, _014339_, _014340_, _014341_, _014342_, _014343_, _014344_, _014345_, _014346_, _014347_, _014348_, _014349_, _014350_, _014351_, _014352_, _014353_, _014354_, _014355_, _014356_, _014357_, _014358_, _014359_, _014360_, _014361_, _014362_, _014363_, _014364_, _014365_, _014366_, _014367_, _014368_, _014369_, _014370_, _014371_, _014372_, _014373_, _014374_, _014375_, _014376_, _014377_, _014378_, _014379_, _014380_, _014381_, _014382_, _014383_, _014384_, _014385_, _014386_, _014387_, _014388_, _014389_, _014390_, _014391_, _014392_, _014393_, _014394_, _014395_, _014396_, _014397_, _014398_, _014399_, _014400_, _014401_, _014402_, _014403_, _014404_, _014405_, _014406_, _014407_, _014408_, _014409_, _014410_, _014411_, _014412_, _014413_, _014414_, _014415_, _014416_, _014417_, _014418_, _014419_, _014420_, _014421_, _014422_, _014423_, _014424_, _014425_, _014426_, _014427_, _014428_, _014429_, _014430_, _014431_, _014432_, _014433_, _014434_, _014435_, _014436_, _014437_, _014438_, _014439_, _014440_, _014441_, _014442_, _014443_, _014444_, _014445_, _014446_, _014447_, _014448_, _014449_, _014450_, _014451_, _014452_, _014453_, _014454_, _014455_, _014456_, _014457_, _014458_, _014459_, _014460_, _014461_, _014462_, _014463_, _014464_, _014465_, _014466_, _014467_, _014468_, _014469_, _014470_, _014471_, _014472_, _014473_, _014474_, _014475_, _014476_, _014477_, _014478_, _014479_, _014480_, _014481_, _014482_, _014483_, _014484_, _014485_, _014486_, _014487_, _014488_, _014489_, _014490_, _014491_, _014492_, _014493_, _014494_, _014495_, _014496_, _014497_, _014498_, _014499_, _014500_, _014501_, _014502_, _014503_, _014504_, _014505_, _014506_, _014507_, _014508_, _014509_, _014510_, _014511_, _014512_, _014513_, _014514_, _014515_, _014516_, _014517_, _014518_, _014519_, _014520_, _014521_, _014522_, _014523_, _014524_, _014525_, _014526_, _014527_, _014528_, _014529_, _014530_, _014531_, _014532_, _014533_, _014534_, _014535_, _014536_, _014537_, _014538_, _014539_, _014540_, _014541_, _014542_, _014543_, _014544_, _014545_, _014546_, _014547_, _014548_, _014549_, _014550_, _014551_, _014552_, _014553_, _014554_, _014555_, _014556_, _014557_, _014558_, _014559_, _014560_, _014561_, _014562_, _014563_, _014564_, _014565_, _014566_, _014567_, _014568_, _014569_, _014570_, _014571_, _014572_, _014573_, _014574_, _014575_, _014576_, _014577_, _014578_, _014579_, _014580_, _014581_, _014582_, _014583_, _014584_, _014585_, _014586_, _014587_, _014588_, _014589_, _014590_, _014591_, _014592_, _014593_, _014594_, _014595_, _014596_, _014597_, _014598_, _014599_, _014600_, _014601_, _014602_, _014603_, _014604_, _014605_, _014606_, _014607_, _014608_, _014609_, _014610_, _014611_, _014612_, _014613_, _014614_, _014615_, _014616_, _014617_, _014618_, _014619_, _014620_, _014621_, _014622_, _014623_, _014624_, _014625_, _014626_, _014627_, _014628_, _014629_, _014630_, _014631_, _014632_, _014633_, _014634_, _014635_, _014636_, _014637_, _014638_, _014639_, _014640_, _014641_, _014642_, _014643_, _014644_, _014645_, _014646_, _014647_, _014648_, _014649_, _014650_, _014651_, _014652_, _014653_, _014654_, _014655_, _014656_, _014657_, _014658_, _014659_, _014660_, _014661_, _014662_, _014663_, _014664_, _014665_, _014666_, _014667_, _014668_, _014669_, _014670_, _014671_, _014672_, _014673_, _014674_, _014675_, _014676_, _014677_, _014678_, _014679_, _014680_, _014681_, _014682_, _014683_, _014684_, _014685_, _014686_, _014687_, _014688_, _014689_, _014690_, _014691_, _014692_, _014693_, _014694_, _014695_, _014696_, _014697_, _014698_, _014699_, _014700_, _014701_, _014702_, _014703_, _014704_, _014705_, _014706_, _014707_, _014708_, _014709_, _014710_, _014711_, _014712_, _014713_, _014714_, _014715_, _014716_, _014717_, _014718_, _014719_, _014720_, _014721_, _014722_, _014723_, _014724_, _014725_, _014726_, _014727_, _014728_, _014729_, _014730_, _014731_, _014732_, _014733_, _014734_, _014735_, _014736_, _014737_, _014738_, _014739_, _014740_, _014741_, _014742_, _014743_, _014744_, _014745_, _014746_, _014747_, _014748_, _014749_, _014750_, _014751_, _014752_, _014753_, _014754_, _014755_, _014756_, _014757_, _014758_, _014759_, _014760_, _014761_, _014762_, _014763_, _014764_, _014765_, _014766_, _014767_, _014768_, _014769_, _014770_, _014771_, _014772_, _014773_, _014774_, _014775_, _014776_, _014777_, _014778_, _014779_, _014780_, _014781_, _014782_, _014783_, _014784_, _014785_, _014786_, _014787_, _014788_, _014789_, _014790_, _014791_, _014792_, _014793_, _014794_, _014795_, _014796_, _014797_, _014798_, _014799_, _014800_, _014801_, _014802_, _014803_, _014804_, _014805_, _014806_, _014807_, _014808_, _014809_, _014810_, _014811_, _014812_, _014813_, _014814_, _014815_, _014816_, _014817_, _014818_, _014819_, _014820_, _014821_, _014822_, _014823_, _014824_, _014825_, _014826_, _014827_, _014828_, _014829_, _014830_, _014831_, _014832_, _014833_, _014834_, _014835_, _014836_, _014837_, _014838_, _014839_, _014840_, _014841_, _014842_, _014843_, _014844_, _014845_, _014846_, _014847_, _014848_, _014849_, _014850_, _014851_, _014852_, _014853_, _014854_, _014855_, _014856_, _014857_, _014858_, _014859_, _014860_, _014861_, _014862_, _014863_, _014864_, _014865_, _014866_, _014867_, _014868_, _014869_, _014870_, _014871_, _014872_, _014873_, _014874_, _014875_, _014876_, _014877_, _014878_, _014879_, _014880_, _014881_, _014882_, _014883_, _014884_, _014885_, _014886_, _014887_, _014888_, _014889_, _014890_, _014891_, _014892_, _014893_, _014894_, _014895_, _014896_, _014897_, _014898_, _014899_, _014900_, _014901_, _014902_, _014903_, _014904_, _014905_, _014906_, _014907_, _014908_, _014909_, _014910_, _014911_, _014912_, _014913_, _014914_, _014915_, _014916_, _014917_, _014918_, _014919_, _014920_, _014921_, _014922_, _014923_, _014924_, _014925_, _014926_, _014927_, _014928_, _014929_, _014930_, _014931_, _014932_, _014933_, _014934_, _014935_, _014936_, _014937_, _014938_, _014939_, _014940_, _014941_, _014942_, _014943_, _014944_, _014945_, _014946_, _014947_, _014948_, _014949_, _014950_, _014951_, _014952_, _014953_, _014954_, _014955_, _014956_, _014957_, _014958_, _014959_, _014960_, _014961_, _014962_, _014963_, _014964_, _014965_, _014966_, _014967_, _014968_, _014969_, _014970_, _014971_, _014972_, _014973_, _014974_, _014975_, _014976_, _014977_, _014978_, _014979_, _014980_, _014981_, _014982_, _014983_, _014984_, _014985_, _014986_, _014987_, _014988_, _014989_, _014990_, _014991_, _014992_, _014993_, _014994_, _014995_, _014996_, _014997_, _014998_, _014999_, _015000_, _015001_, _015002_, _015003_, _015004_, _015005_, _015006_, _015007_, _015008_, _015009_, _015010_, _015011_, _015012_, _015013_, _015014_, _015015_, _015016_, _015017_, _015018_, _015019_, _015020_, _015021_, _015022_, _015023_, _015024_, _015025_, _015026_, _015027_, _015028_, _015029_, _015030_, _015031_, _015032_, _015033_, _015034_, _015035_, _015036_, _015037_, _015038_, _015039_, _015040_, _015041_, _015042_, _015043_, _015044_, _015045_, _015046_, _015047_, _015048_, _015049_, _015050_, _015051_, _015052_, _015053_, _015054_, _015055_, _015056_, _015057_, _015058_, _015059_, _015060_, _015061_, _015062_, _015063_, _015064_, _015065_, _015066_, _015067_, _015068_, _015069_, _015070_, _015071_, _015072_, _015073_, _015074_, _015075_, _015076_, _015077_, _015078_, _015079_, _015080_, _015081_, _015082_, _015083_, _015084_, _015085_, _015086_, _015087_, _015088_, _015089_, _015090_, _015091_, _015092_, _015093_, _015094_, _015095_, _015096_, _015097_, _015098_, _015099_, _015100_, _015101_, _015102_, _015103_, _015104_, _015105_, _015106_, _015107_, _015108_, _015109_, _015110_, _015111_, _015112_, _015113_, _015114_, _015115_, _015116_, _015117_, _015118_, _015119_, _015120_, _015121_, _015122_, _015123_, _015124_, _015125_, _015126_, _015127_, _015128_, _015129_, _015130_, _015131_, _015132_, _015133_, _015134_, _015135_, _015136_, _015137_, _015138_, _015139_, _015140_, _015141_, _015142_, _015143_, _015144_, _015145_, _015146_, _015147_, _015148_, _015149_, _015150_, _015151_, _015152_, _015153_, _015154_, _015155_, _015156_, _015157_, _015158_, _015159_, _015160_, _015161_, _015162_, _015163_, _015164_, _015165_, _015166_, _015167_, _015168_, _015169_, _015170_, _015171_, _015172_, _015173_, _015174_, _015175_, _015176_, _015177_, _015178_, _015179_, _015180_, _015181_, _015182_, _015183_, _015184_, _015185_, _015186_, _015187_, _015188_, _015189_, _015190_, _015191_, _015192_, _015193_, _015194_, _015195_, _015196_, _015197_, _015198_, _015199_, _015200_, _015201_, _015202_, _015203_, _015204_, _015205_, _015206_, _015207_, _015208_, _015209_, _015210_, _015211_, _015212_, _015213_, _015214_, _015215_, _015216_, _015217_, _015218_, _015219_, _015220_, _015221_, _015222_, _015223_, _015224_, _015225_, _015226_, _015227_, _015228_, _015229_, _015230_, _015231_, _015232_, _015233_, _015234_, _015235_, _015236_, _015237_, _015238_, _015239_, _015240_, _015241_, _015242_, _015243_, _015244_, _015245_, _015246_, _015247_, _015248_, _015249_, _015250_, _015251_, _015252_, _015253_, _015254_, _015255_, _015256_, _015257_, _015258_, _015259_, _015260_, _015261_, _015262_, _015263_, _015264_, _015265_, _015266_, _015267_, _015268_, _015269_, _015270_, _015271_, _015272_, _015273_, _015274_, _015275_, _015276_, _015277_, _015278_, _015279_, _015280_, _015281_, _015282_, _015283_, _015284_, _015285_, _015286_, _015287_, _015288_, _015289_, _015290_, _015291_, _015292_, _015293_, _015294_, _015295_, _015296_, _015297_, _015298_, _015299_, _015300_, _015301_, _015302_, _015303_, _015304_, _015305_, _015306_, _015307_, _015308_, _015309_, _015310_, _015311_, _015312_, _015313_, _015314_, _015315_, _015316_, _015317_, _015318_, _015319_, _015320_, _015321_, _015322_, _015323_, _015324_, _015325_, _015326_, _015327_, _015328_, _015329_, _015330_, _015331_, _015332_, _015333_, _015334_, _015335_, _015336_, _015337_, _015338_, _015339_, _015340_, _015341_, _015342_, _015343_, _015344_, _015345_, _015346_, _015347_, _015348_, _015349_, _015350_, _015351_, _015352_, _015353_, _015354_, _015355_, _015356_, _015357_, _015358_, _015359_, _015360_, _015361_, _015362_, _015363_, _015364_, _015365_, _015366_, _015367_, _015368_, _015369_, _015370_, _015371_, _015372_, _015373_, _015374_, _015375_, _015376_, _015377_, _015378_, _015379_, _015380_, _015381_, _015382_, _015383_, _015384_, _015385_, _015386_, _015387_, _015388_, _015389_, _015390_, _015391_, _015392_, _015393_, _015394_, _015395_, _015396_, _015397_, _015398_, _015399_, _015400_, _015401_, _015402_, _015403_, _015404_, _015405_, _015406_, _015407_, _015408_, _015409_, _015410_, _015411_, _015412_, _015413_, _015414_, _015415_, _015416_, _015417_, _015418_, _015419_, _015420_, _015421_, _015422_, _015423_, _015424_, _015425_, _015426_, _015427_, _015428_, _015429_, _015430_, _015431_, _015432_, _015433_, _015434_, _015435_, _015436_, _015437_, _015438_, _015439_, _015440_, _015441_, _015442_, _015443_, _015444_, _015445_, _015446_, _015447_, _015448_, _015449_, _015450_, _015451_, _015452_, _015453_, _015454_, _015455_, _015456_, _015457_, _015458_, _015459_, _015460_, _015461_, _015462_, _015463_, _015464_, _015465_, _015466_, _015467_, _015468_, _015469_, _015470_, _015471_, _015472_, _015473_, _015474_, _015475_, _015476_, _015477_, _015478_, _015479_, _015480_, _015481_, _015482_, _015483_, _015484_, _015485_, _015486_, _015487_, _015488_, _015489_, _015490_, _015491_, _015492_, _015493_, _015494_, _015495_, _015496_, _015497_, _015498_, _015499_, _015500_, _015501_, _015502_, _015503_, _015504_, _015505_, _015506_, _015507_, _015508_, _015509_, _015510_, _015511_, _015512_, _015513_, _015514_, _015515_, _015516_, _015517_, _015518_, _015519_, _015520_, _015521_, _015522_, _015523_, _015524_, _015525_, _015526_, _015527_, _015528_, _015529_, _015530_, _015531_, _015532_, _015533_, _015534_, _015535_, _015536_, _015537_, _015538_, _015539_, _015540_, _015541_, _015542_, _015543_, _015544_, _015545_, _015546_, _015547_, _015548_, _015549_, _015550_, _015551_, _015552_, _015553_, _015554_, _015555_, _015556_, _015557_, _015558_, _015559_, _015560_, _015561_, _015562_, _015563_, _015564_, _015565_, _015566_, _015567_, _015568_, _015569_, _015570_, _015571_, _015572_, _015573_, _015574_, _015575_, _015576_, _015577_, _015578_, _015579_, _015580_, _015581_, _015582_, _015583_, _015584_, _015585_, _015586_, _015587_, _015588_, _015589_, _015590_, _015591_, _015592_, _015593_, _015594_, _015595_, _015596_, _015597_, _015598_, _015599_, _015600_, _015601_, _015602_, _015603_, _015604_, _015605_, _015606_, _015607_, _015608_, _015609_, _015610_, _015611_, _015612_, _015613_, _015614_, _015615_, _015616_, _015617_, _015618_, _015619_, _015620_, _015621_, _015622_, _015623_, _015624_, _015625_, _015626_, _015627_, _015628_, _015629_, _015630_, _015631_, _015632_, _015633_, _015634_, _015635_, _015636_, _015637_, _015638_, _015639_, _015640_, _015641_, _015642_, _015643_, _015644_, _015645_, _015646_, _015647_, _015648_, _015649_, _015650_, _015651_, _015652_, _015653_, _015654_, _015655_, _015656_, _015657_, _015658_, _015659_, _015660_, _015661_, _015662_, _015663_, _015664_, _015665_, _015666_, _015667_, _015668_, _015669_, _015670_, _015671_, _015672_, _015673_, _015674_, _015675_, _015676_, _015677_, _015678_, _015679_, _015680_, _015681_, _015682_, _015683_, _015684_, _015685_, _015686_, _015687_, _015688_, _015689_, _015690_, _015691_, _015692_, _015693_, _015694_, _015695_, _015696_, _015697_, _015698_, _015699_, _015700_, _015701_, _015702_, _015703_, _015704_, _015705_, _015706_, _015707_, _015708_, _015709_, _015710_, _015711_, _015712_, _015713_, _015714_, _015715_, _015716_, _015717_, _015718_, _015719_, _015720_, _015721_, _015722_, _015723_, _015724_, _015725_, _015726_, _015727_, _015728_, _015729_, _015730_, _015731_, _015732_, _015733_, _015734_, _015735_, _015736_, _015737_, _015738_, _015739_, _015740_, _015741_, _015742_, _015743_, _015744_, _015745_, _015746_, _015747_, _015748_, _015749_, _015750_, _015751_, _015752_, _015753_, _015754_, _015755_, _015756_, _015757_, _015758_, _015759_, _015760_, _015761_, _015762_, _015763_, _015764_, _015765_, _015766_, _015767_, _015768_, _015769_, _015770_, _015771_, _015772_, _015773_, _015774_, _015775_, _015776_, _015777_, _015778_, _015779_, _015780_, _015781_, _015782_, _015783_, _015784_, _015785_, _015786_, _015787_, _015788_, _015789_, _015790_, _015791_, _015792_, _015793_, _015794_, _015795_, _015796_, _015797_, _015798_, _015799_, _015800_, _015801_, _015802_, _015803_, _015804_, _015805_, _015806_, _015807_, _015808_, _015809_, _015810_, _015811_, _015812_, _015813_, _015814_, _015815_, _015816_, _015817_, _015818_, _015819_, _015820_, _015821_, _015822_, _015823_, _015824_, _015825_, _015826_, _015827_, _015828_, _015829_, _015830_, _015831_, _015832_, _015833_, _015834_, _015835_, _015836_, _015837_, _015838_, _015839_, _015840_, _015841_, _015842_, _015843_, _015844_, _015845_, _015846_, _015847_, _015848_, _015849_, _015850_, _015851_, _015852_, _015853_, _015854_, _015855_, _015856_, _015857_, _015858_, _015859_, _015860_, _015861_, _015862_, _015863_, _015864_, _015865_, _015866_, _015867_, _015868_, _015869_, _015870_, _015871_, _015872_, _015873_, _015874_, _015875_, _015876_, _015877_, _015878_, _015879_, _015880_, _015881_, _015882_, _015883_, _015884_, _015885_, _015886_, _015887_, _015888_, _015889_, _015890_, _015891_, _015892_, _015893_, _015894_, _015895_, _015896_, _015897_, _015898_, _015899_, _015900_, _015901_, _015902_, _015903_, _015904_, _015905_, _015906_, _015907_, _015908_, _015909_, _015910_, _015911_, _015912_, _015913_, _015914_, _015915_, _015916_, _015917_, _015918_, _015919_, _015920_, _015921_, _015922_, _015923_, _015924_, _015925_, _015926_, _015927_, _015928_, _015929_, _015930_, _015931_, _015932_, _015933_, _015934_, _015935_, _015936_, _015937_, _015938_, _015939_, _015940_, _015941_, _015942_, _015943_, _015944_, _015945_, _015946_, _015947_, _015948_, _015949_, _015950_, _015951_, _015952_, _015953_, _015954_, _015955_, _015956_, _015957_, _015958_, _015959_, _015960_, _015961_, _015962_, _015963_, _015964_, _015965_, _015966_, _015967_, _015968_, _015969_, _015970_, _015971_, _015972_, _015973_, _015974_, _015975_, _015976_, _015977_, _015978_, _015979_, _015980_, _015981_, _015982_, _015983_, _015984_, _015985_, _015986_, _015987_, _015988_, _015989_, _015990_, _015991_, _015992_, _015993_, _015994_, _015995_, _015996_, _015997_, _015998_, _015999_, _016000_, _016001_, _016002_, _016003_, _016004_, _016005_, _016006_, _016007_, _016008_, _016009_, _016010_, _016011_, _016012_, _016013_, _016014_, _016015_, _016016_, _016017_, _016018_, _016019_, _016020_, _016021_, _016022_, _016023_, _016024_, _016025_, _016026_, _016027_, _016028_, _016029_, _016030_, _016031_, _016032_, _016033_, _016034_, _016035_, _016036_, _016037_, _016038_, _016039_, _016040_, _016041_, _016042_, _016043_, _016044_, _016045_, _016046_, _016047_, _016048_, _016049_, _016050_, _016051_, _016052_, _016053_, _016054_, _016055_, _016056_, _016057_, _016058_, _016059_, _016060_, _016061_, _016062_, _016063_, _016064_, _016065_, _016066_, _016067_, _016068_, _016069_, _016070_, _016071_, _016072_, _016073_, _016074_, _016075_, _016076_, _016077_, _016078_, _016079_, _016080_, _016081_, _016082_, _016083_, _016084_, _016085_, _016086_, _016087_, _016088_, _016089_, _016090_, _016091_, _016092_, _016093_, _016094_, _016095_, _016096_, _016097_, _016098_, _016099_, _016100_, _016101_, _016102_, _016103_, _016104_, _016105_, _016106_, _016107_, _016108_, _016109_, _016110_, _016111_, _016112_, _016113_, _016114_, _016115_, _016116_, _016117_, _016118_, _016119_, _016120_, _016121_, _016122_, _016123_, _016124_, _016125_, _016126_, _016127_, _016128_, _016129_, _016130_, _016131_, _016132_, _016133_, _016134_, _016135_, _016136_, _016137_, _016138_, _016139_, _016140_, _016141_, _016142_, _016143_, _016144_, _016145_, _016146_, _016147_, _016148_, _016149_, _016150_, _016151_, _016152_, _016153_, _016154_, _016155_, _016156_, _016157_, _016158_, _016159_, _016160_, _016161_, _016162_, _016163_, _016164_, _016165_, _016166_, _016167_, _016168_, _016169_, _016170_, _016171_, _016172_, _016173_, _016174_, _016175_, _016176_, _016177_, _016178_, _016179_, _016180_, _016181_, _016182_, _016183_, _016184_, _016185_, _016186_, _016187_, _016188_, _016189_, _016190_, _016191_, _016192_, _016193_, _016194_, _016195_, _016196_, _016197_, _016198_, _016199_, _016200_, _016201_, _016202_, _016203_, _016204_, _016205_, _016206_, _016207_, _016208_, _016209_, _016210_, _016211_, _016212_, _016213_, _016214_, _016215_, _016216_, _016217_, _016218_, _016219_, _016220_, _016221_, _016222_, _016223_, _016224_, _016225_, _016226_, _016227_, _016228_, _016229_, _016230_, _016231_, _016232_, _016233_, _016234_, _016235_, _016236_, _016237_, _016238_, _016239_, _016240_, _016241_, _016242_, _016243_, _016244_, _016245_, _016246_, _016247_, _016248_, _016249_, _016250_, _016251_, _016252_, _016253_, _016254_, _016255_, _016256_, _016257_, _016258_, _016259_, _016260_, _016261_, _016262_, _016263_, _016264_, _016265_, _016266_, _016267_, _016268_, _016269_, _016270_, _016271_, _016272_, _016273_, _016274_, _016275_, _016276_, _016277_, _016278_, _016279_, _016280_, _016281_, _016282_, _016283_, _016284_, _016285_, _016286_, _016287_, _016288_, _016289_, _016290_, _016291_, _016292_, _016293_, _016294_, _016295_, _016296_, _016297_, _016298_, _016299_, _016300_, _016301_, _016302_, _016303_, _016304_, _016305_, _016306_, _016307_, _016308_, _016309_, _016310_, _016311_, _016312_, _016313_, _016314_, _016315_, _016316_, _016317_, _016318_, _016319_, _016320_, _016321_, _016322_, _016323_, _016324_, _016325_, _016326_, _016327_, _016328_, _016329_, _016330_, _016331_, _016332_, _016333_, _016334_, _016335_, _016336_, _016337_, _016338_, _016339_, _016340_, _016341_, _016342_, _016343_, _016344_, _016345_, _016346_, _016347_, _016348_, _016349_, _016350_, _016351_, _016352_, _016353_, _016354_, _016355_, _016356_, _016357_, _016358_, _016359_, _016360_, _016361_, _016362_, _016363_, _016364_, _016365_, _016366_, _016367_, _016368_, _016369_, _016370_, _016371_, _016372_, _016373_, _016374_, _016375_, _016376_, _016377_, _016378_, _016379_, _016380_, _016381_, _016382_, _016383_, _016384_, _016385_, _016386_, _016387_, _016388_, _016389_, _016390_, _016391_, _016392_, _016393_, _016394_, _016395_, _016396_, _016397_, _016398_, _016399_, _016400_, _016401_, _016402_, _016403_, _016404_, _016405_, _016406_, _016407_, _016408_, _016409_, _016410_, _016411_, _016412_, _016413_, _016414_, _016415_, _016416_, _016417_, _016418_, _016419_, _016420_, _016421_, _016422_, _016423_, _016424_, _016425_, _016426_, _016427_, _016428_, _016429_, _016430_, _016431_, _016432_, _016433_, _016434_, _016435_, _016436_, _016437_, _016438_, _016439_, _016440_, _016441_, _016442_, _016443_, _016444_, _016445_, _016446_, _016447_, _016448_, _016449_, _016450_, _016451_, _016452_, _016453_, _016454_, _016455_, _016456_, _016457_, _016458_, _016459_, _016460_, _016461_, _016462_, _016463_, _016464_, _016465_, _016466_, _016467_, _016468_, _016469_, _016470_, _016471_, _016472_, _016473_, _016474_, _016475_, _016476_, _016477_, _016478_, _016479_, _016480_, _016481_, _016482_, _016483_, _016484_, _016485_, _016486_, _016487_, _016488_, _016489_, _016490_, _016491_, _016492_, _016493_, _016494_, _016495_, _016496_, _016497_, _016498_, _016499_, _016500_, _016501_, _016502_, _016503_, _016504_, _016505_, _016506_, _016507_, _016508_, _016509_, _016510_, _016511_, _016512_, _016513_, _016514_, _016515_, _016516_, _016517_, _016518_, _016519_, _016520_, _016521_, _016522_, _016523_, _016524_, _016525_, _016526_, _016527_, _016528_, _016529_, _016530_, _016531_, _016532_, _016533_, _016534_, _016535_, _016536_, _016537_, _016538_, _016539_, _016540_, _016541_, _016542_, _016543_, _016544_, _016545_, _016546_, _016547_, _016548_, _016549_, _016550_, _016551_, _016552_, _016553_, _016554_, _016555_, _016556_, _016557_, _016558_, _016559_, _016560_, _016561_, _016562_, _016563_, _016564_, _016565_, _016566_, _016567_, _016568_, _016569_, _016570_, _016571_, _016572_, _016573_, _016574_, _016575_, _016576_, _016577_, _016578_, _016579_, _016580_, _016581_, _016582_, _016583_, _016584_, _016585_, _016586_, _016587_, _016588_, _016589_, _016590_, _016591_, _016592_, _016593_, _016594_, _016595_, _016596_, _016597_, _016598_, _016599_, _016600_, _016601_, _016602_, _016603_, _016604_, _016605_, _016606_, _016607_, _016608_, _016609_, _016610_, _016611_, _016612_, _016613_, _016614_, _016615_, _016616_, _016617_, _016618_, _016619_, _016620_, _016621_, _016622_, _016623_, _016624_, _016625_, _016626_, _016627_, _016628_, _016629_, _016630_, _016631_, _016632_, _016633_, _016634_, _016635_, _016636_, _016637_, _016638_, _016639_, _016640_, _016641_, _016642_, _016643_, _016644_, _016645_, _016646_, _016647_, _016648_, _016649_, _016650_, _016651_, _016652_, _016653_, _016654_, _016655_, _016656_, _016657_, _016658_, _016659_, _016660_, _016661_, _016662_, _016663_, _016664_, _016665_, _016666_, _016667_, _016668_, _016669_, _016670_, _016671_, _016672_, _016673_, _016674_, _016675_, _016676_, _016677_, _016678_, _016679_, _016680_, _016681_, _016682_, _016683_, _016684_, _016685_, _016686_, _016687_, _016688_, _016689_, _016690_, _016691_, _016692_, _016693_, _016694_, _016695_, _016696_, _016697_, _016698_, _016699_, _016700_, _016701_, _016702_, _016703_, _016704_, _016705_, _016706_, _016707_, _016708_, _016709_, _016710_, _016711_, _016712_, _016713_, _016714_, _016715_, _016716_, _016717_, _016718_, _016719_, _016720_, _016721_, _016722_, _016723_, _016724_, _016725_, _016726_, _016727_, _016728_, _016729_, _016730_, _016731_, _016732_, _016733_, _016734_, _016735_, _016736_, _016737_, _016738_, _016739_, _016740_, _016741_, _016742_, _016743_, _016744_, _016745_, _016746_, _016747_, _016748_, _016749_, _016750_, _016751_, _016752_, _016753_, _016754_, _016755_, _016756_, _016757_, _016758_, _016759_, _016760_, _016761_, _016762_, _016763_, _016764_, _016765_, _016766_, _016767_, _016768_, _016769_, _016770_, _016771_, _016772_, _016773_, _016774_, _016775_, _016776_, _016777_, _016778_, _016779_, _016780_, _016781_, _016782_, _016783_, _016784_, _016785_, _016786_, _016787_, _016788_, _016789_, _016790_, _016791_, _016792_, _016793_, _016794_, _016795_, _016796_, _016797_, _016798_, _016799_, _016800_, _016801_, _016802_, _016803_, _016804_, _016805_, _016806_, _016807_, _016808_, _016809_, _016810_, _016811_, _016812_, _016813_, _016814_, _016815_, _016816_, _016817_, _016818_, _016819_, _016820_, _016821_, _016822_, _016823_, _016824_, _016825_, _016826_, _016827_, _016828_, _016829_, _016830_, _016831_, _016832_, _016833_, _016834_, _016835_, _016836_, _016837_, _016838_, _016839_, _016840_, _016841_, _016842_, _016843_, _016844_, _016845_, _016846_, _016847_, _016848_, _016849_, _016850_, _016851_, _016852_, _016853_, _016854_, _016855_, _016856_, _016857_, _016858_, _016859_, _016860_, _016861_, _016862_, _016863_, _016864_, _016865_, _016866_, _016867_, _016868_, _016869_, _016870_, _016871_, _016872_, _016873_, _016874_, _016875_, _016876_, _016877_, _016878_, _016879_, _016880_, _016881_, _016882_, _016883_, _016884_, _016885_, _016886_, _016887_, _016888_, _016889_, _016890_, _016891_, _016892_, _016893_, _016894_, _016895_, _016896_, _016897_, _016898_, _016899_, _016900_, _016901_, _016902_, _016903_, _016904_, _016905_, _016906_, _016907_, _016908_, _016909_, _016910_, _016911_, _016912_, _016913_, _016914_, _016915_, _016916_, _016917_, _016918_, _016919_, _016920_, _016921_, _016922_, _016923_, _016924_, _016925_, _016926_, _016927_, _016928_, _016929_, _016930_, _016931_, _016932_, _016933_, _016934_, _016935_, _016936_, _016937_, _016938_, _016939_, _016940_, _016941_, _016942_, _016943_, _016944_, _016945_, _016946_, _016947_, _016948_, _016949_, _016950_, _016951_, _016952_, _016953_, _016954_, _016955_, _016956_, _016957_, _016958_, _016959_, _016960_, _016961_, _016962_, _016963_, _016964_, _016965_, _016966_, _016967_, _016968_, _016969_, _016970_, _016971_, _016972_, _016973_, _016974_, _016975_, _016976_, _016977_, _016978_, _016979_, _016980_, _016981_, _016982_, _016983_, _016984_, _016985_, _016986_, _016987_, _016988_, _016989_, _016990_, _016991_, _016992_, _016993_, _016994_, _016995_, _016996_, _016997_, _016998_, _016999_, _017000_, _017001_, _017002_, _017003_, _017004_, _017005_, _017006_, _017007_, _017008_, _017009_, _017010_, _017011_, _017012_, _017013_, _017014_, _017015_, _017016_, _017017_, _017018_, _017019_, _017020_, _017021_, _017022_, _017023_, _017024_, _017025_, _017026_, _017027_, _017028_, _017029_, _017030_, _017031_, _017032_, _017033_, _017034_, _017035_, _017036_, _017037_, _017038_, _017039_, _017040_, _017041_, _017042_, _017043_, _017044_, _017045_, _017046_, _017047_, _017048_, _017049_, _017050_, _017051_, _017052_, _017053_, _017054_, _017055_, _017056_, _017057_, _017058_, _017059_, _017060_, _017061_, _017062_, _017063_, _017064_, _017065_, _017066_, _017067_, _017068_, _017069_, _017070_, _017071_, _017072_, _017073_, _017074_, _017075_, _017076_, _017077_, _017078_, _017079_, _017080_, _017081_, _017082_, _017083_, _017084_, _017085_, _017086_, _017087_, _017088_, _017089_, _017090_, _017091_, _017092_, _017093_, _017094_, _017095_, _017096_, _017097_, _017098_, _017099_, _017100_, _017101_, _017102_, _017103_, _017104_, _017105_, _017106_, _017107_, _017108_, _017109_, _017110_, _017111_, _017112_, _017113_, _017114_, _017115_, _017116_, _017117_, _017118_, _017119_, _017120_, _017121_, _017122_, _017123_, _017124_, _017125_, _017126_, _017127_, _017128_, _017129_, _017130_, _017131_, _017132_, _017133_, _017134_, _017135_, _017136_, _017137_, _017138_, _017139_, _017140_, _017141_, _017142_, _017143_, _017144_, _017145_, _017146_, _017147_, _017148_, _017149_, _017150_, _017151_, _017152_, _017153_, _017154_, _017155_, _017156_, _017157_, _017158_, _017159_, _017160_, _017161_, _017162_, _017163_, _017164_, _017165_, _017166_, _017167_, _017168_, _017169_, _017170_, _017171_, _017172_, _017173_, _017174_, _017175_, _017176_, _017177_, _017178_, _017179_, _017180_, _017181_, _017182_, _017183_, _017184_, _017185_, _017186_, _017187_, _017188_, _017189_, _017190_, _017191_, _017192_, _017193_, _017194_, _017195_, _017196_, _017197_, _017198_, _017199_, _017200_, _017201_, _017202_, _017203_, _017204_, _017205_, _017206_, _017207_, _017208_, _017209_, _017210_, _017211_, _017212_, _017213_, _017214_, _017215_, _017216_, _017217_, _017218_, _017219_, _017220_, _017221_, _017222_, _017223_, _017224_, _017225_, _017226_, _017227_, _017228_, _017229_, _017230_, _017231_, _017232_, _017233_, _017234_, _017235_, _017236_, _017237_, _017238_, _017239_, _017240_, _017241_, _017242_, _017243_, _017244_, _017245_, _017246_, _017247_, _017248_, _017249_, _017250_, _017251_, _017252_, _017253_, _017254_, _017255_, _017256_, _017257_, _017258_, _017259_, _017260_, _017261_, _017262_, _017263_, _017264_, _017265_, _017266_, _017267_, _017268_, _017269_, _017270_, _017271_, _017272_, _017273_, _017274_, _017275_, _017276_, _017277_, _017278_, _017279_, _017280_, _017281_, _017282_, _017283_, _017284_, _017285_, _017286_, _017287_, _017288_, _017289_, _017290_, _017291_, _017292_, _017293_, _017294_, _017295_, _017296_, _017297_, _017298_, _017299_, _017300_, _017301_, _017302_, _017303_, _017304_, _017305_, _017306_, _017307_, _017308_, _017309_, _017310_, _017311_, _017312_, _017313_, _017314_, _017315_, _017316_, _017317_, _017318_, _017319_, _017320_, _017321_, _017322_, _017323_, _017324_, _017325_, _017326_, _017327_, _017328_, _017329_, _017330_, _017331_, _017332_, _017333_, _017334_, _017335_, _017336_, _017337_, _017338_, _017339_, _017340_, _017341_, _017342_, _017343_, _017344_, _017345_, _017346_, _017347_, _017348_, _017349_, _017350_, _017351_, _017352_, _017353_, _017354_, _017355_, _017356_, _017357_, _017358_, _017359_, _017360_, _017361_, _017362_, _017363_, _017364_, _017365_, _017366_, _017367_, _017368_, _017369_, _017370_, _017371_, _017372_, _017373_, _017374_, _017375_, _017376_, _017377_, _017378_, _017379_, _017380_, _017381_, _017382_, _017383_, _017384_, _017385_, _017386_, _017387_, _017388_, _017389_, _017390_, _017391_, _017392_, _017393_, _017394_, _017395_, _017396_, _017397_, _017398_, _017399_, _017400_, _017401_, _017402_, _017403_, _017404_, _017405_, _017406_, _017407_, _017408_, _017409_, _017410_, _017411_, _017412_, _017413_, _017414_, _017415_, _017416_, _017417_, _017418_, _017419_, _017420_, _017421_, _017422_, _017423_, _017424_, _017425_, _017426_, _017427_, _017428_, _017429_, _017430_, _017431_, _017432_, _017433_, _017434_, _017435_, _017436_, _017437_, _017438_, _017439_, _017440_, _017441_, _017442_, _017443_, _017444_, _017445_, _017446_, _017447_, _017448_, _017449_, _017450_, _017451_, _017452_, _017453_, _017454_, _017455_, _017456_, _017457_, _017458_, _017459_, _017460_, _017461_, _017462_, _017463_, _017464_, _017465_, _017466_, _017467_, _017468_, _017469_, _017470_, _017471_, _017472_, _017473_, _017474_, _017475_, _017476_, _017477_, _017478_, _017479_, _017480_, _017481_, _017482_, _017483_, _017484_, _017485_, _017486_, _017487_, _017488_, _017489_, _017490_, _017491_, _017492_, _017493_, _017494_, _017495_, _017496_, _017497_, _017498_, _017499_, _017500_, _017501_, _017502_, _017503_, _017504_, _017505_, _017506_, _017507_, _017508_, _017509_, _017510_, _017511_, _017512_, _017513_, _017514_, _017515_, _017516_, _017517_, _017518_, _017519_, _017520_, _017521_, _017522_, _017523_, _017524_, _017525_, _017526_, _017527_, _017528_, _017529_, _017530_, _017531_, _017532_, _017533_, _017534_, _017535_, _017536_, _017537_, _017538_, _017539_, _017540_, _017541_, _017542_, _017543_, _017544_, _017545_, _017546_, _017547_, _017548_, _017549_, _017550_, _017551_, _017552_, _017553_, _017554_, _017555_, _017556_, _017557_, _017558_, _017559_, _017560_, _017561_, _017562_, _017563_, _017564_, _017565_, _017566_, _017567_, _017568_, _017569_, _017570_, _017571_, _017572_, _017573_, _017574_, _017575_, _017576_, _017577_, _017578_, _017579_, _017580_, _017581_, _017582_, _017583_, _017584_, _017585_, _017586_, _017587_, _017588_, _017589_, _017590_, _017591_, _017592_, _017593_, _017594_, _017595_, _017596_, _017597_, _017598_, _017599_, _017600_, _017601_, _017602_, _017603_, _017604_, _017605_, _017606_, _017607_, _017608_, _017609_, _017610_, _017611_, _017612_, _017613_, _017614_, _017615_, _017616_, _017617_, _017618_, _017619_, _017620_, _017621_, _017622_, _017623_, _017624_, _017625_, _017626_, _017627_, _017628_, _017629_, _017630_, _017631_, _017632_, _017633_, _017634_, _017635_, _017636_, _017637_, _017638_, _017639_, _017640_, _017641_, _017642_, _017643_, _017644_, _017645_, _017646_, _017647_, _017648_, _017649_, _017650_, _017651_, _017652_, _017653_, _017654_, _017655_, _017656_, _017657_, _017658_, _017659_, _017660_, _017661_, _017662_, _017663_, _017664_, _017665_, _017666_, _017667_, _017668_, _017669_, _017670_, _017671_, _017672_, _017673_, _017674_, _017675_, _017676_, _017677_, _017678_, _017679_, _017680_, _017681_, _017682_, _017683_, _017684_, _017685_, _017686_, _017687_, _017688_, _017689_, _017690_, _017691_, _017692_, _017693_, _017694_, _017695_, _017696_, _017697_, _017698_, _017699_, _017700_, _017701_, _017702_, _017703_, _017704_, _017705_, _017706_, _017707_, _017708_, _017709_, _017710_, _017711_, _017712_, _017713_, _017714_, _017715_, _017716_, _017717_, _017718_, _017719_, _017720_, _017721_, _017722_, _017723_, _017724_, _017725_, _017726_, _017727_, _017728_, _017729_, _017730_, _017731_, _017732_, _017733_, _017734_, _017735_, _017736_, _017737_, _017738_, _017739_, _017740_, _017741_, _017742_, _017743_, _017744_, _017745_, _017746_, _017747_, _017748_, _017749_, _017750_, _017751_, _017752_, _017753_, _017754_, _017755_, _017756_, _017757_, _017758_, _017759_, _017760_, _017761_, _017762_, _017763_, _017764_, _017765_, _017766_, _017767_, _017768_, _017769_, _017770_, _017771_, _017772_, _017773_, _017774_, _017775_, _017776_, _017777_, _017778_, _017779_, _017780_, _017781_, _017782_, _017783_, _017784_, _017785_, _017786_, _017787_, _017788_, _017789_, _017790_, _017791_, _017792_, _017793_, _017794_, _017795_, _017796_, _017797_, _017798_, _017799_, _017800_, _017801_, _017802_, _017803_, _017804_, _017805_, _017806_, _017807_, _017808_, _017809_, _017810_, _017811_, _017812_, _017813_, _017814_, _017815_, _017816_, _017817_, _017818_, _017819_, _017820_, _017821_, _017822_, _017823_, _017824_, _017825_, _017826_, _017827_, _017828_, _017829_, _017830_, _017831_, _017832_, _017833_, _017834_, _017835_, _017836_, _017837_, _017838_, _017839_, _017840_, _017841_, _017842_, _017843_, _017844_, _017845_, _017846_, _017847_, _017848_, _017849_, _017850_, _017851_, _017852_, _017853_, _017854_, _017855_, _017856_, _017857_, _017858_, _017859_, _017860_, _017861_, _017862_, _017863_, _017864_, _017865_, _017866_, _017867_, _017868_, _017869_, _017870_, _017871_, _017872_, _017873_, _017874_, _017875_, _017876_, _017877_, _017878_, _017879_, _017880_, _017881_, _017882_, _017883_, _017884_, _017885_, _017886_, _017887_, _017888_, _017889_, _017890_, _017891_, _017892_, _017893_, _017894_, _017895_, _017896_, _017897_, _017898_, _017899_, _017900_, _017901_, _017902_, _017903_, _017904_, _017905_, _017906_, _017907_, _017908_, _017909_, _017910_, _017911_, _017912_, _017913_, _017914_, _017915_, _017916_, _017917_, _017918_, _017919_, _017920_, _017921_, _017922_, _017923_, _017924_, _017925_, _017926_, _017927_, _017928_, _017929_, _017930_, _017931_, _017932_, _017933_, _017934_, _017935_, _017936_, _017937_, _017938_, _017939_, _017940_, _017941_, _017942_, _017943_, _017944_, _017945_, _017946_, _017947_, _017948_, _017949_, _017950_, _017951_, _017952_, _017953_, _017954_, _017955_, _017956_, _017957_, _017958_, _017959_, _017960_, _017961_, _017962_, _017963_, _017964_, _017965_, _017966_, _017967_, _017968_, _017969_, _017970_, _017971_, _017972_, _017973_, _017974_, _017975_, _017976_, _017977_, _017978_, _017979_, _017980_, _017981_, _017982_, _017983_, _017984_, _017985_, _017986_, _017987_, _017988_, _017989_, _017990_, _017991_, _017992_, _017993_, _017994_, _017995_, _017996_, _017997_, _017998_, _017999_, _018000_, _018001_, _018002_, _018003_, _018004_, _018005_, _018006_, _018007_, _018008_, _018009_, _018010_, _018011_, _018012_, _018013_, _018014_, _018015_, _018016_, _018017_, _018018_, _018019_, _018020_, _018021_, _018022_, _018023_, _018024_, _018025_, _018026_, _018027_, _018028_, _018029_, _018030_, _018031_, _018032_, _018033_, _018034_, _018035_, _018036_, _018037_, _018038_, _018039_, _018040_, _018041_, _018042_, _018043_, _018044_, _018045_, _018046_, _018047_, _018048_, _018049_, _018050_, _018051_, _018052_, _018053_, _018054_, _018055_, _018056_, _018057_, _018058_, _018059_, _018060_, _018061_, _018062_, _018063_, _018064_, _018065_, _018066_, _018067_, _018068_, _018069_, _018070_, _018071_, _018072_, _018073_, _018074_, _018075_, _018076_, _018077_, _018078_, _018079_, _018080_, _018081_, _018082_, _018083_, _018084_, _018085_, _018086_, _018087_, _018088_, _018089_, _018090_, _018091_, _018092_, _018093_, _018094_, _018095_, _018096_, _018097_, _018098_, _018099_, _018100_, _018101_, _018102_, _018103_, _018104_, _018105_, _018106_, _018107_, _018108_, _018109_, _018110_, _018111_, _018112_, _018113_, _018114_, _018115_, _018116_, _018117_, _018118_, _018119_, _018120_, _018121_, _018122_, _018123_, _018124_, _018125_, _018126_, _018127_, _018128_, _018129_, _018130_, _018131_, _018132_, _018133_, _018134_, _018135_, _018136_, _018137_, _018138_, _018139_, _018140_, _018141_, _018142_, _018143_, _018144_, _018145_, _018146_, _018147_, _018148_, _018149_, _018150_, _018151_, _018152_, _018153_, _018154_, _018155_, _018156_, _018157_, _018158_, _018159_, _018160_, _018161_, _018162_, _018163_, _018164_, _018165_, _018166_, _018167_, _018168_, _018169_, _018170_, _018171_, _018172_, _018173_, _018174_, _018175_, _018176_, _018177_, _018178_, _018179_, _018180_, _018181_, _018182_, _018183_, _018184_, _018185_, _018186_, _018187_, _018188_, _018189_, _018190_, _018191_, _018192_, _018193_, _018194_, _018195_, _018196_, _018197_, _018198_, _018199_, _018200_, _018201_, _018202_, _018203_, _018204_, _018205_, _018206_, _018207_, _018208_, _018209_, _018210_, _018211_, _018212_, _018213_, _018214_, _018215_, _018216_, _018217_, _018218_, _018219_, _018220_, _018221_, _018222_, _018223_, _018224_, _018225_, _018226_, _018227_, _018228_, _018229_, _018230_, _018231_, _018232_, _018233_, _018234_, _018235_, _018236_, _018237_, _018238_, _018239_, _018240_, _018241_, _018242_, _018243_, _018244_, _018245_, _018246_, _018247_, _018248_, _018249_, _018250_, _018251_, _018252_, _018253_, _018254_, _018255_, _018256_, _018257_, _018258_, _018259_, _018260_, _018261_, _018262_, _018263_, _018264_, _018265_, _018266_, _018267_, _018268_, _018269_, _018270_, _018271_, _018272_, _018273_, _018274_, _018275_, _018276_, _018277_, _018278_, _018279_, _018280_, _018281_, _018282_, _018283_, _018284_, _018285_, _018286_, _018287_, _018288_, _018289_, _018290_, _018291_, _018292_, _018293_, _018294_, _018295_, _018296_, _018297_, _018298_, _018299_, _018300_, _018301_, _018302_, _018303_, _018304_, _018305_, _018306_, _018307_, _018308_, _018309_, _018310_, _018311_, _018312_, _018313_, _018314_, _018315_, _018316_, _018317_, _018318_, _018319_, _018320_, _018321_, _018322_, _018323_, _018324_, _018325_, _018326_, _018327_, _018328_, _018329_, _018330_, _018331_, _018332_, _018333_, _018334_, _018335_, _018336_, _018337_, _018338_, _018339_, _018340_, _018341_, _018342_, _018343_, _018344_, _018345_, _018346_, _018347_, _018348_, _018349_, _018350_, _018351_, _018352_, _018353_, _018354_, _018355_, _018356_, _018357_, _018358_, _018359_, _018360_, _018361_, _018362_, _018363_, _018364_, _018365_, _018366_, _018367_, _018368_, _018369_, _018370_, _018371_, _018372_, _018373_, _018374_, _018375_, _018376_, _018377_, _018378_, _018379_, _018380_, _018381_, _018382_, _018383_, _018384_, _018385_, _018386_, _018387_, _018388_, _018389_, _018390_, _018391_, _018392_, _018393_, _018394_, _018395_, _018396_, _018397_, _018398_, _018399_, _018400_, _018401_, _018402_, _018403_, _018404_, _018405_, _018406_, _018407_, _018408_, _018409_, _018410_, _018411_, _018412_, _018413_, _018414_, _018415_, _018416_, _018417_, _018418_, _018419_, _018420_, _018421_, _018422_, _018423_, _018424_, _018425_, _018426_, _018427_, _018428_, _018429_, _018430_, _018431_, _018432_, _018433_, _018434_, _018435_, _018436_, _018437_, _018438_, _018439_, _018440_, _018441_, _018442_, _018443_, _018444_, _018445_, _018446_, _018447_, _018448_, _018449_, _018450_, _018451_, _018452_, _018453_, _018454_, _018455_, _018456_, _018457_, _018458_, _018459_, _018460_, _018461_, _018462_, _018463_, _018464_, _018465_, _018466_, _018467_, _018468_, _018469_, _018470_, _018471_, _018472_, _018473_, _018474_, _018475_, _018476_, _018477_, _018478_, _018479_, _018480_, _018481_, _018482_, _018483_, _018484_, _018485_, _018486_, _018487_, _018488_, _018489_, _018490_, _018491_, _018492_, _018493_, _018494_, _018495_, _018496_, _018497_, _018498_, _018499_, _018500_, _018501_, _018502_, _018503_, _018504_, _018505_, _018506_, _018507_, _018508_, _018509_, _018510_, _018511_, _018512_, _018513_, _018514_, _018515_, _018516_, _018517_, _018518_, _018519_, _018520_, _018521_, _018522_, _018523_, _018524_, _018525_, _018526_, _018527_, _018528_, _018529_, _018530_, _018531_, _018532_, _018533_, _018534_, _018535_, _018536_, _018537_, _018538_, _018539_, _018540_, _018541_, _018542_, _018543_, _018544_, _018545_, _018546_, _018547_, _018548_, _018549_, _018550_, _018551_, _018552_, _018553_, _018554_, _018555_, _018556_, _018557_, _018558_, _018559_, _018560_, _018561_, _018562_, _018563_, _018564_, _018565_, _018566_, _018567_, _018568_, _018569_, _018570_, _018571_, _018572_, _018573_, _018574_, _018575_, _018576_, _018577_, _018578_, _018579_, _018580_, _018581_, _018582_, _018583_, _018584_, _018585_, _018586_, _018587_, _018588_, _018589_, _018590_, _018591_, _018592_, _018593_, _018594_, _018595_, _018596_, _018597_, _018598_, _018599_, _018600_, _018601_, _018602_, _018603_, _018604_, _018605_, _018606_, _018607_, _018608_, _018609_, _018610_, _018611_, _018612_, _018613_, _018614_, _018615_, _018616_, _018617_, _018618_, _018619_, _018620_, _018621_, _018622_, _018623_, _018624_, _018625_, _018626_, _018627_, _018628_, _018629_, _018630_, _018631_, _018632_, _018633_, _018634_, _018635_, _018636_, _018637_, _018638_, _018639_, _018640_, _018641_, _018642_, _018643_, _018644_, _018645_, _018646_, _018647_, _018648_, _018649_, _018650_, _018651_, _018652_, _018653_, _018654_, _018655_, _018656_, _018657_, _018658_, _018659_, _018660_, _018661_, _018662_, _018663_, _018664_, _018665_, _018666_, _018667_, _018668_, _018669_, _018670_, _018671_, _018672_, _018673_, _018674_, _018675_, _018676_, _018677_, _018678_, _018679_, _018680_, _018681_, _018682_, _018683_, _018684_, _018685_, _018686_, _018687_, _018688_, _018689_, _018690_, _018691_, _018692_, _018693_, _018694_, _018695_, _018696_, _018697_, _018698_, _018699_, _018700_, _018701_, _018702_, _018703_, _018704_, _018705_, _018706_, _018707_, _018708_, _018709_, _018710_, _018711_, _018712_, _018713_, _018714_, _018715_, _018716_, _018717_, _018718_, _018719_, _018720_, _018721_, _018722_, _018723_, _018724_, _018725_, _018726_, _018727_, _018728_, _018729_, _018730_, _018731_, _018732_, _018733_, _018734_, _018735_, _018736_, _018737_, _018738_, _018739_, _018740_, _018741_, _018742_, _018743_, _018744_, _018745_, _018746_, _018747_, _018748_, _018749_, _018750_, _018751_, _018752_, _018753_, _018754_, _018755_, _018756_, _018757_, _018758_, _018759_, _018760_, _018761_, _018762_, _018763_, _018764_, _018765_, _018766_, _018767_, _018768_, _018769_, _018770_, _018771_, _018772_, _018773_, _018774_, _018775_, _018776_, _018777_, _018778_, _018779_, _018780_, _018781_, _018782_, _018783_, _018784_, _018785_, _018786_, _018787_, _018788_, _018789_, _018790_, _018791_, _018792_, _018793_, _018794_, _018795_, _018796_, _018797_, _018798_, _018799_, _018800_, _018801_, _018802_, _018803_, _018804_, _018805_, _018806_, _018807_, _018808_, _018809_, _018810_, _018811_, _018812_, _018813_, _018814_, _018815_, _018816_, _018817_, _018818_, _018819_, _018820_, _018821_, _018822_, _018823_, _018824_, _018825_, _018826_, _018827_, _018828_, _018829_, _018830_, _018831_, _018832_, _018833_, _018834_, _018835_, _018836_, _018837_, _018838_, _018839_, _018840_, _018841_, _018842_, _018843_, _018844_, _018845_, _018846_, _018847_, _018848_, _018849_, _018850_, _018851_, _018852_, _018853_, _018854_, _018855_, _018856_, _018857_, _018858_, _018859_, _018860_, _018861_, _018862_, _018863_, _018864_, _018865_, _018866_, _018867_, _018868_, _018869_, _018870_, _018871_, _018872_, _018873_, _018874_, _018875_, _018876_, _018877_, _018878_, _018879_, _018880_, _018881_, _018882_, _018883_, _018884_, _018885_, _018886_, _018887_, _018888_, _018889_, _018890_, _018891_, _018892_, _018893_, _018894_, _018895_, _018896_, _018897_, _018898_, _018899_, _018900_, _018901_, _018902_, _018903_, _018904_, _018905_, _018906_, _018907_, _018908_, _018909_, _018910_, _018911_, _018912_, _018913_, _018914_, _018915_, _018916_, _018917_, _018918_, _018919_, _018920_, _018921_, _018922_, _018923_, _018924_, _018925_, _018926_, _018927_, _018928_, _018929_, _018930_, _018931_, _018932_, _018933_, _018934_, _018935_, _018936_, _018937_, _018938_, _018939_, _018940_, _018941_, _018942_, _018943_, _018944_, _018945_, _018946_, _018947_, _018948_, _018949_, _018950_, _018951_, _018952_, _018953_, _018954_, _018955_, _018956_, _018957_, _018958_, _018959_, _018960_, _018961_, _018962_, _018963_, _018964_, _018965_, _018966_, _018967_, _018968_, _018969_, _018970_, _018971_, _018972_, _018973_, _018974_, _018975_, _018976_, _018977_, _018978_, _018979_, _018980_, _018981_, _018982_, _018983_, _018984_, _018985_, _018986_, _018987_, _018988_, _018989_, _018990_, _018991_, _018992_, _018993_, _018994_, _018995_, _018996_, _018997_, _018998_, _018999_, _019000_, _019001_, _019002_, _019003_, _019004_, _019005_, _019006_, _019007_, _019008_, _019009_, _019010_, _019011_, _019012_, _019013_, _019014_, _019015_, _019016_, _019017_, _019018_, _019019_, _019020_, _019021_, _019022_, _019023_, _019024_, _019025_, _019026_, _019027_, _019028_, _019029_, _019030_, _019031_, _019032_, _019033_, _019034_, _019035_, _019036_, _019037_, _019038_, _019039_, _019040_, _019041_, _019042_, _019043_, _019044_, _019045_, _019046_, _019047_, _019048_, _019049_, _019050_, _019051_, _019052_, _019053_, _019054_, _019055_, _019056_, _019057_, _019058_, _019059_, _019060_, _019061_, _019062_, _019063_, _019064_, _019065_, _019066_, _019067_, _019068_, _019069_, _019070_, _019071_, _019072_, _019073_, _019074_, _019075_, _019076_, _019077_, _019078_, _019079_, _019080_, _019081_, _019082_, _019083_, _019084_, _019085_, _019086_, _019087_, _019088_, _019089_, _019090_, _019091_, _019092_, _019093_, _019094_, _019095_, _019096_, _019097_, _019098_, _019099_, _019100_, _019101_, _019102_, _019103_, _019104_, _019105_, _019106_, _019107_, _019108_, _019109_, _019110_, _019111_, _019112_, _019113_, _019114_, _019115_, _019116_, _019117_, _019118_, _019119_, _019120_, _019121_, _019122_, _019123_, _019124_, _019125_, _019126_, _019127_, _019128_, _019129_, _019130_, _019131_, _019132_, _019133_, _019134_, _019135_, _019136_, _019137_, _019138_, _019139_, _019140_, _019141_, _019142_, _019143_, _019144_, _019145_, _019146_, _019147_, _019148_, _019149_, _019150_, _019151_, _019152_, _019153_, _019154_, _019155_, _019156_, _019157_, _019158_, _019159_, _019160_, _019161_, _019162_, _019163_, _019164_, _019165_, _019166_, _019167_, _019168_, _019169_, _019170_, _019171_, _019172_, _019173_, _019174_, _019175_, _019176_, _019177_, _019178_, _019179_, _019180_, _019181_, _019182_, _019183_, _019184_, _019185_, _019186_, _019187_, _019188_, _019189_, _019190_, _019191_, _019192_, _019193_, _019194_, _019195_, _019196_, _019197_, _019198_, _019199_, _019200_, _019201_, _019202_, _019203_, _019204_, _019205_, _019206_, _019207_, _019208_, _019209_, _019210_, _019211_, _019212_, _019213_, _019214_, _019215_, _019216_, _019217_, _019218_, _019219_, _019220_, _019221_, _019222_, _019223_, _019224_, _019225_, _019226_, _019227_, _019228_, _019229_, _019230_, _019231_, _019232_, _019233_, _019234_, _019235_, _019236_, _019237_, _019238_, _019239_, _019240_, _019241_, _019242_, _019243_, _019244_, _019245_, _019246_, _019247_, _019248_, _019249_, _019250_, _019251_, _019252_, _019253_, _019254_, _019255_, _019256_, _019257_, _019258_, _019259_, _019260_, _019261_, _019262_, _019263_, _019264_, _019265_, _019266_, _019267_, _019268_, _019269_, _019270_, _019271_, _019272_, _019273_, _019274_, _019275_, _019276_, _019277_, _019278_, _019279_, _019280_, _019281_, _019282_, _019283_, _019284_, _019285_, _019286_, _019287_, _019288_, _019289_, _019290_, _019291_, _019292_, _019293_, _019294_, _019295_, _019296_, _019297_, _019298_, _019299_, _019300_, _019301_, _019302_, _019303_, _019304_, _019305_, _019306_, _019307_, _019308_, _019309_, _019310_, _019311_, _019312_, _019313_, _019314_, _019315_, _019316_, _019317_, _019318_, _019319_, _019320_, _019321_, _019322_, _019323_, _019324_, _019325_, _019326_, _019327_, _019328_, _019329_, _019330_, _019331_, _019332_, _019333_, _019334_, _019335_, _019336_, _019337_, _019338_, _019339_, _019340_, _019341_, _019342_, _019343_, _019344_, _019345_, _019346_, _019347_, _019348_, _019349_, _019350_, _019351_, _019352_, _019353_, _019354_, _019355_, _019356_, _019357_, _019358_, _019359_, _019360_, _019361_, _019362_, _019363_, _019364_, _019365_, _019366_, _019367_, _019368_, _019369_, _019370_, _019371_, _019372_, _019373_, _019374_, _019375_, _019376_, _019377_, _019378_, _019379_, _019380_, _019381_, _019382_, _019383_, _019384_, _019385_, _019386_, _019387_, _019388_, _019389_, _019390_, _019391_, _019392_, _019393_, _019394_, _019395_, _019396_, _019397_, _019398_, _019399_, _019400_, _019401_, _019402_, _019403_, _019404_, _019405_, _019406_, _019407_, _019408_, _019409_, _019410_, _019411_, _019412_, _019413_, _019414_, _019415_, _019416_, _019417_, _019418_, _019419_, _019420_, _019421_, _019422_, _019423_, _019424_, _019425_, _019426_, _019427_, _019428_, _019429_, _019430_, _019431_, _019432_, _019433_, _019434_, _019435_, _019436_, _019437_, _019438_, _019439_, _019440_, _019441_, _019442_, _019443_, _019444_, _019445_, _019446_, _019447_, _019448_, _019449_, _019450_, _019451_, _019452_, _019453_, _019454_, _019455_, _019456_, _019457_, _019458_, _019459_, _019460_, _019461_, _019462_, _019463_, _019464_, _019465_, _019466_, _019467_, _019468_, _019469_, _019470_, _019471_, _019472_, _019473_, _019474_, _019475_, _019476_, _019477_, _019478_, _019479_, _019480_, _019481_, _019482_, _019483_, _019484_, _019485_, _019486_, _019487_, _019488_, _019489_, _019490_, _019491_, _019492_, _019493_, _019494_, _019495_, _019496_, _019497_, _019498_, _019499_, _019500_, _019501_, _019502_, _019503_, _019504_, _019505_, _019506_, _019507_, _019508_, _019509_, _019510_, _019511_, _019512_, _019513_, _019514_, _019515_, _019516_, _019517_, _019518_, _019519_, _019520_, _019521_, _019522_, _019523_, _019524_, _019525_, _019526_, _019527_, _019528_, _019529_, _019530_, _019531_, _019532_, _019533_, _019534_, _019535_, _019536_, _019537_, _019538_, _019539_, _019540_, _019541_, _019542_, _019543_, _019544_, _019545_, _019546_, _019547_, _019548_, _019549_, _019550_, _019551_, _019552_, _019553_, _019554_, _019555_, _019556_, _019557_, _019558_, _019559_, _019560_, _019561_, _019562_, _019563_, _019564_, _019565_, _019566_, _019567_, _019568_, _019569_, _019570_, _019571_, _019572_, _019573_, _019574_, _019575_, _019576_, _019577_, _019578_, _019579_, _019580_, _019581_, _019582_, _019583_, _019584_, _019585_, _019586_, _019587_, _019588_, _019589_, _019590_, _019591_, _019592_, _019593_, _019594_, _019595_, _019596_, _019597_, _019598_, _019599_, _019600_, _019601_, _019602_, _019603_, _019604_, _019605_, _019606_, _019607_, _019608_, _019609_, _019610_, _019611_, _019612_, _019613_, _019614_, _019615_, _019616_, _019617_, _019618_, _019619_, _019620_, _019621_, _019622_, _019623_, _019624_, _019625_, _019626_, _019627_, _019628_, _019629_, _019630_, _019631_, _019632_, _019633_, _019634_, _019635_, _019636_, _019637_, _019638_, _019639_, _019640_, _019641_, _019642_, _019643_, _019644_, _019645_, _019646_, _019647_, _019648_, _019649_, _019650_, _019651_, _019652_, _019653_, _019654_, _019655_, _019656_, _019657_, _019658_, _019659_, _019660_, _019661_, _019662_, _019663_, _019664_, _019665_, _019666_, _019667_, _019668_, _019669_, _019670_, _019671_, _019672_, _019673_, _019674_, _019675_, _019676_, _019677_, _019678_, _019679_, _019680_, _019681_, _019682_, _019683_, _019684_, _019685_, _019686_, _019687_, _019688_, _019689_, _019690_, _019691_, _019692_, _019693_, _019694_, _019695_, _019696_, _019697_, _019698_, _019699_, _019700_, _019701_, _019702_, _019703_, _019704_, _019705_, _019706_, _019707_, _019708_, _019709_, _019710_, _019711_, _019712_, _019713_, _019714_, _019715_, _019716_, _019717_, _019718_, _019719_, _019720_, _019721_, _019722_, _019723_, _019724_, _019725_, _019726_, _019727_, _019728_, _019729_, _019730_, _019731_, _019732_, _019733_, _019734_, _019735_, _019736_, _019737_, _019738_, _019739_, _019740_, _019741_, _019742_, _019743_, _019744_, _019745_, _019746_, _019747_, _019748_, _019749_, _019750_, _019751_, _019752_, _019753_, _019754_, _019755_, _019756_, _019757_, _019758_, _019759_, _019760_, _019761_, _019762_, _019763_, _019764_, _019765_, _019766_, _019767_, _019768_, _019769_, _019770_, _019771_, _019772_, _019773_, _019774_, _019775_, _019776_, _019777_, _019778_, _019779_, _019780_, _019781_, _019782_, _019783_, _019784_, _019785_, _019786_, _019787_, _019788_, _019789_, _019790_, _019791_, _019792_, _019793_, _019794_, _019795_, _019796_, _019797_, _019798_, _019799_, _019800_, _019801_, _019802_, _019803_, _019804_, _019805_, _019806_, _019807_, _019808_, _019809_, _019810_, _019811_, _019812_, _019813_, _019814_, _019815_, _019816_, _019817_, _019818_, _019819_, _019820_, _019821_, _019822_, _019823_, _019824_, _019825_, _019826_, _019827_, _019828_, _019829_, _019830_, _019831_, _019832_, _019833_, _019834_, _019835_, _019836_, _019837_, _019838_, _019839_, _019840_, _019841_, _019842_, _019843_, _019844_, _019845_, _019846_, _019847_, _019848_, _019849_, _019850_, _019851_, _019852_, _019853_, _019854_, _019855_, _019856_, _019857_, _019858_, _019859_, _019860_, _019861_, _019862_, _019863_, _019864_, _019865_, _019866_, _019867_, _019868_, _019869_, _019870_, _019871_, _019872_, _019873_, _019874_, _019875_, _019876_, _019877_, _019878_, _019879_, _019880_, _019881_, _019882_, _019883_, _019884_, _019885_, _019886_, _019887_, _019888_, _019889_, _019890_, _019891_, _019892_, _019893_, _019894_, _019895_, _019896_, _019897_, _019898_, _019899_, _019900_, _019901_, _019902_, _019903_, _019904_, _019905_, _019906_, _019907_, _019908_, _019909_, _019910_, _019911_, _019912_, _019913_, _019914_, _019915_, _019916_, _019917_, _019918_, _019919_, _019920_, _019921_, _019922_, _019923_, _019924_, _019925_, _019926_, _019927_, _019928_, _019929_, _019930_, _019931_, _019932_, _019933_, _019934_, _019935_, _019936_, _019937_, _019938_, _019939_, _019940_, _019941_, _019942_, _019943_, _019944_, _019945_, _019946_, _019947_, _019948_, _019949_, _019950_, _019951_, _019952_, _019953_, _019954_, _019955_, _019956_, _019957_, _019958_, _019959_, _019960_, _019961_, _019962_, _019963_, _019964_, _019965_, _019966_, _019967_, _019968_, _019969_, _019970_, _019971_, _019972_, _019973_, _019974_, _019975_, _019976_, _019977_, _019978_, _019979_, _019980_, _019981_, _019982_, _019983_, _019984_, _019985_, _019986_, _019987_, _019988_, _019989_, _019990_, _019991_, _019992_, _019993_, _019994_, _019995_, _019996_, _019997_, _019998_, _019999_, _020000_, _020001_, _020002_, _020003_, _020004_, _020005_, _020006_, _020007_, _020008_, _020009_, _020010_, _020011_, _020012_, _020013_, _020014_, _020015_, _020016_, _020017_, _020018_, _020019_, _020020_, _020021_, _020022_, _020023_, _020024_, _020025_, _020026_, _020027_, _020028_, _020029_, _020030_, _020031_, _020032_, _020033_, _020034_, _020035_, _020036_, _020037_, _020038_, _020039_, _020040_, _020041_, _020042_, _020043_, _020044_, _020045_, _020046_, _020047_, _020048_, _020049_, _020050_, _020051_, _020052_, _020053_, _020054_, _020055_, _020056_, _020057_, _020058_, _020059_, _020060_, _020061_, _020062_, _020063_, _020064_, _020065_, _020066_, _020067_, _020068_, _020069_, _020070_, _020071_, _020072_, _020073_, _020074_, _020075_, _020076_, _020077_, _020078_, _020079_, _020080_, _020081_, _020082_, _020083_, _020084_, _020085_, _020086_, _020087_, _020088_, _020089_, _020090_, _020091_, _020092_, _020093_, _020094_, _020095_, _020096_, _020097_, _020098_, _020099_, _020100_, _020101_, _020102_, _020103_, _020104_, _020105_, _020106_, _020107_, _020108_, _020109_, _020110_, _020111_, _020112_, _020113_, _020114_, _020115_, _020116_, _020117_, _020118_, _020119_, _020120_, _020121_, _020122_, _020123_, _020124_, _020125_, _020126_, _020127_, _020128_, _020129_, _020130_, _020131_, _020132_, _020133_, _020134_, _020135_, _020136_, _020137_, _020138_, _020139_, _020140_, _020141_, _020142_, _020143_, _020144_, _020145_, _020146_, _020147_, _020148_, _020149_, _020150_, _020151_, _020152_, _020153_, _020154_, _020155_, _020156_, _020157_, _020158_, _020159_, _020160_, _020161_, _020162_, _020163_, _020164_, _020165_, _020166_, _020167_, _020168_, _020169_, _020170_, _020171_, _020172_, _020173_, _020174_, _020175_, _020176_, _020177_, _020178_, _020179_, _020180_, _020181_, _020182_, _020183_, _020184_, _020185_, _020186_, _020187_, _020188_, _020189_, _020190_, _020191_, _020192_, _020193_, _020194_, _020195_, _020196_, _020197_, _020198_, _020199_, _020200_, _020201_, _020202_, _020203_, _020204_, _020205_, _020206_, _020207_, _020208_, _020209_, _020210_, _020211_, _020212_, _020213_, _020214_, _020215_, _020216_, _020217_, _020218_, _020219_, _020220_, _020221_, _020222_, _020223_, _020224_, _020225_, _020226_, _020227_, _020228_, _020229_, _020230_, _020231_, _020232_, _020233_, _020234_, _020235_, _020236_, _020237_, _020238_, _020239_, _020240_, _020241_, _020242_, _020243_, _020244_, _020245_, _020246_, _020247_, _020248_, _020249_, _020250_, _020251_, _020252_, _020253_, _020254_, _020255_, _020256_, _020257_, _020258_, _020259_, _020260_, _020261_, _020262_, _020263_, _020264_, _020265_, _020266_, _020267_, _020268_, _020269_, _020270_, _020271_, _020272_, _020273_, _020274_, _020275_, _020276_, _020277_, _020278_, _020279_, _020280_, _020281_, _020282_, _020283_, _020284_, _020285_, _020286_, _020287_, _020288_, _020289_, _020290_, _020291_, _020292_, _020293_, _020294_, _020295_, _020296_, _020297_, _020298_, _020299_, _020300_, _020301_, _020302_, _020303_, _020304_, _020305_, _020306_, _020307_, _020308_, _020309_, _020310_, _020311_, _020312_, _020313_, _020314_, _020315_, _020316_, _020317_, _020318_, _020319_, _020320_, _020321_, _020322_, _020323_, _020324_, _020325_, _020326_, _020327_, _020328_, _020329_, _020330_, _020331_, _020332_, _020333_, _020334_, _020335_, _020336_, _020337_, _020338_, _020339_, _020340_, _020341_, _020342_, _020343_, _020344_, _020345_, _020346_, _020347_, _020348_, _020349_, _020350_, _020351_, _020352_, _020353_, _020354_, _020355_, _020356_, _020357_, _020358_, _020359_, _020360_, _020361_, _020362_, _020363_, _020364_, _020365_, _020366_, _020367_, _020368_, _020369_, _020370_, _020371_, _020372_, _020373_, _020374_, _020375_, _020376_, _020377_, _020378_, _020379_, _020380_, _020381_, _020382_, _020383_, _020384_, _020385_, _020386_, _020387_, _020388_, _020389_, _020390_, _020391_, _020392_, _020393_, _020394_, _020395_, _020396_, _020397_, _020398_, _020399_, _020400_, _020401_, _020402_, _020403_, _020404_, _020405_, _020406_, _020407_, _020408_, _020409_, _020410_, _020411_, _020412_, _020413_, _020414_, _020415_, _020416_, _020417_, _020418_, _020419_, _020420_, _020421_, _020422_, _020423_, _020424_, _020425_, _020426_, _020427_, _020428_, _020429_, _020430_, _020431_, _020432_, _020433_, _020434_, _020435_, _020436_, _020437_, _020438_, _020439_, _020440_, _020441_, _020442_, _020443_, _020444_, _020445_, _020446_, _020447_, _020448_, _020449_, _020450_, _020451_, _020452_, _020453_, _020454_, _020455_, _020456_, _020457_, _020458_, _020459_, _020460_, _020461_, _020462_, _020463_, _020464_, _020465_, _020466_, _020467_, _020468_, _020469_, _020470_, _020471_, _020472_, _020473_, _020474_, _020475_, _020476_, _020477_, _020478_, _020479_, _020480_, _020481_, _020482_, _020483_, _020484_, _020485_, _020486_, _020487_, _020488_, _020489_, _020490_, _020491_, _020492_, _020493_, _020494_, _020495_, _020496_, _020497_, _020498_, _020499_, _020500_, _020501_, _020502_, _020503_, _020504_, _020505_, _020506_, _020507_, _020508_, _020509_, _020510_, _020511_, _020512_, _020513_, _020514_, _020515_, _020516_, _020517_, _020518_, _020519_, _020520_, _020521_, _020522_, _020523_, _020524_, _020525_, _020526_, _020527_, _020528_, _020529_, _020530_, _020531_, _020532_, _020533_, _020534_, _020535_, _020536_, _020537_, _020538_, _020539_, _020540_, _020541_, _020542_, _020543_, _020544_, _020545_, _020546_, _020547_, _020548_, _020549_, _020550_, _020551_, _020552_, _020553_, _020554_, _020555_, _020556_, _020557_, _020558_, _020559_, _020560_, _020561_, _020562_, _020563_, _020564_, _020565_, _020566_, _020567_, _020568_, _020569_, _020570_, _020571_, _020572_, _020573_, _020574_, _020575_, _020576_, _020577_, _020578_, _020579_, _020580_, _020581_, _020582_, _020583_, _020584_, _020585_, _020586_, _020587_, _020588_, _020589_, _020590_, _020591_, _020592_, _020593_, _020594_, _020595_, _020596_, _020597_, _020598_, _020599_, _020600_, _020601_, _020602_, _020603_, _020604_, _020605_, _020606_, _020607_, _020608_, _020609_, _020610_, _020611_, _020612_, _020613_, _020614_, _020615_, _020616_, _020617_, _020618_, _020619_, _020620_, _020621_, _020622_, _020623_, _020624_, _020625_, _020626_, _020627_, _020628_, _020629_, _020630_, _020631_, _020632_, _020633_, _020634_, _020635_, _020636_, _020637_, _020638_, _020639_, _020640_, _020641_, _020642_, _020643_, _020644_, _020645_, _020646_, _020647_, _020648_, _020649_, _020650_, _020651_, _020652_, _020653_, _020654_, _020655_, _020656_, _020657_, _020658_, _020659_, _020660_, _020661_, _020662_, _020663_, _020664_, _020665_, _020666_, _020667_, _020668_, _020669_, _020670_, _020671_, _020672_, _020673_, _020674_, _020675_, _020676_, _020677_, _020678_, _020679_, _020680_, _020681_, _020682_, _020683_, _020684_, _020685_, _020686_, _020687_, _020688_, _020689_, _020690_, _020691_, _020692_, _020693_, _020694_, _020695_, _020696_, _020697_, _020698_, _020699_, _020700_, _020701_, _020702_, _020703_, _020704_, _020705_, _020706_, _020707_, _020708_, _020709_, _020710_, _020711_, _020712_, _020713_, _020714_, _020715_, _020716_, _020717_, _020718_, _020719_, _020720_, _020721_, _020722_, _020723_, _020724_, _020725_, _020726_, _020727_, _020728_, _020729_, _020730_, _020731_, _020732_, _020733_, _020734_, _020735_, _020736_, _020737_, _020738_, _020739_, _020740_, _020741_, _020742_, _020743_, _020744_, _020745_, _020746_, _020747_, _020748_, _020749_, _020750_, _020751_, _020752_, _020753_, _020754_, _020755_, _020756_, _020757_, _020758_, _020759_, _020760_, _020761_, _020762_, _020763_, _020764_, _020765_, _020766_, _020767_, _020768_, _020769_, _020770_, _020771_, _020772_, _020773_, _020774_, _020775_, _020776_, _020777_, _020778_, _020779_, _020780_, _020781_, _020782_, _020783_, _020784_, _020785_, _020786_, _020787_, _020788_, _020789_, _020790_, _020791_, _020792_, _020793_, _020794_, _020795_, _020796_, _020797_, _020798_, _020799_, _020800_, _020801_, _020802_, _020803_, _020804_, _020805_, _020806_, _020807_, _020808_, _020809_, _020810_, _020811_, _020812_, _020813_, _020814_, _020815_, _020816_, _020817_, _020818_, _020819_, _020820_, _020821_, _020822_, _020823_, _020824_, _020825_, _020826_, _020827_, _020828_, _020829_, _020830_, _020831_, _020832_, _020833_, _020834_, _020835_, _020836_, _020837_, _020838_, _020839_, _020840_, _020841_, _020842_, _020843_, _020844_, _020845_, _020846_, _020847_, _020848_, _020849_, _020850_, _020851_, _020852_, _020853_, _020854_, _020855_, _020856_, _020857_, _020858_, _020859_, _020860_, _020861_, _020862_, _020863_, _020864_, _020865_, _020866_, _020867_, _020868_, _020869_, _020870_, _020871_, _020872_, _020873_, _020874_, _020875_, _020876_, _020877_, _020878_, _020879_, _020880_, _020881_, _020882_, _020883_, _020884_, _020885_, _020886_, _020887_, _020888_, _020889_, _020890_, _020891_, _020892_, _020893_, _020894_, _020895_, _020896_, _020897_, _020898_, _020899_, _020900_, _020901_, _020902_, _020903_, _020904_, _020905_, _020906_, _020907_, _020908_, _020909_, _020910_, _020911_, _020912_, _020913_, _020914_, _020915_, _020916_, _020917_, _020918_, _020919_, _020920_, _020921_, _020922_, _020923_, _020924_, _020925_, _020926_, _020927_, _020928_, _020929_, _020930_, _020931_, _020932_, _020933_, _020934_, _020935_, _020936_, _020937_, _020938_, _020939_, _020940_, _020941_, _020942_, _020943_, _020944_, _020945_, _020946_, _020947_, _020948_, _020949_, _020950_, _020951_, _020952_, _020953_, _020954_, _020955_, _020956_, _020957_, _020958_, _020959_, _020960_, _020961_, _020962_, _020963_, _020964_, _020965_, _020966_, _020967_, _020968_, _020969_, _020970_, _020971_, _020972_, _020973_, _020974_, _020975_, _020976_, _020977_, _020978_, _020979_, _020980_, _020981_, _020982_, _020983_, _020984_, _020985_, _020986_, _020987_, _020988_, _020989_, _020990_, _020991_, _020992_, _020993_, _020994_, _020995_, _020996_, _020997_, _020998_, _020999_, _021000_, _021001_, _021002_, _021003_, _021004_, _021005_, _021006_, _021007_, _021008_, _021009_, _021010_, _021011_, _021012_, _021013_, _021014_, _021015_, _021016_, _021017_, _021018_, _021019_, _021020_, _021021_, _021022_, _021023_, _021024_, _021025_, _021026_, _021027_, _021028_, _021029_, _021030_, _021031_, _021032_, _021033_, _021034_, _021035_, _021036_, _021037_, _021038_, _021039_, _021040_, _021041_, _021042_, _021043_, _021044_, _021045_, _021046_, _021047_, _021048_, _021049_, _021050_, _021051_, _021052_, _021053_, _021054_, _021055_, _021056_, _021057_, _021058_, _021059_, _021060_, _021061_, _021062_, _021063_, _021064_, _021065_, _021066_, _021067_, _021068_, _021069_, _021070_, _021071_, _021072_, _021073_, _021074_, _021075_, _021076_, _021077_, _021078_, _021079_, _021080_, _021081_, _021082_, _021083_, _021084_, _021085_, _021086_, _021087_, _021088_, _021089_, _021090_, _021091_, _021092_, _021093_, _021094_, _021095_, _021096_, _021097_, _021098_, _021099_, _021100_, _021101_, _021102_, _021103_, _021104_, _021105_, _021106_, _021107_, _021108_, _021109_, _021110_, _021111_, _021112_, _021113_, _021114_, _021115_, _021116_, _021117_, _021118_, _021119_, _021120_, _021121_, _021122_, _021123_, _021124_, _021125_, _021126_, _021127_, _021128_, _021129_, _021130_, _021131_, _021132_, _021133_, _021134_, _021135_, _021136_, _021137_, _021138_, _021139_, _021140_, _021141_, _021142_, _021143_, _021144_, _021145_, _021146_, _021147_, _021148_, _021149_, _021150_, _021151_, _021152_, _021153_, _021154_, _021155_, _021156_, _021157_, _021158_, _021159_, _021160_, _021161_, _021162_, _021163_, _021164_, _021165_, _021166_, _021167_, _021168_, _021169_, _021170_, _021171_, _021172_, _021173_, _021174_, _021175_, _021176_, _021177_, _021178_, _021179_, _021180_, _021181_, _021182_, _021183_, _021184_, _021185_, _021186_, _021187_, _021188_, _021189_, _021190_, _021191_, _021192_, _021193_, _021194_, _021195_, _021196_, _021197_, _021198_, _021199_, _021200_, _021201_, _021202_, _021203_, _021204_, _021205_, _021206_, _021207_, _021208_, _021209_, _021210_, _021211_, _021212_, _021213_, _021214_, _021215_, _021216_, _021217_, _021218_, _021219_, _021220_, _021221_, _021222_, _021223_, _021224_, _021225_, _021226_, _021227_, _021228_, _021229_, _021230_, _021231_, _021232_, _021233_, _021234_, _021235_, _021236_, _021237_, _021238_, _021239_, _021240_, _021241_, _021242_, _021243_, _021244_, _021245_, _021246_, _021247_, _021248_, _021249_, _021250_, _021251_, _021252_, _021253_, _021254_, _021255_, _021256_, _021257_, _021258_, _021259_, _021260_, _021261_, _021262_, _021263_, _021264_, _021265_, _021266_, _021267_, _021268_, _021269_, _021270_, _021271_, _021272_, _021273_, _021274_, _021275_, _021276_, _021277_, _021278_, _021279_, _021280_, _021281_, _021282_, _021283_, _021284_, _021285_, _021286_, _021287_, _021288_, _021289_, _021290_, _021291_, _021292_, _021293_, _021294_, _021295_, _021296_, _021297_, _021298_, _021299_, _021300_, _021301_, _021302_, _021303_, _021304_, _021305_, _021306_, _021307_, _021308_, _021309_, _021310_, _021311_, _021312_, _021313_, _021314_, _021315_, _021316_, _021317_, _021318_, _021319_, _021320_, _021321_, _021322_, _021323_, _021324_, _021325_, _021326_, _021327_, _021328_, _021329_, _021330_, _021331_, _021332_, _021333_, _021334_, _021335_, _021336_, _021337_, _021338_, _021339_, _021340_, _021341_, _021342_, _021343_, _021344_, _021345_, _021346_, _021347_, _021348_, _021349_, _021350_, _021351_, _021352_, _021353_, _021354_, _021355_, _021356_, _021357_, _021358_, _021359_, _021360_, _021361_, _021362_, _021363_, _021364_, _021365_, _021366_, _021367_, _021368_, _021369_, _021370_, _021371_, _021372_, _021373_, _021374_, _021375_, _021376_, _021377_, _021378_, _021379_, _021380_, _021381_, _021382_, _021383_, _021384_, _021385_, _021386_, _021387_, _021388_, _021389_, _021390_, _021391_, _021392_, _021393_, _021394_, _021395_, _021396_, _021397_, _021398_, _021399_, _021400_, _021401_, _021402_, _021403_, _021404_, _021405_, _021406_, _021407_, _021408_, _021409_, _021410_, _021411_, _021412_, _021413_, _021414_, _021415_, _021416_, _021417_, _021418_, _021419_, _021420_, _021421_, _021422_, _021423_, _021424_, _021425_, _021426_, _021427_, _021428_, _021429_, _021430_, _021431_, _021432_, _021433_, _021434_, _021435_, _021436_, _021437_, _021438_, _021439_, _021440_, _021441_, _021442_, _021443_, _021444_, _021445_, _021446_, _021447_, _021448_, _021449_, _021450_, _021451_, _021452_, _021453_, _021454_, _021455_, _021456_, _021457_, _021458_, _021459_, _021460_, _021461_, _021462_, _021463_, _021464_, _021465_, _021466_, _021467_, _021468_, _021469_, _021470_, _021471_, _021472_, _021473_, _021474_, _021475_, _021476_, _021477_, _021478_, _021479_, _021480_, _021481_, _021482_, _021483_, _021484_, _021485_, _021486_, _021487_, _021488_, _021489_, _021490_, _021491_, _021492_, _021493_, _021494_, _021495_, _021496_, _021497_, _021498_, _021499_, _021500_, _021501_, _021502_, _021503_, _021504_, _021505_, _021506_, _021507_, _021508_, _021509_, _021510_, _021511_, _021512_, _021513_, _021514_, _021515_, _021516_, _021517_, _021518_, _021519_, _021520_, _021521_, _021522_, _021523_, _021524_, _021525_, _021526_, _021527_, _021528_, _021529_, _021530_, _021531_, _021532_, _021533_, _021534_, _021535_, _021536_, _021537_, _021538_, _021539_, _021540_, _021541_, _021542_, _021543_, _021544_, _021545_, _021546_, _021547_, _021548_, _021549_, _021550_, _021551_, _021552_, _021553_, _021554_, _021555_, _021556_, _021557_, _021558_, _021559_, _021560_, _021561_, _021562_, _021563_, _021564_, _021565_, _021566_, _021567_, _021568_, _021569_, _021570_, _021571_, _021572_, _021573_, _021574_, _021575_, _021576_, _021577_, _021578_, _021579_, _021580_, _021581_, _021582_, _021583_, _021584_, _021585_, _021586_, _021587_, _021588_, _021589_, _021590_, _021591_, _021592_, _021593_, _021594_, _021595_, _021596_, _021597_, _021598_, _021599_, _021600_, _021601_, _021602_, _021603_, _021604_, _021605_, _021606_, _021607_, _021608_, _021609_, _021610_, _021611_, _021612_, _021613_, _021614_, _021615_, _021616_, _021617_, _021618_, _021619_, _021620_, _021621_, _021622_, _021623_, _021624_, _021625_, _021626_, _021627_, _021628_, _021629_, _021630_, _021631_, _021632_, _021633_, _021634_, _021635_, _021636_, _021637_, _021638_, _021639_, _021640_, _021641_, _021642_, _021643_, _021644_, _021645_, _021646_, _021647_, _021648_, _021649_, _021650_, _021651_, _021652_, _021653_, _021654_, _021655_, _021656_, _021657_, _021658_, _021659_, _021660_, _021661_, _021662_, _021663_, _021664_, _021665_, _021666_, _021667_, _021668_, _021669_, _021670_, _021671_, _021672_, _021673_, _021674_, _021675_, _021676_, _021677_, _021678_, _021679_, _021680_, _021681_, _021682_, _021683_, _021684_, _021685_, _021686_, _021687_, _021688_, _021689_, _021690_, _021691_, _021692_, _021693_, _021694_, _021695_, _021696_, _021697_, _021698_, _021699_, _021700_, _021701_, _021702_, _021703_, _021704_, _021705_, _021706_, _021707_, _021708_, _021709_, _021710_, _021711_, _021712_, _021713_, _021714_, _021715_, _021716_, _021717_, _021718_, _021719_, _021720_, _021721_, _021722_, _021723_, _021724_, _021725_, _021726_, _021727_, _021728_, _021729_, _021730_, _021731_, _021732_, _021733_, _021734_, _021735_, _021736_, _021737_, _021738_, _021739_, _021740_, _021741_, _021742_, _021743_, _021744_, _021745_, _021746_, _021747_, _021748_, _021749_, _021750_, _021751_, _021752_, _021753_, _021754_, _021755_, _021756_, _021757_, _021758_, _021759_, _021760_, _021761_, _021762_, _021763_, _021764_, _021765_, _021766_, _021767_, _021768_, _021769_, _021770_, _021771_, _021772_, _021773_, _021774_, _021775_, _021776_, _021777_, _021778_, _021779_, _021780_, _021781_, _021782_, _021783_, _021784_, _021785_, _021786_, _021787_, _021788_, _021789_, _021790_, _021791_, _021792_, _021793_, _021794_, _021795_, _021796_, _021797_, _021798_, _021799_, _021800_, _021801_, _021802_, _021803_, _021804_, _021805_, _021806_, _021807_, _021808_, _021809_, _021810_, _021811_, _021812_, _021813_, _021814_, _021815_, _021816_, _021817_, _021818_, _021819_, _021820_, _021821_, _021822_, _021823_, _021824_, _021825_, _021826_, _021827_, _021828_, _021829_, _021830_, _021831_, _021832_, _021833_, _021834_, _021835_, _021836_, _021837_, _021838_, _021839_, _021840_, _021841_, _021842_, _021843_, _021844_, _021845_, _021846_, _021847_, _021848_, _021849_, _021850_, _021851_, _021852_, _021853_, _021854_, _021855_, _021856_, _021857_, _021858_, _021859_, _021860_, _021861_, _021862_, _021863_, _021864_, _021865_, _021866_, _021867_, _021868_, _021869_, _021870_, _021871_, _021872_, _021873_, _021874_, _021875_, _021876_, _021877_, _021878_, _021879_, _021880_, _021881_, _021882_, _021883_, _021884_, _021885_, _021886_, _021887_, _021888_, _021889_, _021890_, _021891_, _021892_, _021893_, _021894_, _021895_, _021896_, _021897_, _021898_, _021899_, _021900_, _021901_, _021902_, _021903_, _021904_, _021905_, _021906_, _021907_, _021908_, _021909_, _021910_, _021911_, _021912_, _021913_, _021914_, _021915_, _021916_, _021917_, _021918_, _021919_, _021920_, _021921_, _021922_, _021923_, _021924_, _021925_, _021926_, _021927_, _021928_, _021929_, _021930_, _021931_, _021932_, _021933_, _021934_, _021935_, _021936_, _021937_, _021938_, _021939_, _021940_, _021941_, _021942_, _021943_, _021944_, _021945_, _021946_, _021947_, _021948_, _021949_, _021950_, _021951_, _021952_, _021953_, _021954_, _021955_, _021956_, _021957_, _021958_, _021959_, _021960_, _021961_, _021962_, _021963_, _021964_, _021965_, _021966_, _021967_, _021968_, _021969_, _021970_, _021971_, _021972_, _021973_, _021974_, _021975_, _021976_, _021977_, _021978_, _021979_, _021980_, _021981_, _021982_, _021983_, _021984_, _021985_, _021986_, _021987_, _021988_, _021989_, _021990_, _021991_, _021992_, _021993_, _021994_, _021995_, _021996_, _021997_, _021998_, _021999_, _022000_, _022001_, _022002_, _022003_, _022004_, _022005_, _022006_, _022007_, _022008_, _022009_, _022010_, _022011_, _022012_, _022013_, _022014_, _022015_, _022016_, _022017_, _022018_, _022019_, _022020_, _022021_, _022022_, _022023_, _022024_, _022025_, _022026_, _022027_, _022028_, _022029_, _022030_, _022031_, _022032_, _022033_, _022034_, _022035_, _022036_, _022037_, _022038_, _022039_, _022040_, _022041_, _022042_, _022043_, _022044_, _022045_, _022046_, _022047_, _022048_, _022049_, _022050_, _022051_, _022052_, _022053_, _022054_, _022055_, _022056_, _022057_, _022058_, _022059_, _022060_, _022061_, _022062_, _022063_, _022064_, _022065_, _022066_, _022067_, _022068_, _022069_, _022070_, _022071_, _022072_, _022073_, _022074_, _022075_, _022076_, _022077_, _022078_, _022079_, _022080_, _022081_, _022082_, _022083_, _022084_, _022085_, _022086_, _022087_, _022088_, _022089_, _022090_, _022091_, _022092_, _022093_, _022094_, _022095_, _022096_, _022097_, _022098_, _022099_, _022100_, _022101_, _022102_, _022103_, _022104_, _022105_, _022106_, _022107_, _022108_, _022109_, _022110_, _022111_, _022112_, _022113_, _022114_, _022115_, _022116_, _022117_, _022118_, _022119_, _022120_, _022121_, _022122_, _022123_, _022124_, _022125_, _022126_, _022127_, _022128_, _022129_, _022130_, _022131_, _022132_, _022133_, _022134_, _022135_, _022136_, _022137_, _022138_, _022139_, _022140_, _022141_, _022142_, _022143_, _022144_, _022145_, _022146_, _022147_, _022148_, _022149_, _022150_, _022151_, _022152_, _022153_, _022154_, _022155_, _022156_, _022157_, _022158_, _022159_, _022160_, _022161_, _022162_, _022163_, _022164_, _022165_, _022166_, _022167_, _022168_, _022169_, _022170_, _022171_, _022172_, _022173_, _022174_, _022175_, _022176_, _022177_, _022178_, _022179_, _022180_, _022181_, _022182_, _022183_, _022184_, _022185_, _022186_, _022187_, _022188_, _022189_, _022190_, _022191_, _022192_, _022193_, _022194_, _022195_, _022196_, _022197_, _022198_, _022199_, _022200_, _022201_, _022202_, _022203_, _022204_, _022205_, _022206_, _022207_, _022208_, _022209_, _022210_, _022211_, _022212_, _022213_, _022214_, _022215_, _022216_, _022217_, _022218_, _022219_, _022220_, _022221_, _022222_, _022223_, _022224_, _022225_, _022226_, _022227_, _022228_, _022229_, _022230_, _022231_, _022232_, _022233_, _022234_, _022235_, _022236_, _022237_, _022238_, _022239_, _022240_, _022241_, _022242_, _022243_, _022244_, _022245_, _022246_, _022247_, _022248_, _022249_, _022250_, _022251_, _022252_, _022253_, _022254_, _022255_, _022256_, _022257_, _022258_, _022259_, _022260_, _022261_, _022262_, _022263_, _022264_, _022265_, _022266_, _022267_, _022268_, _022269_, _022270_, _022271_, _022272_, _022273_, _022274_, _022275_, _022276_, _022277_, _022278_, _022279_, _022280_, _022281_, _022282_, _022283_, _022284_, _022285_, _022286_, _022287_, _022288_, _022289_, _022290_, _022291_, _022292_, _022293_, _022294_, _022295_, _022296_, _022297_, _022298_, _022299_, _022300_, _022301_, _022302_, _022303_, _022304_, _022305_, _022306_, _022307_, _022308_, _022309_, _022310_, _022311_, _022312_, _022313_, _022314_, _022315_, _022316_, _022317_, _022318_, _022319_, _022320_, _022321_, _022322_, _022323_, _022324_, _022325_, _022326_, _022327_, _022328_, _022329_, _022330_, _022331_, _022332_, _022333_, _022334_, _022335_, _022336_, _022337_, _022338_, _022339_, _022340_, _022341_, _022342_, _022343_, _022344_, _022345_, _022346_, _022347_, _022348_, _022349_, _022350_, _022351_, _022352_, _022353_, _022354_, _022355_, _022356_, _022357_, _022358_, _022359_, _022360_, _022361_, _022362_, _022363_, _022364_, _022365_, _022366_, _022367_, _022368_, _022369_, _022370_, _022371_, _022372_, _022373_, _022374_, _022375_, _022376_, _022377_, _022378_, _022379_, _022380_, _022381_, _022382_, _022383_, _022384_, _022385_, _022386_, _022387_, _022388_, _022389_, _022390_, _022391_, _022392_, _022393_, _022394_, _022395_, _022396_, _022397_, _022398_, _022399_, _022400_, _022401_, _022402_, _022403_, _022404_, _022405_, _022406_, _022407_, _022408_, _022409_, _022410_, _022411_, _022412_, _022413_, _022414_, _022415_, _022416_, _022417_, _022418_, _022419_, _022420_, _022421_, _022422_, _022423_, _022424_, _022425_, _022426_, _022427_, _022428_, _022429_, _022430_, _022431_, _022432_, _022433_, _022434_, _022435_, _022436_, _022437_, _022438_, _022439_, _022440_, _022441_, _022442_, _022443_, _022444_, _022445_, _022446_, _022447_, _022448_, _022449_, _022450_, _022451_, _022452_, _022453_, _022454_, _022455_, _022456_, _022457_, _022458_, _022459_, _022460_, _022461_, _022462_, _022463_, _022464_, _022465_, _022466_, _022467_, _022468_, _022469_, _022470_, _022471_, _022472_, _022473_, _022474_, _022475_, _022476_, _022477_, _022478_, _022479_, _022480_, _022481_, _022482_, _022483_, _022484_, _022485_, _022486_, _022487_, _022488_, _022489_, _022490_, _022491_, _022492_, _022493_, _022494_, _022495_, _022496_, _022497_, _022498_, _022499_, _022500_, _022501_, _022502_, _022503_, _022504_, _022505_, _022506_, _022507_, _022508_, _022509_, _022510_, _022511_, _022512_, _022513_, _022514_, _022515_, _022516_, _022517_, _022518_, _022519_, _022520_, _022521_, _022522_, _022523_, _022524_, _022525_, _022526_, _022527_, _022528_, _022529_, _022530_, _022531_, _022532_, _022533_, _022534_, _022535_, _022536_, _022537_, _022538_, _022539_, _022540_, _022541_, _022542_, _022543_, _022544_, _022545_, _022546_, _022547_, _022548_, _022549_, _022550_, _022551_, _022552_, _022553_, _022554_, _022555_, _022556_, _022557_, _022558_, _022559_, _022560_, _022561_, _022562_, _022563_, _022564_, _022565_, _022566_, _022567_, _022568_, _022569_, _022570_, _022571_, _022572_, _022573_, _022574_, _022575_, _022576_, _022577_, _022578_, _022579_, _022580_, _022581_, _022582_, _022583_, _022584_, _022585_, _022586_, _022587_, _022588_, _022589_, _022590_, _022591_, _022592_, _022593_, _022594_, _022595_, _022596_, _022597_, _022598_, _022599_, _022600_, _022601_, _022602_, _022603_, _022604_, _022605_, _022606_, _022607_, _022608_, _022609_, _022610_, _022611_, _022612_, _022613_, _022614_, _022615_, _022616_, _022617_, _022618_, _022619_, _022620_, _022621_, _022622_, _022623_, _022624_, _022625_, _022626_, _022627_, _022628_, _022629_, _022630_, _022631_, _022632_, _022633_, _022634_, _022635_, _022636_, _022637_, _022638_, _022639_, _022640_, _022641_, _022642_, _022643_, _022644_, _022645_, _022646_, _022647_, _022648_, _022649_, _022650_, _022651_, _022652_, _022653_, _022654_, _022655_, _022656_, _022657_, _022658_, _022659_, _022660_, _022661_, _022662_, _022663_, _022664_, _022665_, _022666_, _022667_, _022668_, _022669_, _022670_, _022671_, _022672_, _022673_, _022674_, _022675_, _022676_, _022677_, _022678_, _022679_, _022680_, _022681_, _022682_, _022683_, _022684_, _022685_, _022686_, _022687_, _022688_, _022689_, _022690_, _022691_, _022692_, _022693_, _022694_, _022695_, _022696_, _022697_, _022698_, _022699_, _022700_, _022701_, _022702_, _022703_, _022704_, _022705_, _022706_, _022707_, _022708_, _022709_, _022710_, _022711_, _022712_, _022713_, _022714_, _022715_, _022716_, _022717_, _022718_, _022719_, _022720_, _022721_, _022722_, _022723_, _022724_, _022725_, _022726_, _022727_, _022728_, _022729_, _022730_, _022731_, _022732_, _022733_, _022734_, _022735_, _022736_, _022737_, _022738_, _022739_, _022740_, _022741_, _022742_, _022743_, _022744_, _022745_, _022746_, _022747_, _022748_, _022749_, _022750_, _022751_, _022752_, _022753_, _022754_, _022755_, _022756_, _022757_, _022758_, _022759_, _022760_, _022761_, _022762_, _022763_, _022764_, _022765_, _022766_, _022767_, _022768_, _022769_, _022770_, _022771_, _022772_, _022773_, _022774_, _022775_, _022776_, _022777_, _022778_, _022779_, _022780_, _022781_, _022782_, _022783_, _022784_, _022785_, _022786_, _022787_, _022788_, _022789_, _022790_, _022791_, _022792_, _022793_, _022794_, _022795_, _022796_, _022797_, _022798_, _022799_, _022800_, _022801_, _022802_, _022803_, _022804_, _022805_, _022806_, _022807_, _022808_, _022809_, _022810_, _022811_, _022812_, _022813_, _022814_, _022815_, _022816_, _022817_, _022818_, _022819_, _022820_, _022821_, _022822_, _022823_, _022824_, _022825_, _022826_, _022827_, _022828_, _022829_, _022830_, _022831_, _022832_, _022833_, _022834_, _022835_, _022836_, _022837_, _022838_, _022839_, _022840_, _022841_, _022842_, _022843_, _022844_, _022845_, _022846_, _022847_, _022848_, _022849_, _022850_, _022851_, _022852_, _022853_, _022854_, _022855_, _022856_, _022857_, _022858_, _022859_, _022860_, _022861_, _022862_, _022863_, _022864_, _022865_, _022866_, _022867_, _022868_, _022869_, _022870_, _022871_, _022872_, _022873_, _022874_, _022875_, _022876_, _022877_, _022878_, _022879_, _022880_, _022881_, _022882_, _022883_, _022884_, _022885_, _022886_, _022887_, _022888_, _022889_, _022890_, _022891_, _022892_, _022893_, _022894_, _022895_, _022896_, _022897_, _022898_, _022899_, _022900_, _022901_, _022902_, _022903_, _022904_, _022905_, _022906_, _022907_, _022908_, _022909_, _022910_, _022911_, _022912_, _022913_, _022914_, _022915_, _022916_, _022917_, _022918_, _022919_, _022920_, _022921_, _022922_, _022923_, _022924_, _022925_, _022926_, _022927_, _022928_, _022929_, _022930_, _022931_, _022932_, _022933_, _022934_, _022935_, _022936_, _022937_, _022938_, _022939_, _022940_, _022941_, _022942_, _022943_, _022944_, _022945_, _022946_, _022947_, _022948_, _022949_, _022950_, _022951_, _022952_, _022953_, _022954_, _022955_, _022956_, _022957_, _022958_, _022959_, _022960_, _022961_, _022962_, _022963_, _022964_, _022965_, _022966_, _022967_, _022968_, _022969_, _022970_, _022971_, _022972_, _022973_, _022974_, _022975_, _022976_, _022977_, _022978_, _022979_, _022980_, _022981_, _022982_, _022983_, _022984_, _022985_, _022986_, _022987_, _022988_, _022989_, _022990_, _022991_, _022992_, _022993_, _022994_, _022995_, _022996_, _022997_, _022998_, _022999_, _023000_, _023001_, _023002_, _023003_, _023004_, _023005_, _023006_, _023007_, _023008_, _023009_, _023010_, _023011_, _023012_, _023013_, _023014_, _023015_, _023016_, _023017_, _023018_, _023019_, _023020_, _023021_, _023022_, _023023_, _023024_, _023025_, _023026_, _023027_, _023028_, _023029_, _023030_, _023031_, _023032_, _023033_, _023034_, _023035_, _023036_, _023037_, _023038_, _023039_, _023040_, _023041_, _023042_, _023043_, _023044_, _023045_, _023046_, _023047_, _023048_, _023049_, _023050_, _023051_, _023052_, _023053_, _023054_, _023055_, _023056_, _023057_, _023058_, _023059_, _023060_, _023061_, _023062_, _023063_, _023064_, _023065_, _023066_, _023067_, _023068_, _023069_, _023070_, _023071_, _023072_, _023073_, _023074_, _023075_, _023076_, _023077_, _023078_, _023079_, _023080_, _023081_, _023082_, _023083_, _023084_, _023085_, _023086_, _023087_, _023088_, _023089_, _023090_, _023091_, _023092_, _023093_, _023094_, _023095_, _023096_, _023097_, _023098_, _023099_, _023100_, _023101_, _023102_, _023103_, _023104_, _023105_, _023106_, _023107_, _023108_, _023109_, _023110_, _023111_, _023112_, _023113_, _023114_, _023115_, _023116_, _023117_, _023118_, _023119_, _023120_, _023121_, _023122_, _023123_, _023124_, _023125_, _023126_, _023127_, _023128_, _023129_, _023130_, _023131_, _023132_, _023133_, _023134_, _023135_, _023136_, _023137_, _023138_, _023139_, _023140_, _023141_, _023142_, _023143_, _023144_, _023145_, _023146_, _023147_, _023148_, _023149_, _023150_, _023151_, _023152_, _023153_, _023154_, _023155_, _023156_, _023157_, _023158_, _023159_, _023160_, _023161_, _023162_, _023163_, _023164_, _023165_, _023166_, _023167_, _023168_, _023169_, _023170_, _023171_, _023172_, _023173_, _023174_, _023175_, _023176_, _023177_, _023178_, _023179_, _023180_, _023181_, _023182_, _023183_, _023184_, _023185_, _023186_, _023187_, _023188_, _023189_, _023190_, _023191_, _023192_, _023193_, _023194_, _023195_, _023196_, _023197_, _023198_, _023199_, _023200_, _023201_, _023202_, _023203_, _023204_, _023205_, _023206_, _023207_, _023208_, _023209_, _023210_, _023211_, _023212_, _023213_, _023214_, _023215_, _023216_, _023217_, _023218_, _023219_, _023220_, _023221_, _023222_, _023223_, _023224_, _023225_, _023226_, _023227_, _023228_, _023229_, _023230_, _023231_, _023232_, _023233_, _023234_, _023235_, _023236_, _023237_, _023238_, _023239_, _023240_, _023241_, _023242_, _023243_, _023244_, _023245_, _023246_, _023247_, _023248_, _023249_, _023250_, _023251_, _023252_, _023253_, _023254_, _023255_, _023256_, _023257_, _023258_, _023259_, _023260_, _023261_, _023262_, _023263_, _023264_, _023265_, _023266_, _023267_, _023268_, _023269_, _023270_, _023271_, _023272_, _023273_, _023274_, _023275_, _023276_, _023277_, _023278_, _023279_, _023280_, _023281_, _023282_, _023283_, _023284_, _023285_, _023286_, _023287_, _023288_, _023289_, _023290_, _023291_, _023292_, _023293_, _023294_, _023295_, _023296_, _023297_, _023298_, _023299_, _023300_, _023301_, _023302_, _023303_, _023304_, _023305_, _023306_, _023307_, _023308_, _023309_, _023310_, _023311_, _023312_, _023313_, _023314_, _023315_, _023316_, _023317_, _023318_, _023319_, _023320_, _023321_, _023322_, _023323_, _023324_, _023325_, _023326_, _023327_, _023328_, _023329_, _023330_, _023331_, _023332_, _023333_, _023334_, _023335_, _023336_, _023337_, _023338_, _023339_, _023340_, _023341_, _023342_, _023343_, _023344_, _023345_, _023346_, _023347_, _023348_, _023349_, _023350_, _023351_, _023352_, _023353_, _023354_, _023355_, _023356_, _023357_, _023358_, _023359_, _023360_, _023361_, _023362_, _023363_, _023364_, _023365_, _023366_, _023367_, _023368_, _023369_, _023370_, _023371_, _023372_, _023373_, _023374_, _023375_, _023376_, _023377_, _023378_, _023379_, _023380_, _023381_, _023382_, _023383_, _023384_, _023385_, _023386_, _023387_, _023388_, _023389_, _023390_, _023391_, _023392_, _023393_, _023394_, _023395_, _023396_, _023397_, _023398_, _023399_, _023400_, _023401_, _023402_, _023403_, _023404_, _023405_, _023406_, _023407_, _023408_, _023409_, _023410_, _023411_, _023412_, _023413_, _023414_, _023415_, _023416_, _023417_, _023418_, _023419_, _023420_, _023421_, _023422_, _023423_, _023424_, _023425_, _023426_, _023427_, _023428_, _023429_, _023430_, _023431_, _023432_, _023433_, _023434_, _023435_, _023436_, _023437_, _023438_, _023439_, _023440_, _023441_, _023442_, _023443_, _023444_, _023445_, _023446_, _023447_, _023448_, _023449_, _023450_, _023451_, _023452_, _023453_, _023454_, _023455_, _023456_, _023457_, _023458_, _023459_, _023460_, _023461_, _023462_, _023463_, _023464_, _023465_, _023466_, _023467_, _023468_, _023469_, _023470_, _023471_, _023472_, _023473_, _023474_, _023475_, _023476_, _023477_, _023478_, _023479_, _023480_, _023481_, _023482_, _023483_, _023484_, _023485_, _023486_, _023487_, _023488_, _023489_, _023490_, _023491_, _023492_, _023493_, _023494_, _023495_, _023496_, _023497_, _023498_, _023499_, _023500_, _023501_, _023502_, _023503_, _023504_, _023505_, _023506_, _023507_, _023508_, _023509_, _023510_, _023511_, _023512_, _023513_, _023514_, _023515_, _023516_, _023517_, _023518_, _023519_, _023520_, _023521_, _023522_, _023523_, _023524_, _023525_, _023526_, _023527_, _023528_, _023529_, _023530_, _023531_, _023532_, _023533_, _023534_, _023535_, _023536_, _023537_, _023538_, _023539_, _023540_, _023541_, _023542_, _023543_, _023544_, _023545_, _023546_, _023547_, _023548_, _023549_, _023550_, _023551_, _023552_, _023553_, _023554_, _023555_, _023556_, _023557_, _023558_, _023559_, _023560_, _023561_, _023562_, _023563_, _023564_, _023565_, _023566_, _023567_, _023568_, _023569_, _023570_, _023571_, _023572_, _023573_, _023574_, _023575_, _023576_, _023577_, _023578_, _023579_, _023580_, _023581_, _023582_, _023583_, _023584_, _023585_, _023586_, _023587_, _023588_, _023589_, _023590_, _023591_, _023592_, _023593_, _023594_, _023595_, _023596_, _023597_, _023598_, _023599_, _023600_, _023601_, _023602_, _023603_, _023604_, _023605_, _023606_, _023607_, _023608_, _023609_, _023610_, _023611_, _023612_, _023613_, _023614_, _023615_, _023616_, _023617_, _023618_, _023619_, _023620_, _023621_, _023622_, _023623_, _023624_, _023625_, _023626_, _023627_, _023628_, _023629_, _023630_, _023631_, _023632_, _023633_, _023634_, _023635_, _023636_, _023637_, _023638_, _023639_, _023640_, _023641_, _023642_, _023643_, _023644_, _023645_, _023646_, _023647_, _023648_, _023649_, _023650_, _023651_, _023652_, _023653_, _023654_, _023655_, _023656_, _023657_, _023658_, _023659_, _023660_, _023661_, _023662_, _023663_, _023664_, _023665_, _023666_, _023667_, _023668_, _023669_, _023670_, _023671_, _023672_, _023673_, _023674_, _023675_, _023676_, _023677_, _023678_, _023679_, _023680_, _023681_, _023682_, _023683_, _023684_, _023685_, _023686_, _023687_, _023688_, _023689_, _023690_, _023691_, _023692_, _023693_, _023694_, _023695_, _023696_, _023697_, _023698_, _023699_, _023700_, _023701_, _023702_, _023703_, _023704_, _023705_, _023706_, _023707_, _023708_, _023709_, _023710_, _023711_, _023712_, _023713_, _023714_, _023715_, _023716_, _023717_, _023718_, _023719_, _023720_, _023721_, _023722_, _023723_, _023724_, _023725_, _023726_, _023727_, _023728_, _023729_, _023730_, _023731_, _023732_, _023733_, _023734_, _023735_, _023736_, _023737_, _023738_, _023739_, _023740_, _023741_, _023742_, _023743_, _023744_, _023745_, _023746_, _023747_, _023748_, _023749_, _023750_, _023751_, _023752_, _023753_, _023754_, _023755_, _023756_, _023757_, _023758_, _023759_, _023760_, _023761_, _023762_, _023763_, _023764_, _023765_, _023766_, _023767_, _023768_, _023769_, _023770_, _023771_, _023772_, _023773_, _023774_, _023775_, _023776_, _023777_, _023778_, _023779_, _023780_, _023781_, _023782_, _023783_, _023784_, _023785_, _023786_, _023787_, _023788_, _023789_, _023790_, _023791_, _023792_, _023793_, _023794_, _023795_, _023796_, _023797_, _023798_, _023799_, _023800_, _023801_, _023802_, _023803_, _023804_, _023805_, _023806_, _023807_, _023808_, _023809_, _023810_, _023811_, _023812_, _023813_, _023814_, _023815_, _023816_, _023817_, _023818_, _023819_, _023820_, _023821_, _023822_, _023823_, _023824_, _023825_, _023826_, _023827_, _023828_, _023829_, _023830_, _023831_, _023832_, _023833_, _023834_, _023835_, _023836_, _023837_, _023838_, _023839_, _023840_, _023841_, _023842_, _023843_, _023844_, _023845_, _023846_, _023847_, _023848_, _023849_, _023850_, _023851_, _023852_, _023853_, _023854_, _023855_, _023856_, _023857_, _023858_, _023859_, _023860_, _023861_, _023862_, _023863_, _023864_, _023865_, _023866_, _023867_, _023868_, _023869_, _023870_, _023871_, _023872_, _023873_, _023874_, _023875_, _023876_, _023877_, _023878_, _023879_, _023880_, _023881_, _023882_, _023883_, _023884_, _023885_, _023886_, _023887_, _023888_, _023889_, _023890_, _023891_, _023892_, _023893_, _023894_, _023895_, _023896_, _023897_, _023898_, _023899_, _023900_, _023901_, _023902_, _023903_, _023904_, _023905_, _023906_, _023907_, _023908_, _023909_, _023910_, _023911_, _023912_, _023913_, _023914_, _023915_, _023916_, _023917_, _023918_, _023919_, _023920_, _023921_, _023922_, _023923_, _023924_, _023925_, _023926_, _023927_, _023928_, _023929_, _023930_, _023931_, _023932_, _023933_, _023934_, _023935_, _023936_, _023937_, _023938_, _023939_, _023940_, _023941_, _023942_, _023943_, _023944_, _023945_, _023946_, _023947_, _023948_, _023949_, _023950_, _023951_, _023952_, _023953_, _023954_, _023955_, _023956_, _023957_, _023958_, _023959_, _023960_, _023961_, _023962_, _023963_, _023964_, _023965_, _023966_, _023967_, _023968_, _023969_, _023970_, _023971_, _023972_, _023973_, _023974_, _023975_, _023976_, _023977_, _023978_, _023979_, _023980_, _023981_, _023982_, _023983_, _023984_, _023985_, _023986_, _023987_, _023988_, _023989_, _023990_, _023991_, _023992_, _023993_, _023994_, _023995_, _023996_, _023997_, _023998_, _023999_, _024000_, _024001_, _024002_, _024003_, _024004_, _024005_, _024006_, _024007_, _024008_, _024009_, _024010_, _024011_, _024012_, _024013_, _024014_, _024015_, _024016_, _024017_, _024018_, _024019_, _024020_, _024021_, _024022_, _024023_, _024024_, _024025_, _024026_, _024027_, _024028_, _024029_, _024030_, _024031_, _024032_, _024033_, _024034_, _024035_, _024036_, _024037_, _024038_, _024039_, _024040_, _024041_, _024042_, _024043_, _024044_, _024045_, _024046_, _024047_, _024048_, _024049_, _024050_, _024051_, _024052_, _024053_, _024054_, _024055_, _024056_, _024057_, _024058_, _024059_, _024060_, _024061_, _024062_, _024063_, _024064_, _024065_, _024066_, _024067_, _024068_, _024069_, _024070_, _024071_, _024072_, _024073_, _024074_, _024075_, _024076_, _024077_, _024078_, _024079_, _024080_, _024081_, _024082_, _024083_, _024084_, _024085_, _024086_, _024087_, _024088_, _024089_, _024090_, _024091_, _024092_, _024093_, _024094_, _024095_, _024096_, _024097_, _024098_, _024099_, _024100_, _024101_, _024102_, _024103_, _024104_, _024105_, _024106_, _024107_, _024108_, _024109_, _024110_, _024111_, _024112_, _024113_, _024114_, _024115_, _024116_, _024117_, _024118_, _024119_, _024120_, _024121_, _024122_, _024123_, _024124_, _024125_, _024126_, _024127_, _024128_, _024129_, _024130_, _024131_, _024132_, _024133_, _024134_, _024135_, _024136_, _024137_, _024138_, _024139_, _024140_, _024141_, _024142_, _024143_, _024144_, _024145_, _024146_, _024147_, _024148_, _024149_, _024150_, _024151_, _024152_, _024153_, _024154_, _024155_, _024156_, _024157_, _024158_, _024159_, _024160_, _024161_, _024162_, _024163_, _024164_, _024165_, _024166_, _024167_, _024168_, _024169_, _024170_, _024171_, _024172_, _024173_, _024174_, _024175_, _024176_, _024177_, _024178_, _024179_, _024180_, _024181_, _024182_, _024183_, _024184_, _024185_, _024186_, _024187_, _024188_, _024189_, _024190_, _024191_, _024192_, _024193_, _024194_, _024195_, _024196_, _024197_, _024198_, _024199_, _024200_, _024201_, _024202_, _024203_, _024204_, _024205_, _024206_, _024207_, _024208_, _024209_, _024210_, _024211_, _024212_, _024213_, _024214_, _024215_, _024216_, _024217_, _024218_, _024219_, _024220_, _024221_, _024222_, _024223_, _024224_, _024225_, _024226_, _024227_, _024228_, _024229_, _024230_, _024231_, _024232_, _024233_, _024234_, _024235_, _024236_, _024237_, _024238_, _024239_, _024240_, _024241_, _024242_, _024243_, _024244_, _024245_, _024246_, _024247_, _024248_, _024249_, _024250_, _024251_, _024252_, _024253_, _024254_, _024255_, _024256_, _024257_, _024258_, _024259_, _024260_, _024261_, _024262_, _024263_, _024264_, _024265_, _024266_, _024267_, _024268_, _024269_, _024270_, _024271_, _024272_, _024273_, _024274_, _024275_, _024276_, _024277_, _024278_, _024279_, _024280_, _024281_, _024282_, _024283_, _024284_, _024285_, _024286_, _024287_, _024288_, _024289_, _024290_, _024291_, _024292_, _024293_, _024294_, _024295_, _024296_, _024297_, _024298_, _024299_, _024300_, _024301_, _024302_, _024303_, _024304_, _024305_, _024306_, _024307_, _024308_, _024309_, _024310_, _024311_, _024312_, _024313_, _024314_, _024315_, _024316_, _024317_, _024318_, _024319_, _024320_, _024321_, _024322_, _024323_, _024324_, _024325_, _024326_, _024327_, _024328_, _024329_, _024330_, _024331_, _024332_, _024333_, _024334_, _024335_, _024336_, _024337_, _024338_, _024339_, _024340_, _024341_, _024342_, _024343_, _024344_, _024345_, _024346_, _024347_, _024348_, _024349_, _024350_, _024351_, _024352_, _024353_, _024354_, _024355_, _024356_, _024357_, _024358_, _024359_, _024360_, _024361_, _024362_, _024363_, _024364_, _024365_, _024366_, _024367_, _024368_, _024369_, _024370_, _024371_, _024372_, _024373_, _024374_, _024375_, _024376_, _024377_, _024378_, _024379_, _024380_, _024381_, _024382_, _024383_, _024384_, _024385_, _024386_, _024387_, _024388_, _024389_, _024390_, _024391_, _024392_, _024393_, _024394_, _024395_, _024396_, _024397_, _024398_, _024399_, _024400_, _024401_, _024402_, _024403_, _024404_, _024405_, _024406_, _024407_, _024408_, _024409_, _024410_, _024411_, _024412_, _024413_, _024414_, _024415_, _024416_, _024417_, _024418_, _024419_, _024420_, _024421_, _024422_, _024423_, _024424_, _024425_, _024426_, _024427_, _024428_, _024429_, _024430_, _024431_, _024432_, _024433_, _024434_, _024435_, _024436_, _024437_, _024438_, _024439_, _024440_, _024441_, _024442_, _024443_, _024444_, _024445_, _024446_, _024447_, _024448_, _024449_, _024450_, _024451_, _024452_, _024453_, _024454_, _024455_, _024456_, _024457_, _024458_, _024459_, _024460_, _024461_, _024462_, _024463_, _024464_, _024465_, _024466_, _024467_, _024468_, _024469_, _024470_, _024471_, _024472_, _024473_, _024474_, _024475_, _024476_, _024477_, _024478_, _024479_, _024480_, _024481_, _024482_, _024483_, _024484_, _024485_, _024486_, _024487_, _024488_, _024489_, _024490_, _024491_, _024492_, _024493_, _024494_, _024495_, _024496_, _024497_, _024498_, _024499_, _024500_, _024501_, _024502_, _024503_, _024504_, _024505_, _024506_, _024507_, _024508_, _024509_, _024510_, _024511_, _024512_, _024513_, _024514_, _024515_, _024516_, _024517_, _024518_, _024519_, _024520_, _024521_, _024522_, _024523_, _024524_, _024525_, _024526_, _024527_, _024528_, _024529_, _024530_, _024531_, _024532_, _024533_, _024534_, _024535_, _024536_, _024537_, _024538_, _024539_, _024540_, _024541_, _024542_, _024543_, _024544_, _024545_, _024546_, _024547_, _024548_, _024549_, _024550_, _024551_, _024552_, _024553_, _024554_, _024555_, _024556_, _024557_, _024558_, _024559_, _024560_, _024561_, _024562_, _024563_, _024564_, _024565_, _024566_, _024567_, _024568_, _024569_, _024570_, _024571_, _024572_, _024573_, _024574_, _024575_, _024576_, _024577_, _024578_, _024579_, _024580_, _024581_, _024582_, _024583_, _024584_, _024585_, _024586_, _024587_, _024588_, _024589_, _024590_, _024591_, _024592_, _024593_, _024594_, _024595_, _024596_, _024597_, _024598_, _024599_, _024600_, _024601_, _024602_, _024603_, _024604_, _024605_, _024606_, _024607_, _024608_, _024609_, _024610_, _024611_, _024612_, _024613_, _024614_, _024615_, _024616_, _024617_, _024618_, _024619_, _024620_, _024621_, _024622_, _024623_, _024624_, _024625_, _024626_, _024627_, _024628_, _024629_, _024630_, _024631_, _024632_, _024633_, _024634_, _024635_, _024636_, _024637_, _024638_, _024639_, _024640_, _024641_, _024642_, _024643_, _024644_, _024645_, _024646_, _024647_, _024648_, _024649_, _024650_, _024651_, _024652_, _024653_, _024654_, _024655_, _024656_, _024657_, _024658_, _024659_, _024660_, _024661_, _024662_, _024663_, _024664_, _024665_, _024666_, _024667_, _024668_, _024669_, _024670_, _024671_, _024672_, _024673_, _024674_, _024675_, _024676_, _024677_, _024678_, _024679_, _024680_, _024681_, _024682_, _024683_, _024684_, _024685_, _024686_, _024687_, _024688_, _024689_, _024690_, _024691_, _024692_, _024693_, _024694_, _024695_, _024696_, _024697_, _024698_, _024699_, _024700_, _024701_, _024702_, _024703_, _024704_, _024705_, _024706_, _024707_, _024708_, _024709_, _024710_, _024711_, _024712_, _024713_, _024714_, _024715_, _024716_, _024717_, _024718_, _024719_, _024720_, _024721_, _024722_, _024723_, _024724_, _024725_, _024726_, _024727_, _024728_, _024729_, _024730_, _024731_, _024732_, _024733_, _024734_, _024735_, _024736_, _024737_, _024738_, _024739_, _024740_, _024741_, _024742_, _024743_, _024744_, _024745_, _024746_, _024747_, _024748_, _024749_, _024750_, _024751_, _024752_, _024753_, _024754_, _024755_, _024756_, _024757_, _024758_, _024759_, _024760_, _024761_, _024762_, _024763_, _024764_, _024765_, _024766_, _024767_, _024768_, _024769_, _024770_, _024771_, _024772_, _024773_, _024774_, _024775_, _024776_, _024777_, _024778_, _024779_, _024780_, _024781_, _024782_, _024783_, _024784_, _024785_, _024786_, _024787_, _024788_, _024789_, _024790_, _024791_, _024792_, _024793_, _024794_, _024795_, _024796_, _024797_, _024798_, _024799_, _024800_, _024801_, _024802_, _024803_, _024804_, _024805_, _024806_, _024807_, _024808_, _024809_, _024810_, _024811_, _024812_, _024813_, _024814_, _024815_, _024816_, _024817_, _024818_, _024819_, _024820_, _024821_, _024822_, _024823_, _024824_, _024825_, _024826_, _024827_, _024828_, _024829_, _024830_, _024831_, _024832_, _024833_, _024834_, _024835_, _024836_, _024837_, _024838_, _024839_, _024840_, _024841_, _024842_, _024843_, _024844_, _024845_, _024846_, _024847_, _024848_, _024849_, _024850_, _024851_, _024852_, _024853_, _024854_, _024855_, _024856_, _024857_, _024858_, _024859_, _024860_, _024861_, _024862_, _024863_, _024864_, _024865_, _024866_, _024867_, _024868_, _024869_, _024870_, _024871_, _024872_, _024873_, _024874_, _024875_, _024876_, _024877_, _024878_, _024879_, _024880_, _024881_, _024882_, _024883_, _024884_, _024885_, _024886_, _024887_, _024888_, _024889_, _024890_, _024891_, _024892_, _024893_, _024894_, _024895_, _024896_, _024897_, _024898_, _024899_, _024900_, _024901_, _024902_, _024903_, _024904_, _024905_, _024906_, _024907_, _024908_, _024909_, _024910_, _024911_, _024912_, _024913_, _024914_, _024915_, _024916_, _024917_, _024918_, _024919_, _024920_, _024921_, _024922_, _024923_, _024924_, _024925_, _024926_, _024927_, _024928_, _024929_, _024930_, _024931_, _024932_, _024933_, _024934_, _024935_, _024936_, _024937_, _024938_, _024939_, _024940_, _024941_, _024942_, _024943_, _024944_, _024945_, _024946_, _024947_, _024948_, _024949_, _024950_, _024951_, _024952_, _024953_, _024954_, _024955_, _024956_, _024957_, _024958_, _024959_, _024960_, _024961_, _024962_, _024963_, _024964_, _024965_, _024966_, _024967_, _024968_, _024969_, _024970_, _024971_, _024972_, _024973_, _024974_, _024975_, _024976_, _024977_, _024978_, _024979_, _024980_, _024981_, _024982_, _024983_, _024984_, _024985_, _024986_, _024987_, _024988_, _024989_, _024990_, _024991_, _024992_, _024993_, _024994_, _024995_, _024996_, _024997_, _024998_, _024999_, _025000_, _025001_, _025002_, _025003_, _025004_, _025005_, _025006_, _025007_, _025008_, _025009_, _025010_, _025011_, _025012_, _025013_, _025014_, _025015_, _025016_, _025017_, _025018_, _025019_, _025020_, _025021_, _025022_, _025023_, _025024_, _025025_, _025026_, _025027_, _025028_, _025029_, _025030_, _025031_, _025032_, _025033_, _025034_, _025035_, _025036_, _025037_, _025038_, _025039_, _025040_, _025041_, _025042_, _025043_, _025044_, _025045_, _025046_, _025047_, _025048_, _025049_, _025050_, _025051_, _025052_, _025053_, _025054_, _025055_, _025056_, _025057_, _025058_, _025059_, _025060_, _025061_, _025062_, _025063_, _025064_, _025065_, _025066_, _025067_, _025068_, _025069_, _025070_, _025071_, _025072_, _025073_, _025074_, _025075_, _025076_, _025077_, _025078_, _025079_, _025080_, _025081_, _025082_, _025083_, _025084_, _025085_, _025086_, _025087_, _025088_, _025089_, _025090_, _025091_, _025092_, _025093_, _025094_, _025095_, _025096_, _025097_, _025098_, _025099_, _025100_, _025101_, _025102_, _025103_, _025104_, _025105_, _025106_, _025107_, _025108_, _025109_, _025110_, _025111_, _025112_, _025113_, _025114_, _025115_, _025116_, _025117_, _025118_, _025119_, _025120_, _025121_, _025122_, _025123_, _025124_, _025125_, _025126_, _025127_, _025128_, _025129_, _025130_, _025131_, _025132_, _025133_, _025134_, _025135_, _025136_, _025137_, _025138_, _025139_, _025140_, _025141_, _025142_, _025143_, _025144_, _025145_, _025146_, _025147_, _025148_, _025149_, _025150_, _025151_, _025152_, _025153_, _025154_, _025155_, _025156_, _025157_, _025158_, _025159_, _025160_, _025161_, _025162_, _025163_, _025164_, _025165_, _025166_, _025167_, _025168_, _025169_, _025170_, _025171_, _025172_, _025173_, _025174_, _025175_, _025176_, _025177_, _025178_, _025179_, _025180_, _025181_, _025182_, _025183_, _025184_, _025185_, _025186_, _025187_, _025188_, _025189_, _025190_, _025191_, _025192_, _025193_, _025194_, _025195_, _025196_, _025197_, _025198_, _025199_, _025200_, _025201_, _025202_, _025203_, _025204_, _025205_, _025206_, _025207_, _025208_, _025209_, _025210_, _025211_, _025212_, _025213_, _025214_, _025215_, _025216_, _025217_, _025218_, _025219_, _025220_, _025221_, _025222_, _025223_, _025224_, _025225_, _025226_, _025227_, _025228_, _025229_, _025230_, _025231_, _025232_, _025233_, _025234_, _025235_, _025236_, _025237_, _025238_, _025239_, _025240_, _025241_, _025242_, _025243_, _025244_, _025245_, _025246_, _025247_, _025248_, _025249_, _025250_, _025251_, _025252_, _025253_, _025254_, _025255_, _025256_, _025257_, _025258_, _025259_, _025260_, _025261_, _025262_, _025263_, _025264_, _025265_, _025266_, _025267_, _025268_, _025269_, _025270_, _025271_, _025272_, _025273_, _025274_, _025275_, _025276_, _025277_, _025278_, _025279_, _025280_, _025281_, _025282_, _025283_, _025284_, _025285_, _025286_, _025287_, _025288_, _025289_, _025290_, _025291_, _025292_, _025293_, _025294_, _025295_, _025296_, _025297_, _025298_, _025299_, _025300_, _025301_, _025302_, _025303_, _025304_, _025305_, _025306_, _025307_, _025308_, _025309_, _025310_, _025311_, _025312_, _025313_, _025314_, _025315_, _025316_, _025317_, _025318_, _025319_, _025320_, _025321_, _025322_, _025323_, _025324_, _025325_, _025326_, _025327_, _025328_, _025329_, _025330_, _025331_, _025332_, _025333_, _025334_, _025335_, _025336_, _025337_, _025338_, _025339_, _025340_, _025341_, _025342_, _025343_, _025344_, _025345_, _025346_, _025347_, _025348_, _025349_, _025350_, _025351_, _025352_, _025353_, _025354_, _025355_, _025356_, _025357_, _025358_, _025359_, _025360_, _025361_, _025362_, _025363_, _025364_, _025365_, _025366_, _025367_, _025368_, _025369_, _025370_, _025371_, _025372_, _025373_, _025374_, _025375_, _025376_, _025377_, _025378_, _025379_, _025380_, _025381_, _025382_, _025383_, _025384_, _025385_, _025386_, _025387_, _025388_, _025389_, _025390_, _025391_, _025392_, _025393_, _025394_, _025395_, _025396_, _025397_, _025398_, _025399_, _025400_, _025401_, _025402_, _025403_, _025404_, _025405_, _025406_, _025407_, _025408_, _025409_, _025410_, _025411_, _025412_, _025413_, _025414_, _025415_, _025416_, _025417_, _025418_, _025419_, _025420_, _025421_, _025422_, _025423_, _025424_, _025425_, _025426_, _025427_, _025428_, _025429_, _025430_, _025431_, _025432_, _025433_, _025434_, _025435_, _025436_, _025437_, _025438_, _025439_, _025440_, _025441_, _025442_, _025443_, _025444_, _025445_, _025446_, _025447_, _025448_, _025449_, _025450_, _025451_, _025452_, _025453_, _025454_, _025455_, _025456_, _025457_, _025458_, _025459_, _025460_, _025461_, _025462_, _025463_, _025464_, _025465_, _025466_, _025467_, _025468_, _025469_, _025470_, _025471_, _025472_, _025473_, _025474_, _025475_, _025476_, _025477_, _025478_, _025479_, _025480_, _025481_, _025482_, _025483_, _025484_, _025485_, _025486_, _025487_, _025488_, _025489_, _025490_, _025491_, _025492_, _025493_, _025494_, _025495_, _025496_, _025497_, _025498_, _025499_, _025500_, _025501_, _025502_, _025503_, _025504_, _025505_, _025506_, _025507_, _025508_, _025509_, _025510_, _025511_, _025512_, _025513_, _025514_, _025515_, _025516_, _025517_, _025518_, _025519_, _025520_, _025521_, _025522_, _025523_, _025524_, _025525_, _025526_, _025527_, _025528_, _025529_, _025530_, _025531_, _025532_, _025533_, _025534_, _025535_, _025536_, _025537_, _025538_, _025539_, _025540_, _025541_, _025542_, _025543_, _025544_, _025545_, _025546_, _025547_, _025548_, _025549_, _025550_, _025551_, _025552_, _025553_, _025554_, _025555_, _025556_, _025557_, _025558_, _025559_, _025560_, _025561_, _025562_, _025563_, _025564_, _025565_, _025566_, _025567_, _025568_, _025569_, _025570_, _025571_, _025572_, _025573_, _025574_, _025575_, _025576_, _025577_, _025578_, _025579_, _025580_, _025581_, _025582_, _025583_, _025584_, _025585_, _025586_, _025587_, _025588_, _025589_, _025590_, _025591_, _025592_, _025593_, _025594_, _025595_, _025596_, _025597_, _025598_, _025599_, _025600_, _025601_, _025602_, _025603_, _025604_, _025605_, _025606_, _025607_, _025608_, _025609_, _025610_, _025611_, _025612_, _025613_, _025614_, _025615_, _025616_, _025617_, _025618_, _025619_, _025620_, _025621_, _025622_, _025623_, _025624_, _025625_, _025626_, _025627_, _025628_, _025629_, _025630_, _025631_, _025632_, _025633_, _025634_, _025635_, _025636_, _025637_, _025638_, _025639_, _025640_, _025641_, _025642_, _025643_, _025644_, _025645_, _025646_, _025647_, _025648_, _025649_, _025650_, _025651_, _025652_, _025653_, _025654_, _025655_, _025656_, _025657_, _025658_, _025659_, _025660_, _025661_, _025662_, _025663_, _025664_, _025665_, _025666_, _025667_, _025668_, _025669_, _025670_, _025671_, _025672_, _025673_, _025674_, _025675_, _025676_, _025677_, _025678_, _025679_, _025680_, _025681_, _025682_, _025683_, _025684_, _025685_, _025686_, _025687_, _025688_, _025689_, _025690_, _025691_, _025692_, _025693_, _025694_, _025695_, _025696_, _025697_, _025698_, _025699_, _025700_, _025701_, _025702_, _025703_, _025704_, _025705_, _025706_, _025707_, _025708_, _025709_, _025710_, _025711_, _025712_, _025713_, _025714_, _025715_, _025716_, _025717_, _025718_, _025719_, _025720_, _025721_, _025722_, _025723_, _025724_, _025725_, _025726_, _025727_, _025728_, _025729_, _025730_, _025731_, _025732_, _025733_, _025734_, _025735_, _025736_, _025737_, _025738_, _025739_, _025740_, _025741_, _025742_, _025743_, _025744_, _025745_, _025746_, _025747_, _025748_, _025749_, _025750_, _025751_, _025752_, _025753_, _025754_, _025755_, _025756_, _025757_, _025758_, _025759_, _025760_, _025761_, _025762_, _025763_, _025764_, _025765_, _025766_, _025767_, _025768_, _025769_, _025770_, _025771_, _025772_, _025773_, _025774_, _025775_, _025776_, _025777_, _025778_, _025779_, _025780_, _025781_, _025782_, _025783_, _025784_, _025785_, _025786_, _025787_, _025788_, _025789_, _025790_, _025791_, _025792_, _025793_, _025794_, _025795_, _025796_, _025797_, _025798_, _025799_, _025800_, _025801_, _025802_, _025803_, _025804_, _025805_, _025806_, _025807_, _025808_, _025809_, _025810_, _025811_, _025812_, _025813_, _025814_, _025815_, _025816_, _025817_, _025818_, _025819_, _025820_, _025821_, _025822_, _025823_, _025824_, _025825_, _025826_, _025827_, _025828_, _025829_, _025830_, _025831_, _025832_, _025833_, _025834_, _025835_, _025836_, _025837_, _025838_, _025839_, _025840_, _025841_, _025842_, _025843_, _025844_, _025845_, _025846_, _025847_, _025848_, _025849_, _025850_, _025851_, _025852_, _025853_, _025854_, _025855_, _025856_, _025857_, _025858_, _025859_, _025860_, _025861_, _025862_, _025863_, _025864_, _025865_, _025866_, _025867_, _025868_, _025869_, _025870_, _025871_, _025872_, _025873_, _025874_, _025875_, _025876_, _025877_, _025878_, _025879_, _025880_, _025881_, _025882_, _025883_, _025884_, _025885_, _025886_, _025887_, _025888_, _025889_, _025890_, _025891_, _025892_, _025893_, _025894_, _025895_, _025896_, _025897_, _025898_, _025899_, _025900_, _025901_, _025902_, _025903_, _025904_, _025905_, _025906_, _025907_, _025908_, _025909_, _025910_, _025911_, _025912_, _025913_, _025914_, _025915_, _025916_, _025917_, _025918_, _025919_, _025920_, _025921_, _025922_, _025923_, _025924_, _025925_, _025926_, _025927_, _025928_, _025929_, _025930_, _025931_, _025932_, _025933_, _025934_, _025935_, _025936_, _025937_, _025938_, _025939_, _025940_, _025941_, _025942_, _025943_, _025944_, _025945_, _025946_, _025947_, _025948_, _025949_, _025950_, _025951_, _025952_, _025953_, _025954_, _025955_, _025956_, _025957_, _025958_, _025959_, _025960_, _025961_, _025962_, _025963_, _025964_, _025965_, _025966_, _025967_, _025968_, _025969_, _025970_, _025971_, _025972_, _025973_, _025974_, _025975_, _025976_, _025977_, _025978_, _025979_, _025980_, _025981_, _025982_, _025983_, _025984_, _025985_, _025986_, _025987_, _025988_, _025989_, _025990_, _025991_, _025992_, _025993_, _025994_, _025995_, _025996_, _025997_, _025998_, _025999_, _026000_, _026001_, _026002_, _026003_, _026004_, _026005_, _026006_, _026007_, _026008_, _026009_, _026010_, _026011_, _026012_, _026013_, _026014_, _026015_, _026016_, _026017_, _026018_, _026019_, _026020_, _026021_, _026022_, _026023_, _026024_, _026025_, _026026_, _026027_, _026028_, _026029_, _026030_, _026031_, _026032_, _026033_, _026034_, _026035_, _026036_, _026037_, _026038_, _026039_, _026040_, _026041_, _026042_, _026043_, _026044_, _026045_, _026046_, _026047_, _026048_, _026049_, _026050_, _026051_, _026052_, _026053_, _026054_, _026055_, _026056_, _026057_, _026058_, _026059_, _026060_, _026061_, _026062_, _026063_, _026064_, _026065_, _026066_, _026067_, _026068_, _026069_, _026070_, _026071_, _026072_, _026073_, _026074_, _026075_, _026076_, _026077_, _026078_, _026079_, _026080_, _026081_, _026082_, _026083_, _026084_, _026085_, _026086_, _026087_, _026088_, _026089_, _026090_, _026091_, _026092_, _026093_, _026094_, _026095_, _026096_, _026097_, _026098_, _026099_, _026100_, _026101_, _026102_, _026103_, _026104_, _026105_, _026106_, _026107_, _026108_, _026109_, _026110_, _026111_, _026112_, _026113_, _026114_, _026115_, _026116_, _026117_, _026118_, _026119_, _026120_, _026121_, _026122_, _026123_, _026124_, _026125_, _026126_, _026127_, _026128_, _026129_, _026130_, _026131_, _026132_, _026133_, _026134_, _026135_, _026136_, _026137_, _026138_, _026139_, _026140_, _026141_, _026142_, _026143_, _026144_, _026145_, _026146_, _026147_, _026148_, _026149_, _026150_, _026151_, _026152_, _026153_, _026154_, _026155_, _026156_, _026157_, _026158_, _026159_, _026160_, _026161_, _026162_, _026163_, _026164_, _026165_, _026166_, _026167_, _026168_, _026169_, _026170_, _026171_, _026172_, _026173_, _026174_, _026175_, _026176_, _026177_, _026178_, _026179_, _026180_, _026181_, _026182_, _026183_, _026184_, _026185_, _026186_, _026187_, _026188_, _026189_, _026190_, _026191_, _026192_, _026193_, _026194_, _026195_, _026196_, _026197_, _026198_, _026199_, _026200_, _026201_, _026202_, _026203_, _026204_, _026205_, _026206_, _026207_, _026208_, _026209_, _026210_, _026211_, _026212_, _026213_, _026214_, _026215_, _026216_, _026217_, _026218_, _026219_, _026220_, _026221_, _026222_, _026223_, _026224_, _026225_, _026226_, _026227_, _026228_, _026229_, _026230_, _026231_, _026232_, _026233_, _026234_, _026235_, _026236_, _026237_, _026238_, _026239_, _026240_, _026241_, _026242_, _026243_, _026244_, _026245_, _026246_, _026247_, _026248_, _026249_, _026250_, _026251_, _026252_, _026253_, _026254_, _026255_, _026256_, _026257_, _026258_, _026259_, _026260_, _026261_, _026262_, _026263_, _026264_, _026265_, _026266_, _026267_, _026268_, _026269_, _026270_, _026271_, _026272_, _026273_, _026274_, _026275_, _026276_, _026277_, _026278_, _026279_, _026280_, _026281_, _026282_, _026283_, _026284_, _026285_, _026286_, _026287_, _026288_, _026289_, _026290_, _026291_, _026292_, _026293_, _026294_, _026295_, _026296_, _026297_, _026298_, _026299_, _026300_, _026301_, _026302_, _026303_, _026304_, _026305_, _026306_, _026307_, _026308_, _026309_, _026310_, _026311_, _026312_, _026313_, _026314_, _026315_, _026316_, _026317_, _026318_, _026319_, _026320_, _026321_, _026322_, _026323_, _026324_, _026325_, _026326_, _026327_, _026328_, _026329_, _026330_, _026331_, _026332_, _026333_, _026334_, _026335_, _026336_, _026337_, _026338_, _026339_, _026340_, _026341_, _026342_, _026343_, _026344_, _026345_, _026346_, _026347_, _026348_, _026349_, _026350_, _026351_, _026352_, _026353_, _026354_, _026355_, _026356_, _026357_, _026358_, _026359_, _026360_, _026361_, _026362_, _026363_, _026364_, _026365_, _026366_, _026367_, _026368_, _026369_, _026370_, _026371_, _026372_, _026373_, _026374_, _026375_, _026376_, _026377_, _026378_, _026379_, _026380_, _026381_, _026382_, _026383_, _026384_, _026385_, _026386_, _026387_, _026388_, _026389_, _026390_, _026391_, _026392_, _026393_, _026394_, _026395_, _026396_, _026397_, _026398_, _026399_, _026400_, _026401_, _026402_, _026403_, _026404_, _026405_, _026406_, _026407_, _026408_, _026409_, _026410_, _026411_, _026412_, _026413_, _026414_, _026415_, _026416_, _026417_, _026418_, _026419_, _026420_, _026421_, _026422_, _026423_, _026424_, _026425_, _026426_, _026427_, _026428_, _026429_, _026430_, _026431_, _026432_, _026433_, _026434_, _026435_, _026436_, _026437_, _026438_, _026439_, _026440_, _026441_, _026442_, _026443_, _026444_, _026445_, _026446_, _026447_, _026448_, _026449_, _026450_, _026451_, _026452_, _026453_, _026454_, _026455_, _026456_, _026457_, _026458_, _026459_, _026460_, _026461_, _026462_, _026463_, _026464_, _026465_, _026466_, _026467_, _026468_, _026469_, _026470_, _026471_, _026472_, _026473_, _026474_, _026475_, _026476_, _026477_, _026478_, _026479_, _026480_, _026481_, _026482_, _026483_, _026484_, _026485_, _026486_, _026487_, _026488_, _026489_, _026490_, _026491_, _026492_, _026493_, _026494_, _026495_, _026496_, _026497_, _026498_, _026499_, _026500_, _026501_, _026502_, _026503_, _026504_, _026505_, _026506_, _026507_, _026508_, _026509_, _026510_, _026511_, _026512_, _026513_, _026514_, _026515_, _026516_, _026517_, _026518_, _026519_, _026520_, _026521_, _026522_, _026523_, _026524_, _026525_, _026526_, _026527_, _026528_, _026529_, _026530_, _026531_, _026532_, _026533_, _026534_, _026535_, _026536_, _026537_, _026538_, _026539_, _026540_, _026541_, _026542_, _026543_, _026544_, _026545_, _026546_, _026547_, _026548_, _026549_, _026550_, _026551_, _026552_, _026553_, _026554_, _026555_, _026556_, _026557_, _026558_, _026559_, _026560_, _026561_, _026562_, _026563_, _026564_, _026565_, _026566_, _026567_, _026568_, _026569_, _026570_, _026571_, _026572_, _026573_, _026574_, _026575_, _026576_, _026577_, _026578_, _026579_, _026580_, _026581_, _026582_, _026583_, _026584_, _026585_, _026586_, _026587_, _026588_, _026589_, _026590_, _026591_, _026592_, _026593_, _026594_, _026595_, _026596_, _026597_, _026598_, _026599_, _026600_, _026601_, _026602_, _026603_, _026604_, _026605_, _026606_, _026607_, _026608_, _026609_, _026610_, _026611_, _026612_, _026613_, _026614_, _026615_, _026616_, _026617_, _026618_, _026619_, _026620_, _026621_, _026622_, _026623_, _026624_, _026625_, _026626_, _026627_, _026628_, _026629_, _026630_, _026631_, _026632_, _026633_, _026634_, _026635_, _026636_, _026637_, _026638_, _026639_, _026640_, _026641_, _026642_, _026643_, _026644_, _026645_, _026646_, _026647_, _026648_, _026649_, _026650_, _026651_, _026652_, _026653_, _026654_, _026655_, _026656_, _026657_, _026658_, _026659_, _026660_, _026661_, _026662_, _026663_, _026664_, _026665_, _026666_, _026667_, _026668_, _026669_, _026670_, _026671_, _026672_, _026673_, _026674_, _026675_, _026676_, _026677_, _026678_, _026679_, _026680_, _026681_, _026682_, _026683_, _026684_, _026685_, _026686_, _026687_, _026688_, _026689_, _026690_, _026691_, _026692_, _026693_, _026694_, _026695_, _026696_, _026697_, _026698_, _026699_, _026700_, _026701_, _026702_, _026703_, _026704_, _026705_, _026706_, _026707_, _026708_, _026709_, _026710_, _026711_, _026712_, _026713_, _026714_, _026715_, _026716_, _026717_, _026718_, _026719_, _026720_, _026721_, _026722_, _026723_, _026724_, _026725_, _026726_, _026727_, _026728_, _026729_, _026730_, _026731_, _026732_, _026733_, _026734_, _026735_, _026736_, _026737_, _026738_, _026739_, _026740_, _026741_, _026742_, _026743_, _026744_, _026745_, _026746_, _026747_, _026748_, _026749_, _026750_, _026751_, _026752_, _026753_, _026754_, _026755_, _026756_, _026757_, _026758_, _026759_, _026760_, _026761_, _026762_, _026763_, _026764_, _026765_, _026766_, _026767_, _026768_, _026769_, _026770_, _026771_, _026772_, _026773_, _026774_, _026775_, _026776_, _026777_, _026778_, _026779_, _026780_, _026781_, _026782_, _026783_, _026784_, _026785_, _026786_, _026787_, _026788_, _026789_, _026790_, _026791_, _026792_, _026793_, _026794_, _026795_, _026796_, _026797_, _026798_, _026799_, _026800_, _026801_, _026802_, _026803_, _026804_, _026805_, _026806_, _026807_, _026808_, _026809_, _026810_, _026811_, _026812_, _026813_, _026814_, _026815_, _026816_, _026817_, _026818_, _026819_, _026820_, _026821_, _026822_, _026823_, _026824_, _026825_, _026826_, _026827_, _026828_, _026829_, _026830_, _026831_, _026832_, _026833_, _026834_, _026835_, _026836_, _026837_, _026838_, _026839_, _026840_, _026841_, _026842_, _026843_, _026844_, _026845_, _026846_, _026847_, _026848_, _026849_, _026850_, _026851_, _026852_, _026853_, _026854_, _026855_, _026856_, _026857_, _026858_, _026859_, _026860_, _026861_, _026862_, _026863_, _026864_, _026865_, _026866_, _026867_, _026868_, _026869_, _026870_, _026871_, _026872_, _026873_, _026874_, _026875_, _026876_, _026877_, _026878_, _026879_, _026880_, _026881_, _026882_, _026883_, _026884_, _026885_, _026886_, _026887_, _026888_, _026889_, _026890_, _026891_, _026892_, _026893_, _026894_, _026895_, _026896_, _026897_, _026898_, _026899_, _026900_, _026901_, _026902_, _026903_, _026904_, _026905_, _026906_, _026907_, _026908_, _026909_, _026910_, _026911_, _026912_, _026913_, _026914_, _026915_, _026916_, _026917_, _026918_, _026919_, _026920_, _026921_, _026922_, _026923_, _026924_, _026925_, _026926_, _026927_, _026928_, _026929_, _026930_, _026931_, _026932_, _026933_, _026934_, _026935_, _026936_, _026937_, _026938_, _026939_, _026940_, _026941_, _026942_, _026943_, _026944_, _026945_, _026946_, _026947_, _026948_, _026949_, _026950_, _026951_, _026952_, _026953_, _026954_, _026955_, _026956_, _026957_, _026958_, _026959_, _026960_, _026961_, _026962_, _026963_, _026964_, _026965_, _026966_, _026967_, _026968_, _026969_, _026970_, _026971_, _026972_, _026973_, _026974_, _026975_, _026976_, _026977_, _026978_, _026979_, _026980_, _026981_, _026982_, _026983_, _026984_, _026985_, _026986_, _026987_, _026988_, _026989_, _026990_, _026991_, _026992_, _026993_, _026994_, _026995_, _026996_, _026997_, _026998_, _026999_, _027000_, _027001_, _027002_, _027003_, _027004_, _027005_, _027006_, _027007_, _027008_, _027009_, _027010_, _027011_, _027012_, _027013_, _027014_, _027015_, _027016_, _027017_, _027018_, _027019_, _027020_, _027021_, _027022_, _027023_, _027024_, _027025_, _027026_, _027027_, _027028_, _027029_, _027030_, _027031_, _027032_, _027033_, _027034_, _027035_, _027036_, _027037_, _027038_, _027039_, _027040_, _027041_, _027042_, _027043_, _027044_, _027045_, _027046_, _027047_, _027048_, _027049_, _027050_, _027051_, _027052_, _027053_, _027054_, _027055_, _027056_, _027057_, _027058_, _027059_, _027060_, _027061_, _027062_, _027063_, _027064_, _027065_, _027066_, _027067_, _027068_, _027069_, _027070_, _027071_, _027072_, _027073_, _027074_, _027075_, _027076_, _027077_, _027078_, _027079_, _027080_, _027081_, _027082_, _027083_, _027084_, _027085_, _027086_, _027087_, _027088_, _027089_, _027090_, _027091_, _027092_, _027093_, _027094_, _027095_, _027096_, _027097_, _027098_, _027099_, _027100_, _027101_, _027102_, _027103_, _027104_, _027105_, _027106_, _027107_, _027108_, _027109_, _027110_, _027111_, _027112_, _027113_, _027114_, _027115_, _027116_, _027117_, _027118_, _027119_, _027120_, _027121_, _027122_, _027123_, _027124_, _027125_, _027126_, _027127_, _027128_, _027129_, _027130_, _027131_, _027132_, _027133_, _027134_, _027135_, _027136_, _027137_, _027138_, _027139_, _027140_, _027141_, _027142_, _027143_, _027144_, _027145_, _027146_, _027147_, _027148_, _027149_, _027150_, _027151_, _027152_, _027153_, _027154_, _027155_, _027156_, _027157_, _027158_, _027159_, _027160_, _027161_, _027162_, _027163_, _027164_, _027165_, _027166_, _027167_, _027168_, _027169_, _027170_, _027171_, _027172_, _027173_, _027174_, _027175_, _027176_, _027177_, _027178_, _027179_, _027180_, _027181_, _027182_, _027183_, _027184_, _027185_, _027186_, _027187_, _027188_, _027189_, _027190_, _027191_, _027192_, _027193_, _027194_, _027195_, _027196_, _027197_, _027198_, _027199_, _027200_, _027201_, _027202_, _027203_, _027204_, _027205_, _027206_, _027207_, _027208_, _027209_, _027210_, _027211_, _027212_, _027213_, _027214_, _027215_, _027216_, _027217_, _027218_, _027219_, _027220_, _027221_, _027222_, _027223_, _027224_, _027225_, _027226_, _027227_, _027228_, _027229_, _027230_, _027231_, _027232_, _027233_, _027234_, _027235_, _027236_, _027237_, _027238_, _027239_, _027240_, _027241_, _027242_, _027243_, _027244_, _027245_, _027246_, _027247_, _027248_, _027249_, _027250_, _027251_, _027252_, _027253_, _027254_, _027255_, _027256_, _027257_, _027258_, _027259_, _027260_, _027261_, _027262_, _027263_, _027264_, _027265_, _027266_, _027267_, _027268_, _027269_, _027270_, _027271_, _027272_, _027273_, _027274_, _027275_, _027276_, _027277_, _027278_, _027279_, _027280_, _027281_, _027282_, _027283_, _027284_, _027285_, _027286_, _027287_, _027288_, _027289_, _027290_, _027291_, _027292_, _027293_, _027294_, _027295_, _027296_, _027297_, _027298_, _027299_, _027300_, _027301_, _027302_, _027303_, _027304_, _027305_, _027306_, _027307_, _027308_, _027309_, _027310_, _027311_, _027312_, _027313_, _027314_, _027315_, _027316_, _027317_, _027318_, _027319_, _027320_, _027321_, _027322_, _027323_, _027324_, _027325_, _027326_, _027327_, _027328_, _027329_, _027330_, _027331_, _027332_, _027333_, _027334_, _027335_, _027336_, _027337_, _027338_, _027339_, _027340_, _027341_, _027342_, _027343_, _027344_, _027345_, _027346_, _027347_, _027348_, _027349_, _027350_, _027351_, _027352_, _027353_, _027354_, _027355_, _027356_, _027357_, _027358_, _027359_, _027360_, _027361_, _027362_, _027363_, _027364_, _027365_, _027366_, _027367_, _027368_, _027369_, _027370_, _027371_, _027372_, _027373_, _027374_, _027375_, _027376_, _027377_, _027378_, _027379_, _027380_, _027381_, _027382_, _027383_, _027384_, _027385_, _027386_, _027387_, _027388_, _027389_, _027390_, _027391_, _027392_, _027393_, _027394_, _027395_, _027396_, _027397_, _027398_, _027399_, _027400_, _027401_, _027402_, _027403_, _027404_, _027405_, _027406_, _027407_, _027408_, _027409_, _027410_, _027411_, _027412_, _027413_, _027414_, _027415_, _027416_, _027417_, _027418_, _027419_, _027420_, _027421_, _027422_, _027423_, _027424_, _027425_, _027426_, _027427_, _027428_, _027429_, _027430_, _027431_, _027432_, _027433_, _027434_, _027435_, _027436_, _027437_, _027438_, _027439_, _027440_, _027441_, _027442_, _027443_, _027444_, _027445_, _027446_, _027447_, _027448_, _027449_, _027450_, _027451_, _027452_, _027453_, _027454_, _027455_, _027456_, _027457_, _027458_, _027459_, _027460_, _027461_, _027462_, _027463_, _027464_, _027465_, _027466_, _027467_, _027468_, _027469_, _027470_, _027471_, _027472_, _027473_, _027474_, _027475_, _027476_, _027477_, _027478_, _027479_, _027480_, _027481_, _027482_, _027483_, _027484_, _027485_, _027486_, _027487_, _027488_, _027489_, _027490_, _027491_, _027492_, _027493_, _027494_, _027495_, _027496_, _027497_, _027498_, _027499_, _027500_, _027501_, _027502_, _027503_, _027504_, _027505_, _027506_, _027507_, _027508_, _027509_, _027510_, _027511_, _027512_, _027513_, _027514_, _027515_, _027516_, _027517_, _027518_, _027519_, _027520_, _027521_, _027522_, _027523_, _027524_, _027525_, _027526_, _027527_, _027528_, _027529_, _027530_, _027531_, _027532_, _027533_, _027534_, _027535_, _027536_, _027537_, _027538_, _027539_, _027540_, _027541_, _027542_, _027543_, _027544_, _027545_, _027546_, _027547_, _027548_, _027549_, _027550_, _027551_, _027552_, _027553_, _027554_, _027555_, _027556_, _027557_, _027558_, _027559_, _027560_, _027561_, _027562_, _027563_, _027564_, _027565_, _027566_, _027567_, _027568_, _027569_, _027570_, _027571_, _027572_, _027573_, _027574_, _027575_, _027576_, _027577_, _027578_, _027579_, _027580_, _027581_, _027582_, _027583_, _027584_, _027585_, _027586_, _027587_, _027588_, _027589_, _027590_, _027591_, _027592_, _027593_, _027594_, _027595_, _027596_, _027597_, _027598_, _027599_, _027600_, _027601_, _027602_, _027603_, _027604_, _027605_, _027606_, _027607_, _027608_, _027609_, _027610_, _027611_, _027612_, _027613_, _027614_, _027615_, _027616_, _027617_, _027618_, _027619_, _027620_, _027621_, _027622_, _027623_, _027624_, _027625_, _027626_, _027627_, _027628_, _027629_, _027630_, _027631_, _027632_, _027633_, _027634_, _027635_, _027636_, _027637_, _027638_, _027639_, _027640_, _027641_, _027642_, _027643_, _027644_, _027645_, _027646_, _027647_, _027648_, _027649_, _027650_, _027651_, _027652_, _027653_, _027654_, _027655_, _027656_, _027657_, _027658_, _027659_, _027660_, _027661_, _027662_, _027663_, _027664_, _027665_, _027666_, _027667_, _027668_, _027669_, _027670_, _027671_, _027672_, _027673_, _027674_, _027675_, _027676_, _027677_, _027678_, _027679_, _027680_, _027681_, _027682_, _027683_, _027684_, _027685_, _027686_, _027687_, _027688_, _027689_, _027690_, _027691_, _027692_, _027693_, _027694_, _027695_, _027696_, _027697_, _027698_, _027699_, _027700_, _027701_, _027702_, _027703_, _027704_, _027705_, _027706_, _027707_, _027708_, _027709_, _027710_, _027711_, _027712_, _027713_, _027714_, _027715_, _027716_, _027717_, _027718_, _027719_, _027720_, _027721_, _027722_, _027723_, _027724_, _027725_, _027726_, _027727_, _027728_, _027729_, _027730_, _027731_, _027732_, _027733_, _027734_, _027735_, _027736_, _027737_, _027738_, _027739_, _027740_, _027741_, _027742_, _027743_, _027744_, _027745_, _027746_, _027747_, _027748_, _027749_, _027750_, _027751_, _027752_, _027753_, _027754_, _027755_, _027756_, _027757_, _027758_, _027759_, _027760_, _027761_, _027762_, _027763_, _027764_, _027765_, _027766_, _027767_, _027768_, _027769_, _027770_, _027771_, _027772_, _027773_, _027774_, _027775_, _027776_, _027777_, _027778_, _027779_, _027780_, _027781_, _027782_, _027783_, _027784_, _027785_, _027786_, _027787_, _027788_, _027789_, _027790_, _027791_, _027792_, _027793_, _027794_, _027795_, _027796_, _027797_, _027798_, _027799_, _027800_, _027801_, _027802_, _027803_, _027804_, _027805_, _027806_, _027807_, _027808_, _027809_, _027810_, _027811_, _027812_, _027813_, _027814_, _027815_, _027816_, _027817_, _027818_, _027819_, _027820_, _027821_, _027822_, _027823_, _027824_, _027825_, _027826_, _027827_, _027828_, _027829_, _027830_, _027831_, _027832_, _027833_, _027834_, _027835_, _027836_, _027837_, _027838_, _027839_, _027840_, _027841_, _027842_, _027843_, _027844_, _027845_, _027846_, _027847_, _027848_, _027849_, _027850_, _027851_, _027852_, _027853_, _027854_, _027855_, _027856_, _027857_, _027858_, _027859_, _027860_, _027861_, _027862_, _027863_, _027864_, _027865_, _027866_, _027867_, _027868_, _027869_, _027870_, _027871_, _027872_, _027873_, _027874_, _027875_, _027876_, _027877_, _027878_, _027879_, _027880_, _027881_, _027882_, _027883_, _027884_, _027885_, _027886_, _027887_, _027888_, _027889_, _027890_, _027891_, _027892_, _027893_, _027894_, _027895_, _027896_, _027897_, _027898_, _027899_, _027900_, _027901_, _027902_, _027903_, _027904_, _027905_, _027906_, _027907_, _027908_, _027909_, _027910_, _027911_, _027912_, _027913_, _027914_, _027915_, _027916_, _027917_, _027918_, _027919_, _027920_, _027921_, _027922_, _027923_, _027924_, _027925_, _027926_, _027927_, _027928_, _027929_, _027930_, _027931_, _027932_, _027933_, _027934_, _027935_, _027936_, _027937_, _027938_, _027939_, _027940_, _027941_, _027942_, _027943_, _027944_, _027945_, _027946_, _027947_, _027948_, _027949_, _027950_, _027951_, _027952_, _027953_, _027954_, _027955_, _027956_, _027957_, _027958_, _027959_, _027960_, _027961_, _027962_, _027963_, _027964_, _027965_, _027966_, _027967_, _027968_, _027969_, _027970_, _027971_, _027972_, _027973_, _027974_, _027975_, _027976_, _027977_, _027978_, _027979_, _027980_, _027981_, _027982_, _027983_, _027984_, _027985_, _027986_, _027987_, _027988_, _027989_, _027990_, _027991_, _027992_, _027993_, _027994_, _027995_, _027996_, _027997_, _027998_, _027999_, _028000_, _028001_, _028002_, _028003_, _028004_, _028005_, _028006_, _028007_, _028008_, _028009_, _028010_, _028011_, _028012_, _028013_, _028014_, _028015_, _028016_, _028017_, _028018_, _028019_, _028020_, _028021_, _028022_, _028023_, _028024_, _028025_, _028026_, _028027_, _028028_, _028029_, _028030_, _028031_, _028032_, _028033_, _028034_, _028035_, _028036_, _028037_, _028038_, _028039_, _028040_, _028041_, _028042_, _028043_, _028044_, _028045_, _028046_, _028047_, _028048_, _028049_, _028050_, _028051_, _028052_, _028053_, _028054_, _028055_, _028056_, _028057_, _028058_, _028059_, _028060_, _028061_, _028062_, _028063_, _028064_, _028065_, _028066_, _028067_, _028068_, _028069_, _028070_, _028071_, _028072_, _028073_, _028074_, _028075_, _028076_, _028077_, _028078_, _028079_, _028080_, _028081_, _028082_, _028083_, _028084_, _028085_, _028086_, _028087_, _028088_, _028089_, _028090_, _028091_, _028092_, _028093_, _028094_, _028095_, _028096_, _028097_, _028098_, _028099_, _028100_, _028101_, _028102_, _028103_, _028104_, _028105_, _028106_, _028107_, _028108_, _028109_, _028110_, _028111_, _028112_, _028113_, _028114_, _028115_, _028116_, _028117_, _028118_, _028119_, _028120_, _028121_, _028122_, _028123_, _028124_, _028125_, _028126_, _028127_, _028128_, _028129_, _028130_, _028131_, _028132_, _028133_, _028134_, _028135_, _028136_, _028137_, _028138_, _028139_, _028140_, _028141_, _028142_, _028143_, _028144_, _028145_, _028146_, _028147_, _028148_, _028149_, _028150_, _028151_, _028152_, _028153_, _028154_, _028155_, _028156_, _028157_, _028158_, _028159_, _028160_, _028161_, _028162_, _028163_, _028164_, _028165_, _028166_, _028167_, _028168_, _028169_, _028170_, _028171_, _028172_, _028173_, _028174_, _028175_, _028176_, _028177_, _028178_, _028179_, _028180_, _028181_, _028182_, _028183_, _028184_, _028185_, _028186_, _028187_, _028188_, _028189_, _028190_, _028191_, _028192_, _028193_, _028194_, _028195_, _028196_, _028197_, _028198_, _028199_, _028200_, _028201_, _028202_, _028203_, _028204_, _028205_, _028206_, _028207_, _028208_, _028209_, _028210_, _028211_, _028212_, _028213_, _028214_, _028215_, _028216_, _028217_, _028218_, _028219_, _028220_, _028221_, _028222_, _028223_, _028224_, _028225_, _028226_, _028227_, _028228_, _028229_, _028230_, _028231_, _028232_, _028233_, _028234_, _028235_, _028236_, _028237_, _028238_, _028239_, _028240_, _028241_, _028242_, _028243_, _028244_, _028245_, _028246_, _028247_, _028248_, _028249_, _028250_, _028251_, _028252_, _028253_, _028254_, _028255_, _028256_, _028257_, _028258_, _028259_, _028260_, _028261_, _028262_, _028263_, _028264_, _028265_, _028266_, _028267_, _028268_, _028269_, _028270_, _028271_, _028272_, _028273_, _028274_, _028275_, _028276_, _028277_, _028278_, _028279_, _028280_, _028281_, _028282_, _028283_, _028284_, _028285_, _028286_, _028287_, _028288_, _028289_, _028290_, _028291_, _028292_, _028293_, _028294_, _028295_, _028296_, _028297_, _028298_, _028299_, _028300_, _028301_, _028302_, _028303_, _028304_, _028305_, _028306_, _028307_, _028308_, _028309_, _028310_, _028311_, _028312_, _028313_, _028314_, _028315_, _028316_, _028317_, _028318_, _028319_, _028320_, _028321_, _028322_, _028323_, _028324_, _028325_, _028326_, _028327_, _028328_, _028329_, _028330_, _028331_, _028332_, _028333_, _028334_, _028335_, _028336_, _028337_, _028338_, _028339_, _028340_, _028341_, _028342_, _028343_, _028344_, _028345_, _028346_, _028347_, _028348_, _028349_, _028350_, _028351_, _028352_, _028353_, _028354_, _028355_, _028356_, _028357_, _028358_, _028359_, _028360_, _028361_, _028362_, _028363_, _028364_, _028365_, _028366_, _028367_, _028368_, _028369_, _028370_, _028371_, _028372_, _028373_, _028374_, _028375_, _028376_, _028377_, _028378_, _028379_, _028380_, _028381_, _028382_, _028383_, _028384_, _028385_, _028386_, _028387_, _028388_, _028389_, _028390_, _028391_, _028392_, _028393_, _028394_, _028395_, _028396_, _028397_, _028398_, _028399_, _028400_, _028401_, _028402_, _028403_, _028404_, _028405_, _028406_, _028407_, _028408_, _028409_, _028410_, _028411_, _028412_, _028413_, _028414_, _028415_, _028416_, _028417_, _028418_, _028419_, _028420_, _028421_, _028422_, _028423_, _028424_, _028425_, _028426_, _028427_, _028428_, _028429_, _028430_, _028431_, _028432_, _028433_, _028434_, _028435_, _028436_, _028437_, _028438_, _028439_, _028440_, _028441_, _028442_, _028443_, _028444_, _028445_, _028446_, _028447_, _028448_, _028449_, _028450_, _028451_, _028452_, _028453_, _028454_, _028455_, _028456_, _028457_, _028458_, _028459_, _028460_, _028461_, _028462_, _028463_, _028464_, _028465_, _028466_, _028467_, _028468_, _028469_, _028470_, _028471_, _028472_, _028473_, _028474_, _028475_, _028476_, _028477_, _028478_, _028479_, _028480_, _028481_, _028482_, _028483_, _028484_, _028485_, _028486_, _028487_, _028488_, _028489_, _028490_, _028491_, _028492_, _028493_, _028494_, _028495_, _028496_, _028497_, _028498_, _028499_, _028500_, _028501_, _028502_, _028503_, _028504_, _028505_, _028506_, _028507_, _028508_, _028509_, _028510_, _028511_, _028512_, _028513_, _028514_, _028515_, _028516_, _028517_, _028518_, _028519_, _028520_, _028521_, _028522_, _028523_, _028524_, _028525_, _028526_, _028527_, _028528_, _028529_, _028530_, _028531_, _028532_, _028533_, _028534_, _028535_, _028536_, _028537_, _028538_, _028539_, _028540_, _028541_, _028542_, _028543_, _028544_, _028545_, _028546_, _028547_, _028548_, _028549_, _028550_, _028551_, _028552_, _028553_, _028554_, _028555_, _028556_, _028557_, _028558_, _028559_, _028560_, _028561_, _028562_, _028563_, _028564_, _028565_, _028566_, _028567_, _028568_, _028569_, _028570_, _028571_, _028572_, _028573_, _028574_, _028575_, _028576_, _028577_, _028578_, _028579_, _028580_, _028581_, _028582_, _028583_, _028584_, _028585_, _028586_, _028587_, _028588_, _028589_, _028590_, _028591_, _028592_, _028593_, _028594_, _028595_, _028596_, _028597_, _028598_, _028599_, _028600_, _028601_, _028602_, _028603_, _028604_, _028605_, _028606_, _028607_, _028608_, _028609_, _028610_, _028611_, _028612_, _028613_, _028614_, _028615_, _028616_, _028617_, _028618_, _028619_, _028620_, _028621_, _028622_, _028623_, _028624_, _028625_, _028626_, _028627_, _028628_, _028629_, _028630_, _028631_, _028632_, _028633_, _028634_, _028635_, _028636_, _028637_, _028638_, _028639_, _028640_, _028641_, _028642_, _028643_, _028644_, _028645_, _028646_, _028647_, _028648_, _028649_, _028650_, _028651_, _028652_, _028653_, _028654_, _028655_, _028656_, _028657_, _028658_, _028659_, _028660_, _028661_, _028662_, _028663_, _028664_, _028665_, _028666_, _028667_, _028668_, _028669_, _028670_, _028671_, _028672_, _028673_, _028674_, _028675_, _028676_, _028677_, _028678_, _028679_, _028680_, _028681_, _028682_, _028683_, _028684_, _028685_, _028686_, _028687_, _028688_, _028689_, _028690_, _028691_, _028692_, _028693_, _028694_, _028695_, _028696_, _028697_, _028698_, _028699_, _028700_, _028701_, _028702_, _028703_, _028704_, _028705_, _028706_, _028707_, _028708_, _028709_, _028710_, _028711_, _028712_, _028713_, _028714_, _028715_, _028716_, _028717_, _028718_, _028719_, _028720_, _028721_, _028722_, _028723_, _028724_, _028725_, _028726_, _028727_, _028728_, _028729_, _028730_, _028731_, _028732_, _028733_, _028734_, _028735_, _028736_, _028737_, _028738_, _028739_, _028740_, _028741_, _028742_, _028743_, _028744_, _028745_, _028746_, _028747_, _028748_, _028749_, _028750_, _028751_, _028752_, _028753_, _028754_, _028755_, _028756_, _028757_, _028758_, _028759_, _028760_, _028761_, _028762_, _028763_, _028764_, _028765_, _028766_, _028767_, _028768_, _028769_, _028770_, _028771_, _028772_, _028773_, _028774_, _028775_, _028776_, _028777_, _028778_, _028779_, _028780_, _028781_, _028782_, _028783_, _028784_, _028785_, _028786_, _028787_, _028788_, _028789_, _028790_, _028791_, _028792_, _028793_, _028794_, _028795_, _028796_, _028797_, _028798_, _028799_, _028800_, _028801_, _028802_, _028803_, _028804_, _028805_, _028806_, _028807_, _028808_, _028809_, _028810_, _028811_, _028812_, _028813_, _028814_, _028815_, _028816_, _028817_, _028818_, _028819_, _028820_, _028821_, _028822_, _028823_, _028824_, _028825_, _028826_, _028827_, _028828_, _028829_, _028830_, _028831_, _028832_, _028833_, _028834_, _028835_, _028836_, _028837_, _028838_, _028839_, _028840_, _028841_, _028842_, _028843_, _028844_, _028845_, _028846_, _028847_, _028848_, _028849_, _028850_, _028851_, _028852_, _028853_, _028854_, _028855_, _028856_, _028857_, _028858_, _028859_, _028860_, _028861_, _028862_, _028863_, _028864_, _028865_, _028866_, _028867_, _028868_, _028869_, _028870_, _028871_, _028872_, _028873_, _028874_, _028875_, _028876_, _028877_, _028878_, _028879_, _028880_, _028881_, _028882_, _028883_, _028884_, _028885_, _028886_, _028887_, _028888_, _028889_, _028890_, _028891_, _028892_, _028893_, _028894_, _028895_, _028896_, _028897_, _028898_, _028899_, _028900_, _028901_, _028902_, _028903_, _028904_, _028905_, _028906_, _028907_, _028908_, _028909_, _028910_, _028911_, _028912_, _028913_, _028914_, _028915_, _028916_, _028917_, _028918_, _028919_, _028920_, _028921_, _028922_, _028923_, _028924_, _028925_, _028926_, _028927_, _028928_, _028929_, _028930_, _028931_, _028932_, _028933_, _028934_, _028935_, _028936_, _028937_, _028938_, _028939_, _028940_, _028941_, _028942_, _028943_, _028944_, _028945_, _028946_, _028947_, _028948_, _028949_, _028950_, _028951_, _028952_, _028953_, _028954_, _028955_, _028956_, _028957_, _028958_, _028959_, _028960_, _028961_, _028962_, _028963_, _028964_, _028965_, _028966_, _028967_, _028968_, _028969_, _028970_, _028971_, _028972_, _028973_, _028974_, _028975_, _028976_, _028977_, _028978_, _028979_, _028980_, _028981_, _028982_, _028983_, _028984_, _028985_, _028986_, _028987_, _028988_, _028989_, _028990_, _028991_, _028992_, _028993_, _028994_, _028995_, _028996_, _028997_, _028998_, _028999_, _029000_, _029001_, _029002_, _029003_, _029004_, _029005_, _029006_, _029007_, _029008_, _029009_, _029010_, _029011_, _029012_, _029013_, _029014_, _029015_, _029016_, _029017_, _029018_, _029019_, _029020_, _029021_, _029022_, _029023_, _029024_, _029025_, _029026_, _029027_, _029028_, _029029_, _029030_, _029031_, _029032_, _029033_, _029034_, _029035_, _029036_, _029037_, _029038_, _029039_, _029040_, _029041_, _029042_, _029043_, _029044_, _029045_, _029046_, _029047_, _029048_, _029049_, _029050_, _029051_, _029052_, _029053_, _029054_, _029055_, _029056_, _029057_, _029058_, _029059_, _029060_, _029061_, _029062_, _029063_, _029064_, _029065_, _029066_, _029067_, _029068_, _029069_, _029070_, _029071_, _029072_, _029073_, _029074_, _029075_, _029076_, _029077_, _029078_, _029079_, _029080_, _029081_, _029082_, _029083_, _029084_, _029085_, _029086_, _029087_, _029088_, _029089_, _029090_, _029091_, _029092_, _029093_, _029094_, _029095_, _029096_, _029097_, _029098_, _029099_, _029100_, _029101_, _029102_, _029103_, _029104_, _029105_, _029106_, _029107_, _029108_, _029109_, _029110_, _029111_, _029112_, _029113_, _029114_, _029115_, _029116_, _029117_, _029118_, _029119_, _029120_, _029121_, _029122_, _029123_, _029124_, _029125_, _029126_, _029127_, _029128_, _029129_, _029130_, _029131_, _029132_, _029133_, _029134_, _029135_, _029136_, _029137_, _029138_, _029139_, _029140_, _029141_, _029142_, _029143_, _029144_, _029145_, _029146_, _029147_, _029148_, _029149_, _029150_, _029151_, _029152_, _029153_, _029154_, _029155_, _029156_, _029157_, _029158_, _029159_, _029160_, _029161_, _029162_, _029163_, _029164_, _029165_, _029166_, _029167_, _029168_, _029169_, _029170_, _029171_, _029172_, _029173_, _029174_, _029175_, _029176_, _029177_, _029178_, _029179_, _029180_, _029181_, _029182_, _029183_, _029184_, _029185_, _029186_, _029187_, _029188_, _029189_, _029190_, _029191_, _029192_, _029193_, _029194_, _029195_, _029196_, _029197_, _029198_, _029199_, _029200_, _029201_, _029202_, _029203_, _029204_, _029205_, _029206_, _029207_, _029208_, _029209_, _029210_, _029211_, _029212_, _029213_, _029214_, _029215_, _029216_, _029217_, _029218_, _029219_, _029220_, _029221_, _029222_, _029223_, _029224_, _029225_, _029226_, _029227_, _029228_, _029229_, _029230_, _029231_, _029232_, _029233_, _029234_, _029235_, _029236_, _029237_, _029238_, _029239_, _029240_, _029241_, _029242_, _029243_, _029244_, _029245_, _029246_, _029247_, _029248_, _029249_, _029250_, _029251_, _029252_, _029253_, _029254_, _029255_, _029256_, _029257_, _029258_, _029259_, _029260_, _029261_, _029262_, _029263_, _029264_, _029265_, _029266_, _029267_, _029268_, _029269_, _029270_, _029271_, _029272_, _029273_, _029274_, _029275_, _029276_, _029277_, _029278_, _029279_, _029280_, _029281_, _029282_, _029283_, _029284_, _029285_, _029286_, _029287_, _029288_, _029289_, _029290_, _029291_, _029292_, _029293_, _029294_, _029295_, _029296_, _029297_, _029298_, _029299_, _029300_, _029301_, _029302_, _029303_, _029304_, _029305_, _029306_, _029307_, _029308_, _029309_, _029310_, _029311_, _029312_, _029313_, _029314_, _029315_, _029316_, _029317_, _029318_, _029319_, _029320_, _029321_, _029322_, _029323_, _029324_, _029325_, _029326_, _029327_, _029328_, _029329_, _029330_, _029331_, _029332_, _029333_, _029334_, _029335_, _029336_, _029337_, _029338_, _029339_, _029340_, _029341_, _029342_, _029343_, _029344_, _029345_, _029346_, _029347_, _029348_, _029349_, _029350_, _029351_, _029352_, _029353_, _029354_, _029355_, _029356_, _029357_, _029358_, _029359_, _029360_, _029361_, _029362_, _029363_, _029364_, _029365_, _029366_, _029367_, _029368_, _029369_, _029370_, _029371_, _029372_, _029373_, _029374_, _029375_, _029376_, _029377_, _029378_, _029379_, _029380_, _029381_, _029382_, _029383_, _029384_, _029385_, _029386_, _029387_, _029388_, _029389_, _029390_, _029391_, _029392_, _029393_, _029394_, _029395_, _029396_, _029397_, _029398_, _029399_, _029400_, _029401_, _029402_, _029403_, _029404_, _029405_, _029406_, _029407_, _029408_, _029409_, _029410_, _029411_, _029412_, _029413_, _029414_, _029415_, _029416_, _029417_, _029418_, _029419_, _029420_, _029421_, _029422_, _029423_, _029424_, _029425_, _029426_, _029427_, _029428_, _029429_, _029430_, _029431_, _029432_, _029433_, _029434_, _029435_, _029436_, _029437_, _029438_, _029439_, _029440_, _029441_, _029442_, _029443_, _029444_, _029445_, _029446_, _029447_, _029448_, _029449_, _029450_, _029451_, _029452_, _029453_, _029454_, _029455_, _029456_, _029457_, _029458_, _029459_, _029460_, _029461_, _029462_, _029463_, _029464_, _029465_, _029466_, _029467_, _029468_, _029469_, _029470_, _029471_, _029472_, _029473_, _029474_, _029475_, _029476_, _029477_, _029478_, _029479_, _029480_, _029481_, _029482_, _029483_, _029484_, _029485_, _029486_, _029487_, _029488_, _029489_, _029490_, _029491_, _029492_, _029493_, _029494_, _029495_, _029496_, _029497_, _029498_, _029499_, _029500_, _029501_, _029502_, _029503_, _029504_, _029505_, _029506_, _029507_, _029508_, _029509_, _029510_, _029511_, _029512_, _029513_, _029514_, _029515_, _029516_, _029517_, _029518_, _029519_, _029520_, _029521_, _029522_, _029523_, _029524_, _029525_, _029526_, _029527_, _029528_, _029529_, _029530_, _029531_, _029532_, _029533_, _029534_, _029535_, _029536_, _029537_, _029538_, _029539_, _029540_, _029541_, _029542_, _029543_, _029544_, _029545_, _029546_, _029547_, _029548_, _029549_, _029550_, _029551_, _029552_, _029553_, _029554_, _029555_, _029556_, _029557_, _029558_, _029559_, _029560_, _029561_, _029562_, _029563_, _029564_, _029565_, _029566_, _029567_, _029568_, _029569_, _029570_, _029571_, _029572_, _029573_, _029574_, _029575_, _029576_, _029577_, _029578_, _029579_, _029580_, _029581_, _029582_, _029583_, _029584_, _029585_, _029586_, _029587_, _029588_, _029589_, _029590_, _029591_, _029592_, _029593_, _029594_, _029595_, _029596_, _029597_, _029598_, _029599_, _029600_, _029601_, _029602_, _029603_, _029604_, _029605_, _029606_, _029607_, _029608_, _029609_, _029610_, _029611_, _029612_, _029613_, _029614_, _029615_, _029616_, _029617_, _029618_, _029619_, _029620_, _029621_, _029622_, _029623_, _029624_, _029625_, _029626_, _029627_, _029628_, _029629_, _029630_, _029631_, _029632_, _029633_, _029634_, _029635_, _029636_, _029637_, _029638_, _029639_, _029640_, _029641_, _029642_, _029643_, _029644_, _029645_, _029646_, _029647_, _029648_, _029649_, _029650_, _029651_, _029652_, _029653_, _029654_, _029655_, _029656_, _029657_, _029658_, _029659_, _029660_, _029661_, _029662_, _029663_, _029664_, _029665_, _029666_, _029667_, _029668_, _029669_, _029670_, _029671_, _029672_, _029673_, _029674_, _029675_, _029676_, _029677_, _029678_, _029679_, _029680_, _029681_, _029682_, _029683_, _029684_, _029685_, _029686_, _029687_, _029688_, _029689_, _029690_, _029691_, _029692_, _029693_, _029694_, _029695_, _029696_, _029697_, _029698_, _029699_, _029700_, _029701_, _029702_, _029703_, _029704_, _029705_, _029706_, _029707_, _029708_, _029709_, _029710_, _029711_, _029712_, _029713_, _029714_, _029715_, _029716_, _029717_, _029718_, _029719_, _029720_, _029721_, _029722_, _029723_, _029724_, _029725_, _029726_, _029727_, _029728_, _029729_, _029730_, _029731_, _029732_, _029733_, _029734_, _029735_, _029736_, _029737_, _029738_, _029739_, _029740_, _029741_, _029742_, _029743_, _029744_, _029745_, _029746_, _029747_, _029748_, _029749_, _029750_, _029751_, _029752_, _029753_, _029754_, _029755_, _029756_, _029757_, _029758_, _029759_, _029760_, _029761_, _029762_, _029763_, _029764_, _029765_, _029766_, _029767_, _029768_, _029769_, _029770_, _029771_, _029772_, _029773_, _029774_, _029775_, _029776_, _029777_, _029778_, _029779_, _029780_, _029781_, _029782_, _029783_, _029784_, _029785_, _029786_, _029787_, _029788_, _029789_, _029790_, _029791_, _029792_, _029793_, _029794_, _029795_, _029796_, _029797_, _029798_, _029799_, _029800_, _029801_, _029802_, _029803_, _029804_, _029805_, _029806_, _029807_, _029808_, _029809_, _029810_, _029811_, _029812_, _029813_, _029814_, _029815_, _029816_, _029817_, _029818_, _029819_, _029820_, _029821_, _029822_, _029823_, _029824_, _029825_, _029826_, _029827_, _029828_, _029829_, _029830_, _029831_, _029832_, _029833_, _029834_, _029835_, _029836_, _029837_, _029838_, _029839_, _029840_, _029841_, _029842_, _029843_, _029844_, _029845_, _029846_, _029847_, _029848_, _029849_, _029850_, _029851_, _029852_, _029853_, _029854_, _029855_, _029856_, _029857_, _029858_, _029859_, _029860_, _029861_, _029862_, _029863_, _029864_, _029865_, _029866_, _029867_, _029868_, _029869_, _029870_, _029871_, _029872_, _029873_, _029874_, _029875_, _029876_, _029877_, _029878_, _029879_, _029880_, _029881_, _029882_, _029883_, _029884_, _029885_, _029886_, _029887_, _029888_, _029889_, _029890_, _029891_, _029892_, _029893_, _029894_, _029895_, _029896_, _029897_, _029898_, _029899_, _029900_, _029901_, _029902_, _029903_, _029904_, _029905_, _029906_, _029907_, _029908_, _029909_, _029910_, _029911_, _029912_, _029913_, _029914_, _029915_, _029916_, _029917_, _029918_, _029919_, _029920_, _029921_, _029922_, _029923_, _029924_, _029925_, _029926_, _029927_, _029928_, _029929_, _029930_, _029931_, _029932_, _029933_, _029934_, _029935_, _029936_, _029937_, _029938_, _029939_, _029940_, _029941_, _029942_, _029943_, _029944_, _029945_, _029946_, _029947_, _029948_, _029949_, _029950_, _029951_, _029952_, _029953_, _029954_, _029955_, _029956_, _029957_, _029958_, _029959_, _029960_, _029961_, _029962_, _029963_, _029964_, _029965_, _029966_, _029967_, _029968_, _029969_, _029970_, _029971_, _029972_, _029973_, _029974_, _029975_, _029976_, _029977_, _029978_, _029979_, _029980_, _029981_, _029982_, _029983_, _029984_, _029985_, _029986_, _029987_, _029988_, _029989_, _029990_, _029991_, _029992_, _029993_, _029994_, _029995_, _029996_, _029997_, _029998_, _029999_, _030000_, _030001_, _030002_, _030003_, _030004_, _030005_, _030006_, _030007_, _030008_, _030009_, _030010_, _030011_, _030012_, _030013_, _030014_, _030015_, _030016_, _030017_, _030018_, _030019_, _030020_, _030021_, _030022_, _030023_, _030024_, _030025_, _030026_, _030027_, _030028_, _030029_, _030030_, _030031_, _030032_, _030033_, _030034_, _030035_, _030036_, _030037_, _030038_, _030039_, _030040_, _030041_, _030042_, _030043_, _030044_, _030045_, _030046_, _030047_, _030048_, _030049_, _030050_, _030051_, _030052_, _030053_, _030054_, _030055_, _030056_, _030057_, _030058_, _030059_, _030060_, _030061_, _030062_, _030063_, _030064_, _030065_, _030066_, _030067_, _030068_, _030069_, _030070_, _030071_, _030072_, _030073_, _030074_, _030075_, _030076_, _030077_, _030078_, _030079_, _030080_, _030081_, _030082_, _030083_, _030084_, _030085_, _030086_, _030087_, _030088_, _030089_, _030090_, _030091_, _030092_, _030093_, _030094_, _030095_, _030096_, _030097_, _030098_, _030099_, _030100_, _030101_, _030102_, _030103_, _030104_, _030105_, _030106_, _030107_, _030108_, _030109_, _030110_, _030111_, _030112_, _030113_, _030114_, _030115_, _030116_, _030117_, _030118_, _030119_, _030120_, _030121_, _030122_, _030123_, _030124_, _030125_, _030126_, _030127_, _030128_, _030129_, _030130_, _030131_, _030132_, _030133_, _030134_, _030135_, _030136_, _030137_, _030138_, _030139_, _030140_, _030141_, _030142_, _030143_, _030144_, _030145_, _030146_, _030147_, _030148_, _030149_, _030150_, _030151_, _030152_, _030153_, _030154_, _030155_, _030156_, _030157_, _030158_, _030159_, _030160_, _030161_, _030162_, _030163_, _030164_, _030165_, _030166_, _030167_, _030168_, _030169_, _030170_, _030171_, _030172_, _030173_, _030174_, _030175_, _030176_, _030177_, _030178_, _030179_, _030180_, _030181_, _030182_, _030183_, _030184_, _030185_, _030186_, _030187_, _030188_, _030189_, _030190_, _030191_, _030192_, _030193_, _030194_, _030195_, _030196_, _030197_, _030198_, _030199_, _030200_, _030201_, _030202_, _030203_, _030204_, _030205_, _030206_, _030207_, _030208_, _030209_, _030210_, _030211_, _030212_, _030213_, _030214_, _030215_, _030216_, _030217_, _030218_, _030219_, _030220_, _030221_, _030222_, _030223_, _030224_, _030225_, _030226_, _030227_, _030228_, _030229_, _030230_, _030231_, _030232_, _030233_, _030234_, _030235_, _030236_, _030237_, _030238_, _030239_, _030240_, _030241_, _030242_, _030243_, _030244_, _030245_, _030246_, _030247_, _030248_, _030249_, _030250_, _030251_, _030252_, _030253_, _030254_, _030255_, _030256_, _030257_, _030258_, _030259_, _030260_, _030261_, _030262_, _030263_, _030264_, _030265_, _030266_, _030267_, _030268_, _030269_, _030270_, _030271_, _030272_, _030273_, _030274_, _030275_, _030276_, _030277_, _030278_, _030279_, _030280_, _030281_, _030282_, _030283_, _030284_, _030285_, _030286_, _030287_, _030288_, _030289_, _030290_, _030291_, _030292_, _030293_, _030294_, _030295_, _030296_, _030297_, _030298_, _030299_, _030300_, _030301_, _030302_, _030303_, _030304_, _030305_, _030306_, _030307_, _030308_, _030309_, _030310_, _030311_, _030312_, _030313_, _030314_, _030315_, _030316_, _030317_, _030318_, _030319_, _030320_, _030321_, _030322_, _030323_, _030324_, _030325_, _030326_, _030327_, _030328_, _030329_, _030330_, _030331_, _030332_, _030333_, _030334_, _030335_, _030336_, _030337_, _030338_, _030339_, _030340_, _030341_, _030342_, _030343_, _030344_, _030345_, _030346_, _030347_, _030348_, _030349_, _030350_, _030351_, _030352_, _030353_, _030354_, _030355_, _030356_, _030357_, _030358_, _030359_, _030360_, _030361_, _030362_, _030363_, _030364_, _030365_, _030366_, _030367_, _030368_, _030369_, _030370_, _030371_, _030372_, _030373_, _030374_, _030375_, _030376_, _030377_, _030378_, _030379_, _030380_, _030381_, _030382_, _030383_, _030384_, _030385_, _030386_, _030387_, _030388_, _030389_, _030390_, _030391_, _030392_, _030393_, _030394_, _030395_, _030396_, _030397_, _030398_, _030399_, _030400_, _030401_, _030402_, _030403_, _030404_, _030405_, _030406_, _030407_, _030408_, _030409_, _030410_, _030411_, _030412_, _030413_, _030414_, _030415_, _030416_, _030417_, _030418_, _030419_, _030420_, _030421_, _030422_, _030423_, _030424_, _030425_, _030426_, _030427_, _030428_, _030429_, _030430_, _030431_, _030432_, _030433_, _030434_, _030435_, _030436_, _030437_, _030438_, _030439_, _030440_, _030441_, _030442_, _030443_, _030444_, _030445_, _030446_, _030447_, _030448_, _030449_, _030450_, _030451_, _030452_, _030453_, _030454_, _030455_, _030456_, _030457_, _030458_, _030459_, _030460_, _030461_, _030462_, _030463_, _030464_, _030465_, _030466_, _030467_, _030468_, _030469_, _030470_, _030471_, _030472_, _030473_, _030474_, _030475_, _030476_, _030477_, _030478_, _030479_, _030480_, _030481_, _030482_, _030483_, _030484_, _030485_, _030486_, _030487_, _030488_, _030489_, _030490_, _030491_, _030492_, _030493_, _030494_, _030495_, _030496_, _030497_, _030498_, _030499_, _030500_, _030501_, _030502_, _030503_, _030504_, _030505_, _030506_, _030507_, _030508_, _030509_, _030510_, _030511_, _030512_, _030513_, _030514_, _030515_, _030516_, _030517_, _030518_, _030519_, _030520_, _030521_, _030522_, _030523_, _030524_, _030525_, _030526_, _030527_, _030528_, _030529_, _030530_, _030531_, _030532_, _030533_, _030534_, _030535_, _030536_, _030537_, _030538_, _030539_, _030540_, _030541_, _030542_, _030543_, _030544_, _030545_, _030546_, _030547_, _030548_, _030549_, _030550_, _030551_, _030552_, _030553_, _030554_, _030555_, _030556_, _030557_, _030558_, _030559_, _030560_, _030561_, _030562_, _030563_, _030564_, _030565_, _030566_, _030567_, _030568_, _030569_, _030570_, _030571_, _030572_, _030573_, _030574_, _030575_, _030576_, _030577_, _030578_, _030579_, _030580_, _030581_, _030582_, _030583_, _030584_, _030585_, _030586_, _030587_, _030588_, _030589_, _030590_, _030591_, _030592_, _030593_, _030594_, _030595_, _030596_, _030597_, _030598_, _030599_, _030600_, _030601_, _030602_, _030603_, _030604_, _030605_, _030606_, _030607_, _030608_, _030609_, _030610_, _030611_, _030612_, _030613_, _030614_, _030615_, _030616_, _030617_, _030618_, _030619_, _030620_, _030621_, _030622_, _030623_, _030624_, _030625_, _030626_, _030627_, _030628_, _030629_, _030630_, _030631_, _030632_, _030633_, _030634_, _030635_, _030636_, _030637_, _030638_, _030639_, _030640_, _030641_, _030642_, _030643_, _030644_, _030645_, _030646_, _030647_, _030648_, _030649_, _030650_, _030651_, _030652_, _030653_, _030654_, _030655_, _030656_, _030657_, _030658_, _030659_, _030660_, _030661_, _030662_, _030663_, _030664_, _030665_, _030666_, _030667_, _030668_, _030669_, _030670_, _030671_, _030672_, _030673_, _030674_, _030675_, _030676_, _030677_, _030678_, _030679_, _030680_, _030681_, _030682_, _030683_, _030684_, _030685_, _030686_, _030687_, _030688_, _030689_, _030690_, _030691_, _030692_, _030693_, _030694_, _030695_, _030696_, _030697_, _030698_, _030699_, _030700_, _030701_, _030702_, _030703_, _030704_, _030705_, _030706_, _030707_, _030708_, _030709_, _030710_, _030711_, _030712_, _030713_, _030714_, _030715_, _030716_, _030717_, _030718_, _030719_, _030720_, _030721_, _030722_, _030723_, _030724_, _030725_, _030726_, _030727_, _030728_, _030729_, _030730_, _030731_, _030732_, _030733_, _030734_, _030735_, _030736_, _030737_, _030738_, _030739_, _030740_, _030741_, _030742_, _030743_, _030744_, _030745_, _030746_, _030747_, _030748_, _030749_, _030750_, _030751_, _030752_, _030753_, _030754_, _030755_, _030756_, _030757_, _030758_, _030759_, _030760_, _030761_, _030762_, _030763_, _030764_, _030765_, _030766_, _030767_, _030768_, _030769_, _030770_, _030771_, _030772_, _030773_, _030774_, _030775_, _030776_, _030777_, _030778_, _030779_, _030780_, _030781_, _030782_, _030783_, _030784_, _030785_, _030786_, _030787_, _030788_, _030789_, _030790_, _030791_, _030792_, _030793_, _030794_, _030795_, _030796_, _030797_, _030798_, _030799_, _030800_, _030801_, _030802_, _030803_, _030804_, _030805_, _030806_, _030807_, _030808_, _030809_, _030810_, _030811_, _030812_, _030813_, _030814_, _030815_, _030816_, _030817_, _030818_, _030819_, _030820_, _030821_, _030822_, _030823_, _030824_, _030825_, _030826_, _030827_, _030828_, _030829_, _030830_, _030831_, _030832_, _030833_, _030834_, _030835_, _030836_, _030837_, _030838_, _030839_, _030840_, _030841_, _030842_, _030843_, _030844_, _030845_, _030846_, _030847_, _030848_, _030849_, _030850_, _030851_, _030852_, _030853_, _030854_, _030855_, _030856_, _030857_, _030858_, _030859_, _030860_, _030861_, _030862_, _030863_, _030864_, _030865_, _030866_, _030867_, _030868_, _030869_, _030870_, _030871_, _030872_, _030873_, _030874_, _030875_, _030876_, _030877_, _030878_, _030879_, _030880_, _030881_, _030882_, _030883_, _030884_, _030885_, _030886_, _030887_, _030888_, _030889_, _030890_, _030891_, _030892_, _030893_, _030894_, _030895_, _030896_, _030897_, _030898_, _030899_, _030900_, _030901_, _030902_, _030903_, _030904_, _030905_, _030906_, _030907_, _030908_, _030909_, _030910_, _030911_, _030912_, _030913_, _030914_, _030915_, _030916_, _030917_, _030918_, _030919_, _030920_, _030921_, _030922_, _030923_, _030924_, _030925_, _030926_, _030927_, _030928_, _030929_, _030930_, _030931_, _030932_, _030933_, _030934_, _030935_, _030936_, _030937_, _030938_, _030939_, _030940_, _030941_, _030942_, _030943_, _030944_, _030945_, _030946_, _030947_, _030948_, _030949_, _030950_, _030951_, _030952_, _030953_, _030954_, _030955_, _030956_, _030957_, _030958_, _030959_, _030960_, _030961_, _030962_, _030963_, _030964_, _030965_, _030966_, _030967_, _030968_, _030969_, _030970_, _030971_, _030972_, _030973_, _030974_, _030975_, _030976_, _030977_, _030978_, _030979_, _030980_, _030981_, _030982_, _030983_, _030984_, _030985_, _030986_, _030987_, _030988_, _030989_, _030990_, _030991_, _030992_, _030993_, _030994_, _030995_, _030996_, _030997_, _030998_, _030999_, _031000_, _031001_, _031002_, _031003_, _031004_, _031005_, _031006_, _031007_, _031008_, _031009_, _031010_, _031011_, _031012_, _031013_, _031014_, _031015_, _031016_, _031017_, _031018_, _031019_, _031020_, _031021_, _031022_, _031023_, _031024_, _031025_, _031026_, _031027_, _031028_, _031029_, _031030_, _031031_, _031032_, _031033_, _031034_, _031035_, _031036_, _031037_, _031038_, _031039_, _031040_, _031041_, _031042_, _031043_, _031044_, _031045_, _031046_, _031047_, _031048_, _031049_, _031050_, _031051_, _031052_, _031053_, _031054_, _031055_, _031056_, _031057_, _031058_, _031059_, _031060_, _031061_, _031062_, _031063_, _031064_, _031065_, _031066_, _031067_, _031068_, _031069_, _031070_, _031071_, _031072_, _031073_, _031074_, _031075_, _031076_, _031077_, _031078_, _031079_, _031080_, _031081_, _031082_, _031083_, _031084_, _031085_, _031086_, _031087_, _031088_, _031089_, _031090_, _031091_, _031092_, _031093_, _031094_, _031095_, _031096_, _031097_, _031098_, _031099_, _031100_, _031101_, _031102_, _031103_, _031104_, _031105_, _031106_, _031107_, _031108_, _031109_, _031110_, _031111_, _031112_, _031113_, _031114_, _031115_, _031116_, _031117_, _031118_, _031119_, _031120_, _031121_, _031122_, _031123_, _031124_, _031125_, _031126_, _031127_, _031128_, _031129_, _031130_, _031131_, _031132_, _031133_, _031134_, _031135_, _031136_, _031137_, _031138_, _031139_, _031140_, _031141_, _031142_, _031143_, _031144_, _031145_, _031146_, _031147_, _031148_, _031149_, _031150_, _031151_, _031152_, _031153_, _031154_, _031155_, _031156_, _031157_, _031158_, _031159_, _031160_, _031161_, _031162_, _031163_, _031164_, _031165_, _031166_, _031167_, _031168_, _031169_, _031170_, _031171_, _031172_, _031173_, _031174_, _031175_, _031176_, _031177_, _031178_, _031179_, _031180_, _031181_, _031182_, _031183_, _031184_, _031185_, _031186_, _031187_, _031188_, _031189_, _031190_, _031191_, _031192_, _031193_, _031194_, _031195_, _031196_, _031197_, _031198_, _031199_, _031200_, _031201_, _031202_, _031203_, _031204_, _031205_, _031206_, _031207_, _031208_, _031209_, _031210_, _031211_, _031212_, _031213_, _031214_, _031215_, _031216_, _031217_, _031218_, _031219_, _031220_, _031221_, _031222_, _031223_, _031224_, _031225_, _031226_, _031227_, _031228_, _031229_, _031230_, _031231_, _031232_, _031233_, _031234_, _031235_, _031236_, _031237_, _031238_, _031239_, _031240_, _031241_, _031242_, _031243_, _031244_, _031245_, _031246_, _031247_, _031248_, _031249_, _031250_, _031251_, _031252_, _031253_, _031254_, _031255_, _031256_, _031257_, _031258_, _031259_, _031260_, _031261_, _031262_, _031263_, _031264_, _031265_, _031266_, _031267_, _031268_, _031269_, _031270_, _031271_, _031272_, _031273_, _031274_, _031275_, _031276_, _031277_, _031278_, _031279_, _031280_, _031281_, _031282_, _031283_, _031284_, _031285_, _031286_, _031287_, _031288_, _031289_, _031290_, _031291_, _031292_, _031293_, _031294_, _031295_, _031296_, _031297_, _031298_, _031299_, _031300_, _031301_, _031302_, _031303_, _031304_, _031305_, _031306_, _031307_, _031308_, _031309_, _031310_, _031311_, _031312_, _031313_, _031314_, _031315_, _031316_, _031317_, _031318_, _031319_, _031320_, _031321_, _031322_, _031323_, _031324_, _031325_, _031326_, _031327_, _031328_, _031329_, _031330_, _031331_, _031332_, _031333_, _031334_, _031335_, _031336_, _031337_, _031338_, _031339_, _031340_, _031341_, _031342_, _031343_, _031344_, _031345_, _031346_, _031347_, _031348_, _031349_, _031350_, _031351_, _031352_, _031353_, _031354_, _031355_, _031356_, _031357_, _031358_, _031359_, _031360_, _031361_, _031362_, _031363_, _031364_, _031365_, _031366_, _031367_, _031368_, _031369_, _031370_, _031371_, _031372_, _031373_, _031374_, _031375_, _031376_, _031377_, _031378_, _031379_, _031380_, _031381_, _031382_, _031383_, _031384_, _031385_, _031386_, _031387_, _031388_, _031389_, _031390_, _031391_, _031392_, _031393_, _031394_, _031395_, _031396_, _031397_, _031398_, _031399_, _031400_, _031401_, _031402_, _031403_, _031404_, _031405_, _031406_, _031407_, _031408_, _031409_, _031410_, _031411_, _031412_, _031413_, _031414_, _031415_, _031416_, _031417_, _031418_, _031419_, _031420_, _031421_, _031422_, _031423_, _031424_, _031425_, _031426_, _031427_, _031428_, _031429_, _031430_, _031431_, _031432_, _031433_, _031434_, _031435_, _031436_, _031437_, _031438_, _031439_, _031440_, _031441_, _031442_, _031443_, _031444_, _031445_, _031446_, _031447_, _031448_, _031449_, _031450_, _031451_, _031452_, _031453_, _031454_, _031455_, _031456_, _031457_, _031458_, _031459_, _031460_, _031461_, _031462_, _031463_, _031464_, _031465_, _031466_, _031467_, _031468_, _031469_, _031470_, _031471_, _031472_, _031473_, _031474_, _031475_, _031476_, _031477_, _031478_, _031479_, _031480_, _031481_, _031482_, _031483_, _031484_, _031485_, _031486_, _031487_, _031488_, _031489_, _031490_, _031491_, _031492_, _031493_, _031494_, _031495_, _031496_, _031497_, _031498_, _031499_, _031500_, _031501_, _031502_, _031503_, _031504_, _031505_, _031506_, _031507_, _031508_, _031509_, _031510_, _031511_, _031512_, _031513_, _031514_, _031515_, _031516_, _031517_, _031518_, _031519_, _031520_, _031521_, _031522_, _031523_, _031524_, _031525_, _031526_, _031527_, _031528_, _031529_, _031530_, _031531_, _031532_, _031533_, _031534_, _031535_, _031536_, _031537_, _031538_, _031539_, _031540_, _031541_, _031542_, _031543_, _031544_, _031545_, _031546_, _031547_, _031548_, _031549_, _031550_, _031551_, _031552_, _031553_, _031554_, _031555_, _031556_, _031557_, _031558_, _031559_, _031560_, _031561_, _031562_, _031563_, _031564_, _031565_, _031566_, _031567_, _031568_, _031569_, _031570_, _031571_, _031572_, _031573_, _031574_, _031575_, _031576_, _031577_, _031578_, _031579_, _031580_, _031581_, _031582_, _031583_, _031584_, _031585_, _031586_, _031587_, _031588_, _031589_, _031590_, _031591_, _031592_, _031593_, _031594_, _031595_, _031596_, _031597_, _031598_, _031599_, _031600_, _031601_, _031602_, _031603_, _031604_, _031605_, _031606_, _031607_, _031608_, _031609_, _031610_, _031611_, _031612_, _031613_, _031614_, _031615_, _031616_, _031617_, _031618_, _031619_, _031620_, _031621_, _031622_, _031623_, _031624_, _031625_, _031626_, _031627_, _031628_, _031629_, _031630_, _031631_, _031632_, _031633_, _031634_, _031635_, _031636_, _031637_, _031638_, _031639_, _031640_, _031641_, _031642_, _031643_, _031644_, _031645_, _031646_, _031647_, _031648_, _031649_, _031650_, _031651_, _031652_, _031653_, _031654_, _031655_, _031656_, _031657_, _031658_, _031659_, _031660_, _031661_, _031662_, _031663_, _031664_, _031665_, _031666_, _031667_, _031668_, _031669_, _031670_, _031671_, _031672_, _031673_, _031674_, _031675_, _031676_, _031677_, _031678_, _031679_, _031680_, _031681_, _031682_, _031683_, _031684_, _031685_, _031686_, _031687_, _031688_, _031689_, _031690_, _031691_, _031692_, _031693_, _031694_, _031695_, _031696_, _031697_, _031698_, _031699_, _031700_, _031701_, _031702_, _031703_, _031704_, _031705_, _031706_, _031707_, _031708_, _031709_, _031710_, _031711_, _031712_, _031713_, _031714_, _031715_, _031716_, _031717_, _031718_, _031719_, _031720_, _031721_, _031722_, _031723_, _031724_, _031725_, _031726_, _031727_, _031728_, _031729_, _031730_, _031731_, _031732_, _031733_, _031734_, _031735_, _031736_, _031737_, _031738_, _031739_, _031740_, _031741_, _031742_, _031743_, _031744_, _031745_, _031746_, _031747_, _031748_, _031749_, _031750_, _031751_, _031752_, _031753_, _031754_, _031755_, _031756_, _031757_, _031758_, _031759_, _031760_, _031761_, _031762_, _031763_, _031764_, _031765_, _031766_, _031767_, _031768_, _031769_, _031770_, _031771_, _031772_, _031773_, _031774_, _031775_, _031776_, _031777_, _031778_, _031779_, _031780_, _031781_, _031782_, _031783_, _031784_, _031785_, _031786_, _031787_, _031788_, _031789_, _031790_, _031791_, _031792_, _031793_, _031794_, _031795_, _031796_, _031797_, _031798_, _031799_, _031800_, _031801_, _031802_, _031803_, _031804_, _031805_, _031806_, _031807_, _031808_, _031809_, _031810_, _031811_, _031812_, _031813_, _031814_, _031815_, _031816_, _031817_, _031818_, _031819_, _031820_, _031821_, _031822_, _031823_, _031824_, _031825_, _031826_, _031827_, _031828_, _031829_, _031830_, _031831_, _031832_, _031833_, _031834_, _031835_, _031836_, _031837_, _031838_, _031839_, _031840_, _031841_, _031842_, _031843_, _031844_, _031845_, _031846_, _031847_, _031848_, _031849_, _031850_, _031851_, _031852_, _031853_, _031854_, _031855_, _031856_, _031857_, _031858_, _031859_, _031860_, _031861_, _031862_, _031863_, _031864_, _031865_, _031866_, _031867_, _031868_, _031869_, _031870_, _031871_, _031872_, _031873_, _031874_, _031875_, _031876_, _031877_, _031878_, _031879_, _031880_, _031881_, _031882_, _031883_, _031884_, _031885_, _031886_, _031887_, _031888_, _031889_, _031890_, _031891_, _031892_, _031893_, _031894_, _031895_, _031896_, _031897_, _031898_, _031899_, _031900_, _031901_, _031902_, _031903_, _031904_, _031905_, _031906_, _031907_, _031908_, _031909_, _031910_, _031911_, _031912_, _031913_, _031914_, _031915_, _031916_, _031917_, _031918_, _031919_, _031920_, _031921_, _031922_, _031923_, _031924_, _031925_, _031926_, _031927_, _031928_, _031929_, _031930_, _031931_, _031932_, _031933_, _031934_, _031935_, _031936_, _031937_, _031938_, _031939_, _031940_, _031941_, _031942_, _031943_, _031944_, _031945_, _031946_, _031947_, _031948_, _031949_, _031950_, _031951_, _031952_, _031953_, _031954_, _031955_, _031956_, _031957_, _031958_, _031959_, _031960_, _031961_, _031962_, _031963_, _031964_, _031965_, _031966_, _031967_, _031968_, _031969_, _031970_, _031971_, _031972_, _031973_, _031974_, _031975_, _031976_, _031977_, _031978_, _031979_, _031980_, _031981_, _031982_, _031983_, _031984_, _031985_, _031986_, _031987_, _031988_, _031989_, _031990_, _031991_, _031992_, _031993_, _031994_, _031995_, _031996_, _031997_, _031998_, _031999_, _032000_, _032001_, _032002_, _032003_, _032004_, _032005_, _032006_, _032007_, _032008_, _032009_, _032010_, _032011_, _032012_, _032013_, _032014_, _032015_, _032016_, _032017_, _032018_, _032019_, _032020_, _032021_, _032022_, _032023_, _032024_, _032025_, _032026_, _032027_, _032028_, _032029_, _032030_, _032031_, _032032_, _032033_, _032034_, _032035_, _032036_, _032037_, _032038_, _032039_, _032040_, _032041_, _032042_, _032043_, _032044_, _032045_, _032046_, _032047_, _032048_, _032049_, _032050_, _032051_, _032052_, _032053_, _032054_, _032055_, _032056_, _032057_, _032058_, _032059_, _032060_, _032061_, _032062_, _032063_, _032064_, _032065_, _032066_, _032067_, _032068_, _032069_, _032070_, _032071_, _032072_, _032073_, _032074_, _032075_, _032076_, _032077_, _032078_, _032079_, _032080_, _032081_, _032082_, _032083_, _032084_, _032085_, _032086_, _032087_, _032088_, _032089_, _032090_, _032091_, _032092_, _032093_, _032094_, _032095_, _032096_, _032097_, _032098_, _032099_, _032100_, _032101_, _032102_, _032103_, _032104_, _032105_, _032106_, _032107_, _032108_, _032109_, _032110_, _032111_, _032112_, _032113_, _032114_, _032115_, _032116_, _032117_, _032118_, _032119_, _032120_, _032121_, _032122_, _032123_, _032124_, _032125_, _032126_, _032127_, _032128_, _032129_, _032130_, _032131_, _032132_, _032133_, _032134_, _032135_, _032136_, _032137_, _032138_, _032139_, _032140_, _032141_, _032142_, _032143_, _032144_, _032145_, _032146_, _032147_, _032148_, _032149_, _032150_, _032151_, _032152_, _032153_, _032154_, _032155_, _032156_, _032157_, _032158_, _032159_, _032160_, _032161_, _032162_, _032163_, _032164_, _032165_, _032166_, _032167_, _032168_, _032169_, _032170_, _032171_, _032172_, _032173_, _032174_, _032175_, _032176_, _032177_, _032178_, _032179_, _032180_, _032181_, _032182_, _032183_, _032184_, _032185_, _032186_, _032187_, _032188_, _032189_, _032190_, _032191_, _032192_, _032193_, _032194_, _032195_, _032196_, _032197_, _032198_, _032199_, _032200_, _032201_, _032202_, _032203_, _032204_, _032205_, _032206_, _032207_, _032208_, _032209_, _032210_, _032211_, _032212_, _032213_, _032214_, _032215_, _032216_, _032217_, _032218_, _032219_, _032220_, _032221_, _032222_, _032223_, _032224_, _032225_, _032226_, _032227_, _032228_, _032229_, _032230_, _032231_, _032232_, _032233_, _032234_, _032235_, _032236_, _032237_, _032238_, _032239_, _032240_, _032241_, _032242_, _032243_, _032244_, _032245_, _032246_, _032247_, _032248_, _032249_, _032250_, _032251_, _032252_, _032253_, _032254_, _032255_, _032256_, _032257_, _032258_, _032259_, _032260_, _032261_, _032262_, _032263_, _032264_, _032265_, _032266_, _032267_, _032268_, _032269_, _032270_, _032271_, _032272_, _032273_, _032274_, _032275_, _032276_, _032277_, _032278_, _032279_, _032280_, _032281_, _032282_, _032283_, _032284_, _032285_, _032286_, _032287_, _032288_, _032289_, _032290_, _032291_, _032292_, _032293_, _032294_, _032295_, _032296_, _032297_, _032298_, _032299_, _032300_, _032301_, _032302_, _032303_, _032304_, _032305_, _032306_, _032307_, _032308_, _032309_, _032310_, _032311_, _032312_, _032313_, _032314_, _032315_, _032316_, _032317_, _032318_, _032319_, _032320_, _032321_, _032322_, _032323_, _032324_, _032325_, _032326_, _032327_, _032328_, _032329_, _032330_, _032331_, _032332_, _032333_, _032334_, _032335_, _032336_, _032337_, _032338_, _032339_, _032340_, _032341_, _032342_, _032343_, _032344_, _032345_, _032346_, _032347_, _032348_, _032349_, _032350_, _032351_, _032352_, _032353_, _032354_, _032355_, _032356_, _032357_, _032358_, _032359_, _032360_, _032361_, _032362_, _032363_, _032364_, _032365_, _032366_, _032367_, _032368_, _032369_, _032370_, _032371_, _032372_, _032373_, _032374_, _032375_, _032376_, _032377_, _032378_, _032379_, _032380_, _032381_, _032382_, _032383_, _032384_, _032385_, _032386_, _032387_, _032388_, _032389_, _032390_, _032391_, _032392_, _032393_, _032394_, _032395_, _032396_, _032397_, _032398_, _032399_, _032400_, _032401_, _032402_, _032403_, _032404_, _032405_, _032406_, _032407_, _032408_, _032409_, _032410_, _032411_, _032412_, _032413_, _032414_, _032415_, _032416_, _032417_, _032418_, _032419_, _032420_, _032421_, _032422_, _032423_, _032424_, _032425_, _032426_, _032427_, _032428_, _032429_, _032430_, _032431_, _032432_, _032433_, _032434_, _032435_, _032436_, _032437_, _032438_, _032439_, _032440_, _032441_, _032442_, _032443_, _032444_, _032445_, _032446_, _032447_, _032448_, _032449_, _032450_, _032451_, _032452_, _032453_, _032454_, _032455_, _032456_, _032457_, _032458_, _032459_, _032460_, _032461_, _032462_, _032463_, _032464_, _032465_, _032466_, _032467_, _032468_, _032469_, _032470_, _032471_, _032472_, _032473_, _032474_, _032475_, _032476_, _032477_, _032478_, _032479_, _032480_, _032481_, _032482_, _032483_, _032484_, _032485_, _032486_, _032487_, _032488_, _032489_, _032490_, _032491_, _032492_, _032493_, _032494_, _032495_, _032496_, _032497_, _032498_, _032499_, _032500_, _032501_, _032502_, _032503_, _032504_, _032505_, _032506_, _032507_, _032508_, _032509_, _032510_, _032511_, _032512_, _032513_, _032514_, _032515_, _032516_, _032517_, _032518_, _032519_, _032520_, _032521_, _032522_, _032523_, _032524_, _032525_, _032526_, _032527_, _032528_, _032529_, _032530_, _032531_, _032532_, _032533_, _032534_, _032535_, _032536_, _032537_, _032538_, _032539_, _032540_, _032541_, _032542_, _032543_, _032544_, _032545_, _032546_, _032547_, _032548_, _032549_, _032550_, _032551_, _032552_, _032553_, _032554_, _032555_, _032556_, _032557_, _032558_, _032559_, _032560_, _032561_, _032562_, _032563_, _032564_, _032565_, _032566_, _032567_, _032568_, _032569_, _032570_, _032571_, _032572_, _032573_, _032574_, _032575_, _032576_, _032577_, _032578_, _032579_, _032580_, _032581_, _032582_, _032583_, _032584_, _032585_, _032586_, _032587_, _032588_, _032589_, _032590_, _032591_, _032592_, _032593_, _032594_, _032595_, _032596_, _032597_, _032598_, _032599_, _032600_, _032601_, _032602_, _032603_, _032604_, _032605_, _032606_, _032607_, _032608_, _032609_, _032610_, _032611_, _032612_, _032613_, _032614_, _032615_, _032616_, _032617_, _032618_, _032619_, _032620_, _032621_, _032622_, _032623_, _032624_, _032625_, _032626_, _032627_, _032628_, _032629_, _032630_, _032631_, _032632_, _032633_, _032634_, _032635_, _032636_, _032637_, _032638_, _032639_, _032640_, _032641_, _032642_, _032643_, _032644_, _032645_, _032646_, _032647_, _032648_, _032649_, _032650_, _032651_, _032652_, _032653_, _032654_, _032655_, _032656_, _032657_, _032658_, _032659_, _032660_, _032661_, _032662_, _032663_, _032664_, _032665_, _032666_, _032667_, _032668_, _032669_, _032670_, _032671_, _032672_, _032673_, _032674_, _032675_, _032676_, _032677_, _032678_, _032679_, _032680_, _032681_, _032682_, _032683_, _032684_, _032685_, _032686_, _032687_, _032688_, _032689_, _032690_, _032691_, _032692_, _032693_, _032694_, _032695_, _032696_, _032697_, _032698_, _032699_, _032700_, _032701_, _032702_, _032703_, _032704_, _032705_, _032706_, _032707_, _032708_, _032709_, _032710_, _032711_, _032712_, _032713_, _032714_, _032715_, _032716_, _032717_, _032718_, _032719_, _032720_, _032721_, _032722_, _032723_, _032724_, _032725_, _032726_, _032727_, _032728_, _032729_, _032730_, _032731_, _032732_, _032733_, _032734_, _032735_, _032736_, _032737_, _032738_, _032739_, _032740_, _032741_, _032742_, _032743_, _032744_, _032745_, _032746_, _032747_, _032748_, _032749_, _032750_, _032751_, _032752_, _032753_, _032754_, _032755_, _032756_, _032757_, _032758_, _032759_, _032760_, _032761_, _032762_, _032763_, _032764_, _032765_, _032766_, _032767_, _032768_, _032769_, _032770_, _032771_, _032772_, _032773_, _032774_, _032775_, _032776_, _032777_, _032778_, _032779_, _032780_, _032781_, _032782_, _032783_, _032784_, _032785_, _032786_, _032787_, _032788_, _032789_, _032790_, _032791_, _032792_, _032793_, _032794_, _032795_, _032796_, _032797_, _032798_, _032799_, _032800_, _032801_, _032802_, _032803_, _032804_, _032805_, _032806_, _032807_, _032808_, _032809_, _032810_, _032811_, _032812_, _032813_, _032814_, _032815_, _032816_, _032817_, _032818_, _032819_, _032820_, _032821_, _032822_, _032823_, _032824_, _032825_, _032826_, _032827_, _032828_, _032829_, _032830_, _032831_, _032832_, _032833_, _032834_, _032835_, _032836_, _032837_, _032838_, _032839_, _032840_, _032841_, _032842_, _032843_, _032844_, _032845_, _032846_, _032847_, _032848_, _032849_, _032850_, _032851_, _032852_, _032853_, _032854_, _032855_, _032856_, _032857_, _032858_, _032859_, _032860_, _032861_, _032862_, _032863_, _032864_, _032865_, _032866_, _032867_, _032868_, _032869_, _032870_, _032871_, _032872_, _032873_, _032874_, _032875_, _032876_, _032877_, _032878_, _032879_, _032880_, _032881_, _032882_, _032883_, _032884_, _032885_, _032886_, _032887_, _032888_, _032889_, _032890_, _032891_, _032892_, _032893_, _032894_, _032895_, _032896_, _032897_, _032898_, _032899_, _032900_, _032901_, _032902_, _032903_, _032904_, _032905_, _032906_, _032907_, _032908_, _032909_, _032910_, _032911_, _032912_, _032913_, _032914_, _032915_, _032916_, _032917_, _032918_, _032919_, _032920_, _032921_, _032922_, _032923_, _032924_, _032925_, _032926_, _032927_, _032928_, _032929_, _032930_, _032931_, _032932_, _032933_, _032934_, _032935_, _032936_, _032937_, _032938_, _032939_, _032940_, _032941_, _032942_, _032943_, _032944_, _032945_, _032946_, _032947_, _032948_, _032949_, _032950_, _032951_, _032952_, _032953_, _032954_, _032955_, _032956_, _032957_, _032958_, _032959_, _032960_, _032961_, _032962_, _032963_, _032964_, _032965_, _032966_, _032967_, _032968_, _032969_, _032970_, _032971_, _032972_, _032973_, _032974_, _032975_, _032976_, _032977_, _032978_, _032979_, _032980_, _032981_, _032982_, _032983_, _032984_, _032985_, _032986_, _032987_, _032988_, _032989_, _032990_, _032991_, _032992_, _032993_, _032994_, _032995_, _032996_, _032997_, _032998_, _032999_, _033000_, _033001_, _033002_, _033003_, _033004_, _033005_, _033006_, _033007_, _033008_, _033009_, _033010_, _033011_, _033012_, _033013_, _033014_, _033015_, _033016_, _033017_, _033018_, _033019_, _033020_, _033021_, _033022_, _033023_, _033024_, _033025_, _033026_, _033027_, _033028_, _033029_, _033030_, _033031_, _033032_, _033033_, _033034_, _033035_, _033036_, _033037_, _033038_, _033039_, _033040_, _033041_, _033042_, _033043_, _033044_, _033045_, _033046_, _033047_, _033048_, _033049_, _033050_, _033051_, _033052_, _033053_, _033054_, _033055_, _033056_, _033057_, _033058_, _033059_, _033060_, _033061_, _033062_, _033063_, _033064_, _033065_, _033066_, _033067_, _033068_, _033069_, _033070_, _033071_, _033072_, _033073_, _033074_, _033075_, _033076_, _033077_, _033078_, _033079_, _033080_, _033081_, _033082_, _033083_, _033084_, _033085_, _033086_, _033087_, _033088_, _033089_, _033090_, _033091_, _033092_, _033093_, _033094_, _033095_, _033096_, _033097_, _033098_, _033099_, _033100_, _033101_, _033102_, _033103_, _033104_, _033105_, _033106_, _033107_, _033108_, _033109_, _033110_, _033111_, _033112_, _033113_, _033114_, _033115_, _033116_, _033117_, _033118_, _033119_, _033120_, _033121_, _033122_, _033123_, _033124_, _033125_, _033126_, _033127_, _033128_, _033129_, _033130_, _033131_, _033132_, _033133_, _033134_, _033135_, _033136_, _033137_, _033138_, _033139_, _033140_, _033141_, _033142_, _033143_, _033144_, _033145_, _033146_, _033147_, _033148_, _033149_, _033150_, _033151_, _033152_, _033153_, _033154_, _033155_, _033156_, _033157_, _033158_, _033159_, _033160_, _033161_, _033162_, _033163_, _033164_, _033165_, _033166_, _033167_, _033168_, _033169_, _033170_, _033171_, _033172_, _033173_, _033174_, _033175_, _033176_, _033177_, _033178_, _033179_, _033180_, _033181_, _033182_, _033183_, _033184_, _033185_, _033186_, _033187_, _033188_, _033189_, _033190_, _033191_, _033192_, _033193_, _033194_, _033195_, _033196_, _033197_, _033198_, _033199_, _033200_, _033201_, _033202_, _033203_, _033204_, _033205_, _033206_, _033207_, _033208_, _033209_, _033210_, _033211_, _033212_, _033213_, _033214_, _033215_, _033216_, _033217_, _033218_, _033219_, _033220_, _033221_, _033222_, _033223_, _033224_, _033225_, _033226_, _033227_, _033228_, _033229_, _033230_, _033231_, _033232_, _033233_, _033234_, _033235_, _033236_, _033237_, _033238_, _033239_, _033240_, _033241_, _033242_, _033243_, _033244_, _033245_, _033246_, _033247_, _033248_, _033249_, _033250_, _033251_, _033252_, _033253_, _033254_, _033255_, _033256_, _033257_, _033258_, _033259_, _033260_, _033261_, _033262_, _033263_, _033264_, _033265_, _033266_, _033267_, _033268_, _033269_, _033270_, _033271_, _033272_, _033273_, _033274_, _033275_, _033276_, _033277_, _033278_, _033279_, _033280_, _033281_, _033282_, _033283_, _033284_, _033285_, _033286_, _033287_, _033288_, _033289_, _033290_, _033291_, _033292_, _033293_, _033294_, _033295_, _033296_, _033297_, _033298_, _033299_, _033300_, _033301_, _033302_, _033303_, _033304_, _033305_, _033306_, _033307_, _033308_, _033309_, _033310_, _033311_, _033312_, _033313_, _033314_, _033315_, _033316_, _033317_, _033318_, _033319_, _033320_, _033321_, _033322_, _033323_, _033324_, _033325_, _033326_, _033327_, _033328_, _033329_, _033330_, _033331_, _033332_, _033333_, _033334_, _033335_, _033336_, _033337_, _033338_, _033339_, _033340_, _033341_, _033342_, _033343_, _033344_, _033345_, _033346_, _033347_, _033348_, _033349_, _033350_, _033351_, _033352_, _033353_, _033354_, _033355_, _033356_, _033357_, _033358_, _033359_, _033360_, _033361_, _033362_, _033363_, _033364_, _033365_, _033366_, _033367_, _033368_, _033369_, _033370_, _033371_, _033372_, _033373_, _033374_, _033375_, _033376_, _033377_, _033378_, _033379_, _033380_, _033381_, _033382_, _033383_, _033384_, _033385_, _033386_, _033387_, _033388_, _033389_, _033390_, _033391_, _033392_, _033393_, _033394_, _033395_, _033396_, _033397_, _033398_, _033399_, _033400_, _033401_, _033402_, _033403_, _033404_, _033405_, _033406_, _033407_, _033408_, _033409_, _033410_, _033411_, _033412_, _033413_, _033414_, _033415_, _033416_, _033417_, _033418_, _033419_, _033420_, _033421_, _033422_, _033423_, _033424_, _033425_, _033426_, _033427_, _033428_, _033429_, _033430_, _033431_, _033432_, _033433_, _033434_, _033435_, _033436_, _033437_, _033438_, _033439_, _033440_, _033441_, _033442_, _033443_, _033444_, _033445_, _033446_, _033447_, _033448_, _033449_, _033450_, _033451_, _033452_, _033453_, _033454_, _033455_, _033456_, _033457_, _033458_, _033459_, _033460_, _033461_, _033462_, _033463_, _033464_, _033465_, _033466_, _033467_, _033468_, _033469_, _033470_, _033471_, _033472_, _033473_, _033474_, _033475_, _033476_, _033477_, _033478_, _033479_, _033480_, _033481_, _033482_, _033483_, _033484_, _033485_, _033486_, _033487_, _033488_, _033489_, _033490_, _033491_, _033492_, _033493_, _033494_, _033495_, _033496_, _033497_, _033498_, _033499_, _033500_, _033501_, _033502_, _033503_, _033504_, _033505_, _033506_, _033507_, _033508_, _033509_, _033510_, _033511_, _033512_, _033513_, _033514_, _033515_, _033516_, _033517_, _033518_, _033519_, _033520_, _033521_, _033522_, _033523_, _033524_, _033525_, _033526_, _033527_, _033528_, _033529_, _033530_, _033531_, _033532_, _033533_, _033534_, _033535_, _033536_, _033537_, _033538_, _033539_, _033540_, _033541_, _033542_, _033543_, _033544_, _033545_, _033546_, _033547_, _033548_, _033549_, _033550_, _033551_, _033552_, _033553_, _033554_, _033555_, _033556_, _033557_, _033558_, _033559_, _033560_, _033561_, _033562_, _033563_, _033564_, _033565_, _033566_, _033567_, _033568_, _033569_, _033570_, _033571_, _033572_, _033573_, _033574_, _033575_, _033576_, _033577_, _033578_, _033579_, _033580_, _033581_, _033582_, _033583_, _033584_, _033585_, _033586_, _033587_, _033588_, _033589_, _033590_, _033591_, _033592_, _033593_, _033594_, _033595_, _033596_, _033597_, _033598_, _033599_, _033600_, _033601_, _033602_, _033603_, _033604_, _033605_, _033606_, _033607_, _033608_, _033609_, _033610_, _033611_, _033612_, _033613_, _033614_, _033615_, _033616_, _033617_, _033618_, _033619_, _033620_, _033621_, _033622_, _033623_, _033624_, _033625_, _033626_, _033627_, _033628_, _033629_, _033630_, _033631_, _033632_, _033633_, _033634_, _033635_, _033636_, _033637_, _033638_, _033639_, _033640_, _033641_, _033642_, _033643_, _033644_, _033645_, _033646_, _033647_, _033648_, _033649_, _033650_, _033651_, _033652_, _033653_, _033654_, _033655_, _033656_, _033657_, _033658_, _033659_, _033660_, _033661_, _033662_, _033663_, _033664_, _033665_, _033666_, _033667_, _033668_, _033669_, _033670_, _033671_, _033672_, _033673_, _033674_, _033675_, _033676_, _033677_, _033678_, _033679_, _033680_, _033681_, _033682_, _033683_, _033684_, _033685_, _033686_, _033687_, _033688_, _033689_, _033690_, _033691_, _033692_, _033693_, _033694_, _033695_, _033696_, _033697_, _033698_, _033699_, _033700_, _033701_, _033702_, _033703_, _033704_, _033705_, _033706_, _033707_, _033708_, _033709_, _033710_, _033711_, _033712_, _033713_, _033714_, _033715_, _033716_, _033717_, _033718_, _033719_, _033720_, _033721_, _033722_, _033723_, _033724_, _033725_, _033726_, _033727_, _033728_, _033729_, _033730_, _033731_, _033732_, _033733_, _033734_, _033735_, _033736_, _033737_, _033738_, _033739_, _033740_, _033741_, _033742_, _033743_, _033744_, _033745_, _033746_, _033747_, _033748_, _033749_, _033750_, _033751_, _033752_, _033753_, _033754_, _033755_, _033756_, _033757_, _033758_, _033759_, _033760_, _033761_, _033762_, _033763_, _033764_, _033765_, _033766_, _033767_, _033768_, _033769_, _033770_, _033771_, _033772_, _033773_, _033774_, _033775_, _033776_, _033777_, _033778_, _033779_, _033780_, _033781_, _033782_, _033783_, _033784_, _033785_, _033786_, _033787_, _033788_, _033789_, _033790_, _033791_, _033792_, _033793_, _033794_, _033795_, _033796_, _033797_, _033798_, _033799_, _033800_, _033801_, _033802_, _033803_, _033804_, _033805_, _033806_, _033807_, _033808_, _033809_, _033810_, _033811_, _033812_, _033813_, _033814_, _033815_, _033816_, _033817_, _033818_, _033819_, _033820_, _033821_, _033822_, _033823_, _033824_, _033825_, _033826_, _033827_, _033828_, _033829_, _033830_, _033831_, _033832_, _033833_, _033834_, _033835_, _033836_, _033837_, _033838_, _033839_, _033840_, _033841_, _033842_, _033843_, _033844_, _033845_, _033846_, _033847_, _033848_, _033849_, _033850_, _033851_, _033852_, _033853_, _033854_, _033855_, _033856_, _033857_, _033858_, _033859_, _033860_, _033861_, _033862_, _033863_, _033864_, _033865_, _033866_, _033867_, _033868_, _033869_, _033870_, _033871_, _033872_, _033873_, _033874_, _033875_, _033876_, _033877_, _033878_, _033879_, _033880_, _033881_, _033882_, _033883_, _033884_, _033885_, _033886_, _033887_, _033888_, _033889_, _033890_, _033891_, _033892_, _033893_, _033894_, _033895_, _033896_, _033897_, _033898_, _033899_, _033900_, _033901_, _033902_, _033903_, _033904_, _033905_, _033906_, _033907_, _033908_, _033909_, _033910_, _033911_, _033912_, _033913_, _033914_, _033915_, _033916_, _033917_, _033918_, _033919_, _033920_, _033921_, _033922_, _033923_, _033924_, _033925_, _033926_, _033927_, _033928_, _033929_, _033930_, _033931_, _033932_, _033933_, _033934_, _033935_, _033936_, _033937_, _033938_, _033939_, _033940_, _033941_, _033942_, _033943_, _033944_, _033945_, _033946_, _033947_, _033948_, _033949_, _033950_, _033951_, _033952_, _033953_, _033954_, _033955_, _033956_, _033957_, _033958_, _033959_, _033960_, _033961_, _033962_, _033963_, _033964_, _033965_, _033966_, _033967_, _033968_, _033969_, _033970_, _033971_, _033972_, _033973_, _033974_, _033975_, _033976_, _033977_, _033978_, _033979_, _033980_, _033981_, _033982_, _033983_, _033984_, _033985_, _033986_, _033987_, _033988_, _033989_, _033990_, _033991_, _033992_, _033993_, _033994_, _033995_, _033996_, _033997_, _033998_, _033999_, _034000_, _034001_, _034002_, _034003_, _034004_, _034005_, _034006_, _034007_, _034008_, _034009_, _034010_, _034011_, _034012_, _034013_, _034014_, _034015_, _034016_, _034017_, _034018_, _034019_, _034020_, _034021_, _034022_, _034023_, _034024_, _034025_, _034026_, _034027_, _034028_, _034029_, _034030_, _034031_, _034032_, _034033_, _034034_, _034035_, _034036_, _034037_, _034038_, _034039_, _034040_, _034041_, _034042_, _034043_, _034044_, _034045_, _034046_, _034047_, _034048_, _034049_, _034050_, _034051_, _034052_, _034053_, _034054_, _034055_, _034056_, _034057_, _034058_, _034059_, _034060_, _034061_, _034062_, _034063_, _034064_, _034065_, _034066_, _034067_, _034068_, _034069_, _034070_, _034071_, _034072_, _034073_, _034074_, _034075_, _034076_, _034077_, _034078_, _034079_, _034080_, _034081_, _034082_, _034083_, _034084_, _034085_, _034086_, _034087_, _034088_, _034089_, _034090_, _034091_, _034092_, _034093_, _034094_, _034095_, _034096_, _034097_, _034098_, _034099_, _034100_, _034101_, _034102_, _034103_, _034104_, _034105_, _034106_, _034107_, _034108_, _034109_, _034110_, _034111_, _034112_, _034113_, _034114_, _034115_, _034116_, _034117_, _034118_, _034119_, _034120_, _034121_, _034122_, _034123_, _034124_, _034125_, _034126_, _034127_, _034128_, _034129_, _034130_, _034131_, _034132_, _034133_, _034134_, _034135_, _034136_, _034137_, _034138_, _034139_, _034140_, _034141_, _034142_, _034143_, _034144_, _034145_, _034146_, _034147_, _034148_, _034149_, _034150_, _034151_, _034152_, _034153_, _034154_, _034155_, _034156_, _034157_, _034158_, _034159_, _034160_, _034161_, _034162_, _034163_, _034164_, _034165_, _034166_, _034167_, _034168_, _034169_, _034170_, _034171_, _034172_, _034173_, _034174_, _034175_, _034176_, _034177_, _034178_, _034179_, _034180_, _034181_, _034182_, _034183_, _034184_, _034185_, _034186_, _034187_, _034188_, _034189_, _034190_, _034191_, _034192_, _034193_, _034194_, _034195_, _034196_, _034197_, _034198_, _034199_, _034200_, _034201_, _034202_, _034203_, _034204_, _034205_, _034206_, _034207_, _034208_, _034209_, _034210_, _034211_, _034212_, _034213_, _034214_, _034215_, _034216_, _034217_, _034218_, _034219_, _034220_, _034221_, _034222_, _034223_, _034224_, _034225_, _034226_, _034227_, _034228_, _034229_, _034230_, _034231_, _034232_, _034233_, _034234_, _034235_, _034236_, _034237_, _034238_, _034239_, _034240_, _034241_, _034242_, _034243_, _034244_, _034245_, _034246_, _034247_, _034248_, _034249_, _034250_, _034251_, _034252_, _034253_, _034254_, _034255_, _034256_, _034257_, _034258_, _034259_, _034260_, _034261_, _034262_, _034263_, _034264_, _034265_, _034266_, _034267_, _034268_, _034269_, _034270_, _034271_, _034272_, _034273_, _034274_, _034275_, _034276_, _034277_, _034278_, _034279_, _034280_, _034281_, _034282_, _034283_, _034284_, _034285_, _034286_, _034287_, _034288_, _034289_, _034290_, _034291_, _034292_, _034293_, _034294_, _034295_, _034296_, _034297_, _034298_, _034299_, _034300_, _034301_, _034302_, _034303_, _034304_, _034305_, _034306_, _034307_, _034308_, _034309_, _034310_, _034311_, _034312_, _034313_, _034314_, _034315_, _034316_, _034317_, _034318_, _034319_, _034320_, _034321_, _034322_, _034323_, _034324_, _034325_, _034326_, _034327_, _034328_, _034329_, _034330_, _034331_, _034332_, _034333_, _034334_, _034335_, _034336_, _034337_, _034338_, _034339_, _034340_, _034341_, _034342_, _034343_, _034344_, _034345_, _034346_, _034347_, _034348_, _034349_, _034350_, _034351_, _034352_, _034353_, _034354_, _034355_, _034356_, _034357_, _034358_, _034359_, _034360_, _034361_, _034362_, _034363_, _034364_, _034365_, _034366_, _034367_, _034368_, _034369_, _034370_, _034371_, _034372_, _034373_, _034374_, _034375_, _034376_, _034377_, _034378_, _034379_, _034380_, _034381_, _034382_, _034383_, _034384_, _034385_, _034386_, _034387_, _034388_, _034389_, _034390_, _034391_, _034392_, _034393_, _034394_, _034395_, _034396_, _034397_, _034398_, _034399_, _034400_, _034401_, _034402_, _034403_, _034404_, _034405_, _034406_, _034407_, _034408_, _034409_, _034410_, _034411_, _034412_, _034413_, _034414_, _034415_, _034416_, _034417_, _034418_, _034419_, _034420_, _034421_, _034422_, _034423_, _034424_, _034425_, _034426_, _034427_, _034428_, _034429_, _034430_, _034431_, _034432_, _034433_, _034434_, _034435_, _034436_, _034437_, _034438_, _034439_, _034440_, _034441_, _034442_, _034443_, _034444_, _034445_, _034446_, _034447_, _034448_, _034449_, _034450_, _034451_, _034452_, _034453_, _034454_, _034455_, _034456_, _034457_, _034458_, _034459_, _034460_, _034461_, _034462_, _034463_, _034464_, _034465_, _034466_, _034467_, _034468_, _034469_, _034470_, _034471_, _034472_, _034473_, _034474_, _034475_, _034476_, _034477_, _034478_, _034479_, _034480_, _034481_, _034482_, _034483_, _034484_, _034485_, _034486_, _034487_, _034488_, _034489_, _034490_, _034491_, _034492_, _034493_, _034494_, _034495_, _034496_, _034497_, _034498_, _034499_, _034500_, _034501_, _034502_, _034503_, _034504_, _034505_, _034506_, _034507_, _034508_, _034509_, _034510_, _034511_, _034512_, _034513_, _034514_, _034515_, _034516_, _034517_, _034518_, _034519_, _034520_, _034521_, _034522_, _034523_, _034524_, _034525_, _034526_, _034527_, _034528_, _034529_, _034530_, _034531_, _034532_, _034533_, _034534_, _034535_, _034536_, _034537_, _034538_, _034539_, _034540_, _034541_, _034542_, _034543_, _034544_, _034545_, _034546_, _034547_, _034548_, _034549_, _034550_, _034551_, _034552_, _034553_, _034554_, _034555_, _034556_, _034557_, _034558_, _034559_, _034560_, _034561_, _034562_, _034563_, _034564_, _034565_, _034566_, _034567_, _034568_, _034569_, _034570_, _034571_, _034572_, _034573_, _034574_, _034575_, _034576_, _034577_, _034578_, _034579_, _034580_, _034581_, _034582_, _034583_, _034584_, _034585_, _034586_, _034587_, _034588_, _034589_, _034590_, _034591_, _034592_, _034593_, _034594_, _034595_, _034596_, _034597_, _034598_, _034599_, _034600_, _034601_, _034602_, _034603_, _034604_, _034605_, _034606_, _034607_, _034608_, _034609_, _034610_, _034611_, _034612_, _034613_, _034614_, _034615_, _034616_, _034617_, _034618_, _034619_, _034620_, _034621_, _034622_, _034623_, _034624_, _034625_, _034626_, _034627_, _034628_, _034629_, _034630_, _034631_, _034632_, _034633_, _034634_, _034635_, _034636_, _034637_, _034638_, _034639_, _034640_, _034641_, _034642_, _034643_, _034644_, _034645_, _034646_, _034647_, _034648_, _034649_, _034650_, _034651_, _034652_, _034653_, _034654_, _034655_, _034656_, _034657_, _034658_, _034659_, _034660_, _034661_, _034662_, _034663_, _034664_, _034665_, _034666_, _034667_, _034668_, _034669_, _034670_, _034671_, _034672_, _034673_, _034674_, _034675_, _034676_, _034677_, _034678_, _034679_, _034680_, _034681_, _034682_, _034683_, _034684_, _034685_, _034686_, _034687_, _034688_, _034689_, _034690_, _034691_, _034692_, _034693_, _034694_, _034695_, _034696_, _034697_, _034698_, _034699_, _034700_, _034701_, _034702_, _034703_, _034704_, _034705_, _034706_, _034707_, _034708_, _034709_, _034710_, _034711_, _034712_, _034713_, _034714_, _034715_, _034716_, _034717_, _034718_, _034719_, _034720_, _034721_, _034722_, _034723_, _034724_, _034725_, _034726_, _034727_, _034728_, _034729_, _034730_, _034731_, _034732_, _034733_, _034734_, _034735_, _034736_, _034737_, _034738_, _034739_, _034740_, _034741_, _034742_, _034743_, _034744_, _034745_, _034746_, _034747_, _034748_, _034749_, _034750_, _034751_, _034752_, _034753_, _034754_, _034755_, _034756_, _034757_, _034758_, _034759_, _034760_, _034761_, _034762_, _034763_, _034764_, _034765_, _034766_, _034767_, _034768_, _034769_, _034770_, _034771_, _034772_, _034773_, _034774_, _034775_, _034776_, _034777_, _034778_, _034779_, _034780_, _034781_, _034782_, _034783_, _034784_, _034785_, _034786_, _034787_, _034788_, _034789_, _034790_, _034791_, _034792_, _034793_, _034794_, _034795_, _034796_, _034797_, _034798_, _034799_, _034800_, _034801_, _034802_, _034803_, _034804_, _034805_, _034806_, _034807_, _034808_, _034809_, _034810_, _034811_, _034812_, _034813_, _034814_, _034815_, _034816_, _034817_, _034818_, _034819_, _034820_, _034821_, _034822_, _034823_, _034824_, _034825_, _034826_, _034827_, _034828_, _034829_, _034830_, _034831_, _034832_, _034833_, _034834_, _034835_, _034836_, _034837_, _034838_, _034839_, _034840_, _034841_, _034842_, _034843_, _034844_, _034845_, _034846_, _034847_, _034848_, _034849_, _034850_, _034851_, _034852_, _034853_, _034854_, _034855_, _034856_, _034857_, _034858_, _034859_, _034860_, _034861_, _034862_, _034863_, _034864_, _034865_, _034866_, _034867_, _034868_, _034869_, _034870_, _034871_, _034872_, _034873_, _034874_, _034875_, _034876_, _034877_, _034878_, _034879_, _034880_, _034881_, _034882_, _034883_, _034884_, _034885_, _034886_, _034887_, _034888_, _034889_, _034890_, _034891_, _034892_, _034893_, _034894_, _034895_, _034896_, _034897_, _034898_, _034899_, _034900_, _034901_, _034902_, _034903_, _034904_, _034905_, _034906_, _034907_, _034908_, _034909_, _034910_, _034911_, _034912_, _034913_, _034914_, _034915_, _034916_, _034917_, _034918_, _034919_, _034920_, _034921_, _034922_, _034923_, _034924_, _034925_, _034926_, _034927_, _034928_, _034929_, _034930_, _034931_, _034932_, _034933_, _034934_, _034935_, _034936_, _034937_, _034938_, _034939_, _034940_, _034941_, _034942_, _034943_, _034944_, _034945_, _034946_, _034947_, _034948_, _034949_, _034950_, _034951_, _034952_, _034953_, _034954_, _034955_, _034956_, _034957_, _034958_, _034959_, _034960_, _034961_, _034962_, _034963_, _034964_, _034965_, _034966_, _034967_, _034968_, _034969_, _034970_, _034971_, _034972_, _034973_, _034974_, _034975_, _034976_, _034977_, _034978_, _034979_, _034980_, _034981_, _034982_, _034983_, _034984_, _034985_, _034986_, _034987_, _034988_, _034989_, _034990_, _034991_, _034992_, _034993_, _034994_, _034995_, _034996_, _034997_, _034998_, _034999_, _035000_, _035001_, _035002_, _035003_, _035004_, _035005_, _035006_, _035007_, _035008_, _035009_, _035010_, _035011_, _035012_, _035013_, _035014_, _035015_, _035016_, _035017_, _035018_, _035019_, _035020_, _035021_, _035022_, _035023_, _035024_, _035025_, _035026_, _035027_, _035028_, _035029_, _035030_, _035031_, _035032_, _035033_, _035034_, _035035_, _035036_, _035037_, _035038_, _035039_, _035040_, _035041_, _035042_, _035043_, _035044_, _035045_, _035046_, _035047_, _035048_, _035049_, _035050_, _035051_, _035052_, _035053_, _035054_, _035055_, _035056_, _035057_, _035058_, _035059_, _035060_, _035061_, _035062_, _035063_, _035064_, _035065_, _035066_, _035067_, _035068_, _035069_, _035070_, _035071_, _035072_, _035073_, _035074_, _035075_, _035076_, _035077_, _035078_, _035079_, _035080_, _035081_, _035082_, _035083_, _035084_, _035085_, _035086_, _035087_, _035088_, _035089_, _035090_, _035091_, _035092_, _035093_, _035094_, _035095_, _035096_, _035097_, _035098_, _035099_, _035100_, _035101_, _035102_, _035103_, _035104_, _035105_, _035106_, _035107_, _035108_, _035109_, _035110_, _035111_, _035112_, _035113_, _035114_, _035115_, _035116_, _035117_, _035118_, _035119_, _035120_, _035121_, _035122_, _035123_, _035124_, _035125_, _035126_, _035127_, _035128_, _035129_, _035130_, _035131_, _035132_, _035133_, _035134_, _035135_, _035136_, _035137_, _035138_, _035139_, _035140_, _035141_, _035142_, _035143_, _035144_, _035145_, _035146_, _035147_, _035148_, _035149_, _035150_, _035151_, _035152_, _035153_, _035154_, _035155_, _035156_, _035157_, _035158_, _035159_, _035160_, _035161_, _035162_, _035163_, _035164_, _035165_, _035166_, _035167_, _035168_, _035169_, _035170_, _035171_, _035172_, _035173_, _035174_, _035175_, _035176_, _035177_, _035178_, _035179_, _035180_, _035181_, _035182_, _035183_, _035184_, _035185_, _035186_, _035187_, _035188_, _035189_, _035190_, _035191_, _035192_, _035193_, _035194_, _035195_, _035196_, _035197_, _035198_, _035199_, _035200_, _035201_, _035202_, _035203_, _035204_, _035205_, _035206_, _035207_, _035208_, _035209_, _035210_, _035211_, _035212_, _035213_, _035214_, _035215_, _035216_, _035217_, _035218_, _035219_, _035220_, _035221_, _035222_, _035223_, _035224_, _035225_, _035226_, _035227_, _035228_, _035229_, _035230_, _035231_, _035232_, _035233_, _035234_, _035235_, _035236_, _035237_, _035238_, _035239_, _035240_, _035241_, _035242_, _035243_, _035244_, _035245_, _035246_, _035247_, _035248_, _035249_, _035250_, _035251_, _035252_, _035253_, _035254_, _035255_, _035256_, _035257_, _035258_, _035259_, _035260_, _035261_, _035262_, _035263_, _035264_, _035265_, _035266_, _035267_, _035268_, _035269_, _035270_, _035271_, _035272_, _035273_, _035274_, _035275_, _035276_, _035277_, _035278_, _035279_, _035280_, _035281_, _035282_, _035283_, _035284_, _035285_, _035286_, _035287_, _035288_, _035289_, _035290_, _035291_, _035292_, _035293_, _035294_, _035295_, _035296_, _035297_, _035298_, _035299_, _035300_, _035301_, _035302_, _035303_, _035304_, _035305_, _035306_, _035307_, _035308_, _035309_, _035310_, _035311_, _035312_, _035313_, _035314_, _035315_, _035316_, _035317_, _035318_, _035319_, _035320_, _035321_, _035322_, _035323_, _035324_, _035325_, _035326_, _035327_, _035328_, _035329_, _035330_, _035331_, _035332_, _035333_, _035334_, _035335_, _035336_, _035337_, _035338_, _035339_, _035340_, _035341_, _035342_, _035343_, _035344_, _035345_, _035346_, _035347_, _035348_, _035349_, _035350_, _035351_, _035352_, _035353_, _035354_, _035355_, _035356_, _035357_, _035358_, _035359_, _035360_, _035361_, _035362_, _035363_, _035364_, _035365_, _035366_, _035367_, _035368_, _035369_, _035370_, _035371_, _035372_, _035373_, _035374_, _035375_, _035376_, _035377_, _035378_, _035379_, _035380_, _035381_, _035382_, _035383_, _035384_, _035385_, _035386_, _035387_, _035388_, _035389_, _035390_, _035391_, _035392_, _035393_, _035394_, _035395_, _035396_, _035397_, _035398_, _035399_, _035400_, _035401_, _035402_, _035403_, _035404_, _035405_, _035406_, _035407_, _035408_, _035409_, _035410_, _035411_, _035412_, _035413_, _035414_, _035415_, _035416_, _035417_, _035418_, _035419_, _035420_, _035421_, _035422_, _035423_, _035424_, _035425_, _035426_, _035427_, _035428_, _035429_, _035430_, _035431_, _035432_, _035433_, _035434_, _035435_, _035436_, _035437_, _035438_, _035439_, _035440_, _035441_, _035442_, _035443_, _035444_, _035445_, _035446_, _035447_, _035448_, _035449_, _035450_, _035451_, _035452_, _035453_, _035454_, _035455_, _035456_, _035457_, _035458_, _035459_, _035460_, _035461_, _035462_, _035463_, _035464_, _035465_, _035466_, _035467_, _035468_, _035469_, _035470_, _035471_, _035472_, _035473_, _035474_, _035475_, _035476_, _035477_, _035478_, _035479_, _035480_, _035481_, _035482_, _035483_, _035484_, _035485_, _035486_, _035487_, _035488_, _035489_, _035490_, _035491_, _035492_, _035493_, _035494_, _035495_, _035496_, _035497_, _035498_, _035499_, _035500_, _035501_, _035502_, _035503_, _035504_, _035505_, _035506_, _035507_, _035508_, _035509_, _035510_, _035511_, _035512_, _035513_, _035514_, _035515_, _035516_, _035517_, _035518_, _035519_, _035520_, _035521_, _035522_, _035523_, _035524_, _035525_, _035526_, _035527_, _035528_, _035529_, _035530_, _035531_, _035532_, _035533_, _035534_, _035535_, _035536_, _035537_, _035538_, _035539_, _035540_, _035541_, _035542_, _035543_, _035544_, _035545_, _035546_, _035547_, _035548_, _035549_, _035550_, _035551_, _035552_, _035553_, _035554_, _035555_, _035556_, _035557_, _035558_, _035559_, _035560_, _035561_, _035562_, _035563_, _035564_, _035565_, _035566_, _035567_, _035568_, _035569_, _035570_, _035571_, _035572_, _035573_, _035574_, _035575_, _035576_, _035577_, _035578_, _035579_, _035580_, _035581_, _035582_, _035583_, _035584_, _035585_, _035586_, _035587_, _035588_, _035589_, _035590_, _035591_, _035592_, _035593_, _035594_, _035595_, _035596_, _035597_, _035598_, _035599_, _035600_, _035601_, _035602_, _035603_, _035604_, _035605_, _035606_, _035607_, _035608_, _035609_, _035610_, _035611_, _035612_, _035613_, _035614_, _035615_, _035616_, _035617_, _035618_, _035619_, _035620_, _035621_, _035622_, _035623_, _035624_, _035625_, _035626_, _035627_, _035628_, _035629_, _035630_, _035631_, _035632_, _035633_, _035634_, _035635_, _035636_, _035637_, _035638_, _035639_, _035640_, _035641_, _035642_, _035643_, _035644_, _035645_, _035646_, _035647_, _035648_, _035649_, _035650_, _035651_, _035652_, _035653_, _035654_, _035655_, _035656_, _035657_, _035658_, _035659_, _035660_, _035661_, _035662_, _035663_, _035664_, _035665_, _035666_, _035667_, _035668_, _035669_, _035670_, _035671_, _035672_, _035673_, _035674_, _035675_, _035676_, _035677_, _035678_, _035679_, _035680_, _035681_, _035682_, _035683_, _035684_, _035685_, _035686_, _035687_, _035688_, _035689_, _035690_, _035691_, _035692_, _035693_, _035694_, _035695_, _035696_, _035697_, _035698_, _035699_, _035700_, _035701_, _035702_, _035703_, _035704_, _035705_, _035706_, _035707_, _035708_, _035709_, _035710_, _035711_, _035712_, _035713_, _035714_, _035715_, _035716_, _035717_, _035718_, _035719_, _035720_, _035721_, _035722_, _035723_, _035724_, _035725_, _035726_, _035727_, _035728_, _035729_, _035730_, _035731_, _035732_, _035733_, _035734_, _035735_, _035736_, _035737_, _035738_, _035739_, _035740_, _035741_, _035742_, _035743_, _035744_, _035745_, _035746_, _035747_, _035748_, _035749_, _035750_, _035751_, _035752_, _035753_, _035754_, _035755_, _035756_, _035757_, _035758_, _035759_, _035760_, _035761_, _035762_, _035763_, _035764_, _035765_, _035766_, _035767_, _035768_, _035769_, _035770_, _035771_, _035772_, _035773_, _035774_, _035775_, _035776_, _035777_, _035778_, _035779_, _035780_, _035781_, _035782_, _035783_, _035784_, _035785_, _035786_, _035787_, _035788_, _035789_, _035790_, _035791_, _035792_, _035793_, _035794_, _035795_, _035796_, _035797_, _035798_, _035799_, _035800_, _035801_, _035802_, _035803_, _035804_, _035805_, _035806_, _035807_, _035808_, _035809_, _035810_, _035811_, _035812_, _035813_, _035814_, _035815_, _035816_, _035817_, _035818_, _035819_, _035820_, _035821_, _035822_, _035823_, _035824_, _035825_, _035826_, _035827_, _035828_, _035829_, _035830_, _035831_, _035832_, _035833_, _035834_, _035835_, _035836_, _035837_, _035838_, _035839_, _035840_, _035841_, _035842_, _035843_, _035844_, _035845_, _035846_, _035847_, _035848_, _035849_, _035850_, _035851_, _035852_, _035853_, _035854_, _035855_, _035856_, _035857_, _035858_, _035859_, _035860_, _035861_, _035862_, _035863_, _035864_, _035865_, _035866_, _035867_, _035868_, _035869_, _035870_, _035871_, _035872_, _035873_, _035874_, _035875_, _035876_, _035877_, _035878_, _035879_, _035880_, _035881_, _035882_, _035883_, _035884_, _035885_, _035886_, _035887_, _035888_, _035889_, _035890_, _035891_, _035892_, _035893_, _035894_, _035895_, _035896_, _035897_, _035898_, _035899_, _035900_, _035901_, _035902_, _035903_, _035904_, _035905_, _035906_, _035907_, _035908_, _035909_, _035910_, _035911_, _035912_, _035913_, _035914_, _035915_, _035916_, _035917_, _035918_, _035919_, _035920_, _035921_, _035922_, _035923_, _035924_, _035925_, _035926_, _035927_, _035928_, _035929_, _035930_, _035931_, _035932_, _035933_, _035934_, _035935_, _035936_, _035937_, _035938_, _035939_, _035940_, _035941_, _035942_, _035943_, _035944_, _035945_, _035946_, _035947_, _035948_, _035949_, _035950_, _035951_, _035952_, _035953_, _035954_, _035955_, _035956_, _035957_, _035958_, _035959_, _035960_, _035961_, _035962_, _035963_, _035964_, _035965_, _035966_, _035967_, _035968_, _035969_, _035970_, _035971_, _035972_, _035973_, _035974_, _035975_, _035976_, _035977_, _035978_, _035979_, _035980_, _035981_, _035982_, _035983_, _035984_, _035985_, _035986_, _035987_, _035988_, _035989_, _035990_, _035991_, _035992_, _035993_, _035994_, _035995_, _035996_, _035997_, _035998_, _035999_, _036000_, _036001_, _036002_, _036003_, _036004_, _036005_, _036006_, _036007_, _036008_, _036009_, _036010_, _036011_, _036012_, _036013_, _036014_, _036015_, _036016_, _036017_, _036018_, _036019_, _036020_, _036021_, _036022_, _036023_, _036024_, _036025_, _036026_, _036027_, _036028_, _036029_, _036030_, _036031_, _036032_, _036033_, _036034_, _036035_, _036036_, _036037_, _036038_, _036039_, _036040_, _036041_, _036042_, _036043_, _036044_, _036045_, _036046_, _036047_, _036048_, _036049_, _036050_, _036051_, _036052_, _036053_, _036054_, _036055_, _036056_, _036057_, _036058_, _036059_, _036060_, _036061_, _036062_, _036063_, _036064_, _036065_, _036066_, _036067_, _036068_, _036069_, _036070_, _036071_, _036072_, _036073_, _036074_, _036075_, _036076_, _036077_, _036078_, _036079_, _036080_, _036081_, _036082_, _036083_, _036084_, _036085_, _036086_, _036087_, _036088_, _036089_, _036090_, _036091_, _036092_, _036093_, _036094_, _036095_, _036096_, _036097_, _036098_, _036099_, _036100_, _036101_, _036102_, _036103_, _036104_, _036105_, _036106_, _036107_, _036108_, _036109_, _036110_, _036111_, _036112_, _036113_, _036114_, _036115_, _036116_, _036117_, _036118_, _036119_, _036120_, _036121_, _036122_, _036123_, _036124_, _036125_, _036126_, _036127_, _036128_, _036129_, _036130_, _036131_, _036132_, _036133_, _036134_, _036135_, _036136_, _036137_, _036138_, _036139_, _036140_, _036141_, _036142_, _036143_, _036144_, _036145_, _036146_, _036147_, _036148_, _036149_, _036150_, _036151_, _036152_, _036153_, _036154_, _036155_, _036156_, _036157_, _036158_, _036159_, _036160_, _036161_, _036162_, _036163_, _036164_, _036165_, _036166_, _036167_, _036168_, _036169_, _036170_, _036171_, _036172_, _036173_, _036174_, _036175_, _036176_, _036177_, _036178_, _036179_, _036180_, _036181_, _036182_, _036183_, _036184_, _036185_, _036186_, _036187_, _036188_, _036189_, _036190_, _036191_, _036192_, _036193_, _036194_, _036195_, _036196_, _036197_, _036198_, _036199_, _036200_, _036201_, _036202_, _036203_, _036204_, _036205_, _036206_, _036207_, _036208_, _036209_, _036210_, _036211_, _036212_, _036213_, _036214_, _036215_, _036216_, _036217_, _036218_, _036219_, _036220_, _036221_, _036222_, _036223_, _036224_, _036225_, _036226_, _036227_, _036228_, _036229_, _036230_, _036231_, _036232_, _036233_, _036234_, _036235_, _036236_, _036237_, _036238_, _036239_, _036240_, _036241_, _036242_, _036243_, _036244_, _036245_, _036246_, _036247_, _036248_, _036249_, _036250_, _036251_, _036252_, _036253_, _036254_, _036255_, _036256_, _036257_, _036258_, _036259_, _036260_, _036261_, _036262_, _036263_, _036264_, _036265_, _036266_, _036267_, _036268_, _036269_, _036270_, _036271_, _036272_, _036273_, _036274_, _036275_, _036276_, _036277_, _036278_, _036279_, _036280_, _036281_, _036282_, _036283_, _036284_, _036285_, _036286_, _036287_, _036288_, _036289_, _036290_, _036291_, _036292_, _036293_, _036294_, _036295_, _036296_, _036297_, _036298_, _036299_, _036300_, _036301_, _036302_, _036303_, _036304_, _036305_, _036306_, _036307_, _036308_, _036309_, _036310_, _036311_, _036312_, _036313_, _036314_, _036315_, _036316_, _036317_, _036318_, _036319_, _036320_, _036321_, _036322_, _036323_, _036324_, _036325_, _036326_, _036327_, _036328_, _036329_, _036330_, _036331_, _036332_, _036333_, _036334_, _036335_, _036336_, _036337_, _036338_, _036339_, _036340_, _036341_, _036342_, _036343_, _036344_, _036345_, _036346_, _036347_, _036348_, _036349_, _036350_, _036351_, _036352_, _036353_, _036354_, _036355_, _036356_, _036357_, _036358_, _036359_, _036360_, _036361_, _036362_, _036363_, _036364_, _036365_, _036366_, _036367_, _036368_, _036369_, _036370_, _036371_, _036372_, _036373_, _036374_, _036375_, _036376_, _036377_, _036378_, _036379_, _036380_, _036381_, _036382_, _036383_, _036384_, _036385_, _036386_, _036387_, _036388_, _036389_, _036390_, _036391_, _036392_, _036393_, _036394_, _036395_, _036396_, _036397_, _036398_, _036399_, _036400_, _036401_, _036402_, _036403_, _036404_, _036405_, _036406_, _036407_, _036408_, _036409_, _036410_, _036411_, _036412_, _036413_, _036414_, _036415_, _036416_, _036417_, _036418_, _036419_, _036420_, _036421_, _036422_, _036423_, _036424_, _036425_, _036426_, _036427_, _036428_, _036429_, _036430_, _036431_, _036432_, _036433_, _036434_, _036435_, _036436_, _036437_, _036438_, _036439_, _036440_, _036441_, _036442_, _036443_, _036444_, _036445_, _036446_, _036447_, _036448_, _036449_, _036450_, _036451_, _036452_, _036453_, _036454_, _036455_, _036456_, _036457_, _036458_, _036459_, _036460_, _036461_, _036462_, _036463_, _036464_, _036465_, _036466_, _036467_, _036468_, _036469_, _036470_, _036471_, _036472_, _036473_, _036474_, _036475_, _036476_, _036477_, _036478_, _036479_, _036480_, _036481_, _036482_, _036483_, _036484_, _036485_, _036486_, _036487_, _036488_, _036489_, _036490_, _036491_, _036492_, _036493_, _036494_, _036495_, _036496_, _036497_, _036498_, _036499_, _036500_, _036501_, _036502_, _036503_, _036504_, _036505_, _036506_, _036507_, _036508_, _036509_, _036510_, _036511_, _036512_, _036513_, _036514_, _036515_, _036516_, _036517_, _036518_, _036519_, _036520_, _036521_, _036522_, _036523_, _036524_, _036525_, _036526_, _036527_, _036528_, _036529_, _036530_, _036531_, _036532_, _036533_, _036534_, _036535_, _036536_, _036537_, _036538_, _036539_, _036540_, _036541_, _036542_, _036543_, _036544_, _036545_, _036546_, _036547_, _036548_, _036549_, _036550_, _036551_, _036552_, _036553_, _036554_, _036555_, _036556_, _036557_, _036558_, _036559_, _036560_, _036561_, _036562_, _036563_, _036564_, _036565_, _036566_, _036567_, _036568_, _036569_, _036570_, _036571_, _036572_, _036573_, _036574_, _036575_, _036576_, _036577_, _036578_, _036579_, _036580_, _036581_, _036582_, _036583_, _036584_, _036585_, _036586_, _036587_, _036588_, _036589_, _036590_, _036591_, _036592_, _036593_, _036594_, _036595_, _036596_, _036597_, _036598_, _036599_, _036600_, _036601_, _036602_, _036603_, _036604_, _036605_, _036606_, _036607_, _036608_, _036609_, _036610_, _036611_, _036612_, _036613_, _036614_, _036615_, _036616_, _036617_, _036618_, _036619_, _036620_, _036621_, _036622_, _036623_, _036624_, _036625_, _036626_, _036627_, _036628_, _036629_, _036630_, _036631_, _036632_, _036633_, _036634_, _036635_, _036636_, _036637_, _036638_, _036639_, _036640_, _036641_, _036642_, _036643_, _036644_, _036645_, _036646_, _036647_, _036648_, _036649_, _036650_, _036651_, _036652_, _036653_, _036654_, _036655_, _036656_, _036657_, _036658_, _036659_, _036660_, _036661_, _036662_, _036663_, _036664_, _036665_, _036666_, _036667_, _036668_, _036669_, _036670_, _036671_, _036672_, _036673_, _036674_, _036675_, _036676_, _036677_, _036678_, _036679_, _036680_, _036681_, _036682_, _036683_, _036684_, _036685_, _036686_, _036687_, _036688_, _036689_, _036690_, _036691_, _036692_, _036693_, _036694_, _036695_, _036696_, _036697_, _036698_, _036699_, _036700_, _036701_, _036702_, _036703_, _036704_, _036705_, _036706_, _036707_, _036708_, _036709_, _036710_, _036711_, _036712_, _036713_, _036714_, _036715_, _036716_, _036717_, _036718_, _036719_, _036720_, _036721_, _036722_, _036723_, _036724_, _036725_, _036726_, _036727_, _036728_, _036729_, _036730_, _036731_, _036732_, _036733_, _036734_, _036735_, _036736_, _036737_, _036738_, _036739_, _036740_, _036741_, _036742_, _036743_, _036744_, _036745_, _036746_, _036747_, _036748_, _036749_, _036750_, _036751_, _036752_, _036753_, _036754_, _036755_, _036756_, _036757_, _036758_, _036759_, _036760_, _036761_, _036762_, _036763_, _036764_, _036765_, _036766_, _036767_, _036768_, _036769_, _036770_, _036771_, _036772_, _036773_, _036774_, _036775_, _036776_, _036777_, _036778_, _036779_, _036780_, _036781_, _036782_, _036783_, _036784_, _036785_, _036786_, _036787_, _036788_, _036789_, _036790_, _036791_, _036792_, _036793_, _036794_, _036795_, _036796_, _036797_, _036798_, _036799_, _036800_, _036801_, _036802_, _036803_, _036804_, _036805_, _036806_, _036807_, _036808_, _036809_, _036810_, _036811_, _036812_, _036813_, _036814_, _036815_, _036816_, _036817_, _036818_, _036819_, _036820_, _036821_, _036822_, _036823_, _036824_, _036825_, _036826_, _036827_, _036828_, _036829_, _036830_, _036831_, _036832_, _036833_, _036834_, _036835_, _036836_, _036837_, _036838_, _036839_, _036840_, _036841_, _036842_, _036843_, _036844_, _036845_, _036846_, _036847_, _036848_, _036849_, _036850_, _036851_, _036852_, _036853_, _036854_, _036855_, _036856_, _036857_, _036858_, _036859_, _036860_, _036861_, _036862_, _036863_, _036864_, _036865_, _036866_, _036867_, _036868_, _036869_, _036870_, _036871_, _036872_, _036873_, _036874_, _036875_, _036876_, _036877_, _036878_, _036879_, _036880_, _036881_, _036882_, _036883_, _036884_, _036885_, _036886_, _036887_, _036888_, _036889_, _036890_, _036891_, _036892_, _036893_, _036894_, _036895_, _036896_, _036897_, _036898_, _036899_, _036900_, _036901_, _036902_, _036903_, _036904_, _036905_, _036906_, _036907_, _036908_, _036909_, _036910_, _036911_, _036912_, _036913_, _036914_, _036915_, _036916_, _036917_, _036918_, _036919_, _036920_, _036921_, _036922_, _036923_, _036924_, _036925_, _036926_, _036927_, _036928_, _036929_, _036930_, _036931_, _036932_, _036933_, _036934_, _036935_, _036936_, _036937_, _036938_, _036939_, _036940_, _036941_, _036942_, _036943_, _036944_, _036945_, _036946_, _036947_, _036948_, _036949_, _036950_, _036951_, _036952_, _036953_, _036954_, _036955_, _036956_, _036957_, _036958_, _036959_, _036960_, _036961_, _036962_, _036963_, _036964_, _036965_, _036966_, _036967_, _036968_, _036969_, _036970_, _036971_, _036972_, _036973_, _036974_, _036975_, _036976_, _036977_, _036978_, _036979_, _036980_, _036981_, _036982_, _036983_, _036984_, _036985_, _036986_, _036987_, _036988_, _036989_, _036990_, _036991_, _036992_, _036993_, _036994_, _036995_, _036996_, _036997_, _036998_, _036999_, _037000_, _037001_, _037002_, _037003_, _037004_, _037005_, _037006_, _037007_, _037008_, _037009_, _037010_, _037011_, _037012_, _037013_, _037014_, _037015_, _037016_, _037017_, _037018_, _037019_, _037020_, _037021_, _037022_, _037023_, _037024_, _037025_, _037026_, _037027_, _037028_, _037029_, _037030_, _037031_, _037032_, _037033_, _037034_, _037035_, _037036_, _037037_, _037038_, _037039_, _037040_, _037041_, _037042_, _037043_, _037044_, _037045_, _037046_, _037047_, _037048_, _037049_, _037050_, _037051_, _037052_, _037053_, _037054_, _037055_, _037056_, _037057_, _037058_, _037059_, _037060_, _037061_, _037062_, _037063_, _037064_, _037065_, _037066_, _037067_, _037068_, _037069_, _037070_, _037071_, _037072_, _037073_, _037074_, _037075_, _037076_, _037077_, _037078_, _037079_, _037080_, _037081_, _037082_, _037083_, _037084_, _037085_, _037086_, _037087_, _037088_, _037089_, _037090_, _037091_, _037092_, _037093_, _037094_, _037095_, _037096_, _037097_, _037098_, _037099_, _037100_, _037101_, _037102_, _037103_, _037104_, _037105_, _037106_, _037107_, _037108_, _037109_, _037110_, _037111_, _037112_, _037113_, _037114_, _037115_, _037116_, _037117_, _037118_, _037119_, _037120_, _037121_, _037122_, _037123_, _037124_, _037125_, _037126_, _037127_, _037128_, _037129_, _037130_, _037131_, _037132_, _037133_, _037134_, _037135_, _037136_, _037137_, _037138_, _037139_, _037140_, _037141_, _037142_, _037143_, _037144_, _037145_, _037146_, _037147_, _037148_, _037149_, _037150_, _037151_, _037152_, _037153_, _037154_, _037155_, _037156_, _037157_, _037158_, _037159_, _037160_, _037161_, _037162_, _037163_, _037164_, _037165_, _037166_, _037167_, _037168_, _037169_, _037170_, _037171_, _037172_, _037173_, _037174_, _037175_, _037176_, _037177_, _037178_, _037179_, _037180_, _037181_, _037182_, _037183_, _037184_, _037185_, _037186_, _037187_, _037188_, _037189_, _037190_, _037191_, _037192_, _037193_, _037194_, _037195_, _037196_, _037197_, _037198_, _037199_, _037200_, _037201_, _037202_, _037203_, _037204_, _037205_, _037206_, _037207_, _037208_, _037209_, _037210_, _037211_, _037212_, _037213_, _037214_, _037215_, _037216_, _037217_, _037218_, _037219_, _037220_, _037221_, _037222_, _037223_, _037224_, _037225_, _037226_, _037227_, _037228_, _037229_, _037230_, _037231_, _037232_, _037233_, _037234_, _037235_, _037236_, _037237_, _037238_, _037239_, _037240_, _037241_, _037242_, _037243_, _037244_, _037245_, _037246_, _037247_, _037248_, _037249_, _037250_, _037251_, _037252_, _037253_, _037254_, _037255_, _037256_, _037257_, _037258_, _037259_, _037260_, _037261_, _037262_, _037263_, _037264_, _037265_, _037266_, _037267_, _037268_, _037269_, _037270_, _037271_, _037272_, _037273_, _037274_, _037275_, _037276_, _037277_, _037278_, _037279_, _037280_, _037281_, _037282_, _037283_, _037284_, _037285_, _037286_, _037287_, _037288_, _037289_, _037290_, _037291_, _037292_, _037293_, _037294_, _037295_, _037296_, _037297_, _037298_, _037299_, _037300_, _037301_, _037302_, _037303_, _037304_, _037305_, _037306_, _037307_, _037308_, _037309_, _037310_, _037311_, _037312_, _037313_, _037314_, _037315_, _037316_, _037317_, _037318_, _037319_, _037320_, _037321_, _037322_, _037323_, _037324_, _037325_, _037326_, _037327_, _037328_, _037329_, _037330_, _037331_, _037332_, _037333_, _037334_, _037335_, _037336_, _037337_, _037338_, _037339_, _037340_, _037341_, _037342_, _037343_, _037344_, _037345_, _037346_, _037347_, _037348_, _037349_, _037350_, _037351_, _037352_, _037353_, _037354_, _037355_, _037356_, _037357_, _037358_, _037359_, _037360_, _037361_, _037362_, _037363_, _037364_, _037365_, _037366_, _037367_, _037368_, _037369_, _037370_, _037371_, _037372_, _037373_, _037374_, _037375_, _037376_, _037377_, _037378_, _037379_, _037380_, _037381_, _037382_, _037383_, _037384_, _037385_, _037386_, _037387_, _037388_, _037389_, _037390_, _037391_, _037392_, _037393_, _037394_, _037395_, _037396_, _037397_, _037398_, _037399_, _037400_, _037401_, _037402_, _037403_, _037404_, _037405_, _037406_, _037407_, _037408_, _037409_, _037410_, _037411_, _037412_, _037413_, _037414_, _037415_, _037416_, _037417_, _037418_, _037419_, _037420_, _037421_, _037422_, _037423_, _037424_, _037425_, _037426_, _037427_, _037428_, _037429_, _037430_, _037431_, _037432_, _037433_, _037434_, _037435_, _037436_, _037437_, _037438_, _037439_, _037440_, _037441_, _037442_, _037443_, _037444_, _037445_, _037446_, _037447_, _037448_, _037449_, _037450_, _037451_, _037452_, _037453_, _037454_, _037455_, _037456_, _037457_, _037458_, _037459_, _037460_, _037461_, _037462_, _037463_, _037464_, _037465_, _037466_, _037467_, _037468_, _037469_, _037470_, _037471_, _037472_, _037473_, _037474_, _037475_, _037476_, _037477_, _037478_, _037479_, _037480_, _037481_, _037482_, _037483_, _037484_, _037485_, _037486_, _037487_, _037488_, _037489_, _037490_, _037491_, _037492_, _037493_, _037494_, _037495_, _037496_, _037497_, _037498_, _037499_, _037500_, _037501_, _037502_, _037503_, _037504_, _037505_, _037506_, _037507_, _037508_, _037509_, _037510_, _037511_, _037512_, _037513_, _037514_, _037515_, _037516_, _037517_, _037518_, _037519_, _037520_, _037521_, _037522_, _037523_, _037524_, _037525_, _037526_, _037527_, _037528_, _037529_, _037530_, _037531_, _037532_, _037533_, _037534_, _037535_, _037536_, _037537_, _037538_, _037539_, _037540_, _037541_, _037542_, _037543_, _037544_, _037545_, _037546_, _037547_, _037548_, _037549_, _037550_, _037551_, _037552_, _037553_, _037554_, _037555_, _037556_, _037557_, _037558_, _037559_, _037560_, _037561_, _037562_, _037563_, _037564_, _037565_, _037566_, _037567_, _037568_, _037569_, _037570_, _037571_, _037572_, _037573_, _037574_, _037575_, _037576_, _037577_, _037578_, _037579_, _037580_, _037581_, _037582_, _037583_, _037584_, _037585_, _037586_, _037587_, _037588_, _037589_, _037590_, _037591_, _037592_, _037593_, _037594_, _037595_, _037596_, _037597_, _037598_, _037599_, _037600_, _037601_, _037602_, _037603_, _037604_, _037605_, _037606_, _037607_, _037608_, _037609_, _037610_, _037611_, _037612_, _037613_, _037614_, _037615_, _037616_, _037617_, _037618_, _037619_, _037620_, _037621_, _037622_, _037623_, _037624_, _037625_, _037626_, _037627_, _037628_, _037629_, _037630_, _037631_, _037632_, _037633_, _037634_, _037635_, _037636_, _037637_, _037638_, _037639_, _037640_, _037641_, _037642_, _037643_, _037644_, _037645_, _037646_, _037647_, _037648_, _037649_, _037650_, _037651_, _037652_, _037653_, _037654_, _037655_, _037656_, _037657_, _037658_, _037659_, _037660_, _037661_, _037662_, _037663_, _037664_, _037665_, _037666_, _037667_, _037668_, _037669_, _037670_, _037671_, _037672_, _037673_, _037674_, _037675_, _037676_, _037677_, _037678_, _037679_, _037680_, _037681_, _037682_, _037683_, _037684_, _037685_, _037686_, _037687_, _037688_, _037689_, _037690_, _037691_, _037692_, _037693_, _037694_, _037695_, _037696_, _037697_, _037698_, _037699_, _037700_, _037701_, _037702_, _037703_, _037704_, _037705_, _037706_, _037707_, _037708_, _037709_, _037710_, _037711_, _037712_, _037713_, _037714_, _037715_, _037716_, _037717_, _037718_, _037719_, _037720_, _037721_, _037722_, _037723_, _037724_, _037725_, _037726_, _037727_, _037728_, _037729_, _037730_, _037731_, _037732_, _037733_, _037734_, _037735_, _037736_, _037737_, _037738_, _037739_, _037740_, _037741_, _037742_, _037743_, _037744_, _037745_, _037746_, _037747_, _037748_, _037749_, _037750_, _037751_, _037752_, _037753_, _037754_, _037755_, _037756_, _037757_, _037758_, _037759_, _037760_, _037761_, _037762_, _037763_, _037764_, _037765_, _037766_, _037767_, _037768_, _037769_, _037770_, _037771_, _037772_, _037773_, _037774_, _037775_, _037776_, _037777_, _037778_, _037779_, _037780_, _037781_, _037782_, _037783_, _037784_, _037785_, _037786_, _037787_, _037788_, _037789_, _037790_, _037791_, _037792_, _037793_, _037794_, _037795_, _037796_, _037797_, _037798_, _037799_, _037800_, _037801_, _037802_, _037803_, _037804_, _037805_, _037806_, _037807_, _037808_, _037809_, _037810_, _037811_, _037812_, _037813_, _037814_, _037815_, _037816_, _037817_, _037818_, _037819_, _037820_, _037821_, _037822_, _037823_, _037824_, _037825_, _037826_, _037827_, _037828_, _037829_, _037830_, _037831_, _037832_, _037833_, _037834_, _037835_, _037836_, _037837_, _037838_, _037839_, _037840_, _037841_, _037842_, _037843_, _037844_, _037845_, _037846_, _037847_, _037848_, _037849_, _037850_, _037851_, _037852_, _037853_, _037854_, _037855_, _037856_, _037857_, _037858_, _037859_, _037860_, _037861_, _037862_, _037863_, _037864_, _037865_, _037866_, _037867_, _037868_, _037869_, _037870_, _037871_, _037872_, _037873_, _037874_, _037875_, _037876_, _037877_, _037878_, _037879_, _037880_, _037881_, _037882_, _037883_, _037884_, _037885_, _037886_, _037887_, _037888_, _037889_, _037890_, _037891_, _037892_, _037893_, _037894_, _037895_, _037896_, _037897_, _037898_, _037899_, _037900_, _037901_, _037902_, _037903_, _037904_, _037905_, _037906_, _037907_, _037908_, _037909_, _037910_, _037911_, _037912_, _037913_, _037914_, _037915_, _037916_, _037917_, _037918_, _037919_, _037920_, _037921_, _037922_, _037923_, _037924_, _037925_, _037926_, _037927_, _037928_, _037929_, _037930_, _037931_, _037932_, _037933_, _037934_, _037935_, _037936_, _037937_, _037938_, _037939_, _037940_, _037941_, _037942_, _037943_, _037944_, _037945_, _037946_, _037947_, _037948_, _037949_, _037950_, _037951_, _037952_, _037953_, _037954_, _037955_, _037956_, _037957_, _037958_, _037959_, _037960_, _037961_, _037962_, _037963_, _037964_, _037965_, _037966_, _037967_, _037968_, _037969_, _037970_, _037971_, _037972_, _037973_, _037974_, _037975_, _037976_, _037977_, _037978_, _037979_, _037980_, _037981_, _037982_, _037983_, _037984_, _037985_, _037986_, _037987_, _037988_, _037989_, _037990_, _037991_, _037992_, _037993_, _037994_, _037995_, _037996_, _037997_, _037998_, _037999_, _038000_, _038001_, _038002_, _038003_, _038004_, _038005_, _038006_, _038007_, _038008_, _038009_, _038010_, _038011_, _038012_, _038013_, _038014_, _038015_, _038016_, _038017_, _038018_, _038019_, _038020_, _038021_, _038022_, _038023_, _038024_, _038025_, _038026_, _038027_, _038028_, _038029_, _038030_, _038031_, _038032_, _038033_, _038034_, _038035_, _038036_, _038037_, _038038_, _038039_, _038040_, _038041_, _038042_, _038043_, _038044_, _038045_, _038046_, _038047_, _038048_, _038049_, _038050_, _038051_, _038052_, _038053_, _038054_, _038055_, _038056_, _038057_, _038058_, _038059_, _038060_, _038061_, _038062_, _038063_, _038064_, _038065_, _038066_, _038067_, _038068_, _038069_, _038070_, _038071_, _038072_, _038073_, _038074_, _038075_, _038076_, _038077_, _038078_, _038079_, _038080_, _038081_, _038082_, _038083_, _038084_, _038085_, _038086_, _038087_, _038088_, _038089_, _038090_, _038091_, _038092_, _038093_, _038094_, _038095_, _038096_, _038097_, _038098_, _038099_, _038100_, _038101_, _038102_, _038103_, _038104_, _038105_, _038106_, _038107_, _038108_, _038109_, _038110_, _038111_, _038112_, _038113_, _038114_, _038115_, _038116_, _038117_, _038118_, _038119_, _038120_, _038121_, _038122_, _038123_, _038124_, _038125_, _038126_, _038127_, _038128_, _038129_, _038130_, _038131_, _038132_, _038133_, _038134_, _038135_, _038136_, _038137_, _038138_, _038139_, _038140_, _038141_, _038142_, _038143_, _038144_, _038145_, _038146_, _038147_, _038148_, _038149_, _038150_, _038151_, _038152_, _038153_, _038154_, _038155_, _038156_, _038157_, _038158_, _038159_, _038160_, _038161_, _038162_, _038163_, _038164_, _038165_, _038166_, _038167_, _038168_, _038169_, _038170_, _038171_, _038172_, _038173_, _038174_, _038175_, _038176_, _038177_, _038178_, _038179_, _038180_, _038181_, _038182_, _038183_, _038184_, _038185_, _038186_, _038187_, _038188_, _038189_, _038190_, _038191_, _038192_, _038193_, _038194_, _038195_, _038196_, _038197_, _038198_, _038199_, _038200_, _038201_, _038202_, _038203_, _038204_, _038205_, _038206_, _038207_, _038208_, _038209_, _038210_, _038211_, _038212_, _038213_, _038214_, _038215_, _038216_, _038217_, _038218_, _038219_, _038220_, _038221_, _038222_, _038223_, _038224_, _038225_, _038226_, _038227_, _038228_, _038229_, _038230_, _038231_, _038232_, _038233_, _038234_, _038235_, _038236_, _038237_, _038238_, _038239_, _038240_, _038241_, _038242_, _038243_, _038244_, _038245_, _038246_, _038247_, _038248_, _038249_, _038250_, _038251_, _038252_, _038253_, _038254_, _038255_, _038256_, _038257_, _038258_, _038259_, _038260_, _038261_, _038262_, _038263_, _038264_, _038265_, _038266_, _038267_, _038268_, _038269_, _038270_, _038271_, _038272_, _038273_, _038274_, _038275_, _038276_, _038277_, _038278_, _038279_, _038280_, _038281_, _038282_, _038283_, _038284_, _038285_, _038286_, _038287_, _038288_, _038289_, _038290_, _038291_, _038292_, _038293_, _038294_, _038295_, _038296_, _038297_, _038298_, _038299_, _038300_, _038301_, _038302_, _038303_, _038304_, _038305_, _038306_, _038307_, _038308_, _038309_, _038310_, _038311_, _038312_, _038313_, _038314_, _038315_, _038316_, _038317_, _038318_, _038319_, _038320_, _038321_, _038322_, _038323_, _038324_, _038325_, _038326_, _038327_, _038328_, _038329_, _038330_, _038331_, _038332_, _038333_, _038334_, _038335_, _038336_, _038337_, _038338_, _038339_, _038340_, _038341_, _038342_, _038343_, _038344_, _038345_, _038346_, _038347_, _038348_, _038349_, _038350_, _038351_, _038352_, _038353_, _038354_, _038355_, _038356_, _038357_, _038358_, _038359_, _038360_, _038361_, _038362_, _038363_, _038364_, _038365_, _038366_, _038367_, _038368_, _038369_, _038370_, _038371_, _038372_, _038373_, _038374_, _038375_, _038376_, _038377_, _038378_, _038379_, _038380_, _038381_, _038382_, _038383_, _038384_, _038385_, _038386_, _038387_, _038388_, _038389_, _038390_, _038391_, _038392_, _038393_, _038394_, _038395_, _038396_, _038397_, _038398_, _038399_, _038400_, _038401_, _038402_, _038403_, _038404_, _038405_, _038406_, _038407_, _038408_, _038409_, _038410_, _038411_, _038412_, _038413_, _038414_, _038415_, _038416_, _038417_, _038418_, _038419_, _038420_, _038421_, _038422_, _038423_, _038424_, _038425_, _038426_, _038427_, _038428_, _038429_, _038430_, _038431_, _038432_, _038433_, _038434_, _038435_, _038436_, _038437_, _038438_, _038439_, _038440_, _038441_, _038442_, _038443_, _038444_, _038445_, _038446_, _038447_, _038448_, _038449_, _038450_, _038451_, _038452_, _038453_, _038454_, _038455_, _038456_, _038457_, _038458_, _038459_, _038460_, _038461_, _038462_, _038463_, _038464_, _038465_, _038466_, _038467_, _038468_, _038469_, _038470_, _038471_, _038472_, _038473_, _038474_, _038475_, _038476_, _038477_, _038478_, _038479_, _038480_, _038481_, _038482_, _038483_, _038484_, _038485_, _038486_, _038487_, _038488_, _038489_, _038490_, _038491_, _038492_, _038493_, _038494_, _038495_, _038496_, _038497_, _038498_, _038499_, _038500_, _038501_, _038502_, _038503_, _038504_, _038505_, _038506_, _038507_, _038508_, _038509_, _038510_, _038511_, _038512_, _038513_, _038514_, _038515_, _038516_, _038517_, _038518_, _038519_, _038520_, _038521_, _038522_, _038523_, _038524_, _038525_, _038526_, _038527_, _038528_, _038529_, _038530_, _038531_, _038532_, _038533_, _038534_, _038535_, _038536_, _038537_, _038538_, _038539_, _038540_, _038541_, _038542_, _038543_, _038544_, _038545_, _038546_, _038547_, _038548_, _038549_, _038550_, _038551_, _038552_, _038553_, _038554_, _038555_, _038556_, _038557_, _038558_, _038559_, _038560_, _038561_, _038562_, _038563_, _038564_, _038565_, _038566_, _038567_, _038568_, _038569_, _038570_, _038571_, _038572_, _038573_, _038574_, _038575_, _038576_, _038577_, _038578_, _038579_, _038580_, _038581_, _038582_, _038583_, _038584_, _038585_, _038586_, _038587_, _038588_, _038589_, _038590_, _038591_, _038592_, _038593_, _038594_, _038595_, _038596_, _038597_, _038598_, _038599_, _038600_, _038601_, _038602_, _038603_, _038604_, _038605_, _038606_, _038607_, _038608_, _038609_, _038610_, _038611_, _038612_, _038613_, _038614_, _038615_, _038616_, _038617_, _038618_, _038619_, _038620_, _038621_, _038622_, _038623_, _038624_, _038625_, _038626_, _038627_, _038628_, _038629_, _038630_, _038631_, _038632_, _038633_, _038634_, _038635_, _038636_, _038637_, _038638_, _038639_, _038640_, _038641_, _038642_, _038643_, _038644_, _038645_, _038646_, _038647_, _038648_, _038649_, _038650_, _038651_, _038652_, _038653_, _038654_, _038655_, _038656_, _038657_, _038658_, _038659_, _038660_, _038661_, _038662_, _038663_, _038664_, _038665_, _038666_, _038667_, _038668_, _038669_, _038670_, _038671_, _038672_, _038673_, _038674_, _038675_, _038676_, _038677_, _038678_, _038679_, _038680_, _038681_, _038682_, _038683_, _038684_, _038685_, _038686_, _038687_, _038688_, _038689_, _038690_, _038691_, _038692_, _038693_, _038694_, _038695_, _038696_, _038697_, _038698_, _038699_, _038700_, _038701_, _038702_, _038703_, _038704_, _038705_, _038706_, _038707_, _038708_, _038709_, _038710_, _038711_, _038712_, _038713_, _038714_, _038715_, _038716_, _038717_, _038718_, _038719_, _038720_, _038721_, _038722_, _038723_, _038724_, _038725_, _038726_, _038727_, _038728_, _038729_, _038730_, _038731_, _038732_, _038733_, _038734_, _038735_, _038736_, _038737_, _038738_, _038739_, _038740_, _038741_, _038742_, _038743_, _038744_, _038745_, _038746_, _038747_, _038748_, _038749_, _038750_, _038751_, _038752_, _038753_, _038754_, _038755_, _038756_, _038757_, _038758_, _038759_, _038760_, _038761_, _038762_, _038763_, _038764_, _038765_, _038766_, _038767_, _038768_, _038769_, _038770_, _038771_, _038772_, _038773_, _038774_, _038775_, _038776_, _038777_, _038778_, _038779_, _038780_, _038781_, _038782_, _038783_, _038784_, _038785_, _038786_, _038787_, _038788_, _038789_, _038790_, _038791_, _038792_, _038793_, _038794_, _038795_, _038796_, _038797_, _038798_, _038799_, _038800_, _038801_, _038802_, _038803_, _038804_, _038805_, _038806_, _038807_, _038808_, _038809_, _038810_, _038811_, _038812_, _038813_, _038814_, _038815_, _038816_, _038817_, _038818_, _038819_, _038820_, _038821_, _038822_, _038823_, _038824_, _038825_, _038826_, _038827_, _038828_, _038829_, _038830_, _038831_, _038832_, _038833_, _038834_, _038835_, _038836_, _038837_, _038838_, _038839_, _038840_, _038841_, _038842_, _038843_, _038844_, _038845_, _038846_, _038847_, _038848_, _038849_, _038850_, _038851_, _038852_, _038853_, _038854_, _038855_, _038856_, _038857_, _038858_, _038859_, _038860_, _038861_, _038862_, _038863_, _038864_, _038865_, _038866_, _038867_, _038868_, _038869_, _038870_, _038871_, _038872_, _038873_, _038874_, _038875_, _038876_, _038877_, _038878_, _038879_, _038880_, _038881_, _038882_, _038883_, _038884_, _038885_, _038886_, _038887_, _038888_, _038889_, _038890_, _038891_, _038892_, _038893_, _038894_, _038895_, _038896_, _038897_, _038898_, _038899_, _038900_, _038901_, _038902_, _038903_, _038904_, _038905_, _038906_, _038907_, _038908_, _038909_, _038910_, _038911_, _038912_, _038913_, _038914_, _038915_, _038916_, _038917_, _038918_, _038919_, _038920_, _038921_, _038922_, _038923_, _038924_, _038925_, _038926_, _038927_, _038928_, _038929_, _038930_, _038931_, _038932_, _038933_, _038934_, _038935_, _038936_, _038937_, _038938_, _038939_, _038940_, _038941_, _038942_, _038943_, _038944_, _038945_, _038946_, _038947_, _038948_, _038949_, _038950_, _038951_, _038952_, _038953_, _038954_, _038955_, _038956_, _038957_, _038958_, _038959_, _038960_, _038961_, _038962_, _038963_, _038964_, _038965_, _038966_, _038967_, _038968_, _038969_, _038970_, _038971_, _038972_, _038973_, _038974_, _038975_, _038976_, _038977_, _038978_, _038979_, _038980_, _038981_, _038982_, _038983_, _038984_, _038985_, _038986_, _038987_, _038988_, _038989_, _038990_, _038991_, _038992_, _038993_, _038994_, _038995_, _038996_, _038997_, _038998_, _038999_, _039000_, _039001_, _039002_, _039003_, _039004_, _039005_, _039006_, _039007_, _039008_, _039009_, _039010_, _039011_, _039012_, _039013_, _039014_, _039015_, _039016_, _039017_, _039018_, _039019_, _039020_, _039021_, _039022_, _039023_, _039024_, _039025_, _039026_, _039027_, _039028_, _039029_, _039030_, _039031_, _039032_, _039033_, _039034_, _039035_, _039036_, _039037_, _039038_, _039039_, _039040_, _039041_, _039042_, _039043_, _039044_, _039045_, _039046_, _039047_, _039048_, _039049_, _039050_, _039051_, _039052_, _039053_, _039054_, _039055_, _039056_, _039057_, _039058_, _039059_, _039060_, _039061_, _039062_, _039063_, _039064_, _039065_, _039066_, _039067_, _039068_, _039069_, _039070_, _039071_, _039072_, _039073_, _039074_, _039075_, _039076_, _039077_, _039078_, _039079_, _039080_, _039081_, _039082_, _039083_, _039084_, _039085_, _039086_, _039087_, _039088_, _039089_, _039090_, _039091_, _039092_, _039093_, _039094_, _039095_, _039096_, _039097_, _039098_, _039099_, _039100_, _039101_, _039102_, _039103_, _039104_, _039105_, _039106_, _039107_, _039108_, _039109_, _039110_, _039111_, _039112_, _039113_, _039114_, _039115_, _039116_, _039117_, _039118_, _039119_, _039120_, _039121_, _039122_, _039123_, _039124_, _039125_, _039126_, _039127_, _039128_, _039129_, _039130_, _039131_, _039132_, _039133_, _039134_, _039135_, _039136_, _039137_, _039138_, _039139_, _039140_, _039141_, _039142_, _039143_, _039144_, _039145_, _039146_, _039147_, _039148_, _039149_, _039150_, _039151_, _039152_, _039153_, _039154_, _039155_, _039156_, _039157_, _039158_, _039159_, _039160_, _039161_, _039162_, _039163_, _039164_, _039165_, _039166_, _039167_, _039168_, _039169_, _039170_, _039171_, _039172_, _039173_, _039174_, _039175_, _039176_, _039177_, _039178_, _039179_, _039180_, _039181_, _039182_, _039183_, _039184_, _039185_, _039186_, _039187_, _039188_, _039189_, _039190_, _039191_, _039192_, _039193_, _039194_, _039195_, _039196_, _039197_, _039198_, _039199_, _039200_, _039201_, _039202_, _039203_, _039204_, _039205_, _039206_, _039207_, _039208_, _039209_, _039210_, _039211_, _039212_, _039213_, _039214_, _039215_, _039216_, _039217_, _039218_, _039219_, _039220_, _039221_, _039222_, _039223_, _039224_, _039225_, _039226_, _039227_, _039228_, _039229_, _039230_, _039231_, _039232_, _039233_, _039234_, _039235_, _039236_, _039237_, _039238_, _039239_, _039240_, _039241_, _039242_, _039243_, _039244_, _039245_, _039246_, _039247_, _039248_, _039249_, _039250_, _039251_, _039252_, _039253_, _039254_, _039255_, _039256_, _039257_, _039258_, _039259_, _039260_, _039261_, _039262_, _039263_, _039264_, _039265_, _039266_, _039267_, _039268_, _039269_, _039270_, _039271_, _039272_, _039273_, _039274_, _039275_, _039276_, _039277_, _039278_, _039279_, _039280_, _039281_, _039282_, _039283_, _039284_, _039285_, _039286_, _039287_, _039288_, _039289_, _039290_, _039291_, _039292_, _039293_, _039294_, _039295_, _039296_, _039297_, _039298_, _039299_, _039300_, _039301_, _039302_, _039303_, _039304_, _039305_, _039306_, _039307_, _039308_, _039309_, _039310_, _039311_, _039312_, _039313_, _039314_, _039315_, _039316_, _039317_, _039318_, _039319_, _039320_, _039321_, _039322_, _039323_, _039324_, _039325_, _039326_, _039327_, _039328_, _039329_, _039330_, _039331_, _039332_, _039333_, _039334_, _039335_, _039336_, _039337_, _039338_, _039339_, _039340_, _039341_, _039342_, _039343_, _039344_, _039345_, _039346_, _039347_, _039348_, _039349_, _039350_, _039351_, _039352_, _039353_, _039354_, _039355_, _039356_, _039357_, _039358_, _039359_, _039360_, _039361_, _039362_, _039363_, _039364_, _039365_, _039366_, _039367_, _039368_, _039369_, _039370_, _039371_, _039372_, _039373_, _039374_, _039375_, _039376_, _039377_, _039378_, _039379_, _039380_, _039381_, _039382_, _039383_, _039384_, _039385_, _039386_, _039387_, _039388_, _039389_, _039390_, _039391_, _039392_, _039393_, _039394_, _039395_, _039396_, _039397_, _039398_, _039399_, _039400_, _039401_, _039402_, _039403_, _039404_, _039405_, _039406_, _039407_, _039408_, _039409_, _039410_, _039411_, _039412_, _039413_, _039414_, _039415_, _039416_, _039417_, _039418_, _039419_, _039420_, _039421_, _039422_, _039423_, _039424_, _039425_, _039426_, _039427_, _039428_, _039429_, _039430_, _039431_, _039432_, _039433_, _039434_, _039435_, _039436_, _039437_, _039438_, _039439_, _039440_, _039441_, _039442_, _039443_, _039444_, _039445_, _039446_, _039447_, _039448_, _039449_, _039450_, _039451_, _039452_, _039453_, _039454_, _039455_, _039456_, _039457_, _039458_, _039459_, _039460_, _039461_, _039462_, _039463_, _039464_, _039465_, _039466_, _039467_, _039468_, _039469_, _039470_, _039471_, _039472_, _039473_, _039474_, _039475_, _039476_, _039477_, _039478_, _039479_, _039480_, _039481_, _039482_, _039483_, _039484_, _039485_, _039486_, _039487_, _039488_, _039489_, _039490_, _039491_, _039492_, _039493_, _039494_, _039495_, _039496_, _039497_, _039498_, _039499_, _039500_, _039501_, _039502_, _039503_, _039504_, _039505_, _039506_, _039507_, _039508_, _039509_, _039510_, _039511_, _039512_, _039513_, _039514_, _039515_, _039516_, _039517_, _039518_, _039519_, _039520_, _039521_, _039522_, _039523_, _039524_, _039525_, _039526_, _039527_, _039528_, _039529_, _039530_, _039531_, _039532_, _039533_, _039534_, _039535_, _039536_, _039537_, _039538_, _039539_, _039540_, _039541_, _039542_, _039543_, _039544_, _039545_, _039546_, _039547_, _039548_, _039549_, _039550_, _039551_, _039552_, _039553_, _039554_, _039555_, _039556_, _039557_, _039558_, _039559_, _039560_, _039561_, _039562_, _039563_, _039564_, _039565_, _039566_, _039567_, _039568_, _039569_, _039570_, _039571_, _039572_, _039573_, _039574_, _039575_, _039576_, _039577_, _039578_, _039579_, _039580_, _039581_, _039582_, _039583_, _039584_, _039585_, _039586_, _039587_, _039588_, _039589_, _039590_, _039591_, _039592_, _039593_, _039594_, _039595_, _039596_, _039597_, _039598_, _039599_, _039600_, _039601_, _039602_, _039603_, _039604_, _039605_, _039606_, _039607_, _039608_, _039609_, _039610_, _039611_, _039612_, _039613_, _039614_, _039615_, _039616_, _039617_, _039618_, _039619_, _039620_, _039621_, _039622_, _039623_, _039624_, _039625_, _039626_, _039627_, _039628_, _039629_, _039630_, _039631_, _039632_, _039633_, _039634_, _039635_, _039636_, _039637_, _039638_, _039639_, _039640_, _039641_, _039642_, _039643_, _039644_, _039645_, _039646_, _039647_, _039648_, _039649_, _039650_, _039651_, _039652_, _039653_, _039654_, _039655_, _039656_, _039657_, _039658_, _039659_, _039660_, _039661_, _039662_, _039663_, _039664_, _039665_, _039666_, _039667_, _039668_, _039669_, _039670_, _039671_, _039672_, _039673_, _039674_, _039675_, _039676_, _039677_, _039678_, _039679_, _039680_, _039681_, _039682_, _039683_, _039684_, _039685_, _039686_, _039687_, _039688_, _039689_, _039690_, _039691_, _039692_, _039693_, _039694_, _039695_, _039696_, _039697_, _039698_, _039699_, _039700_, _039701_, _039702_, _039703_, _039704_, _039705_, _039706_, _039707_, _039708_, _039709_, _039710_, _039711_, _039712_, _039713_, _039714_, _039715_, _039716_, _039717_, _039718_, _039719_, _039720_, _039721_, _039722_, _039723_, _039724_, _039725_, _039726_, _039727_, _039728_, _039729_, _039730_, _039731_, _039732_, _039733_, _039734_, _039735_, _039736_, _039737_, _039738_, _039739_, _039740_, _039741_, _039742_, _039743_, _039744_, _039745_, _039746_, _039747_, _039748_, _039749_, _039750_, _039751_, _039752_, _039753_, _039754_, _039755_, _039756_, _039757_, _039758_, _039759_, _039760_, _039761_, _039762_, _039763_, _039764_, _039765_, _039766_, _039767_, _039768_, _039769_, _039770_, _039771_, _039772_, _039773_, _039774_, _039775_, _039776_, _039777_, _039778_, _039779_, _039780_, _039781_, _039782_, _039783_, _039784_, _039785_, _039786_, _039787_, _039788_, _039789_, _039790_, _039791_, _039792_, _039793_, _039794_, _039795_, _039796_, _039797_, _039798_, _039799_, _039800_, _039801_, _039802_, _039803_, _039804_, _039805_, _039806_, _039807_, _039808_, _039809_, _039810_, _039811_, _039812_, _039813_, _039814_, _039815_, _039816_, _039817_, _039818_, _039819_, _039820_, _039821_, _039822_, _039823_, _039824_, _039825_, _039826_, _039827_, _039828_, _039829_, _039830_, _039831_, _039832_, _039833_, _039834_, _039835_, _039836_, _039837_, _039838_, _039839_, _039840_, _039841_, _039842_, _039843_, _039844_, _039845_, _039846_, _039847_, _039848_, _039849_, _039850_, _039851_, _039852_, _039853_, _039854_, _039855_, _039856_, _039857_, _039858_, _039859_, _039860_, _039861_, _039862_, _039863_, _039864_, _039865_, _039866_, _039867_, _039868_, _039869_, _039870_, _039871_, _039872_, _039873_, _039874_, _039875_, _039876_, _039877_, _039878_, _039879_, _039880_, _039881_, _039882_, _039883_, _039884_, _039885_, _039886_, _039887_, _039888_, _039889_, _039890_, _039891_, _039892_, _039893_, _039894_, _039895_, _039896_, _039897_, _039898_, _039899_, _039900_, _039901_, _039902_, _039903_, _039904_, _039905_, _039906_, _039907_, _039908_, _039909_, _039910_, _039911_, _039912_, _039913_, _039914_, _039915_, _039916_, _039917_, _039918_, _039919_, _039920_, _039921_, _039922_, _039923_, _039924_, _039925_, _039926_, _039927_, _039928_, _039929_, _039930_, _039931_, _039932_, _039933_, _039934_, _039935_, _039936_, _039937_, _039938_, _039939_, _039940_, _039941_, _039942_, _039943_, _039944_, _039945_, _039946_, _039947_, _039948_, _039949_, _039950_, _039951_, _039952_, _039953_, _039954_, _039955_, _039956_, _039957_, _039958_, _039959_, _039960_, _039961_, _039962_, _039963_, _039964_, _039965_, _039966_, _039967_, _039968_, _039969_, _039970_, _039971_, _039972_, _039973_, _039974_, _039975_, _039976_, _039977_, _039978_, _039979_, _039980_, _039981_, _039982_, _039983_, _039984_, _039985_, _039986_, _039987_, _039988_, _039989_, _039990_, _039991_, _039992_, _039993_, _039994_, _039995_, _039996_, _039997_, _039998_, _039999_, _040000_, _040001_, _040002_, _040003_, _040004_, _040005_, _040006_, _040007_, _040008_, _040009_, _040010_, _040011_, _040012_, _040013_, _040014_, _040015_, _040016_, _040017_, _040018_, _040019_, _040020_, _040021_, _040022_, _040023_, _040024_, _040025_, _040026_, _040027_, _040028_, _040029_, _040030_, _040031_, _040032_, _040033_, _040034_, _040035_, _040036_, _040037_, _040038_, _040039_, _040040_, _040041_, _040042_, _040043_, _040044_, _040045_, _040046_, _040047_, _040048_, _040049_, _040050_, _040051_, _040052_, _040053_, _040054_, _040055_, _040056_, _040057_, _040058_, _040059_, _040060_, _040061_, _040062_, _040063_, _040064_, _040065_, _040066_, _040067_, _040068_, _040069_, _040070_, _040071_, _040072_, _040073_, _040074_, _040075_, _040076_, _040077_, _040078_, _040079_, _040080_, _040081_, _040082_, _040083_, _040084_, _040085_, _040086_, _040087_, _040088_, _040089_, _040090_, _040091_, _040092_, _040093_, _040094_, _040095_, _040096_, _040097_, _040098_, _040099_, _040100_, _040101_, _040102_, _040103_, _040104_, _040105_, _040106_, _040107_, _040108_, _040109_, _040110_, _040111_, _040112_, _040113_, _040114_, _040115_, _040116_, _040117_, _040118_, _040119_, _040120_, _040121_, _040122_, _040123_, _040124_, _040125_, _040126_, _040127_, _040128_, _040129_, _040130_, _040131_, _040132_, _040133_, _040134_, _040135_, _040136_, _040137_, _040138_, _040139_, _040140_, _040141_, _040142_, _040143_, _040144_, _040145_, _040146_, _040147_, _040148_, _040149_, _040150_, _040151_, _040152_, _040153_, _040154_, _040155_, _040156_, _040157_, _040158_, _040159_, _040160_, _040161_, _040162_, _040163_, _040164_, _040165_, _040166_, _040167_, _040168_, _040169_, _040170_, _040171_, _040172_, _040173_, _040174_, _040175_, _040176_, _040177_, _040178_, _040179_, _040180_, _040181_, _040182_, _040183_, _040184_, _040185_, _040186_, _040187_, _040188_, _040189_, _040190_, _040191_, _040192_, _040193_, _040194_, _040195_, _040196_, _040197_, _040198_, _040199_, _040200_, _040201_, _040202_, _040203_, _040204_, _040205_, _040206_, _040207_, _040208_, _040209_, _040210_, _040211_, _040212_, _040213_, _040214_, _040215_, _040216_, _040217_, _040218_, _040219_, _040220_, _040221_, _040222_, _040223_, _040224_, _040225_, _040226_, _040227_, _040228_, _040229_, _040230_, _040231_, _040232_, _040233_, _040234_, _040235_, _040236_, _040237_, _040238_, _040239_, _040240_, _040241_, _040242_, _040243_, _040244_, _040245_, _040246_, _040247_, _040248_, _040249_, _040250_, _040251_, _040252_, _040253_, _040254_, _040255_, _040256_, _040257_, _040258_, _040259_, _040260_, _040261_, _040262_, _040263_, _040264_, _040265_, _040266_, _040267_, _040268_, _040269_, _040270_, _040271_, _040272_, _040273_, _040274_, _040275_, _040276_, _040277_, _040278_, _040279_, _040280_, _040281_, _040282_, _040283_, _040284_, _040285_, _040286_, _040287_, _040288_, _040289_, _040290_, _040291_, _040292_, _040293_, _040294_, _040295_, _040296_, _040297_, _040298_, _040299_, _040300_, _040301_, _040302_, _040303_, _040304_, _040305_, _040306_, _040307_, _040308_, _040309_, _040310_, _040311_, _040312_, _040313_, _040314_, _040315_, _040316_, _040317_, _040318_, _040319_, _040320_, _040321_, _040322_, _040323_, _040324_, _040325_, _040326_, _040327_, _040328_, _040329_, _040330_, _040331_, _040332_, _040333_, _040334_, _040335_, _040336_, _040337_, _040338_, _040339_, _040340_, _040341_, _040342_, _040343_, _040344_, _040345_, _040346_, _040347_, _040348_, _040349_, _040350_, _040351_, _040352_, _040353_, _040354_, _040355_, _040356_, _040357_, _040358_, _040359_, _040360_, _040361_, _040362_, _040363_, _040364_, _040365_, _040366_, _040367_, _040368_, _040369_, _040370_, _040371_, _040372_, _040373_, _040374_, _040375_, _040376_, _040377_, _040378_, _040379_, _040380_, _040381_, _040382_, _040383_, _040384_, _040385_, _040386_, _040387_, _040388_, _040389_, _040390_, _040391_, _040392_, _040393_, _040394_, _040395_, _040396_, _040397_, _040398_, _040399_, _040400_, _040401_, _040402_, _040403_, _040404_, _040405_, _040406_, _040407_, _040408_, _040409_, _040410_, _040411_, _040412_, _040413_, _040414_, _040415_, _040416_, _040417_, _040418_, _040419_, _040420_, _040421_, _040422_, _040423_, _040424_, _040425_, _040426_, _040427_, _040428_, _040429_, _040430_, _040431_, _040432_, _040433_, _040434_, _040435_, _040436_, _040437_, _040438_, _040439_, _040440_, _040441_, _040442_, _040443_, _040444_, _040445_, _040446_, _040447_, _040448_, _040449_, _040450_, _040451_, _040452_, _040453_, _040454_, _040455_, _040456_, _040457_, _040458_, _040459_, _040460_, _040461_, _040462_, _040463_, _040464_, _040465_, _040466_, _040467_, _040468_, _040469_, _040470_, _040471_, _040472_, _040473_, _040474_, _040475_, _040476_, _040477_, _040478_, _040479_, _040480_, _040481_, _040482_, _040483_, _040484_, _040485_, _040486_, _040487_, _040488_, _040489_, _040490_, _040491_, _040492_, _040493_, _040494_, _040495_, _040496_, _040497_, _040498_, _040499_, _040500_, _040501_, _040502_, _040503_, _040504_, _040505_, _040506_, _040507_, _040508_, _040509_, _040510_, _040511_, _040512_, _040513_, _040514_, _040515_, _040516_, _040517_, _040518_, _040519_, _040520_, _040521_, _040522_, _040523_, _040524_, _040525_, _040526_, _040527_, _040528_, _040529_, _040530_, _040531_, _040532_, _040533_, _040534_, _040535_, _040536_, _040537_, _040538_, _040539_, _040540_, _040541_, _040542_, _040543_, _040544_, _040545_, _040546_, _040547_, _040548_, _040549_, _040550_, _040551_, _040552_, _040553_, _040554_, _040555_, _040556_, _040557_, _040558_, _040559_, _040560_, _040561_, _040562_, _040563_, _040564_, _040565_, _040566_, _040567_, _040568_, _040569_, _040570_, _040571_, _040572_, _040573_, _040574_, _040575_, _040576_, _040577_, _040578_, _040579_, _040580_, _040581_, _040582_, _040583_, _040584_, _040585_, _040586_, _040587_, _040588_, _040589_, _040590_, _040591_, _040592_, _040593_, _040594_, _040595_, _040596_, _040597_, _040598_, _040599_, _040600_, _040601_, _040602_, _040603_, _040604_, _040605_, _040606_, _040607_, _040608_, _040609_, _040610_, _040611_, _040612_, _040613_, _040614_, _040615_, _040616_, _040617_, _040618_, _040619_, _040620_, _040621_, _040622_, _040623_, _040624_, _040625_, _040626_, _040627_, _040628_, _040629_, _040630_, _040631_, _040632_, _040633_, _040634_, _040635_, _040636_, _040637_, _040638_, _040639_, _040640_, _040641_, _040642_, _040643_, _040644_, _040645_, _040646_, _040647_, _040648_, _040649_, _040650_, _040651_, _040652_, _040653_, _040654_, _040655_, _040656_, _040657_, _040658_, _040659_, _040660_, _040661_, _040662_, _040663_, _040664_, _040665_, _040666_, _040667_, _040668_, _040669_, _040670_, _040671_, _040672_, _040673_, _040674_, _040675_, _040676_, _040677_, _040678_, _040679_, _040680_, _040681_, _040682_, _040683_, _040684_, _040685_, _040686_, _040687_, _040688_, _040689_, _040690_, _040691_, _040692_, _040693_, _040694_, _040695_, _040696_, _040697_, _040698_, _040699_, _040700_, _040701_, _040702_, _040703_, _040704_, _040705_, _040706_, _040707_, _040708_, _040709_, _040710_, _040711_, _040712_, _040713_, _040714_, _040715_, _040716_, _040717_, _040718_, _040719_, _040720_, _040721_, _040722_, _040723_, _040724_, _040725_, _040726_, _040727_, _040728_, _040729_, _040730_, _040731_, _040732_, _040733_, _040734_, _040735_, _040736_, _040737_, _040738_, _040739_, _040740_, _040741_, _040742_, _040743_, _040744_, _040745_, _040746_, _040747_, _040748_, _040749_, _040750_, _040751_, _040752_, _040753_, _040754_, _040755_, _040756_, _040757_, _040758_, _040759_, _040760_, _040761_, _040762_, _040763_, _040764_, _040765_, _040766_, _040767_, _040768_, _040769_, _040770_, _040771_, _040772_, _040773_, _040774_, _040775_, _040776_, _040777_, _040778_, _040779_, _040780_, _040781_, _040782_, _040783_, _040784_, _040785_, _040786_, _040787_, _040788_, _040789_, _040790_, _040791_, _040792_, _040793_, _040794_, _040795_, _040796_, _040797_, _040798_, _040799_, _040800_, _040801_, _040802_, _040803_, _040804_, _040805_, _040806_, _040807_, _040808_, _040809_, _040810_, _040811_, _040812_, _040813_, _040814_, _040815_, _040816_, _040817_, _040818_, _040819_, _040820_, _040821_, _040822_, _040823_, _040824_, _040825_, _040826_, _040827_, _040828_, _040829_, _040830_, _040831_, _040832_, _040833_, _040834_, _040835_, _040836_, _040837_, _040838_, _040839_, _040840_, _040841_, _040842_, _040843_, _040844_, _040845_, _040846_, _040847_, _040848_, _040849_, _040850_, _040851_, _040852_, _040853_, _040854_, _040855_, _040856_, _040857_, _040858_, _040859_, _040860_, _040861_, _040862_, _040863_, _040864_, _040865_, _040866_, _040867_, _040868_, _040869_, _040870_, _040871_, _040872_, _040873_, _040874_, _040875_, _040876_, _040877_, _040878_, _040879_, _040880_, _040881_, _040882_, _040883_, _040884_, _040885_, _040886_, _040887_, _040888_, _040889_, _040890_, _040891_, _040892_, _040893_, _040894_, _040895_, _040896_, _040897_, _040898_, _040899_, _040900_, _040901_, _040902_, _040903_, _040904_, _040905_, _040906_, _040907_, _040908_, _040909_, _040910_, _040911_, _040912_, _040913_, _040914_, _040915_, _040916_, _040917_, _040918_, _040919_, _040920_, _040921_, _040922_, _040923_, _040924_, _040925_, _040926_, _040927_, _040928_, _040929_, _040930_, _040931_, _040932_, _040933_, _040934_, _040935_, _040936_, _040937_, _040938_, _040939_, _040940_, _040941_, _040942_, _040943_, _040944_, _040945_, _040946_, _040947_, _040948_, _040949_, _040950_, _040951_, _040952_, _040953_, _040954_, _040955_, _040956_, _040957_, _040958_, _040959_, _040960_, _040961_, _040962_, _040963_, _040964_, _040965_, _040966_, _040967_, _040968_, _040969_, _040970_, _040971_, _040972_, _040973_, _040974_, _040975_, _040976_, _040977_, _040978_, _040979_, _040980_, _040981_, _040982_, _040983_, _040984_, _040985_, _040986_, _040987_, _040988_, _040989_, _040990_, _040991_, _040992_, _040993_, _040994_, _040995_, _040996_, _040997_, _040998_, _040999_, _041000_, _041001_, _041002_, _041003_, _041004_, _041005_, _041006_, _041007_, _041008_, _041009_, _041010_, _041011_, _041012_, _041013_, _041014_, _041015_, _041016_, _041017_, _041018_, _041019_, _041020_, _041021_, _041022_, _041023_, _041024_, _041025_, _041026_, _041027_, _041028_, _041029_, _041030_, _041031_, _041032_, _041033_, _041034_, _041035_, _041036_, _041037_, _041038_, _041039_, _041040_, _041041_, _041042_, _041043_, _041044_, _041045_, _041046_, _041047_, _041048_, _041049_, _041050_, _041051_, _041052_, _041053_, _041054_, _041055_, _041056_, _041057_, _041058_, _041059_, _041060_, _041061_, _041062_, _041063_, _041064_, _041065_, _041066_, _041067_, _041068_, _041069_, _041070_, _041071_, _041072_, _041073_, _041074_, _041075_, _041076_, _041077_, _041078_, _041079_, _041080_, _041081_, _041082_, _041083_, _041084_, _041085_, _041086_, _041087_, _041088_, _041089_, _041090_, _041091_, _041092_, _041093_, _041094_, _041095_, _041096_, _041097_, _041098_, _041099_, _041100_, _041101_, _041102_, _041103_, _041104_, _041105_, _041106_, _041107_, _041108_, _041109_, _041110_, _041111_, _041112_, _041113_, _041114_, _041115_, _041116_, _041117_, _041118_, _041119_, _041120_, _041121_, _041122_, _041123_, _041124_, _041125_, _041126_, _041127_, _041128_, _041129_, _041130_, _041131_, _041132_, _041133_, _041134_, _041135_, _041136_, _041137_, _041138_, _041139_, _041140_, _041141_, _041142_, _041143_, _041144_, _041145_, _041146_, _041147_, _041148_, _041149_, _041150_, _041151_, _041152_, _041153_, _041154_, _041155_, _041156_, _041157_, _041158_, _041159_, _041160_, _041161_, _041162_, _041163_, _041164_, _041165_, _041166_, _041167_, _041168_, _041169_, _041170_, _041171_, _041172_, _041173_, _041174_, _041175_, _041176_, _041177_, _041178_, _041179_, _041180_, _041181_, _041182_, _041183_, _041184_, _041185_, _041186_, _041187_, _041188_, _041189_, _041190_, _041191_, _041192_, _041193_, _041194_, _041195_, _041196_, _041197_, _041198_, _041199_, _041200_, _041201_, _041202_, _041203_, _041204_, _041205_, _041206_, _041207_, _041208_, _041209_, _041210_, _041211_, _041212_, _041213_, _041214_, _041215_, _041216_, _041217_, _041218_, _041219_, _041220_, _041221_, _041222_, _041223_, _041224_, _041225_, _041226_, _041227_, _041228_, _041229_, _041230_, _041231_, _041232_, _041233_, _041234_, _041235_, _041236_, _041237_, _041238_, _041239_, _041240_, _041241_, _041242_, _041243_, _041244_, _041245_, _041246_, _041247_, _041248_, _041249_, _041250_, _041251_, _041252_, _041253_, _041254_, _041255_, _041256_, _041257_, _041258_, _041259_, _041260_, _041261_, _041262_, _041263_, _041264_, _041265_, _041266_, _041267_, _041268_, _041269_, _041270_, _041271_, _041272_, _041273_, _041274_, _041275_, _041276_, _041277_, _041278_, _041279_, _041280_, _041281_, _041282_, _041283_, _041284_, _041285_, _041286_, _041287_, _041288_, _041289_, _041290_, _041291_, _041292_, _041293_, _041294_, _041295_, _041296_, _041297_, _041298_, _041299_, _041300_, _041301_, _041302_, _041303_, _041304_, _041305_, _041306_, _041307_, _041308_, _041309_, _041310_, _041311_, _041312_, _041313_, _041314_, _041315_, _041316_, _041317_, _041318_, _041319_, _041320_, _041321_, _041322_, _041323_, _041324_, _041325_, _041326_, _041327_, _041328_, _041329_, _041330_, _041331_, _041332_, _041333_, _041334_, _041335_, _041336_, _041337_, _041338_, _041339_, _041340_, _041341_, _041342_, _041343_, _041344_, _041345_, _041346_, _041347_, _041348_, _041349_, _041350_, _041351_, _041352_, _041353_, _041354_, _041355_, _041356_, _041357_, _041358_, _041359_, _041360_, _041361_, _041362_, _041363_, _041364_, _041365_, _041366_, _041367_, _041368_, _041369_, _041370_, _041371_, _041372_, _041373_, _041374_, _041375_, _041376_, _041377_, _041378_, _041379_, _041380_, _041381_, _041382_, _041383_, _041384_, _041385_, _041386_, _041387_, _041388_, _041389_, _041390_, _041391_, _041392_, _041393_, _041394_, _041395_, _041396_, _041397_, _041398_, _041399_, _041400_, _041401_, _041402_, _041403_, _041404_, _041405_, _041406_, _041407_, _041408_, _041409_, _041410_, _041411_, _041412_, _041413_, _041414_, _041415_, _041416_, _041417_, _041418_, _041419_, _041420_, _041421_, _041422_, _041423_, _041424_, _041425_, _041426_, _041427_, _041428_, _041429_, _041430_, _041431_, _041432_, _041433_, _041434_, _041435_, _041436_, _041437_, _041438_, _041439_, _041440_, _041441_, _041442_, _041443_, _041444_, _041445_, _041446_, _041447_, _041448_, _041449_, _041450_, _041451_, _041452_, _041453_, _041454_, _041455_, _041456_, _041457_, _041458_, _041459_, _041460_, _041461_, _041462_, _041463_, _041464_, _041465_, _041466_, _041467_, _041468_, _041469_, _041470_, _041471_, _041472_, _041473_, _041474_, _041475_, _041476_, _041477_, _041478_, _041479_, _041480_, _041481_, _041482_, _041483_, _041484_, _041485_, _041486_, _041487_, _041488_, _041489_, _041490_, _041491_, _041492_, _041493_, _041494_, _041495_, _041496_, _041497_, _041498_, _041499_, _041500_, _041501_, _041502_, _041503_, _041504_, _041505_, _041506_, _041507_, _041508_, _041509_, _041510_, _041511_, _041512_, _041513_, _041514_, _041515_, _041516_, _041517_, _041518_, _041519_, _041520_, _041521_, _041522_, _041523_, _041524_, _041525_, _041526_, _041527_, _041528_, _041529_, _041530_, _041531_, _041532_, _041533_, _041534_, _041535_, _041536_, _041537_, _041538_, _041539_, _041540_, _041541_, _041542_, _041543_, _041544_, _041545_, _041546_, _041547_, _041548_, _041549_, _041550_, _041551_, _041552_, _041553_, _041554_, _041555_, _041556_, _041557_, _041558_, _041559_, _041560_, _041561_, _041562_, _041563_, _041564_, _041565_, _041566_, _041567_, _041568_, _041569_, _041570_, _041571_, _041572_, _041573_, _041574_, _041575_, _041576_, _041577_, _041578_, _041579_, _041580_, _041581_, _041582_, _041583_, _041584_, _041585_, _041586_, _041587_, _041588_, _041589_, _041590_, _041591_, _041592_, _041593_, _041594_, _041595_, _041596_, _041597_, _041598_, _041599_, _041600_, _041601_, _041602_, _041603_, _041604_, _041605_, _041606_, _041607_, _041608_, _041609_, _041610_, _041611_, _041612_, _041613_, _041614_, _041615_, _041616_, _041617_, _041618_, _041619_, _041620_, _041621_, _041622_, _041623_, _041624_, _041625_, _041626_, _041627_, _041628_, _041629_, _041630_, _041631_, _041632_, _041633_, _041634_, _041635_, _041636_, _041637_, _041638_, _041639_, _041640_, _041641_, _041642_, _041643_, _041644_, _041645_, _041646_, _041647_, _041648_, _041649_, _041650_, _041651_, _041652_, _041653_, _041654_, _041655_, _041656_, _041657_, _041658_, _041659_, _041660_, _041661_, _041662_, _041663_, _041664_, _041665_, _041666_, _041667_, _041668_, _041669_, _041670_, _041671_, _041672_, _041673_, _041674_, _041675_, _041676_, _041677_, _041678_, _041679_, _041680_, _041681_, _041682_, _041683_, _041684_, _041685_, _041686_, _041687_, _041688_, _041689_, _041690_, _041691_, _041692_, _041693_, _041694_, _041695_, _041696_, _041697_, _041698_, _041699_, _041700_, _041701_, _041702_, _041703_, _041704_, _041705_, _041706_, _041707_, _041708_, _041709_, _041710_, _041711_, _041712_, _041713_, _041714_, _041715_, _041716_, _041717_, _041718_, _041719_, _041720_, _041721_, _041722_, _041723_, _041724_, _041725_, _041726_, _041727_, _041728_, _041729_, _041730_, _041731_, _041732_, _041733_, _041734_, _041735_, _041736_, _041737_, _041738_, _041739_, _041740_, _041741_, _041742_, _041743_, _041744_, _041745_, _041746_, _041747_, _041748_, _041749_, _041750_, _041751_, _041752_, _041753_, _041754_, _041755_, _041756_, _041757_, _041758_, _041759_, _041760_, _041761_, _041762_, _041763_, _041764_, _041765_, _041766_, _041767_, _041768_, _041769_, _041770_, _041771_, _041772_, _041773_, _041774_, _041775_, _041776_, _041777_, _041778_, _041779_, _041780_, _041781_, _041782_, _041783_, _041784_, _041785_, _041786_, _041787_, _041788_, _041789_, _041790_, _041791_, _041792_, _041793_, _041794_, _041795_, _041796_, _041797_, _041798_, _041799_, _041800_, _041801_, _041802_, _041803_, _041804_, _041805_, _041806_, _041807_, _041808_, _041809_, _041810_, _041811_, _041812_, _041813_, _041814_, _041815_, _041816_, _041817_, _041818_, _041819_, _041820_, _041821_, _041822_, _041823_, _041824_, _041825_, _041826_, _041827_, _041828_, _041829_, _041830_, _041831_, _041832_, _041833_, _041834_, _041835_, _041836_, _041837_, _041838_, _041839_, _041840_, _041841_, _041842_, _041843_, _041844_, _041845_, _041846_, _041847_, _041848_, _041849_, _041850_, _041851_, _041852_, _041853_, _041854_, _041855_, _041856_, _041857_, _041858_, _041859_, _041860_, _041861_, _041862_, _041863_, _041864_, _041865_, _041866_, _041867_, _041868_, _041869_, _041870_, _041871_, _041872_, _041873_, _041874_, _041875_, _041876_, _041877_, _041878_, _041879_, _041880_, _041881_, _041882_, _041883_, _041884_, _041885_, _041886_, _041887_, _041888_, _041889_, _041890_, _041891_, _041892_, _041893_, _041894_, _041895_, _041896_, _041897_, _041898_, _041899_, _041900_, _041901_, _041902_, _041903_, _041904_, _041905_, _041906_, _041907_, _041908_, _041909_, _041910_, _041911_, _041912_, _041913_, _041914_, _041915_, _041916_, _041917_, _041918_, _041919_, _041920_, _041921_, _041922_, _041923_, _041924_, _041925_, _041926_, _041927_, _041928_, _041929_, _041930_, _041931_, _041932_, _041933_, _041934_, _041935_, _041936_, _041937_, _041938_, _041939_, _041940_, _041941_, _041942_, _041943_, _041944_, _041945_, _041946_, _041947_, _041948_, _041949_, _041950_, _041951_, _041952_, _041953_, _041954_, _041955_, _041956_, _041957_, _041958_, _041959_, _041960_, _041961_, _041962_, _041963_, _041964_, _041965_, _041966_, _041967_, _041968_, _041969_, _041970_, _041971_, _041972_, _041973_, _041974_, _041975_, _041976_, _041977_, _041978_, _041979_, _041980_, _041981_, _041982_, _041983_, _041984_, _041985_, _041986_, _041987_, _041988_, _041989_, _041990_, _041991_, _041992_, _041993_, _041994_, _041995_, _041996_, _041997_, _041998_, _041999_, _042000_, _042001_, _042002_, _042003_, _042004_, _042005_, _042006_, _042007_, _042008_, _042009_, _042010_, _042011_, _042012_, _042013_, _042014_, _042015_, _042016_, _042017_, _042018_, _042019_, _042020_, _042021_, _042022_, _042023_, _042024_, _042025_, _042026_, _042027_, _042028_, _042029_, _042030_, _042031_, _042032_, _042033_, _042034_, _042035_, _042036_, _042037_, _042038_, _042039_, _042040_, _042041_, _042042_, _042043_, _042044_, _042045_, _042046_, _042047_, _042048_, _042049_, _042050_, _042051_, _042052_, _042053_, _042054_, _042055_, _042056_, _042057_, _042058_, _042059_, _042060_, _042061_, _042062_, _042063_, _042064_, _042065_, _042066_, _042067_, _042068_, _042069_, _042070_, _042071_, _042072_, _042073_, _042074_, _042075_, _042076_, _042077_, _042078_, _042079_, _042080_, _042081_, _042082_, _042083_, _042084_, _042085_, _042086_, _042087_, _042088_, _042089_, _042090_, _042091_, _042092_, _042093_, _042094_, _042095_, _042096_, _042097_, _042098_, _042099_, _042100_, _042101_, _042102_, _042103_, _042104_, _042105_, _042106_, _042107_, _042108_, _042109_, _042110_, _042111_, _042112_, _042113_, _042114_, _042115_, _042116_, _042117_, _042118_, _042119_, _042120_, _042121_, _042122_, _042123_, _042124_, _042125_, _042126_, _042127_, _042128_, _042129_, _042130_, _042131_, _042132_, _042133_, _042134_, _042135_, _042136_, _042137_, _042138_, _042139_, _042140_, _042141_, _042142_, _042143_, _042144_, _042145_, _042146_, _042147_, _042148_, _042149_, _042150_, _042151_, _042152_, _042153_, _042154_, _042155_, _042156_, _042157_, _042158_, _042159_, _042160_, _042161_, _042162_, _042163_, _042164_, _042165_, _042166_, _042167_, _042168_, _042169_, _042170_, _042171_, _042172_, _042173_, _042174_, _042175_, _042176_, _042177_, _042178_, _042179_, _042180_, _042181_, _042182_, _042183_, _042184_, _042185_, _042186_, _042187_, _042188_, _042189_, _042190_, _042191_, _042192_, _042193_, _042194_, _042195_, _042196_, _042197_, _042198_, _042199_, _042200_, _042201_, _042202_, _042203_, _042204_, _042205_, _042206_, _042207_, _042208_, _042209_, _042210_, _042211_, _042212_, _042213_, _042214_, _042215_, _042216_, _042217_, _042218_, _042219_, _042220_, _042221_, _042222_, _042223_, _042224_, _042225_, _042226_, _042227_, _042228_, _042229_, _042230_, _042231_, _042232_, _042233_, _042234_, _042235_, _042236_, _042237_, _042238_, _042239_, _042240_, _042241_, _042242_, _042243_, _042244_, _042245_, _042246_, _042247_, _042248_, _042249_, _042250_, _042251_, _042252_, _042253_, _042254_, _042255_, _042256_, _042257_, _042258_, _042259_, _042260_, _042261_, _042262_, _042263_, _042264_, _042265_, _042266_, _042267_, _042268_, _042269_, _042270_, _042271_, _042272_, _042273_, _042274_, _042275_, _042276_, _042277_, _042278_, _042279_, _042280_, _042281_, _042282_, _042283_, _042284_, _042285_, _042286_, _042287_, _042288_, _042289_, _042290_, _042291_, _042292_, _042293_, _042294_, _042295_, _042296_, _042297_, _042298_, _042299_, _042300_, _042301_, _042302_, _042303_, _042304_, _042305_, _042306_, _042307_, _042308_, _042309_, _042310_, _042311_, _042312_, _042313_, _042314_, _042315_, _042316_, _042317_, _042318_, _042319_, _042320_, _042321_, _042322_, _042323_, _042324_, _042325_, _042326_, _042327_, _042328_, _042329_, _042330_, _042331_, _042332_, _042333_, _042334_, _042335_, _042336_, _042337_, _042338_, _042339_, _042340_, _042341_, _042342_, _042343_, _042344_, _042345_, _042346_, _042347_, _042348_, _042349_, _042350_, _042351_, _042352_, _042353_, _042354_, _042355_, _042356_, _042357_, _042358_, _042359_, _042360_, _042361_, _042362_, _042363_, _042364_, _042365_, _042366_, _042367_, _042368_, _042369_, _042370_, _042371_, _042372_, _042373_, _042374_, _042375_, _042376_, _042377_, _042378_, _042379_, _042380_, _042381_, _042382_, _042383_, _042384_, _042385_, _042386_, _042387_, _042388_, _042389_, _042390_, _042391_, _042392_, _042393_, _042394_, _042395_, _042396_, _042397_, _042398_, _042399_, _042400_, _042401_, _042402_, _042403_, _042404_, _042405_, _042406_, _042407_, _042408_, _042409_, _042410_, _042411_, _042412_, _042413_, _042414_, _042415_, _042416_, _042417_, _042418_, _042419_, _042420_, _042421_, _042422_, _042423_, _042424_, _042425_, _042426_, _042427_, _042428_, _042429_, _042430_, _042431_, _042432_, _042433_, _042434_, _042435_, _042436_, _042437_, _042438_, _042439_, _042440_, _042441_, _042442_, _042443_, _042444_, _042445_, _042446_, _042447_, _042448_, _042449_, _042450_, _042451_, _042452_, _042453_, _042454_, _042455_, _042456_, _042457_, _042458_, _042459_, _042460_, _042461_, _042462_, _042463_, _042464_, _042465_, _042466_, _042467_, _042468_, _042469_, _042470_, _042471_, _042472_, _042473_, _042474_, _042475_, _042476_, _042477_, _042478_, _042479_, _042480_, _042481_, _042482_, _042483_, _042484_, _042485_, _042486_, _042487_, _042488_, _042489_, _042490_, _042491_, _042492_, _042493_, _042494_, _042495_, _042496_, _042497_, _042498_, _042499_, _042500_, _042501_, _042502_, _042503_, _042504_, _042505_, _042506_, _042507_, _042508_, _042509_, _042510_, _042511_, _042512_, _042513_, _042514_, _042515_, _042516_, _042517_, _042518_, _042519_, _042520_, _042521_, _042522_, _042523_, _042524_, _042525_, _042526_, _042527_, _042528_, _042529_, _042530_, _042531_, _042532_, _042533_, _042534_, _042535_, _042536_, _042537_, _042538_, _042539_, _042540_, _042541_, _042542_, _042543_, _042544_, _042545_, _042546_, _042547_, _042548_, _042549_, _042550_, _042551_, _042552_, _042553_, _042554_, _042555_, _042556_, _042557_, _042558_, _042559_, _042560_, _042561_, _042562_, _042563_, _042564_, _042565_, _042566_, _042567_, _042568_, _042569_, _042570_, _042571_, _042572_, _042573_, _042574_, _042575_, _042576_, _042577_, _042578_, _042579_, _042580_, _042581_, _042582_, _042583_, _042584_, _042585_, _042586_, _042587_, _042588_, _042589_, _042590_, _042591_, _042592_, _042593_, _042594_, _042595_, _042596_, _042597_, _042598_, _042599_, _042600_, _042601_, _042602_, _042603_, _042604_, _042605_, _042606_, _042607_, _042608_, _042609_, _042610_, _042611_, _042612_, _042613_, _042614_, _042615_, _042616_, _042617_, _042618_, _042619_, _042620_, _042621_, _042622_, _042623_, _042624_, _042625_, _042626_, _042627_, _042628_, _042629_, _042630_, _042631_, _042632_, _042633_, _042634_, _042635_, _042636_, _042637_, _042638_, _042639_, _042640_, _042641_, _042642_, _042643_, _042644_, _042645_, _042646_, _042647_, _042648_, _042649_, _042650_, _042651_, _042652_, _042653_, _042654_, _042655_, _042656_, _042657_, _042658_, _042659_, _042660_, _042661_, _042662_, _042663_, _042664_, _042665_, _042666_, _042667_, _042668_, _042669_, _042670_, _042671_, _042672_, _042673_, _042674_, _042675_, _042676_, _042677_, _042678_, _042679_, _042680_, _042681_, _042682_, _042683_, _042684_, _042685_, _042686_, _042687_, _042688_, _042689_, _042690_, _042691_, _042692_, _042693_, _042694_, _042695_, _042696_, _042697_, _042698_, _042699_, _042700_, _042701_, _042702_, _042703_, _042704_, _042705_, _042706_, _042707_, _042708_, _042709_, _042710_, _042711_, _042712_, _042713_, _042714_, _042715_, _042716_, _042717_, _042718_, _042719_, _042720_, _042721_, _042722_, _042723_, _042724_, _042725_, _042726_, _042727_, _042728_, _042729_, _042730_, _042731_, _042732_, _042733_, _042734_, _042735_, _042736_, _042737_, _042738_, _042739_, _042740_, _042741_, _042742_, _042743_, _042744_, _042745_, _042746_, _042747_, _042748_, _042749_, _042750_, _042751_, _042752_, _042753_, _042754_, _042755_, _042756_, _042757_, _042758_, _042759_, _042760_, _042761_, _042762_, _042763_, _042764_, _042765_, _042766_, _042767_, _042768_, _042769_, _042770_, _042771_, _042772_, _042773_, _042774_, _042775_, _042776_, _042777_, _042778_, _042779_, _042780_, _042781_, _042782_, _042783_, _042784_, _042785_, _042786_, _042787_, _042788_, _042789_, _042790_, _042791_, _042792_, _042793_, _042794_, _042795_, _042796_, _042797_, _042798_, _042799_, _042800_, _042801_, _042802_, _042803_, _042804_, _042805_, _042806_, _042807_, _042808_, _042809_, _042810_, _042811_, _042812_, _042813_, _042814_, _042815_, _042816_, _042817_, _042818_, _042819_, _042820_, _042821_, _042822_, _042823_, _042824_, _042825_, _042826_, _042827_, _042828_, _042829_, _042830_, _042831_, _042832_, _042833_, _042834_, _042835_, _042836_, _042837_, _042838_, _042839_, _042840_, _042841_, _042842_, _042843_, _042844_, _042845_, _042846_, _042847_, _042848_, _042849_, _042850_, _042851_, _042852_, _042853_, _042854_, _042855_, _042856_, _042857_, _042858_, _042859_, _042860_, _042861_, _042862_, _042863_, _042864_, _042865_, _042866_, _042867_, _042868_, _042869_, _042870_, _042871_, _042872_, _042873_, _042874_, _042875_, _042876_, _042877_, _042878_, _042879_, _042880_, _042881_, _042882_, _042883_, _042884_, _042885_, _042886_, _042887_, _042888_, _042889_, _042890_, _042891_, _042892_, _042893_, _042894_, _042895_, _042896_, _042897_, _042898_, _042899_, _042900_, _042901_, _042902_, _042903_, _042904_, _042905_, _042906_, _042907_, _042908_, _042909_, _042910_, _042911_, _042912_, _042913_, _042914_, _042915_, _042916_, _042917_, _042918_, _042919_, _042920_, _042921_, _042922_, _042923_, _042924_, _042925_, _042926_, _042927_, _042928_, _042929_, _042930_, _042931_, _042932_, _042933_, _042934_, _042935_, _042936_, _042937_, _042938_, _042939_, _042940_, _042941_, _042942_, _042943_, _042944_, _042945_, _042946_, _042947_, _042948_, _042949_, _042950_, _042951_, _042952_, _042953_, _042954_, _042955_, _042956_, _042957_, _042958_, _042959_, _042960_, _042961_, _042962_, _042963_, _042964_, _042965_, _042966_, _042967_, _042968_, _042969_, _042970_, _042971_, _042972_, _042973_, _042974_, _042975_, _042976_, _042977_, _042978_, _042979_, _042980_, _042981_, _042982_, _042983_, _042984_, _042985_, _042986_, _042987_, _042988_, _042989_, _042990_, _042991_, _042992_, _042993_, _042994_, _042995_, _042996_, _042997_, _042998_, _042999_, _043000_, _043001_, _043002_, _043003_, _043004_, _043005_, _043006_, _043007_, _043008_, _043009_, _043010_, _043011_, _043012_, _043013_, _043014_, _043015_, _043016_, _043017_, _043018_, _043019_, _043020_, _043021_, _043022_, _043023_, _043024_, _043025_, _043026_, _043027_, _043028_, _043029_, _043030_, _043031_, _043032_, _043033_, _043034_, _043035_, _043036_, _043037_, _043038_, _043039_, _043040_, _043041_, _043042_, _043043_, _043044_, _043045_, _043046_, _043047_, _043048_, _043049_, _043050_, _043051_, _043052_, _043053_, _043054_, _043055_, _043056_, _043057_, _043058_, _043059_, _043060_, _043061_, _043062_, _043063_, _043064_, _043065_, _043066_, _043067_, _043068_, _043069_, _043070_, _043071_, _043072_, _043073_, _043074_, _043075_, _043076_, _043077_, _043078_, _043079_, _043080_, _043081_, _043082_, _043083_, _043084_, _043085_, _043086_, _043087_, _043088_, _043089_, _043090_, _043091_, _043092_, _043093_, _043094_, _043095_, _043096_, _043097_, _043098_, _043099_, _043100_, _043101_, _043102_, _043103_, _043104_, _043105_, _043106_, _043107_, _043108_, _043109_, _043110_, _043111_, _043112_, _043113_, _043114_, _043115_, _043116_, _043117_, _043118_, _043119_, _043120_, _043121_, _043122_, _043123_, _043124_, _043125_, _043126_, _043127_, _043128_, _043129_, _043130_, _043131_, _043132_, _043133_, _043134_, _043135_, _043136_, _043137_, _043138_, _043139_, _043140_, _043141_, _043142_, _043143_, _043144_, _043145_, _043146_, _043147_, _043148_, _043149_, _043150_, _043151_, _043152_, _043153_, _043154_, _043155_, _043156_, _043157_, _043158_, _043159_, _043160_, _043161_, _043162_, _043163_, _043164_, _043165_, _043166_, _043167_, _043168_, _043169_, _043170_, _043171_, _043172_, _043173_, _043174_, _043175_, _043176_, _043177_, _043178_, _043179_, _043180_, _043181_, _043182_, _043183_, _043184_, _043185_, _043186_, _043187_, _043188_, _043189_, _043190_, _043191_, _043192_, _043193_, _043194_, _043195_, _043196_, _043197_, _043198_, _043199_, _043200_, _043201_, _043202_, _043203_, _043204_, _043205_, _043206_, _043207_, _043208_, _043209_, _043210_, _043211_, _043212_, _043213_, _043214_, _043215_, _043216_, _043217_, _043218_, _043219_, _043220_, _043221_, _043222_, _043223_, _043224_, _043225_, _043226_, _043227_, _043228_, _043229_, _043230_, _043231_, _043232_, _043233_, _043234_, _043235_, _043236_, _043237_, _043238_, _043239_, _043240_, _043241_, _043242_, _043243_, _043244_, _043245_, _043246_, _043247_, _043248_, _043249_, _043250_, _043251_, _043252_, _043253_, _043254_, _043255_, _043256_, _043257_, _043258_, _043259_, _043260_, _043261_, _043262_, _043263_, _043264_, _043265_, _043266_, _043267_, _043268_, _043269_, _043270_, _043271_, _043272_, _043273_, _043274_, _043275_, _043276_, _043277_, _043278_, _043279_, _043280_, _043281_, _043282_, _043283_, _043284_, _043285_, _043286_, _043287_, _043288_, _043289_, _043290_, _043291_, _043292_, _043293_, _043294_, _043295_, _043296_, _043297_, _043298_, _043299_, _043300_, _043301_, _043302_, _043303_, _043304_, _043305_, _043306_, _043307_, _043308_, _043309_, _043310_, _043311_, _043312_, _043313_, _043314_, _043315_, _043316_, _043317_, _043318_, _043319_, _043320_, _043321_, _043322_, _043323_, _043324_, _043325_, _043326_, _043327_, _043328_, _043329_, _043330_, _043331_, _043332_, _043333_, _043334_, _043335_, _043336_, _043337_, _043338_, _043339_, _043340_, _043341_, _043342_, _043343_, _043344_, _043345_, _043346_, _043347_, _043348_, _043349_, _043350_, _043351_, _043352_, _043353_, _043354_, _043355_, _043356_, _043357_, _043358_, _043359_, _043360_, _043361_, _043362_, _043363_, _043364_, _043365_, _043366_, _043367_, _043368_, _043369_, _043370_, _043371_, _043372_, _043373_, _043374_, _043375_, _043376_, _043377_, _043378_, _043379_, _043380_, _043381_, _043382_, _043383_, _043384_, _043385_, _043386_, _043387_, _043388_, _043389_, _043390_, _043391_, _043392_, _043393_, _043394_, _043395_, _043396_, _043397_, _043398_, _043399_, _043400_, _043401_, _043402_, _043403_, _043404_, _043405_, _043406_, _043407_, _043408_, _043409_, _043410_, _043411_, _043412_, _043413_, _043414_, _043415_, _043416_, _043417_, _043418_, _043419_, _043420_, _043421_, _043422_, _043423_, _043424_, _043425_, _043426_, _043427_, _043428_, _043429_, _043430_, _043431_, _043432_, _043433_, _043434_, _043435_, _043436_, _043437_, _043438_, _043439_, _043440_, _043441_, _043442_, _043443_, _043444_, _043445_, _043446_, _043447_, _043448_, _043449_, _043450_, _043451_, _043452_, _043453_, _043454_, _043455_, _043456_, _043457_, _043458_, _043459_, _043460_, _043461_, _043462_, _043463_, _043464_, _043465_, _043466_, _043467_, _043468_, _043469_, _043470_, _043471_, _043472_, _043473_, _043474_, _043475_, _043476_, _043477_, _043478_, _043479_, _043480_, _043481_, _043482_, _043483_, _043484_, _043485_, _043486_, _043487_, _043488_, _043489_, _043490_, _043491_, _043492_, _043493_, _043494_, _043495_, _043496_, _043497_, _043498_, _043499_, _043500_, _043501_, _043502_, _043503_, _043504_, _043505_, _043506_, _043507_, _043508_, _043509_, _043510_, _043511_, _043512_, _043513_, _043514_, _043515_, _043516_, _043517_, _043518_, _043519_, _043520_, _043521_, _043522_, _043523_, _043524_, _043525_, _043526_, _043527_, _043528_, _043529_, _043530_, _043531_, _043532_, _043533_, _043534_, _043535_, _043536_, _043537_, _043538_, _043539_, _043540_, _043541_, _043542_, _043543_, _043544_, _043545_, _043546_, _043547_, _043548_, _043549_, _043550_, _043551_, _043552_, _043553_, _043554_, _043555_, _043556_, _043557_, _043558_, _043559_, _043560_, _043561_, _043562_, _043563_, _043564_, _043565_, _043566_, _043567_, _043568_, _043569_, _043570_, _043571_, _043572_, _043573_, _043574_, _043575_, _043576_, _043577_, _043578_, _043579_, _043580_, _043581_, _043582_, _043583_, _043584_, _043585_, _043586_, _043587_, _043588_, _043589_, _043590_, _043591_, _043592_, _043593_, _043594_, _043595_, _043596_, _043597_, _043598_, _043599_, _043600_, _043601_, _043602_, _043603_, _043604_, _043605_, _043606_, _043607_, _043608_, _043609_, _043610_, _043611_, _043612_, _043613_, _043614_, _043615_, _043616_, _043617_, _043618_, _043619_, _043620_, _043621_, _043622_, _043623_, _043624_, _043625_, _043626_, _043627_, _043628_, _043629_, _043630_, _043631_, _043632_, _043633_, _043634_, _043635_, _043636_, _043637_, _043638_, _043639_, _043640_, _043641_, _043642_, _043643_, _043644_, _043645_, _043646_, _043647_, _043648_, _043649_, _043650_, _043651_, _043652_, _043653_, _043654_, _043655_, _043656_, _043657_, _043658_, _043659_, _043660_, _043661_, _043662_, _043663_, _043664_, _043665_, _043666_, _043667_, _043668_, _043669_, _043670_, _043671_, _043672_, _043673_, _043674_, _043675_, _043676_, _043677_, _043678_, _043679_, _043680_, _043681_, _043682_, _043683_, _043684_, _043685_, _043686_, _043687_, _043688_, _043689_, _043690_, _043691_, _043692_, _043693_, _043694_, _043695_, _043696_, _043697_, _043698_, _043699_, _043700_, _043701_, _043702_, _043703_, _043704_, _043705_, _043706_, _043707_, _043708_, _043709_, _043710_, _043711_, _043712_, _043713_, _043714_, _043715_, _043716_, _043717_, _043718_, _043719_, _043720_, _043721_, _043722_, _043723_, _043724_, _043725_, _043726_, _043727_, _043728_, _043729_, _043730_, _043731_, _043732_, _043733_, _043734_, _043735_, _043736_, _043737_, _043738_, _043739_, _043740_, _043741_, _043742_, _043743_, _043744_, _043745_, _043746_, _043747_, _043748_, _043749_, _043750_, _043751_, _043752_, _043753_, _043754_, _043755_, _043756_, _043757_, _043758_, _043759_, _043760_, _043761_, _043762_, _043763_, _043764_, _043765_, _043766_, _043767_, _043768_, _043769_, _043770_, _043771_, _043772_, _043773_, _043774_, _043775_, _043776_, _043777_, _043778_, _043779_, _043780_, _043781_, _043782_, _043783_, _043784_, _043785_, _043786_, _043787_, _043788_, _043789_, _043790_, _043791_, _043792_, _043793_, _043794_, _043795_, _043796_, _043797_, _043798_, _043799_, _043800_, _043801_, _043802_, _043803_, _043804_, _043805_, _043806_, _043807_, _043808_, _043809_, _043810_, _043811_, _043812_, _043813_, _043814_, _043815_, _043816_, _043817_, _043818_, _043819_, _043820_, _043821_, _043822_, _043823_, _043824_, _043825_, _043826_, _043827_, _043828_, _043829_, _043830_, _043831_, _043832_, _043833_, _043834_, _043835_, _043836_, _043837_, _043838_, _043839_, _043840_, _043841_, _043842_, _043843_, _043844_, _043845_, _043846_, _043847_, _043848_, _043849_, _043850_, _043851_, _043852_, _043853_, _043854_, _043855_, _043856_, _043857_, _043858_, _043859_, _043860_, _043861_, _043862_, _043863_, _043864_, _043865_, _043866_, _043867_, _043868_, _043869_, _043870_, _043871_, _043872_, _043873_, _043874_, _043875_, _043876_, _043877_, _043878_, _043879_, _043880_, _043881_, _043882_, _043883_, _043884_, _043885_, _043886_, _043887_, _043888_, _043889_, _043890_, _043891_, _043892_, _043893_, _043894_, _043895_, _043896_, _043897_, _043898_, _043899_, _043900_, _043901_, _043902_, _043903_, _043904_, _043905_, _043906_, _043907_, _043908_, _043909_, _043910_, _043911_, _043912_, _043913_, _043914_, _043915_, _043916_, _043917_, _043918_, _043919_, _043920_, _043921_, _043922_, _043923_, _043924_, _043925_, _043926_, _043927_, _043928_, _043929_, _043930_, _043931_, _043932_, _043933_, _043934_, _043935_, _043936_, _043937_, _043938_, _043939_, _043940_, _043941_, _043942_, _043943_, _043944_, _043945_, _043946_, _043947_, _043948_, _043949_, _043950_, _043951_, _043952_, _043953_, _043954_, _043955_, _043956_, _043957_, _043958_, _043959_, _043960_, _043961_, _043962_, _043963_, _043964_, _043965_, _043966_, _043967_, _043968_, _043969_, _043970_, _043971_, _043972_, _043973_, _043974_, _043975_, _043976_, _043977_, _043978_, _043979_, _043980_, _043981_, _043982_, _043983_, _043984_, _043985_, _043986_, _043987_, _043988_, _043989_, _043990_, _043991_, _043992_, _043993_, _043994_, _043995_, _043996_, _043997_, _043998_, _043999_, _044000_, _044001_, _044002_, _044003_, _044004_, _044005_, _044006_, _044007_, _044008_, _044009_, _044010_, _044011_, _044012_, _044013_, _044014_, _044015_, _044016_, _044017_, _044018_, _044019_, _044020_, _044021_, _044022_, _044023_, _044024_, _044025_, _044026_, _044027_, _044028_, _044029_, _044030_, _044031_, _044032_, _044033_, _044034_, _044035_, _044036_, _044037_, _044038_, _044039_, _044040_, _044041_, _044042_, _044043_, _044044_, _044045_, _044046_, _044047_, _044048_, _044049_, _044050_, _044051_, _044052_, _044053_, _044054_, _044055_, _044056_, _044057_, _044058_, _044059_, _044060_, _044061_, _044062_, _044063_, _044064_, _044065_, _044066_, _044067_, _044068_, _044069_, _044070_, _044071_, _044072_, _044073_, _044074_, _044075_, _044076_, _044077_, _044078_, _044079_, _044080_, _044081_, _044082_, _044083_, _044084_, _044085_, _044086_, _044087_, _044088_, _044089_, _044090_, _044091_, _044092_, _044093_, _044094_, _044095_, _044096_, _044097_, _044098_, _044099_, _044100_, _044101_, _044102_, _044103_, _044104_, _044105_, _044106_, _044107_, _044108_, _044109_, _044110_, _044111_, _044112_, _044113_, _044114_, _044115_, _044116_, _044117_, _044118_, _044119_, _044120_, _044121_, _044122_, _044123_, _044124_, _044125_, _044126_, _044127_, _044128_, _044129_, _044130_, _044131_, _044132_, _044133_, _044134_, _044135_, _044136_, _044137_, _044138_, _044139_, _044140_, _044141_, _044142_, _044143_, _044144_, _044145_, _044146_, _044147_, _044148_, _044149_, _044150_, _044151_, _044152_, _044153_, _044154_, _044155_, _044156_, _044157_, _044158_, _044159_, _044160_, _044161_, _044162_, _044163_, _044164_, _044165_, _044166_, _044167_, _044168_, _044169_, _044170_, _044171_, _044172_, _044173_, _044174_, _044175_, _044176_, _044177_, _044178_, _044179_, _044180_, _044181_, _044182_, _044183_, _044184_, _044185_, _044186_, _044187_, _044188_, _044189_, _044190_, _044191_, _044192_, _044193_, _044194_, _044195_, _044196_, _044197_, _044198_, _044199_, _044200_, _044201_, _044202_, _044203_, _044204_, _044205_, _044206_, _044207_, _044208_, _044209_, _044210_, _044211_, _044212_, _044213_, _044214_, _044215_, _044216_, _044217_, _044218_, _044219_, _044220_, _044221_, _044222_, _044223_, _044224_, _044225_, _044226_, _044227_, _044228_, _044229_, _044230_, _044231_, _044232_, _044233_, _044234_, _044235_, _044236_, _044237_, _044238_, _044239_, _044240_, _044241_, _044242_, _044243_, _044244_, _044245_, _044246_, _044247_, _044248_, _044249_, _044250_, _044251_, _044252_, _044253_, _044254_, _044255_, _044256_, _044257_, _044258_, _044259_, _044260_, _044261_, _044262_, _044263_, _044264_, _044265_, _044266_, _044267_, _044268_, _044269_, _044270_, _044271_, _044272_, _044273_, _044274_, _044275_, _044276_, _044277_, _044278_, _044279_, _044280_, _044281_, _044282_, _044283_, _044284_, _044285_, _044286_, _044287_, _044288_, _044289_, _044290_, _044291_, _044292_, _044293_, _044294_, _044295_, _044296_, _044297_, _044298_, _044299_, _044300_, _044301_, _044302_, _044303_, _044304_, _044305_, _044306_, _044307_, _044308_, _044309_, _044310_, _044311_, _044312_, _044313_, _044314_, _044315_, _044316_, _044317_, _044318_, _044319_, _044320_, _044321_, _044322_, _044323_, _044324_, _044325_, _044326_, _044327_, _044328_, _044329_, _044330_, _044331_, _044332_, _044333_, _044334_, _044335_, _044336_, _044337_, _044338_, _044339_, _044340_, _044341_, _044342_, _044343_, _044344_, _044345_, _044346_, _044347_, _044348_, _044349_, _044350_, _044351_, _044352_, _044353_, _044354_, _044355_, _044356_, _044357_, _044358_, _044359_, _044360_, _044361_, _044362_, _044363_, _044364_, _044365_, _044366_, _044367_, _044368_, _044369_, _044370_, _044371_, _044372_, _044373_, _044374_, _044375_, _044376_, _044377_, _044378_, _044379_, _044380_, _044381_, _044382_, _044383_, _044384_, _044385_, _044386_, _044387_, _044388_, _044389_, _044390_, _044391_, _044392_, _044393_, _044394_, _044395_, _044396_, _044397_, _044398_, _044399_, _044400_, _044401_, _044402_, _044403_, _044404_, _044405_, _044406_, _044407_, _044408_, _044409_, _044410_, _044411_, _044412_, _044413_, _044414_, _044415_, _044416_, _044417_, _044418_, _044419_, _044420_, _044421_, _044422_, _044423_, _044424_, _044425_, _044426_, _044427_, _044428_, _044429_, _044430_, _044431_, _044432_, _044433_, _044434_, _044435_, _044436_, _044437_, _044438_, _044439_, _044440_, _044441_, _044442_, _044443_, _044444_, _044445_, _044446_, _044447_, _044448_, _044449_, _044450_, _044451_, _044452_, _044453_, _044454_, _044455_, _044456_, _044457_, _044458_, _044459_, _044460_, _044461_, _044462_, _044463_, _044464_, _044465_, _044466_, _044467_, _044468_, _044469_, _044470_, _044471_, _044472_, _044473_, _044474_, _044475_, _044476_, _044477_, _044478_, _044479_, _044480_, _044481_, _044482_, _044483_, _044484_, _044485_, _044486_, _044487_, _044488_, _044489_, _044490_, _044491_, _044492_, _044493_, _044494_, _044495_, _044496_, _044497_, _044498_, _044499_, _044500_, _044501_, _044502_, _044503_, _044504_, _044505_, _044506_, _044507_, _044508_, _044509_, _044510_, _044511_, _044512_, _044513_, _044514_, _044515_, _044516_, _044517_, _044518_, _044519_, _044520_, _044521_, _044522_, _044523_, _044524_, _044525_, _044526_, _044527_, _044528_, _044529_, _044530_, _044531_, _044532_, _044533_, _044534_, _044535_, _044536_, _044537_, _044538_, _044539_, _044540_, _044541_, _044542_, _044543_, _044544_, _044545_, _044546_, _044547_, _044548_, _044549_, _044550_, _044551_, _044552_, _044553_, _044554_, _044555_, _044556_, _044557_, _044558_, _044559_, _044560_, _044561_, _044562_, _044563_, _044564_, _044565_, _044566_, _044567_, _044568_, _044569_, _044570_, _044571_, _044572_, _044573_, _044574_, _044575_, _044576_, _044577_, _044578_, _044579_, _044580_, _044581_, _044582_, _044583_, _044584_, _044585_, _044586_, _044587_, _044588_, _044589_, _044590_, _044591_, _044592_, _044593_, _044594_, _044595_, _044596_, _044597_, _044598_, _044599_, _044600_, _044601_, _044602_, _044603_, _044604_, _044605_, _044606_, _044607_, _044608_, _044609_, _044610_, _044611_, _044612_, _044613_, _044614_, _044615_, _044616_, _044617_, _044618_, _044619_, _044620_, _044621_, _044622_, _044623_, _044624_, _044625_, _044626_, _044627_, _044628_, _044629_, _044630_, _044631_, _044632_, _044633_, _044634_, _044635_, _044636_, _044637_, _044638_, _044639_, _044640_, _044641_, _044642_, _044643_, _044644_, _044645_, _044646_, _044647_, _044648_, _044649_, _044650_, _044651_, _044652_, _044653_, _044654_, _044655_, _044656_, _044657_, _044658_, _044659_, _044660_, _044661_, _044662_, _044663_, _044664_, _044665_, _044666_, _044667_, _044668_, _044669_, _044670_, _044671_, _044672_, _044673_, _044674_, _044675_, _044676_, _044677_, _044678_, _044679_, _044680_, _044681_, _044682_, _044683_, _044684_, _044685_, _044686_, _044687_, _044688_, _044689_, _044690_, _044691_, _044692_, _044693_, _044694_, _044695_, _044696_, _044697_, _044698_, _044699_, _044700_, _044701_, _044702_, _044703_, _044704_, _044705_, _044706_, _044707_, _044708_, _044709_, _044710_, _044711_, _044712_, _044713_, _044714_, _044715_, _044716_, _044717_, _044718_, _044719_, _044720_, _044721_, _044722_, _044723_, _044724_, _044725_, _044726_, _044727_, _044728_, _044729_, _044730_, _044731_, _044732_, _044733_, _044734_, _044735_, _044736_, _044737_, _044738_, _044739_, _044740_, _044741_, _044742_, _044743_, _044744_, _044745_, _044746_, _044747_, _044748_, _044749_, _044750_, _044751_, _044752_, _044753_, _044754_, _044755_, _044756_, _044757_, _044758_, _044759_, _044760_, _044761_, _044762_, _044763_, _044764_, _044765_, _044766_, _044767_, _044768_, _044769_, _044770_, _044771_, _044772_, _044773_, _044774_, _044775_, _044776_, _044777_, _044778_, _044779_, _044780_, _044781_, _044782_, _044783_, _044784_, _044785_, _044786_, _044787_, _044788_, _044789_, _044790_, _044791_, _044792_, _044793_, _044794_, _044795_, _044796_, _044797_, _044798_, _044799_, _044800_, _044801_, _044802_, _044803_, _044804_, _044805_, _044806_, _044807_, _044808_, _044809_, _044810_, _044811_, _044812_, _044813_, _044814_, _044815_, _044816_, _044817_, _044818_, _044819_, _044820_, _044821_, _044822_, _044823_, _044824_, _044825_, _044826_, _044827_, _044828_, _044829_, _044830_, _044831_, _044832_, _044833_, _044834_, _044835_, _044836_, _044837_, _044838_, _044839_, _044840_, _044841_, _044842_, _044843_, _044844_, _044845_, _044846_, _044847_, _044848_, _044849_, _044850_, _044851_, _044852_, _044853_, _044854_, _044855_, _044856_, _044857_, _044858_, _044859_, _044860_, _044861_, _044862_, _044863_, _044864_, _044865_, _044866_, _044867_, _044868_, _044869_, _044870_, _044871_, _044872_, _044873_, _044874_, _044875_, _044876_, _044877_, _044878_, _044879_, _044880_, _044881_, _044882_, _044883_, _044884_, _044885_, _044886_, _044887_, _044888_, _044889_, _044890_, _044891_, _044892_, _044893_, _044894_, _044895_, _044896_, _044897_, _044898_, _044899_, _044900_, _044901_, _044902_, _044903_, _044904_, _044905_, _044906_, _044907_, _044908_, _044909_, _044910_, _044911_, _044912_, _044913_, _044914_, _044915_, _044916_, _044917_, _044918_, _044919_, _044920_, _044921_, _044922_, _044923_, _044924_, _044925_, _044926_, _044927_, _044928_, _044929_, _044930_, _044931_, _044932_, _044933_, _044934_, _044935_, _044936_, _044937_, _044938_, _044939_, _044940_, _044941_, _044942_, _044943_, _044944_, _044945_, _044946_, _044947_, _044948_, _044949_, _044950_, _044951_, _044952_, _044953_, _044954_, _044955_, _044956_, _044957_, _044958_, _044959_, _044960_, _044961_, _044962_, _044963_, _044964_, _044965_, _044966_, _044967_, _044968_, _044969_, _044970_, _044971_, _044972_, _044973_, _044974_, _044975_, _044976_, _044977_, _044978_, _044979_, _044980_, _044981_, _044982_, _044983_, _044984_, _044985_, _044986_, _044987_, _044988_, _044989_, _044990_, _044991_, _044992_, _044993_, _044994_, _044995_, _044996_, _044997_, _044998_, _044999_, _045000_, _045001_, _045002_, _045003_, _045004_, _045005_, _045006_, _045007_, _045008_, _045009_, _045010_, _045011_, _045012_, _045013_, _045014_, _045015_, _045016_, _045017_, _045018_, _045019_, _045020_, _045021_, _045022_, _045023_, _045024_, _045025_, _045026_, _045027_, _045028_, _045029_, _045030_, _045031_, _045032_, _045033_, _045034_, _045035_, _045036_, _045037_, _045038_, _045039_, _045040_, _045041_, _045042_, _045043_, _045044_, _045045_, _045046_, _045047_, _045048_, _045049_, _045050_, _045051_, _045052_, _045053_, _045054_, _045055_, _045056_, _045057_, _045058_, _045059_, _045060_, _045061_, _045062_, _045063_, _045064_, _045065_, _045066_, _045067_, _045068_, _045069_, _045070_, _045071_, _045072_, _045073_, _045074_, _045075_, _045076_, _045077_, _045078_, _045079_, _045080_, _045081_, _045082_, _045083_, _045084_, _045085_, _045086_, _045087_, _045088_, _045089_, _045090_, _045091_, _045092_, _045093_, _045094_, _045095_, _045096_, _045097_, _045098_, _045099_, _045100_, _045101_, _045102_, _045103_, _045104_, _045105_, _045106_, _045107_, _045108_, _045109_, _045110_, _045111_, _045112_, _045113_, _045114_, _045115_, _045116_, _045117_, _045118_, _045119_, _045120_, _045121_, _045122_, _045123_, _045124_, _045125_, _045126_, _045127_, _045128_, _045129_, _045130_, _045131_, _045132_, _045133_, _045134_, _045135_, _045136_, _045137_, _045138_, _045139_, _045140_, _045141_, _045142_, _045143_, _045144_, _045145_, _045146_, _045147_, _045148_, _045149_, _045150_, _045151_, _045152_, _045153_, _045154_, _045155_, _045156_, _045157_, _045158_, _045159_, _045160_, _045161_, _045162_, _045163_, _045164_, _045165_, _045166_, _045167_, _045168_, _045169_, _045170_, _045171_, _045172_, _045173_, _045174_, _045175_, _045176_, _045177_, _045178_, _045179_, _045180_, _045181_, _045182_, _045183_, _045184_, _045185_, _045186_, _045187_, _045188_, _045189_, _045190_, _045191_, _045192_, _045193_, _045194_, _045195_, _045196_, _045197_, _045198_, _045199_, _045200_, _045201_, _045202_, _045203_, _045204_, _045205_, _045206_, _045207_, _045208_, _045209_, _045210_, _045211_, _045212_, _045213_, _045214_, _045215_, _045216_, _045217_, _045218_, _045219_, _045220_, _045221_, _045222_, _045223_, _045224_, _045225_, _045226_, _045227_, _045228_, _045229_, _045230_, _045231_, _045232_, _045233_, _045234_, _045235_, _045236_, _045237_, _045238_, _045239_, _045240_, _045241_, _045242_, _045243_, _045244_, _045245_, _045246_, _045247_, _045248_, _045249_, _045250_, _045251_, _045252_, _045253_, _045254_, _045255_, _045256_, _045257_, _045258_, _045259_, _045260_, _045261_, _045262_, _045263_, _045264_, _045265_, _045266_, _045267_, _045268_, _045269_, _045270_, _045271_, _045272_, _045273_, _045274_, _045275_, _045276_, _045277_, _045278_, _045279_, _045280_, _045281_, _045282_, _045283_, _045284_, _045285_, _045286_, _045287_, _045288_, _045289_, _045290_, _045291_, _045292_, _045293_, _045294_, _045295_, _045296_, _045297_, _045298_, _045299_, _045300_, _045301_, _045302_, _045303_, _045304_, _045305_, _045306_, _045307_, _045308_, _045309_, _045310_, _045311_, _045312_, _045313_, _045314_, _045315_, _045316_, _045317_, _045318_, _045319_, _045320_, _045321_, _045322_, _045323_, _045324_, _045325_, _045326_, _045327_, _045328_, _045329_, _045330_, _045331_, _045332_, _045333_, _045334_, _045335_, _045336_, _045337_, _045338_, _045339_, _045340_, _045341_, _045342_, _045343_, _045344_, _045345_, _045346_, _045347_, _045348_, _045349_, _045350_, _045351_, _045352_, _045353_, _045354_, _045355_, _045356_, _045357_, _045358_, _045359_, _045360_, _045361_, _045362_, _045363_, _045364_, _045365_, _045366_, _045367_, _045368_, _045369_, _045370_, _045371_, _045372_, _045373_, _045374_, _045375_, _045376_, _045377_, _045378_, _045379_, _045380_, _045381_, _045382_, _045383_, _045384_, _045385_, _045386_, _045387_, _045388_, _045389_, _045390_, _045391_, _045392_, _045393_, _045394_, _045395_, _045396_, _045397_, _045398_, _045399_, _045400_, _045401_, _045402_, _045403_, _045404_, _045405_, _045406_, _045407_, _045408_, _045409_, _045410_, _045411_, _045412_, _045413_, _045414_, _045415_, _045416_, _045417_, _045418_, _045419_, _045420_, _045421_, _045422_, _045423_, _045424_, _045425_, _045426_, _045427_, _045428_, _045429_, _045430_, _045431_, _045432_, _045433_, _045434_, _045435_, _045436_, _045437_, _045438_, _045439_, _045440_, _045441_, _045442_, _045443_, _045444_, _045445_, _045446_, _045447_, _045448_, _045449_, _045450_, _045451_, _045452_, _045453_, _045454_, _045455_, _045456_, _045457_, _045458_, _045459_, _045460_, _045461_, _045462_, _045463_, _045464_, _045465_, _045466_, _045467_, _045468_, _045469_, _045470_, _045471_, _045472_, _045473_, _045474_, _045475_, _045476_, _045477_, _045478_, _045479_, _045480_, _045481_, _045482_, _045483_, _045484_, _045485_, _045486_, _045487_, _045488_, _045489_, _045490_, _045491_, _045492_, _045493_, _045494_, _045495_, _045496_, _045497_, _045498_, _045499_, _045500_, _045501_, _045502_, _045503_, _045504_, _045505_, _045506_, _045507_, _045508_, _045509_, _045510_, _045511_, _045512_, _045513_, _045514_, _045515_, _045516_, _045517_, _045518_, _045519_, _045520_, _045521_, _045522_, _045523_, _045524_, _045525_, _045526_, _045527_, _045528_, _045529_, _045530_, _045531_, _045532_, _045533_, _045534_, _045535_, _045536_, _045537_, _045538_, _045539_, _045540_, _045541_, _045542_, _045543_, _045544_, _045545_, _045546_, _045547_, _045548_, _045549_, _045550_, _045551_, _045552_, _045553_, _045554_, _045555_, _045556_, _045557_, _045558_, _045559_, _045560_, _045561_, _045562_, _045563_, _045564_, _045565_, _045566_, _045567_, _045568_, _045569_, _045570_, _045571_, _045572_, _045573_, _045574_, _045575_, _045576_, _045577_, _045578_, _045579_, _045580_, _045581_, _045582_, _045583_, _045584_, _045585_, _045586_, _045587_, _045588_, _045589_, _045590_, _045591_, _045592_, _045593_, _045594_, _045595_, _045596_, _045597_, _045598_, _045599_, _045600_, _045601_, _045602_, _045603_, _045604_, _045605_, _045606_, _045607_, _045608_, _045609_, _045610_, _045611_, _045612_, _045613_, _045614_, _045615_, _045616_, _045617_, _045618_, _045619_, _045620_, _045621_, _045622_, _045623_, _045624_, _045625_, _045626_, _045627_, _045628_, _045629_, _045630_, _045631_, _045632_, _045633_, _045634_, _045635_, _045636_, _045637_, _045638_, _045639_, _045640_, _045641_, _045642_, _045643_, _045644_, _045645_, _045646_, _045647_, _045648_, _045649_, _045650_, _045651_, _045652_, _045653_, _045654_, _045655_, _045656_, _045657_, _045658_, _045659_, _045660_, _045661_, _045662_, _045663_, _045664_, _045665_, _045666_, _045667_, _045668_, _045669_, _045670_, _045671_, _045672_, _045673_, _045674_, _045675_, _045676_, _045677_, _045678_, _045679_, _045680_, _045681_, _045682_, _045683_, _045684_, _045685_, _045686_, _045687_, _045688_, _045689_, _045690_, _045691_, _045692_, _045693_, _045694_, _045695_, _045696_, _045697_, _045698_, _045699_, _045700_, _045701_, _045702_, _045703_, _045704_, _045705_, _045706_, _045707_, _045708_, _045709_, _045710_, _045711_, _045712_, _045713_, _045714_, _045715_, _045716_, _045717_, _045718_, _045719_, _045720_, _045721_, _045722_, _045723_, _045724_, _045725_, _045726_, _045727_, _045728_, _045729_, _045730_, _045731_, _045732_, _045733_, _045734_, _045735_, _045736_, _045737_, _045738_, _045739_, _045740_, _045741_, _045742_, _045743_, _045744_, _045745_, _045746_, _045747_, _045748_, _045749_, _045750_, _045751_, _045752_, _045753_, _045754_, _045755_, _045756_, _045757_, _045758_, _045759_, _045760_, _045761_, _045762_, _045763_, _045764_, _045765_, _045766_, _045767_, _045768_, _045769_, _045770_, _045771_, _045772_, _045773_, _045774_, _045775_, _045776_, _045777_, _045778_, _045779_, _045780_, _045781_, _045782_, _045783_, _045784_, _045785_, _045786_, _045787_, _045788_, _045789_, _045790_, _045791_, _045792_, _045793_, _045794_, _045795_, _045796_, _045797_, _045798_, _045799_, _045800_, _045801_, _045802_, _045803_, _045804_, _045805_, _045806_, _045807_, _045808_, _045809_, _045810_, _045811_, _045812_, _045813_, _045814_, _045815_, _045816_, _045817_, _045818_, _045819_, _045820_, _045821_, _045822_, _045823_, _045824_, _045825_, _045826_, _045827_, _045828_, _045829_, _045830_, _045831_, _045832_, _045833_, _045834_, _045835_, _045836_, _045837_, _045838_, _045839_, _045840_, _045841_, _045842_, _045843_, _045844_, _045845_, _045846_, _045847_, _045848_, _045849_, _045850_, _045851_, _045852_, _045853_, _045854_, _045855_, _045856_, _045857_, _045858_, _045859_, _045860_, _045861_, _045862_, _045863_, _045864_, _045865_, _045866_, _045867_, _045868_, _045869_, _045870_, _045871_, _045872_, _045873_, _045874_, _045875_, _045876_, _045877_, _045878_, _045879_, _045880_, _045881_, _045882_, _045883_, _045884_, _045885_, _045886_, _045887_, _045888_, _045889_, _045890_, _045891_, _045892_, _045893_, _045894_, _045895_, _045896_, _045897_, _045898_, _045899_, _045900_, _045901_, _045902_, _045903_, _045904_, _045905_, _045906_, _045907_, _045908_, _045909_, _045910_, _045911_, _045912_, _045913_, _045914_, _045915_, _045916_, _045917_, _045918_, _045919_, _045920_, _045921_, _045922_, _045923_, _045924_, _045925_, _045926_, _045927_, _045928_, _045929_, _045930_, _045931_, _045932_, _045933_, _045934_, _045935_, _045936_, _045937_, _045938_, _045939_, _045940_, _045941_, _045942_, _045943_, _045944_, _045945_, _045946_, _045947_, _045948_, _045949_, _045950_, _045951_, _045952_, _045953_, _045954_, _045955_, _045956_, _045957_, _045958_, _045959_, _045960_, _045961_, _045962_, _045963_, _045964_, _045965_, _045966_, _045967_, _045968_, _045969_, _045970_, _045971_, _045972_, _045973_, _045974_, _045975_, _045976_, _045977_, _045978_, _045979_, _045980_, _045981_, _045982_, _045983_, _045984_, _045985_, _045986_, _045987_, _045988_, _045989_, _045990_, _045991_, _045992_, _045993_, _045994_, _045995_, _045996_, _045997_, _045998_, _045999_, _046000_, _046001_, _046002_, _046003_, _046004_, _046005_, _046006_, _046007_, _046008_, _046009_, _046010_, _046011_, _046012_, _046013_, _046014_, _046015_, _046016_, _046017_, _046018_, _046019_, _046020_, _046021_, _046022_, _046023_, _046024_, _046025_, _046026_, _046027_, _046028_, _046029_, _046030_, _046031_, _046032_, _046033_, _046034_, _046035_, _046036_, _046037_, _046038_, _046039_, _046040_, _046041_, _046042_, _046043_, _046044_, _046045_, _046046_, _046047_, _046048_, _046049_, _046050_, _046051_, _046052_, _046053_, _046054_, _046055_, _046056_, _046057_, _046058_, _046059_, _046060_, _046061_, _046062_, _046063_, _046064_, _046065_, _046066_, _046067_, _046068_, _046069_, _046070_, _046071_, _046072_, _046073_, _046074_, _046075_, _046076_, _046077_, _046078_, _046079_, _046080_, _046081_, _046082_, _046083_, _046084_, _046085_, _046086_, _046087_, _046088_, _046089_, _046090_, _046091_, _046092_, _046093_, _046094_, _046095_, _046096_, _046097_, _046098_, _046099_, _046100_, _046101_, _046102_, _046103_, _046104_, _046105_, _046106_, _046107_, _046108_, _046109_, _046110_, _046111_, _046112_, _046113_, _046114_, _046115_, _046116_, _046117_, _046118_, _046119_, _046120_, _046121_, _046122_, _046123_, _046124_, _046125_, _046126_, _046127_, _046128_, _046129_, _046130_, _046131_, _046132_, _046133_, _046134_, _046135_, _046136_, _046137_, _046138_, _046139_, _046140_, _046141_, _046142_, _046143_, _046144_, _046145_, _046146_, _046147_, _046148_, _046149_, _046150_, _046151_, _046152_, _046153_, _046154_, _046155_, _046156_, _046157_, _046158_, _046159_, _046160_, _046161_, _046162_, _046163_, _046164_, _046165_, _046166_, _046167_, _046168_, _046169_, _046170_, _046171_, _046172_, _046173_, _046174_, _046175_, _046176_, _046177_, _046178_, _046179_, _046180_, _046181_, _046182_, _046183_, _046184_, _046185_, _046186_, _046187_, _046188_, _046189_, _046190_, _046191_, _046192_, _046193_, _046194_, _046195_, _046196_, _046197_, _046198_, _046199_, _046200_, _046201_, _046202_, _046203_, _046204_, _046205_, _046206_, _046207_, _046208_, _046209_, _046210_, _046211_, _046212_, _046213_, _046214_, _046215_, _046216_, _046217_, _046218_, _046219_, _046220_, _046221_, _046222_, _046223_, _046224_, _046225_, _046226_, _046227_, _046228_, _046229_, _046230_, _046231_, _046232_, _046233_, _046234_, _046235_, _046236_, _046237_, _046238_, _046239_, _046240_, _046241_, _046242_, _046243_, _046244_, _046245_, _046246_, _046247_, _046248_, _046249_, _046250_, _046251_, _046252_, _046253_, _046254_, _046255_, _046256_, _046257_, _046258_, _046259_, _046260_, _046261_, _046262_, _046263_, _046264_, _046265_, _046266_, _046267_, _046268_, _046269_, _046270_, _046271_, _046272_, _046273_, _046274_, _046275_, _046276_, _046277_, _046278_, _046279_, _046280_, _046281_, _046282_, _046283_, _046284_, _046285_, _046286_, _046287_, _046288_, _046289_, _046290_, _046291_, _046292_, _046293_, _046294_, _046295_, _046296_, _046297_, _046298_, _046299_, _046300_, _046301_, _046302_, _046303_, _046304_, _046305_, _046306_, _046307_, _046308_, _046309_, _046310_, _046311_, _046312_, _046313_, _046314_, _046315_, _046316_, _046317_, _046318_, _046319_, _046320_, _046321_, _046322_, _046323_, _046324_, _046325_, _046326_, _046327_, _046328_, _046329_, _046330_, _046331_, _046332_, _046333_, _046334_, _046335_, _046336_, _046337_, _046338_, _046339_, _046340_, _046341_, _046342_, _046343_, _046344_, _046345_, _046346_, _046347_, _046348_, _046349_, _046350_, _046351_, _046352_, _046353_, _046354_, _046355_, _046356_, _046357_, _046358_, _046359_, _046360_, _046361_, _046362_, _046363_, _046364_, _046365_, _046366_, _046367_, _046368_, _046369_, _046370_, _046371_, _046372_, _046373_, _046374_, _046375_, _046376_, _046377_, _046378_, _046379_, _046380_, _046381_, _046382_, _046383_, _046384_, _046385_, _046386_, _046387_, _046388_, _046389_, _046390_, _046391_, _046392_, _046393_, _046394_, _046395_, _046396_, _046397_, _046398_, _046399_, _046400_, _046401_, _046402_, _046403_, _046404_, _046405_, _046406_, _046407_, _046408_, _046409_, _046410_, _046411_, _046412_, _046413_, _046414_, _046415_, _046416_, _046417_, _046418_, _046419_, _046420_, _046421_, _046422_, _046423_, _046424_, _046425_, _046426_, _046427_, _046428_, _046429_, _046430_, _046431_, _046432_, _046433_, _046434_, _046435_, _046436_, _046437_, _046438_, _046439_, _046440_, _046441_, _046442_, _046443_, _046444_, _046445_, _046446_, _046447_, _046448_, _046449_, _046450_, _046451_, _046452_, _046453_, _046454_, _046455_, _046456_, _046457_, _046458_, _046459_, _046460_, _046461_, _046462_, _046463_, _046464_, _046465_, _046466_, _046467_, _046468_, _046469_, _046470_, _046471_, _046472_, _046473_, _046474_, _046475_, _046476_, _046477_, _046478_, _046479_, _046480_, _046481_, _046482_, _046483_, _046484_, _046485_, _046486_, _046487_, _046488_, _046489_, _046490_, _046491_, _046492_, _046493_, _046494_, _046495_, _046496_, _046497_, _046498_, _046499_, _046500_, _046501_, _046502_, _046503_, _046504_, _046505_, _046506_, _046507_, _046508_, _046509_, _046510_, _046511_, _046512_, _046513_, _046514_, _046515_, _046516_, _046517_, _046518_, _046519_, _046520_, _046521_, _046522_, _046523_, _046524_, _046525_, _046526_, _046527_, _046528_, _046529_, _046530_, _046531_, _046532_, _046533_, _046534_, _046535_, _046536_, _046537_, _046538_, _046539_, _046540_, _046541_, _046542_, _046543_, _046544_, _046545_, _046546_, _046547_, _046548_, _046549_, _046550_, _046551_, _046552_, _046553_, _046554_, _046555_, _046556_, _046557_, _046558_, _046559_, _046560_, _046561_, _046562_, _046563_, _046564_, _046565_, _046566_, _046567_, _046568_, _046569_, _046570_, _046571_, _046572_, _046573_, _046574_, _046575_, _046576_, _046577_, _046578_, _046579_, _046580_, _046581_, _046582_, _046583_, _046584_, _046585_, _046586_, _046587_, _046588_, _046589_, _046590_, _046591_, _046592_, _046593_, _046594_, _046595_, _046596_, _046597_, _046598_, _046599_, _046600_, _046601_, _046602_, _046603_, _046604_, _046605_, _046606_, _046607_, _046608_, _046609_, _046610_, _046611_, _046612_, _046613_, _046614_, _046615_, _046616_, _046617_, _046618_, _046619_, _046620_, _046621_, _046622_, _046623_, _046624_, _046625_, _046626_, _046627_, _046628_, _046629_, _046630_, _046631_, _046632_, _046633_, _046634_, _046635_, _046636_, _046637_, _046638_, _046639_, _046640_, _046641_, _046642_, _046643_, _046644_, _046645_, _046646_, _046647_, _046648_, _046649_, _046650_, _046651_, _046652_, _046653_, _046654_, _046655_, _046656_, _046657_, _046658_, _046659_, _046660_, _046661_, _046662_, _046663_, _046664_, _046665_, _046666_, _046667_, _046668_, _046669_, _046670_, _046671_, _046672_, _046673_, _046674_, _046675_, _046676_, _046677_, _046678_, _046679_, _046680_, _046681_, _046682_, _046683_, _046684_, _046685_, _046686_, _046687_, _046688_, _046689_, _046690_, _046691_, _046692_, _046693_, _046694_, _046695_, _046696_, _046697_, _046698_, _046699_, _046700_, _046701_, _046702_, _046703_, _046704_, _046705_, _046706_, _046707_, _046708_, _046709_, _046710_, _046711_, _046712_, _046713_, _046714_, _046715_, _046716_, _046717_, _046718_, _046719_, _046720_, _046721_, _046722_, _046723_, _046724_, _046725_, _046726_, _046727_, _046728_, _046729_, _046730_, _046731_, _046732_, _046733_, _046734_, _046735_, _046736_, _046737_, _046738_, _046739_, _046740_, _046741_, _046742_, _046743_, _046744_, _046745_, _046746_, _046747_, _046748_, _046749_, _046750_, _046751_, _046752_, _046753_, _046754_, _046755_, _046756_, _046757_, _046758_, _046759_, _046760_, _046761_, _046762_, _046763_, _046764_, _046765_, _046766_, _046767_, _046768_, _046769_, _046770_, _046771_, _046772_, _046773_, _046774_, _046775_, _046776_, _046777_, _046778_, _046779_, _046780_, _046781_, _046782_, _046783_, _046784_, _046785_, _046786_, _046787_, _046788_, _046789_, _046790_, _046791_, _046792_, _046793_, _046794_, _046795_, _046796_, _046797_, _046798_, _046799_, _046800_, _046801_, _046802_, _046803_, _046804_, _046805_, _046806_, _046807_, _046808_, _046809_, _046810_, _046811_, _046812_, _046813_, _046814_, _046815_, _046816_, _046817_, _046818_, _046819_, _046820_, _046821_, _046822_, _046823_, _046824_, _046825_, _046826_, _046827_, _046828_, _046829_, _046830_, _046831_, _046832_, _046833_, _046834_, _046835_, _046836_, _046837_, _046838_, _046839_, _046840_, _046841_, _046842_, _046843_, _046844_, _046845_, _046846_, _046847_, _046848_, _046849_, _046850_, _046851_, _046852_, _046853_, _046854_, _046855_, _046856_, _046857_, _046858_, _046859_, _046860_, _046861_, _046862_, _046863_, _046864_, _046865_, _046866_, _046867_, _046868_, _046869_, _046870_, _046871_, _046872_, _046873_, _046874_, _046875_, _046876_, _046877_, _046878_, _046879_, _046880_, _046881_, _046882_, _046883_, _046884_, _046885_, _046886_, _046887_, _046888_, _046889_, _046890_, _046891_, _046892_, _046893_, _046894_, _046895_, _046896_, _046897_, _046898_, _046899_, _046900_, _046901_, _046902_, _046903_, _046904_, _046905_, _046906_, _046907_, _046908_, _046909_, _046910_, _046911_, _046912_, _046913_, _046914_, _046915_, _046916_, _046917_, _046918_, _046919_, _046920_, _046921_, _046922_, _046923_, _046924_, _046925_, _046926_, _046927_, _046928_, _046929_, _046930_, _046931_, _046932_, _046933_, _046934_, _046935_, _046936_, _046937_, _046938_, _046939_, _046940_, _046941_, _046942_, _046943_, _046944_, _046945_, _046946_, _046947_, _046948_, _046949_, _046950_, _046951_, _046952_, _046953_, _046954_, _046955_, _046956_, _046957_, _046958_, _046959_, _046960_, _046961_, _046962_, _046963_, _046964_, _046965_, _046966_, _046967_, _046968_, _046969_, _046970_, _046971_, _046972_, _046973_, _046974_, _046975_, _046976_, _046977_, _046978_, _046979_, _046980_, _046981_, _046982_, _046983_, _046984_, _046985_, _046986_, _046987_, _046988_, _046989_, _046990_, _046991_, _046992_, _046993_, _046994_, _046995_, _046996_, _046997_, _046998_, _046999_, _047000_, _047001_, _047002_, _047003_, _047004_, _047005_, _047006_, _047007_, _047008_, _047009_, _047010_, _047011_, _047012_, _047013_, _047014_, _047015_, _047016_, _047017_, _047018_, _047019_, _047020_, _047021_, _047022_, _047023_, _047024_, _047025_, _047026_, _047027_, _047028_, _047029_, _047030_, _047031_, _047032_, _047033_, _047034_, _047035_, _047036_, _047037_, _047038_, _047039_, _047040_, _047041_, _047042_, _047043_, _047044_, _047045_, _047046_, _047047_, _047048_, _047049_, _047050_, _047051_, _047052_, _047053_, _047054_, _047055_, _047056_, _047057_, _047058_, _047059_, _047060_, _047061_, _047062_, _047063_, _047064_, _047065_, _047066_, _047067_, _047068_, _047069_, _047070_, _047071_, _047072_, _047073_, _047074_, _047075_, _047076_, _047077_, _047078_, _047079_, _047080_, _047081_, _047082_, _047083_, _047084_, _047085_, _047086_, _047087_, _047088_, _047089_, _047090_, _047091_, _047092_, _047093_, _047094_, _047095_, _047096_, _047097_, _047098_, _047099_, _047100_, _047101_, _047102_, _047103_, _047104_, _047105_, _047106_, _047107_, _047108_, _047109_, _047110_, _047111_, _047112_, _047113_, _047114_, _047115_, _047116_, _047117_, _047118_, _047119_, _047120_, _047121_, _047122_, _047123_, _047124_, _047125_, _047126_, _047127_, _047128_, _047129_, _047130_, _047131_, _047132_, _047133_, _047134_, _047135_, _047136_, _047137_, _047138_, _047139_, _047140_, _047141_, _047142_, _047143_, _047144_, _047145_, _047146_, _047147_, _047148_, _047149_, _047150_, _047151_, _047152_, _047153_, _047154_, _047155_, _047156_, _047157_, _047158_, _047159_, _047160_, _047161_, _047162_, _047163_, _047164_, _047165_, _047166_, _047167_, _047168_, _047169_, _047170_, _047171_, _047172_, _047173_, _047174_, _047175_, _047176_, _047177_, _047178_, _047179_, _047180_, _047181_, _047182_, _047183_, _047184_, _047185_, _047186_, _047187_, _047188_, _047189_, _047190_, _047191_, _047192_, _047193_, _047194_, _047195_, _047196_, _047197_, _047198_, _047199_, _047200_, _047201_, _047202_, _047203_, _047204_, _047205_, _047206_, _047207_, _047208_, _047209_, _047210_, _047211_, _047212_, _047213_, _047214_, _047215_, _047216_, _047217_, _047218_, _047219_, _047220_, _047221_, _047222_, _047223_, _047224_, _047225_, _047226_, _047227_, _047228_, _047229_, _047230_, _047231_, _047232_, _047233_, _047234_, _047235_, _047236_, _047237_, _047238_, _047239_, _047240_, _047241_, _047242_, _047243_, _047244_, _047245_, _047246_, _047247_, _047248_, _047249_, _047250_, _047251_, _047252_, _047253_, _047254_, _047255_, _047256_, _047257_, _047258_, _047259_, _047260_, _047261_, _047262_, _047263_, _047264_, _047265_, _047266_, _047267_, _047268_, _047269_, _047270_, _047271_, _047272_, _047273_, _047274_, _047275_, _047276_, _047277_, _047278_, _047279_, _047280_, _047281_, _047282_, _047283_, _047284_, _047285_, _047286_, _047287_, _047288_, _047289_, _047290_, _047291_, _047292_, _047293_, _047294_, _047295_, _047296_, _047297_, _047298_, _047299_, _047300_, _047301_, _047302_, _047303_, _047304_, _047305_, _047306_, _047307_, _047308_, _047309_, _047310_, _047311_, _047312_, _047313_, _047314_, _047315_, _047316_, _047317_, _047318_, _047319_, _047320_, _047321_, _047322_, _047323_, _047324_, _047325_, _047326_, _047327_, _047328_, _047329_, _047330_, _047331_, _047332_, _047333_, _047334_, _047335_, _047336_, _047337_, _047338_, _047339_, _047340_, _047341_, _047342_, _047343_, _047344_, _047345_, _047346_, _047347_, _047348_, _047349_, _047350_, _047351_, _047352_, _047353_, _047354_, _047355_, _047356_, _047357_, _047358_, _047359_, _047360_, _047361_, _047362_, _047363_, _047364_, _047365_, _047366_, _047367_, _047368_, _047369_, _047370_, _047371_, _047372_, _047373_, _047374_, _047375_, _047376_, _047377_, _047378_, _047379_, _047380_, _047381_, _047382_, _047383_, _047384_, _047385_, _047386_, _047387_, _047388_, _047389_, _047390_, _047391_, _047392_, _047393_, _047394_, _047395_, _047396_, _047397_, _047398_, _047399_, _047400_, _047401_, _047402_, _047403_, _047404_, _047405_, _047406_, _047407_, _047408_, _047409_, _047410_, _047411_, _047412_, _047413_, _047414_, _047415_, _047416_, _047417_, _047418_, _047419_, _047420_, _047421_, _047422_, _047423_, _047424_, _047425_, _047426_, _047427_, _047428_, _047429_, _047430_, _047431_, _047432_, _047433_, _047434_, _047435_, _047436_, _047437_, _047438_, _047439_, _047440_, _047441_, _047442_, _047443_, _047444_, _047445_, _047446_, _047447_, _047448_, _047449_, _047450_, _047451_, _047452_, _047453_, _047454_, _047455_, _047456_, _047457_, _047458_, _047459_, _047460_, _047461_, _047462_, _047463_, _047464_, _047465_, _047466_, _047467_, _047468_, _047469_, _047470_, _047471_, _047472_, _047473_, _047474_, _047475_, _047476_, _047477_, _047478_, _047479_, _047480_, _047481_, _047482_, _047483_, _047484_, _047485_, _047486_, _047487_, _047488_, _047489_, _047490_, _047491_, _047492_, _047493_, _047494_, _047495_, _047496_, _047497_, _047498_, _047499_, _047500_, _047501_, _047502_, _047503_, _047504_, _047505_, _047506_, _047507_, _047508_, _047509_, _047510_, _047511_, _047512_, _047513_, _047514_, _047515_, _047516_, _047517_, _047518_, _047519_, _047520_, _047521_, _047522_, _047523_, _047524_, _047525_, _047526_, _047527_, _047528_, _047529_, _047530_, _047531_, _047532_, _047533_, _047534_, _047535_, _047536_, _047537_, _047538_, _047539_, _047540_, _047541_, _047542_, _047543_, _047544_, _047545_, _047546_, _047547_, _047548_, _047549_, _047550_, _047551_, _047552_, _047553_, _047554_, _047555_, _047556_, _047557_, _047558_, _047559_, _047560_, _047561_, _047562_, _047563_, _047564_, _047565_, _047566_, _047567_, _047568_, _047569_, _047570_, _047571_, _047572_, _047573_, _047574_, _047575_, _047576_, _047577_, _047578_, _047579_, _047580_, _047581_, _047582_, _047583_, _047584_, _047585_, _047586_, _047587_, _047588_, _047589_, _047590_, _047591_, _047592_, _047593_, _047594_, _047595_, _047596_, _047597_, _047598_, _047599_, _047600_, _047601_, _047602_, _047603_, _047604_, _047605_, _047606_, _047607_, _047608_, _047609_, _047610_, _047611_, _047612_, _047613_, _047614_, _047615_, _047616_, _047617_, _047618_, _047619_, _047620_, _047621_, _047622_, _047623_, _047624_, _047625_, _047626_, _047627_, _047628_, _047629_, _047630_, _047631_, _047632_, _047633_, _047634_, _047635_, _047636_, _047637_, _047638_, _047639_, _047640_, _047641_, _047642_, _047643_, _047644_, _047645_, _047646_, _047647_, _047648_, _047649_, _047650_, _047651_, _047652_, _047653_, _047654_, _047655_, _047656_, _047657_, _047658_, _047659_, _047660_, _047661_, _047662_, _047663_, _047664_, _047665_, _047666_, _047667_, _047668_, _047669_, _047670_, _047671_, _047672_, _047673_, _047674_, _047675_, _047676_, _047677_, _047678_, _047679_, _047680_, _047681_, _047682_, _047683_, _047684_, _047685_, _047686_, _047687_, _047688_, _047689_, _047690_, _047691_, _047692_, _047693_, _047694_, _047695_, _047696_, _047697_, _047698_, _047699_, _047700_, _047701_, _047702_, _047703_, _047704_, _047705_, _047706_, _047707_, _047708_, _047709_, _047710_, _047711_, _047712_, _047713_, _047714_, _047715_, _047716_, _047717_, _047718_, _047719_, _047720_, _047721_, _047722_, _047723_, _047724_, _047725_, _047726_, _047727_, _047728_, _047729_, _047730_, _047731_, _047732_, _047733_, _047734_, _047735_, _047736_, _047737_, _047738_, _047739_, _047740_, _047741_, _047742_, _047743_, _047744_, _047745_, _047746_, _047747_, _047748_, _047749_, _047750_, _047751_, _047752_, _047753_, _047754_, _047755_, _047756_, _047757_, _047758_, _047759_, _047760_, _047761_, _047762_, _047763_, _047764_, _047765_, _047766_, _047767_, _047768_, _047769_, _047770_, _047771_, _047772_, _047773_, _047774_, _047775_, _047776_, _047777_, _047778_, _047779_, _047780_, _047781_, _047782_, _047783_, _047784_, _047785_, _047786_, _047787_, _047788_, _047789_, _047790_, _047791_, _047792_, _047793_, _047794_, _047795_, _047796_, _047797_, _047798_, _047799_, _047800_, _047801_, _047802_, _047803_, _047804_, _047805_, _047806_, _047807_, _047808_, _047809_, _047810_, _047811_, _047812_, _047813_, _047814_, _047815_, _047816_, _047817_, _047818_, _047819_, _047820_, _047821_, _047822_, _047823_, _047824_, _047825_, _047826_, _047827_, _047828_, _047829_, _047830_, _047831_, _047832_, _047833_, _047834_, _047835_, _047836_, _047837_, _047838_, _047839_, _047840_, _047841_, _047842_, _047843_, _047844_, _047845_, _047846_, _047847_, _047848_, _047849_, _047850_, _047851_, _047852_, _047853_, _047854_, _047855_, _047856_, _047857_, _047858_, _047859_, _047860_, _047861_, _047862_, _047863_, _047864_, _047865_, _047866_, _047867_, _047868_, _047869_, _047870_, _047871_, _047872_, _047873_, _047874_, _047875_, _047876_, _047877_, _047878_, _047879_, _047880_, _047881_, _047882_, _047883_, _047884_, _047885_, _047886_, _047887_, _047888_, _047889_, _047890_, _047891_, _047892_, _047893_, _047894_, _047895_, _047896_, _047897_, _047898_, _047899_, _047900_, _047901_, _047902_, _047903_, _047904_, _047905_, _047906_, _047907_, _047908_, _047909_, _047910_, _047911_, _047912_, _047913_, _047914_, _047915_, _047916_, _047917_, _047918_, _047919_, _047920_, _047921_, _047922_, _047923_, _047924_, _047925_, _047926_, _047927_, _047928_, _047929_, _047930_, _047931_, _047932_, _047933_, _047934_, _047935_, _047936_, _047937_, _047938_, _047939_, _047940_, _047941_, _047942_, _047943_, _047944_, _047945_, _047946_, _047947_, _047948_, _047949_, _047950_, _047951_, _047952_, _047953_, _047954_, _047955_, _047956_, _047957_, _047958_, _047959_, _047960_, _047961_, _047962_, _047963_, _047964_, _047965_, _047966_, _047967_, _047968_, _047969_, _047970_, _047971_, _047972_, _047973_, _047974_, _047975_, _047976_, _047977_, _047978_, _047979_, _047980_, _047981_, _047982_, _047983_, _047984_, _047985_, _047986_, _047987_, _047988_, _047989_, _047990_, _047991_, _047992_, _047993_, _047994_, _047995_, _047996_, _047997_, _047998_, _047999_, _048000_, _048001_, _048002_, _048003_, _048004_, _048005_, _048006_, _048007_, _048008_, _048009_, _048010_, _048011_, _048012_, _048013_, _048014_, _048015_, _048016_, _048017_, _048018_, _048019_, _048020_, _048021_, _048022_, _048023_, _048024_, _048025_, _048026_, _048027_, _048028_, _048029_, _048030_, _048031_, _048032_, _048033_, _048034_, _048035_, _048036_, _048037_, _048038_, _048039_, _048040_, _048041_, _048042_, _048043_, _048044_, _048045_, _048046_, _048047_, _048048_, _048049_, _048050_, _048051_, _048052_, _048053_, _048054_, _048055_, _048056_, _048057_, _048058_, _048059_, _048060_, _048061_, _048062_, _048063_, _048064_, _048065_, _048066_, _048067_, _048068_, _048069_, _048070_, _048071_, _048072_, _048073_, _048074_, _048075_, _048076_, _048077_, _048078_, _048079_, _048080_, _048081_, _048082_, _048083_, _048084_, _048085_, _048086_, _048087_, _048088_, _048089_, _048090_, _048091_, _048092_, _048093_, _048094_, _048095_, _048096_, _048097_, _048098_, _048099_, _048100_, _048101_, _048102_, _048103_, _048104_, _048105_, _048106_, _048107_, _048108_, _048109_, _048110_, _048111_, _048112_, _048113_, _048114_, _048115_, _048116_, _048117_, _048118_, _048119_, _048120_, _048121_, _048122_, _048123_, _048124_, _048125_, _048126_, _048127_, _048128_, _048129_, _048130_, _048131_, _048132_, _048133_, _048134_, _048135_, _048136_, _048137_, _048138_, _048139_, _048140_, _048141_, _048142_, _048143_, _048144_, _048145_, _048146_, _048147_, _048148_, _048149_, _048150_, _048151_, _048152_, _048153_, _048154_, _048155_, _048156_, _048157_, _048158_, _048159_, _048160_, _048161_, _048162_, _048163_, _048164_, _048165_, _048166_, _048167_, _048168_, _048169_, _048170_, _048171_, _048172_, _048173_, _048174_, _048175_, _048176_, _048177_, _048178_, _048179_, _048180_, _048181_, _048182_, _048183_, _048184_, _048185_, _048186_, _048187_, _048188_, _048189_, _048190_, _048191_, _048192_, _048193_, _048194_, _048195_, _048196_, _048197_, _048198_, _048199_, _048200_, _048201_, _048202_, _048203_, _048204_, _048205_, _048206_, _048207_, _048208_, _048209_, _048210_, _048211_, _048212_, _048213_, _048214_, _048215_, _048216_, _048217_, _048218_, _048219_, _048220_, _048221_, _048222_, _048223_, _048224_, _048225_, _048226_, _048227_, _048228_, _048229_, _048230_, _048231_, _048232_, _048233_, _048234_, _048235_, _048236_, _048237_, _048238_, _048239_, _048240_, _048241_, _048242_, _048243_, _048244_, _048245_, _048246_, _048247_, _048248_, _048249_, _048250_, _048251_, _048252_, _048253_, _048254_, _048255_, _048256_, _048257_, _048258_, _048259_, _048260_, _048261_, _048262_, _048263_, _048264_, _048265_, _048266_, _048267_, _048268_, _048269_, _048270_, _048271_, _048272_, _048273_, _048274_, _048275_, _048276_, _048277_, _048278_, _048279_, _048280_, _048281_, _048282_, _048283_, _048284_, _048285_, _048286_, _048287_, _048288_, _048289_, _048290_, _048291_, _048292_, _048293_, _048294_, _048295_, _048296_, _048297_, _048298_, _048299_, _048300_, _048301_, _048302_, _048303_, _048304_, _048305_, _048306_, _048307_, _048308_, _048309_, _048310_, _048311_, _048312_, _048313_, _048314_, _048315_, _048316_, _048317_, _048318_, _048319_, _048320_, _048321_, _048322_, _048323_, _048324_, _048325_, _048326_, _048327_, _048328_, _048329_, _048330_, _048331_, _048332_, _048333_, _048334_, _048335_, _048336_, _048337_, _048338_, _048339_, _048340_, _048341_, _048342_, _048343_, _048344_, _048345_, _048346_, _048347_, _048348_, _048349_, _048350_, _048351_, _048352_, _048353_, _048354_, _048355_, _048356_, _048357_, _048358_, _048359_, _048360_, _048361_, _048362_, _048363_, _048364_, _048365_, _048366_, _048367_, _048368_, _048369_, _048370_, _048371_, _048372_, _048373_, _048374_, _048375_, _048376_, _048377_, _048378_, _048379_, _048380_, _048381_, _048382_, _048383_, _048384_, _048385_, _048386_, _048387_, _048388_, _048389_, _048390_, _048391_, _048392_, _048393_, _048394_, _048395_, _048396_, _048397_, _048398_, _048399_, _048400_, _048401_, _048402_, _048403_, _048404_, _048405_, _048406_, _048407_, _048408_, _048409_, _048410_, _048411_, _048412_, _048413_, _048414_, _048415_, _048416_, _048417_, _048418_, _048419_, _048420_, _048421_, _048422_, _048423_, _048424_, _048425_, _048426_, _048427_, _048428_, _048429_, _048430_, _048431_, _048432_, _048433_, _048434_, _048435_, _048436_, _048437_, _048438_, _048439_, _048440_, _048441_, _048442_, _048443_, _048444_, _048445_, _048446_, _048447_, _048448_, _048449_, _048450_, _048451_, _048452_, _048453_, _048454_, _048455_, _048456_, _048457_, _048458_, _048459_, _048460_, _048461_, _048462_, _048463_, _048464_, _048465_, _048466_, _048467_, _048468_, _048469_, _048470_, _048471_, _048472_, _048473_, _048474_, _048475_, _048476_, _048477_, _048478_, _048479_, _048480_, _048481_, _048482_, _048483_, _048484_, _048485_, _048486_, _048487_, _048488_, _048489_, _048490_, _048491_, _048492_, _048493_, _048494_, _048495_, _048496_, _048497_, _048498_, _048499_, _048500_, _048501_, _048502_, _048503_, _048504_, _048505_, _048506_, _048507_, _048508_, _048509_, _048510_, _048511_, _048512_, _048513_, _048514_, _048515_, _048516_, _048517_, _048518_, _048519_, _048520_, _048521_, _048522_, _048523_, _048524_, _048525_, _048526_, _048527_, _048528_, _048529_, _048530_, _048531_, _048532_, _048533_, _048534_, _048535_, _048536_, _048537_, _048538_, _048539_, _048540_, _048541_, _048542_, _048543_, _048544_, _048545_, _048546_, _048547_, _048548_, _048549_, _048550_, _048551_, _048552_, _048553_, _048554_, _048555_, _048556_, _048557_, _048558_, _048559_, _048560_, _048561_, _048562_, _048563_, _048564_, _048565_, _048566_, _048567_, _048568_, _048569_, _048570_, _048571_, _048572_, _048573_, _048574_, _048575_, _048576_, _048577_, _048578_, _048579_, _048580_, _048581_, _048582_, _048583_, _048584_, _048585_, _048586_, _048587_, _048588_, _048589_, _048590_, _048591_, _048592_, _048593_, _048594_, _048595_, _048596_, _048597_, _048598_, _048599_, _048600_, _048601_, _048602_, _048603_, _048604_, _048605_, _048606_, _048607_, _048608_, _048609_, _048610_, _048611_, _048612_, _048613_, _048614_, _048615_, _048616_, _048617_, _048618_, _048619_, _048620_, _048621_, _048622_, _048623_, _048624_, _048625_, _048626_, _048627_, _048628_, _048629_, _048630_, _048631_, _048632_, _048633_, _048634_, _048635_, _048636_, _048637_, _048638_, _048639_, _048640_, _048641_, _048642_, _048643_, _048644_, _048645_, _048646_, _048647_, _048648_, _048649_, _048650_, _048651_, _048652_, _048653_, _048654_, _048655_, _048656_, _048657_, _048658_, _048659_, _048660_, _048661_, _048662_, _048663_, _048664_, _048665_, _048666_, _048667_, _048668_, _048669_, _048670_, _048671_, _048672_, _048673_, _048674_, _048675_, _048676_, _048677_, _048678_, _048679_, _048680_, _048681_, _048682_, _048683_, _048684_, _048685_, _048686_, _048687_, _048688_, _048689_, _048690_, _048691_, _048692_, _048693_, _048694_, _048695_, _048696_, _048697_, _048698_, _048699_, _048700_, _048701_, _048702_, _048703_, _048704_, _048705_, _048706_, _048707_, _048708_, _048709_, _048710_, _048711_, _048712_, _048713_, _048714_, _048715_, _048716_, _048717_, _048718_, _048719_, _048720_, _048721_, _048722_, _048723_, _048724_, _048725_, _048726_, _048727_, _048728_, _048729_, _048730_, _048731_, _048732_, _048733_, _048734_, _048735_, _048736_, _048737_, _048738_, _048739_, _048740_, _048741_, _048742_, _048743_, _048744_, _048745_, _048746_, _048747_, _048748_, _048749_, _048750_, _048751_, _048752_, _048753_, _048754_, _048755_, _048756_, _048757_, _048758_, _048759_, _048760_, _048761_, _048762_, _048763_, _048764_, _048765_, _048766_, _048767_, _048768_, _048769_, _048770_, _048771_, _048772_, _048773_, _048774_, _048775_, _048776_, _048777_, _048778_, _048779_, _048780_, _048781_, _048782_, _048783_, _048784_, _048785_, _048786_, _048787_, _048788_, _048789_, _048790_, _048791_, _048792_, _048793_, _048794_, _048795_, _048796_, _048797_, _048798_, _048799_, _048800_, _048801_, _048802_, _048803_, _048804_, _048805_, _048806_, _048807_, _048808_, _048809_, _048810_, _048811_, _048812_, _048813_, _048814_, _048815_, _048816_, _048817_, _048818_, _048819_, _048820_, _048821_, _048822_, _048823_, _048824_, _048825_, _048826_, _048827_, _048828_, _048829_, _048830_, _048831_, _048832_, _048833_, _048834_, _048835_, _048836_, _048837_, _048838_, _048839_, _048840_, _048841_, _048842_, _048843_, _048844_, _048845_, _048846_, _048847_, _048848_, _048849_, _048850_, _048851_, _048852_, _048853_, _048854_, _048855_, _048856_, _048857_, _048858_, _048859_, _048860_, _048861_, _048862_, _048863_, _048864_, _048865_, _048866_, _048867_, _048868_, _048869_, _048870_, _048871_, _048872_, _048873_, _048874_, _048875_, _048876_, _048877_, _048878_, _048879_, _048880_, _048881_, _048882_, _048883_, _048884_, _048885_, _048886_, _048887_, _048888_, _048889_, _048890_, _048891_, _048892_, _048893_, _048894_, _048895_, _048896_, _048897_, _048898_, _048899_, _048900_, _048901_, _048902_, _048903_, _048904_, _048905_, _048906_, _048907_, _048908_, _048909_, _048910_, _048911_, _048912_, _048913_, _048914_, _048915_, _048916_, _048917_, _048918_, _048919_, _048920_, _048921_, _048922_, _048923_, _048924_, _048925_, _048926_, _048927_, _048928_, _048929_, _048930_, _048931_, _048932_, _048933_, _048934_, _048935_, _048936_, _048937_, _048938_, _048939_, _048940_, _048941_, _048942_, _048943_, _048944_, _048945_, _048946_, _048947_, _048948_, _048949_, _048950_, _048951_, _048952_, _048953_, _048954_, _048955_, _048956_, _048957_, _048958_, _048959_, _048960_, _048961_, _048962_, _048963_, _048964_, _048965_, _048966_, _048967_, _048968_, _048969_, _048970_, _048971_, _048972_, _048973_, _048974_, _048975_, _048976_, _048977_, _048978_, _048979_, _048980_, _048981_, _048982_, _048983_, _048984_, _048985_, _048986_, _048987_, _048988_, _048989_, _048990_, _048991_, _048992_, _048993_, _048994_, _048995_, _048996_, _048997_, _048998_, _048999_, _049000_, _049001_, _049002_, _049003_, _049004_, _049005_, _049006_, _049007_, _049008_, _049009_, _049010_, _049011_, _049012_, _049013_, _049014_, _049015_, _049016_, _049017_, _049018_, _049019_, _049020_, _049021_, _049022_, _049023_, _049024_, _049025_, _049026_, _049027_, _049028_, _049029_, _049030_, _049031_, _049032_, _049033_, _049034_, _049035_, _049036_, _049037_, _049038_, _049039_, _049040_, _049041_, _049042_, _049043_, _049044_, _049045_, _049046_, _049047_, _049048_, _049049_, _049050_, _049051_, _049052_, _049053_, _049054_, _049055_, _049056_, _049057_, _049058_, _049059_, _049060_, _049061_, _049062_, _049063_, _049064_, _049065_, _049066_, _049067_, _049068_, _049069_, _049070_, _049071_, _049072_, _049073_, _049074_, _049075_, _049076_, _049077_, _049078_, _049079_, _049080_, _049081_, _049082_, _049083_, _049084_, _049085_, _049086_, _049087_, _049088_, _049089_, _049090_, _049091_, _049092_, _049093_, _049094_, _049095_, _049096_, _049097_, _049098_, _049099_, _049100_, _049101_, _049102_, _049103_, _049104_, _049105_, _049106_, _049107_, _049108_, _049109_, _049110_, _049111_, _049112_, _049113_, _049114_, _049115_, _049116_, _049117_, _049118_, _049119_, _049120_, _049121_, _049122_, _049123_, _049124_, _049125_, _049126_, _049127_, _049128_, _049129_, _049130_, _049131_, _049132_, _049133_, _049134_, _049135_, _049136_, _049137_, _049138_, _049139_, _049140_, _049141_, _049142_, _049143_, _049144_, _049145_, _049146_, _049147_, _049148_, _049149_, _049150_, _049151_, _049152_, _049153_, _049154_, _049155_, _049156_, _049157_, _049158_, _049159_, _049160_, _049161_, _049162_, _049163_, _049164_, _049165_, _049166_, _049167_, _049168_, _049169_, _049170_, _049171_, _049172_, _049173_, _049174_, _049175_, _049176_, _049177_, _049178_, _049179_, _049180_, _049181_, _049182_, _049183_, _049184_, _049185_, _049186_, _049187_, _049188_, _049189_, _049190_, _049191_, _049192_, _049193_, _049194_, _049195_, _049196_, _049197_, _049198_, _049199_, _049200_, _049201_, _049202_, _049203_, _049204_, _049205_, _049206_, _049207_, _049208_, _049209_, _049210_, _049211_, _049212_, _049213_, _049214_, _049215_, _049216_, _049217_, _049218_, _049219_, _049220_, _049221_, _049222_, _049223_, _049224_, _049225_, _049226_, _049227_, _049228_, _049229_, _049230_, _049231_, _049232_, _049233_, _049234_, _049235_, _049236_, _049237_, _049238_, _049239_, _049240_, _049241_, _049242_, _049243_, _049244_, _049245_, _049246_, _049247_, _049248_, _049249_, _049250_, _049251_, _049252_, _049253_, _049254_, _049255_, _049256_, _049257_, _049258_, _049259_, _049260_, _049261_, _049262_, _049263_, _049264_, _049265_, _049266_, _049267_, _049268_, _049269_, _049270_, _049271_, _049272_, _049273_, _049274_, _049275_, _049276_, _049277_, _049278_, _049279_, _049280_, _049281_, _049282_, _049283_, _049284_, _049285_, _049286_, _049287_, _049288_, _049289_, _049290_, _049291_, _049292_, _049293_, _049294_, _049295_, _049296_, _049297_, _049298_, _049299_, _049300_, _049301_, _049302_, _049303_, _049304_, _049305_, _049306_, _049307_, _049308_, _049309_, _049310_, _049311_, _049312_, _049313_, _049314_, _049315_, _049316_, _049317_, _049318_, _049319_, _049320_, _049321_, _049322_, _049323_, _049324_, _049325_, _049326_, _049327_, _049328_, _049329_, _049330_, _049331_, _049332_, _049333_, _049334_, _049335_, _049336_, _049337_, _049338_, _049339_, _049340_, _049341_, _049342_, _049343_, _049344_, _049345_, _049346_, _049347_, _049348_, _049349_, _049350_, _049351_, _049352_, _049353_, _049354_, _049355_, _049356_, _049357_, _049358_, _049359_, _049360_, _049361_, _049362_, _049363_, _049364_, _049365_, _049366_, _049367_, _049368_, _049369_, _049370_, _049371_, _049372_, _049373_, _049374_, _049375_, _049376_, _049377_, _049378_, _049379_, _049380_, _049381_, _049382_, _049383_, _049384_, _049385_, _049386_, _049387_, _049388_, _049389_, _049390_, _049391_, _049392_, _049393_, _049394_, _049395_, _049396_, _049397_, _049398_, _049399_, _049400_, _049401_, _049402_, _049403_, _049404_, _049405_, _049406_, _049407_, _049408_, _049409_, _049410_, _049411_, _049412_, _049413_, _049414_, _049415_, _049416_, _049417_, _049418_, _049419_, _049420_, _049421_, _049422_, _049423_, _049424_, _049425_, _049426_, _049427_, _049428_, _049429_, _049430_, _049431_, _049432_, _049433_, _049434_, _049435_, _049436_, _049437_, _049438_, _049439_, _049440_, _049441_, _049442_, _049443_, _049444_, _049445_, _049446_, _049447_, _049448_, _049449_, _049450_, _049451_, _049452_, _049453_, _049454_, _049455_, _049456_, _049457_, _049458_, _049459_, _049460_, _049461_, _049462_, _049463_, _049464_, _049465_, _049466_, _049467_, _049468_, _049469_, _049470_, _049471_, _049472_, _049473_, _049474_, _049475_, _049476_, _049477_, _049478_, _049479_, _049480_, _049481_, _049482_, _049483_, _049484_, _049485_, _049486_, _049487_, _049488_, _049489_, _049490_, _049491_, _049492_, _049493_, _049494_, _049495_, _049496_, _049497_, _049498_, _049499_, _049500_, _049501_, _049502_, _049503_, _049504_, _049505_, _049506_, _049507_, _049508_, _049509_, _049510_, _049511_, _049512_, _049513_, _049514_, _049515_, _049516_, _049517_, _049518_, _049519_, _049520_, _049521_, _049522_, _049523_, _049524_, _049525_, _049526_, _049527_, _049528_, _049529_, _049530_, _049531_, _049532_, _049533_, _049534_, _049535_, _049536_, _049537_, _049538_, _049539_, _049540_, _049541_, _049542_, _049543_, _049544_, _049545_, _049546_, _049547_, _049548_, _049549_, _049550_, _049551_, _049552_, _049553_, _049554_, _049555_, _049556_, _049557_, _049558_, _049559_, _049560_, _049561_, _049562_, _049563_, _049564_, _049565_, _049566_, _049567_, _049568_, _049569_, _049570_, _049571_, _049572_, _049573_, _049574_, _049575_, _049576_, _049577_, _049578_, _049579_, _049580_, _049581_, _049582_, _049583_, _049584_, _049585_, _049586_, _049587_, _049588_, _049589_, _049590_, _049591_, _049592_, _049593_, _049594_, _049595_, _049596_, _049597_, _049598_, _049599_, _049600_, _049601_, _049602_, _049603_, _049604_, _049605_, _049606_, _049607_, _049608_, _049609_, _049610_, _049611_, _049612_, _049613_, _049614_, _049615_, _049616_, _049617_, _049618_, _049619_, _049620_, _049621_, _049622_, _049623_, _049624_, _049625_, _049626_, _049627_, _049628_, _049629_, _049630_, _049631_, _049632_, _049633_, _049634_, _049635_, _049636_, _049637_, _049638_, _049639_, _049640_, _049641_, _049642_, _049643_, _049644_, _049645_, _049646_, _049647_, _049648_, _049649_, _049650_, _049651_, _049652_, _049653_, _049654_, _049655_, _049656_, _049657_, _049658_, _049659_, _049660_, _049661_, _049662_, _049663_, _049664_, _049665_, _049666_, _049667_, _049668_, _049669_, _049670_, _049671_, _049672_, _049673_, _049674_, _049675_, _049676_, _049677_, _049678_, _049679_, _049680_, _049681_, _049682_, _049683_, _049684_, _049685_, _049686_, _049687_, _049688_, _049689_, _049690_, _049691_, _049692_, _049693_, _049694_, _049695_, _049696_, _049697_, _049698_, _049699_, _049700_, _049701_, _049702_, _049703_, _049704_, _049705_, _049706_, _049707_, _049708_, _049709_, _049710_, _049711_, _049712_, _049713_, _049714_, _049715_, _049716_, _049717_, _049718_, _049719_, _049720_, _049721_, _049722_, _049723_, _049724_, _049725_, _049726_, _049727_, _049728_, _049729_, _049730_, _049731_, _049732_, _049733_, _049734_, _049735_, _049736_, _049737_, _049738_, _049739_, _049740_, _049741_, _049742_, _049743_, _049744_, _049745_, _049746_, _049747_, _049748_, _049749_, _049750_, _049751_, _049752_, _049753_, _049754_, _049755_, _049756_, _049757_, _049758_, _049759_, _049760_, _049761_, _049762_, _049763_, _049764_, _049765_, _049766_, _049767_, _049768_, _049769_, _049770_, _049771_, _049772_, _049773_, _049774_, _049775_, _049776_, _049777_, _049778_, _049779_, _049780_, _049781_, _049782_, _049783_, _049784_, _049785_, _049786_, _049787_, _049788_, _049789_, _049790_, _049791_, _049792_, _049793_, _049794_, _049795_, _049796_, _049797_, _049798_, _049799_, _049800_, _049801_, _049802_, _049803_, _049804_, _049805_, _049806_, _049807_, _049808_, _049809_, _049810_, _049811_, _049812_, _049813_, _049814_, _049815_, _049816_, _049817_, _049818_, _049819_, _049820_, _049821_, _049822_, _049823_, _049824_, _049825_, _049826_, _049827_, _049828_, _049829_, _049830_, _049831_, _049832_, _049833_, _049834_, _049835_, _049836_, _049837_, _049838_, _049839_, _049840_, _049841_, _049842_, _049843_, _049844_, _049845_, _049846_, _049847_, _049848_, _049849_, _049850_, _049851_, _049852_, _049853_, _049854_, _049855_, _049856_, _049857_, _049858_, _049859_, _049860_, _049861_, _049862_, _049863_, _049864_, _049865_, _049866_, _049867_, _049868_, _049869_, _049870_, _049871_, _049872_, _049873_, _049874_, _049875_, _049876_, _049877_, _049878_, _049879_, _049880_, _049881_, _049882_, _049883_, _049884_, _049885_, _049886_, _049887_, _049888_, _049889_, _049890_, _049891_, _049892_, _049893_, _049894_, _049895_, _049896_, _049897_, _049898_, _049899_, _049900_, _049901_, _049902_, _049903_, _049904_, _049905_, _049906_, _049907_, _049908_, _049909_, _049910_, _049911_, _049912_, _049913_, _049914_, _049915_, _049916_, _049917_, _049918_, _049919_, _049920_, _049921_, _049922_, _049923_, _049924_, _049925_, _049926_, _049927_, _049928_, _049929_, _049930_, _049931_, _049932_, _049933_, _049934_, _049935_, _049936_, _049937_, _049938_, _049939_, _049940_, _049941_, _049942_, _049943_, _049944_, _049945_, _049946_, _049947_, _049948_, _049949_, _049950_, _049951_, _049952_, _049953_, _049954_, _049955_, _049956_, _049957_, _049958_, _049959_, _049960_, _049961_, _049962_, _049963_, _049964_, _049965_, _049966_, _049967_, _049968_, _049969_, _049970_, _049971_, _049972_, _049973_, _049974_, _049975_, _049976_, _049977_, _049978_, _049979_, _049980_, _049981_, _049982_, _049983_, _049984_, _049985_, _049986_, _049987_, _049988_, _049989_, _049990_, _049991_, _049992_, _049993_, _049994_, _049995_, _049996_, _049997_, _049998_, _049999_, _050000_, _050001_, _050002_, _050003_, _050004_, _050005_, _050006_, _050007_, _050008_, _050009_, _050010_, _050011_, _050012_, _050013_, _050014_, _050015_, _050016_, _050017_, _050018_, _050019_, _050020_, _050021_, _050022_, _050023_, _050024_, _050025_, _050026_, _050027_, _050028_, _050029_, _050030_, _050031_, _050032_, _050033_, _050034_, _050035_, _050036_, _050037_, _050038_, _050039_, _050040_, _050041_, _050042_, _050043_, _050044_, _050045_, _050046_, _050047_, _050048_, _050049_, _050050_, _050051_, _050052_, _050053_, _050054_, _050055_, _050056_, _050057_, _050058_, _050059_, _050060_, _050061_, _050062_, _050063_, _050064_, _050065_, _050066_, _050067_, _050068_, _050069_, _050070_, _050071_, _050072_, _050073_, _050074_, _050075_, _050076_, _050077_, _050078_, _050079_, _050080_, _050081_, _050082_, _050083_, _050084_, _050085_, _050086_, _050087_, _050088_, _050089_, _050090_, _050091_, _050092_, _050093_, _050094_, _050095_, _050096_, _050097_, _050098_, _050099_, _050100_, _050101_, _050102_, _050103_, _050104_, _050105_, _050106_, _050107_, _050108_, _050109_, _050110_, _050111_, _050112_, _050113_, _050114_, _050115_, _050116_, _050117_, _050118_, _050119_, _050120_, _050121_, _050122_, _050123_, _050124_, _050125_, _050126_, _050127_, _050128_, _050129_, _050130_, _050131_, _050132_, _050133_, _050134_, _050135_, _050136_, _050137_, _050138_, _050139_, _050140_, _050141_, _050142_, _050143_, _050144_, _050145_, _050146_, _050147_, _050148_, _050149_, _050150_, _050151_, _050152_, _050153_, _050154_, _050155_, _050156_, _050157_, _050158_, _050159_, _050160_, _050161_, _050162_, _050163_, _050164_, _050165_, _050166_, _050167_, _050168_, _050169_, _050170_, _050171_, _050172_, _050173_, _050174_, _050175_, _050176_, _050177_, _050178_, _050179_, _050180_, _050181_, _050182_, _050183_, _050184_, _050185_, _050186_, _050187_, _050188_, _050189_, _050190_, _050191_, _050192_, _050193_, _050194_, _050195_, _050196_, _050197_, _050198_, _050199_, _050200_, _050201_, _050202_, _050203_, _050204_, _050205_, _050206_, _050207_, _050208_, _050209_, _050210_, _050211_, _050212_, _050213_, _050214_, _050215_, _050216_, _050217_, _050218_, _050219_, _050220_, _050221_, _050222_, _050223_, _050224_, _050225_, _050226_, _050227_, _050228_, _050229_, _050230_, _050231_, _050232_, _050233_, _050234_, _050235_, _050236_, _050237_, _050238_, _050239_, _050240_, _050241_, _050242_, _050243_, _050244_, _050245_, _050246_, _050247_, _050248_, _050249_, _050250_, _050251_, _050252_, _050253_, _050254_, _050255_, _050256_, _050257_, _050258_, _050259_, _050260_, _050261_, _050262_, _050263_, _050264_, _050265_, _050266_, _050267_, _050268_, _050269_, _050270_, _050271_, _050272_, _050273_, _050274_, _050275_, _050276_, _050277_, _050278_, _050279_, _050280_, _050281_, _050282_, _050283_, _050284_, _050285_, _050286_, _050287_, _050288_, _050289_, _050290_, _050291_, _050292_, _050293_, _050294_, _050295_, _050296_, _050297_, _050298_, _050299_, _050300_, _050301_, _050302_, _050303_, _050304_, _050305_, _050306_, _050307_, _050308_, _050309_, _050310_, _050311_, _050312_, _050313_, _050314_, _050315_, _050316_, _050317_, _050318_, _050319_, _050320_, _050321_, _050322_, _050323_, _050324_, _050325_, _050326_, _050327_, _050328_, _050329_, _050330_, _050331_, _050332_, _050333_, _050334_, _050335_, _050336_, _050337_, _050338_, _050339_, _050340_, _050341_, _050342_, _050343_, _050344_, _050345_, _050346_, _050347_, _050348_, _050349_, _050350_, _050351_, _050352_, _050353_, _050354_, _050355_, _050356_, _050357_, _050358_, _050359_, _050360_, _050361_, _050362_, _050363_, _050364_, _050365_, _050366_, _050367_, _050368_, _050369_, _050370_, _050371_, _050372_, _050373_, _050374_, _050375_, _050376_, _050377_, _050378_, _050379_, _050380_, _050381_, _050382_, _050383_, _050384_, _050385_, _050386_, _050387_, _050388_, _050389_, _050390_, _050391_, _050392_, _050393_, _050394_, _050395_, _050396_, _050397_, _050398_, _050399_, _050400_, _050401_, _050402_, _050403_, _050404_, _050405_, _050406_, _050407_, _050408_, _050409_, _050410_, _050411_, _050412_, _050413_, _050414_, _050415_, _050416_, _050417_, _050418_, _050419_, _050420_, _050421_, _050422_, _050423_, _050424_, _050425_, _050426_, _050427_, _050428_, _050429_, _050430_, _050431_, _050432_, _050433_, _050434_, _050435_, _050436_, _050437_, _050438_, _050439_, _050440_, _050441_, _050442_, _050443_, _050444_, _050445_, _050446_, _050447_, _050448_, _050449_, _050450_, _050451_, _050452_, _050453_, _050454_, _050455_, _050456_, _050457_, _050458_, _050459_, _050460_, _050461_, _050462_, _050463_, _050464_, _050465_, _050466_, _050467_, _050468_, _050469_, _050470_, _050471_, _050472_, _050473_, _050474_, _050475_, _050476_, _050477_, _050478_, _050479_, _050480_, _050481_, _050482_, _050483_, _050484_, _050485_, _050486_, _050487_, _050488_, _050489_, _050490_, _050491_, _050492_, _050493_, _050494_, _050495_, _050496_, _050497_, _050498_, _050499_, _050500_, _050501_, _050502_, _050503_, _050504_, _050505_, _050506_, _050507_, _050508_, _050509_, _050510_, _050511_, _050512_, _050513_, _050514_, _050515_, _050516_, _050517_, _050518_, _050519_, _050520_, _050521_, _050522_, _050523_, _050524_, _050525_, _050526_, _050527_, _050528_, _050529_, _050530_, _050531_, _050532_, _050533_, _050534_, _050535_, _050536_, _050537_, _050538_, _050539_, _050540_, _050541_, _050542_, _050543_, _050544_, _050545_, _050546_, _050547_, _050548_, _050549_, _050550_, _050551_, _050552_, _050553_, _050554_, _050555_, _050556_, _050557_, _050558_, _050559_, _050560_, _050561_, _050562_, _050563_, _050564_, _050565_, _050566_, _050567_, _050568_, _050569_, _050570_, _050571_, _050572_, _050573_, _050574_, _050575_, _050576_, _050577_, _050578_, _050579_, _050580_, _050581_, _050582_, _050583_, _050584_, _050585_, _050586_, _050587_, _050588_, _050589_, _050590_, _050591_, _050592_, _050593_, _050594_, _050595_, _050596_, _050597_, _050598_, _050599_, _050600_, _050601_, _050602_, _050603_, _050604_, _050605_, _050606_, _050607_, _050608_, _050609_, _050610_, _050611_, _050612_, _050613_, _050614_, _050615_, _050616_, _050617_, _050618_, _050619_, _050620_, _050621_, _050622_, _050623_, _050624_, _050625_, _050626_, _050627_, _050628_, _050629_, _050630_, _050631_, _050632_, _050633_, _050634_, _050635_, _050636_, _050637_, _050638_, _050639_, _050640_, _050641_, _050642_, _050643_, _050644_, _050645_, _050646_, _050647_, _050648_, _050649_, _050650_, _050651_, _050652_, _050653_, _050654_, _050655_, _050656_, _050657_, _050658_, _050659_, _050660_, _050661_, _050662_, _050663_, _050664_, _050665_, _050666_, _050667_, _050668_, _050669_, _050670_, _050671_, _050672_, _050673_, _050674_, _050675_, _050676_, _050677_, _050678_, _050679_, _050680_, _050681_, _050682_, _050683_, _050684_, _050685_, _050686_, _050687_, _050688_, _050689_, _050690_, _050691_, _050692_, _050693_, _050694_, _050695_, _050696_, _050697_, _050698_, _050699_, _050700_, _050701_, _050702_, _050703_, _050704_, _050705_, _050706_, _050707_, _050708_, _050709_, _050710_, _050711_, _050712_, _050713_, _050714_, _050715_, _050716_, _050717_, _050718_, _050719_, _050720_, _050721_, _050722_, _050723_, _050724_, _050725_, _050726_, _050727_, _050728_, _050729_, _050730_, _050731_, _050732_, _050733_, _050734_, _050735_, _050736_, _050737_, _050738_, _050739_, _050740_, _050741_, _050742_, _050743_, _050744_, _050745_, _050746_, _050747_, _050748_, _050749_, _050750_, _050751_, _050752_, _050753_, _050754_, _050755_, _050756_, _050757_, _050758_, _050759_, _050760_, _050761_, _050762_, _050763_, _050764_, _050765_, _050766_, _050767_, _050768_, _050769_, _050770_, _050771_, _050772_, _050773_, _050774_, _050775_, _050776_, _050777_, _050778_, _050779_, _050780_, _050781_, _050782_, _050783_, _050784_, _050785_, _050786_, _050787_, _050788_, _050789_, _050790_, _050791_, _050792_, _050793_, _050794_, _050795_, _050796_, _050797_, _050798_, _050799_, _050800_, _050801_, _050802_, _050803_, _050804_, _050805_, _050806_, _050807_, _050808_, _050809_, _050810_, _050811_, _050812_, _050813_, _050814_, _050815_, _050816_, _050817_, _050818_, _050819_, _050820_, _050821_, _050822_, _050823_, _050824_, _050825_, _050826_, _050827_, _050828_, _050829_, _050830_, _050831_, _050832_, _050833_, _050834_, _050835_, _050836_, _050837_, _050838_, _050839_, _050840_, _050841_, _050842_, _050843_, _050844_, _050845_, _050846_, _050847_, _050848_, _050849_, _050850_, _050851_, _050852_, _050853_, _050854_, _050855_, _050856_, _050857_, _050858_, _050859_, _050860_, _050861_, _050862_, _050863_, _050864_, _050865_, _050866_, _050867_, _050868_, _050869_, _050870_, _050871_, _050872_, _050873_, _050874_, _050875_, _050876_, _050877_, _050878_, _050879_, _050880_, _050881_, _050882_, _050883_, _050884_, _050885_, _050886_, _050887_, _050888_, _050889_, _050890_, _050891_, _050892_, _050893_, _050894_, _050895_, _050896_, _050897_, _050898_, _050899_, _050900_, _050901_, _050902_, _050903_, _050904_, _050905_, _050906_, _050907_, _050908_, _050909_, _050910_, _050911_, _050912_, _050913_, _050914_, _050915_, _050916_, _050917_, _050918_, _050919_, _050920_, _050921_, _050922_, _050923_, _050924_, _050925_, _050926_, _050927_, _050928_, _050929_, _050930_, _050931_, _050932_, _050933_, _050934_, _050935_, _050936_, _050937_, _050938_, _050939_, _050940_, _050941_, _050942_, _050943_, _050944_, _050945_, _050946_, _050947_, _050948_, _050949_, _050950_, _050951_, _050952_, _050953_, _050954_, _050955_, _050956_, _050957_, _050958_, _050959_, _050960_, _050961_, _050962_, _050963_, _050964_, _050965_, _050966_, _050967_, _050968_, _050969_, _050970_, _050971_, _050972_, _050973_, _050974_, _050975_, _050976_, _050977_, _050978_, _050979_, _050980_, _050981_, _050982_, _050983_, _050984_, _050985_, _050986_, _050987_, _050988_, _050989_, _050990_, _050991_, _050992_, _050993_, _050994_, _050995_, _050996_, _050997_, _050998_, _050999_, _051000_, _051001_, _051002_, _051003_, _051004_, _051005_, _051006_, _051007_, _051008_, _051009_, _051010_, _051011_, _051012_, _051013_, _051014_, _051015_, _051016_, _051017_, _051018_, _051019_, _051020_, _051021_, _051022_, _051023_, _051024_, _051025_, _051026_, _051027_, _051028_, _051029_, _051030_, _051031_, _051032_, _051033_, _051034_, _051035_, _051036_, _051037_, _051038_, _051039_, _051040_, _051041_, _051042_, _051043_, _051044_, _051045_, _051046_, _051047_, _051048_, _051049_, _051050_, _051051_, _051052_, _051053_, _051054_, _051055_, _051056_, _051057_, _051058_, _051059_, _051060_, _051061_, _051062_, _051063_, _051064_, _051065_, _051066_, _051067_, _051068_, _051069_, _051070_, _051071_, _051072_, _051073_, _051074_, _051075_, _051076_, _051077_, _051078_, _051079_, _051080_, _051081_, _051082_, _051083_, _051084_, _051085_, _051086_, _051087_, _051088_, _051089_, _051090_, _051091_, _051092_, _051093_, _051094_, _051095_, _051096_, _051097_, _051098_, _051099_, _051100_, _051101_, _051102_, _051103_, _051104_, _051105_, _051106_, _051107_, _051108_, _051109_, _051110_, _051111_, _051112_, _051113_, _051114_, _051115_, _051116_, _051117_, _051118_, _051119_, _051120_, _051121_, _051122_, _051123_, _051124_, _051125_, _051126_, _051127_, _051128_, _051129_, _051130_, _051131_, _051132_, _051133_, _051134_, _051135_, _051136_, _051137_, _051138_, _051139_, _051140_, _051141_, _051142_, _051143_, _051144_, _051145_, _051146_, _051147_, _051148_, _051149_, _051150_, _051151_, _051152_, _051153_, _051154_, _051155_, _051156_, _051157_, _051158_, _051159_, _051160_, _051161_, _051162_, _051163_, _051164_, _051165_, _051166_, _051167_, _051168_, _051169_, _051170_, _051171_, _051172_, _051173_, _051174_, _051175_, _051176_, _051177_, _051178_, _051179_, _051180_, _051181_, _051182_, _051183_, _051184_, _051185_, _051186_, _051187_, _051188_, _051189_, _051190_, _051191_, _051192_, _051193_, _051194_, _051195_, _051196_, _051197_, _051198_, _051199_, _051200_, _051201_, _051202_, _051203_, _051204_, _051205_, _051206_, _051207_, _051208_, _051209_, _051210_, _051211_, _051212_, _051213_, _051214_, _051215_, _051216_, _051217_, _051218_, _051219_, _051220_, _051221_, _051222_, _051223_, _051224_, _051225_, _051226_, _051227_, _051228_, _051229_, _051230_, _051231_, _051232_, _051233_, _051234_, _051235_, _051236_, _051237_, _051238_, _051239_, _051240_, _051241_, _051242_, _051243_, _051244_, _051245_, _051246_, _051247_, _051248_, _051249_, _051250_, _051251_, _051252_, _051253_, _051254_, _051255_, _051256_, _051257_, _051258_, _051259_, _051260_, _051261_, _051262_, _051263_, _051264_, _051265_, _051266_, _051267_, _051268_, _051269_, _051270_, _051271_, _051272_, _051273_, _051274_, _051275_, _051276_, _051277_, _051278_, _051279_, _051280_, _051281_, _051282_, _051283_, _051284_, _051285_, _051286_, _051287_, _051288_, _051289_, _051290_, _051291_, _051292_, _051293_, _051294_, _051295_, _051296_, _051297_, _051298_, _051299_, _051300_, _051301_, _051302_, _051303_, _051304_, _051305_, _051306_, _051307_, _051308_, _051309_, _051310_, _051311_, _051312_, _051313_, _051314_, _051315_, _051316_, _051317_, _051318_, _051319_, _051320_, _051321_, _051322_, _051323_, _051324_, _051325_, _051326_, _051327_, _051328_, _051329_, _051330_, _051331_, _051332_, _051333_, _051334_, _051335_, _051336_, _051337_, _051338_, _051339_, _051340_, _051341_, _051342_, _051343_, _051344_, _051345_, _051346_, _051347_, _051348_, _051349_, _051350_, _051351_, _051352_, _051353_, _051354_, _051355_, _051356_, _051357_, _051358_, _051359_, _051360_, _051361_, _051362_, _051363_, _051364_, _051365_, _051366_, _051367_, _051368_, _051369_, _051370_, _051371_, _051372_, _051373_, _051374_, _051375_, _051376_, _051377_, _051378_, _051379_, _051380_, _051381_, _051382_, _051383_, _051384_, _051385_, _051386_, _051387_, _051388_, _051389_, _051390_, _051391_, _051392_, _051393_, _051394_, _051395_, _051396_, _051397_, _051398_, _051399_, _051400_, _051401_, _051402_, _051403_, _051404_, _051405_, _051406_, _051407_, _051408_, _051409_, _051410_, _051411_, _051412_, _051413_, _051414_, _051415_, _051416_, _051417_, _051418_, _051419_, _051420_, _051421_, _051422_, _051423_, _051424_, _051425_, _051426_, _051427_, _051428_, _051429_, _051430_, _051431_, _051432_, _051433_, _051434_, _051435_, _051436_, _051437_, _051438_, _051439_, _051440_, _051441_, _051442_, _051443_, _051444_, _051445_, _051446_, _051447_, _051448_, _051449_, _051450_, _051451_, _051452_, _051453_, _051454_, _051455_, _051456_, _051457_, _051458_, _051459_, _051460_, _051461_, _051462_, _051463_, _051464_, _051465_, _051466_, _051467_, _051468_, _051469_, _051470_, _051471_, _051472_, _051473_, _051474_, _051475_, _051476_, _051477_, _051478_, _051479_, _051480_, _051481_, _051482_, _051483_, _051484_, _051485_, _051486_, _051487_, _051488_, _051489_, _051490_, _051491_, _051492_, _051493_, _051494_, _051495_, _051496_, _051497_, _051498_, _051499_, _051500_, _051501_, _051502_, _051503_, _051504_, _051505_, _051506_, _051507_, _051508_, _051509_, _051510_, _051511_, _051512_, _051513_, _051514_, _051515_, _051516_, _051517_, _051518_, _051519_, _051520_, _051521_, _051522_, _051523_, _051524_, _051525_, _051526_, _051527_, _051528_, _051529_, _051530_, _051531_, _051532_, _051533_, _051534_, _051535_, _051536_, _051537_, _051538_, _051539_, _051540_, _051541_, _051542_, _051543_, _051544_, _051545_, _051546_, _051547_, _051548_, _051549_, _051550_, _051551_, _051552_, _051553_, _051554_, _051555_, _051556_, _051557_, _051558_, _051559_, _051560_, _051561_, _051562_, _051563_, _051564_, _051565_, _051566_, _051567_, _051568_, _051569_, _051570_, _051571_, _051572_, _051573_, _051574_, _051575_, _051576_, _051577_, _051578_, _051579_, _051580_, _051581_, _051582_, _051583_, _051584_, _051585_, _051586_, _051587_, _051588_, _051589_, _051590_, _051591_, _051592_, _051593_, _051594_, _051595_, _051596_, _051597_, _051598_, _051599_, _051600_, _051601_, _051602_, _051603_, _051604_, _051605_, _051606_, _051607_, _051608_, _051609_, _051610_, _051611_, _051612_, _051613_, _051614_, _051615_, _051616_, _051617_, _051618_, _051619_, _051620_, _051621_, _051622_, _051623_, _051624_, _051625_, _051626_, _051627_, _051628_, _051629_, _051630_, _051631_, _051632_, _051633_, _051634_, _051635_, _051636_, _051637_, _051638_, _051639_, _051640_, _051641_, _051642_, _051643_, _051644_, _051645_, _051646_, _051647_, _051648_, _051649_, _051650_, _051651_, _051652_, _051653_, _051654_, _051655_, _051656_, _051657_, _051658_, _051659_, _051660_, _051661_, _051662_, _051663_, _051664_, _051665_, _051666_, _051667_, _051668_, _051669_, _051670_, _051671_, _051672_, _051673_, _051674_, _051675_, _051676_, _051677_, _051678_, _051679_, _051680_, _051681_, _051682_, _051683_, _051684_, _051685_, _051686_, _051687_, _051688_, _051689_, _051690_, _051691_, _051692_, _051693_, _051694_, _051695_, _051696_, _051697_, _051698_, _051699_, _051700_, _051701_, _051702_, _051703_, _051704_, _051705_, _051706_, _051707_, _051708_, _051709_, _051710_, _051711_, _051712_, _051713_, _051714_, _051715_, _051716_, _051717_, _051718_, _051719_, _051720_, _051721_, _051722_, _051723_, _051724_, _051725_, _051726_, _051727_, _051728_, _051729_, _051730_, _051731_, _051732_, _051733_, _051734_, _051735_, _051736_, _051737_, _051738_, _051739_, _051740_, _051741_, _051742_, _051743_, _051744_, _051745_, _051746_, _051747_, _051748_, _051749_, _051750_, _051751_, _051752_, _051753_, _051754_, _051755_, _051756_, _051757_, _051758_, _051759_, _051760_, _051761_, _051762_, _051763_, _051764_, _051765_, _051766_, _051767_, _051768_, _051769_, _051770_, _051771_, _051772_, _051773_, _051774_, _051775_, _051776_, _051777_, _051778_, _051779_, _051780_, _051781_, _051782_, _051783_, _051784_, _051785_, _051786_, _051787_, _051788_, _051789_, _051790_, _051791_, _051792_, _051793_, _051794_, _051795_, _051796_, _051797_, _051798_, _051799_, _051800_, _051801_, _051802_, _051803_, _051804_, _051805_, _051806_, _051807_, _051808_, _051809_, _051810_, _051811_, _051812_, _051813_, _051814_, _051815_, _051816_, _051817_, _051818_, _051819_, _051820_, _051821_, _051822_, _051823_, _051824_, _051825_, _051826_, _051827_, _051828_, _051829_, _051830_, _051831_, _051832_, _051833_, _051834_, _051835_, _051836_, _051837_, _051838_, _051839_, _051840_, _051841_, _051842_, _051843_, _051844_, _051845_, _051846_, _051847_, _051848_, _051849_, _051850_, _051851_, _051852_, _051853_, _051854_, _051855_, _051856_, _051857_, _051858_, _051859_, _051860_, _051861_, _051862_, _051863_, _051864_, _051865_, _051866_, _051867_, _051868_, _051869_, _051870_, _051871_, _051872_, _051873_, _051874_, _051875_, _051876_, _051877_, _051878_, _051879_, _051880_, _051881_, _051882_, _051883_, _051884_, _051885_, _051886_, _051887_, _051888_, _051889_, _051890_, _051891_, _051892_, _051893_, _051894_, _051895_, _051896_, _051897_, _051898_, _051899_, _051900_, _051901_, _051902_, _051903_, _051904_, _051905_, _051906_, _051907_, _051908_, _051909_, _051910_, _051911_, _051912_, _051913_, _051914_, _051915_, _051916_, _051917_, _051918_, _051919_, _051920_, _051921_, _051922_, _051923_, _051924_, _051925_, _051926_, _051927_, _051928_, _051929_, _051930_, _051931_, _051932_, _051933_, _051934_, _051935_, _051936_, _051937_, _051938_, _051939_, _051940_, _051941_, _051942_, _051943_, _051944_, _051945_, _051946_, _051947_, _051948_, _051949_, _051950_, _051951_, _051952_, _051953_, _051954_, _051955_, _051956_, _051957_, _051958_, _051959_, _051960_, _051961_, _051962_, _051963_, _051964_, _051965_, _051966_, _051967_, _051968_, _051969_, _051970_, _051971_, _051972_, _051973_, _051974_, _051975_, _051976_, _051977_, _051978_, _051979_, _051980_, _051981_, _051982_, _051983_, _051984_, _051985_, _051986_, _051987_, _051988_, _051989_, _051990_, _051991_, _051992_, _051993_, _051994_, _051995_, _051996_, _051997_, _051998_, _051999_, _052000_, _052001_, _052002_, _052003_, _052004_, _052005_, _052006_, _052007_, _052008_, _052009_, _052010_, _052011_, _052012_, _052013_, _052014_, _052015_, _052016_, _052017_, _052018_, _052019_, _052020_, _052021_, _052022_, _052023_, _052024_, _052025_, _052026_, _052027_, _052028_, _052029_, _052030_, _052031_, _052032_, _052033_, _052034_, _052035_, _052036_, _052037_, _052038_, _052039_, _052040_, _052041_, _052042_, _052043_, _052044_, _052045_, _052046_, _052047_, _052048_, _052049_, _052050_, _052051_, _052052_, _052053_, _052054_, _052055_, _052056_, _052057_, _052058_, _052059_, _052060_, _052061_, _052062_, _052063_, _052064_, _052065_, _052066_, _052067_, _052068_, _052069_, _052070_, _052071_, _052072_, _052073_, _052074_, _052075_, _052076_, _052077_, _052078_, _052079_, _052080_, _052081_, _052082_, _052083_, _052084_, _052085_, _052086_, _052087_, _052088_, _052089_, _052090_, _052091_, _052092_, _052093_, _052094_, _052095_, _052096_, _052097_, _052098_, _052099_, _052100_, _052101_, _052102_, _052103_, _052104_, _052105_, _052106_, _052107_, _052108_, _052109_, _052110_, _052111_, _052112_, _052113_, _052114_, _052115_, _052116_, _052117_, _052118_, _052119_, _052120_, _052121_, _052122_, _052123_, _052124_, _052125_, _052126_, _052127_, _052128_, _052129_, _052130_, _052131_, _052132_, _052133_, _052134_, _052135_, _052136_, _052137_, _052138_, _052139_, _052140_, _052141_, _052142_, _052143_, _052144_, _052145_, _052146_, _052147_, _052148_, _052149_, _052150_, _052151_, _052152_, _052153_, _052154_, _052155_, _052156_, _052157_, _052158_, _052159_, _052160_, _052161_, _052162_, _052163_, _052164_, _052165_, _052166_, _052167_, _052168_, _052169_, _052170_, _052171_, _052172_, _052173_, _052174_, _052175_, _052176_, _052177_, _052178_, _052179_, _052180_, _052181_, _052182_, _052183_, _052184_, _052185_, _052186_, _052187_, _052188_, _052189_, _052190_, _052191_, _052192_, _052193_, _052194_, _052195_, _052196_, _052197_, _052198_, _052199_, _052200_, _052201_, _052202_, _052203_, _052204_, _052205_, _052206_, _052207_, _052208_, _052209_, _052210_, _052211_, _052212_, _052213_, _052214_, _052215_, _052216_, _052217_, _052218_, _052219_, _052220_, _052221_, _052222_, _052223_, _052224_, _052225_, _052226_, _052227_, _052228_, _052229_, _052230_, _052231_, _052232_, _052233_, _052234_, _052235_, _052236_, _052237_, _052238_, _052239_, _052240_, _052241_, _052242_, _052243_, _052244_, _052245_, _052246_, _052247_, _052248_, _052249_, _052250_, _052251_, _052252_, _052253_, _052254_, _052255_, _052256_, _052257_, _052258_, _052259_, _052260_, _052261_, _052262_, _052263_, _052264_, _052265_, _052266_, _052267_, _052268_, _052269_, _052270_, _052271_, _052272_, _052273_, _052274_, _052275_, _052276_, _052277_, _052278_, _052279_, _052280_, _052281_, _052282_, _052283_, _052284_, _052285_, _052286_, _052287_, _052288_, _052289_, _052290_, _052291_, _052292_, _052293_, _052294_, _052295_, _052296_, _052297_, _052298_, _052299_, _052300_, _052301_, _052302_, _052303_, _052304_, _052305_, _052306_, _052307_, _052308_, _052309_, _052310_, _052311_, _052312_, _052313_, _052314_, _052315_, _052316_, _052317_, _052318_, _052319_, _052320_, _052321_, _052322_, _052323_, _052324_, _052325_, _052326_, _052327_, _052328_, _052329_, _052330_, _052331_, _052332_, _052333_, _052334_, _052335_, _052336_, _052337_, _052338_, _052339_, _052340_, _052341_, _052342_, _052343_, _052344_, _052345_, _052346_, _052347_, _052348_, _052349_, _052350_, _052351_, _052352_, _052353_, _052354_, _052355_, _052356_, _052357_, _052358_, _052359_, _052360_, _052361_, _052362_, _052363_, _052364_, _052365_, _052366_, _052367_, _052368_, _052369_, _052370_, _052371_, _052372_, _052373_, _052374_, _052375_, _052376_, _052377_, _052378_, _052379_, _052380_, _052381_, _052382_, _052383_, _052384_, _052385_, _052386_, _052387_, _052388_, _052389_, _052390_, _052391_, _052392_, _052393_, _052394_, _052395_, _052396_, _052397_, _052398_, _052399_, _052400_, _052401_, _052402_, _052403_, _052404_, _052405_, _052406_, _052407_, _052408_, _052409_, _052410_, _052411_, _052412_, _052413_, _052414_, _052415_, _052416_, _052417_, _052418_, _052419_, _052420_, _052421_, _052422_, _052423_, _052424_, _052425_, _052426_, _052427_, _052428_, _052429_, _052430_, _052431_, _052432_, _052433_, _052434_, _052435_, _052436_, _052437_, _052438_, _052439_, _052440_, _052441_, _052442_, _052443_, _052444_, _052445_, _052446_, _052447_, _052448_, _052449_, _052450_, _052451_, _052452_, _052453_, _052454_, _052455_, _052456_, _052457_, _052458_, _052459_, _052460_, _052461_, _052462_, _052463_, _052464_, _052465_, _052466_, _052467_, _052468_, _052469_, _052470_, _052471_, _052472_, _052473_, _052474_, _052475_, _052476_, _052477_, _052478_, _052479_, _052480_, _052481_, _052482_, _052483_, _052484_, _052485_, _052486_, _052487_, _052488_, _052489_, _052490_, _052491_, _052492_, _052493_, _052494_, _052495_, _052496_, _052497_, _052498_, _052499_, _052500_, _052501_, _052502_, _052503_, _052504_, _052505_, _052506_, _052507_, _052508_, _052509_, _052510_, _052511_, _052512_, _052513_, _052514_, _052515_, _052516_, _052517_, _052518_, _052519_, _052520_, _052521_, _052522_, _052523_, _052524_, _052525_, _052526_, _052527_, _052528_, _052529_, _052530_, _052531_, _052532_, _052533_, _052534_, _052535_, _052536_, _052537_, _052538_, _052539_, _052540_, _052541_, _052542_, _052543_, _052544_, _052545_, _052546_, _052547_, _052548_, _052549_, _052550_, _052551_, _052552_, _052553_, _052554_, _052555_, _052556_, _052557_, _052558_, _052559_, _052560_, _052561_, _052562_, _052563_, _052564_, _052565_, _052566_, _052567_, _052568_, _052569_, _052570_, _052571_, _052572_, _052573_, _052574_, _052575_, _052576_, _052577_, _052578_, _052579_, _052580_, _052581_, _052582_, _052583_, _052584_, _052585_, _052586_, _052587_, _052588_, _052589_, _052590_, _052591_, _052592_, _052593_, _052594_, _052595_, _052596_, _052597_, _052598_, _052599_, _052600_, _052601_, _052602_, _052603_, _052604_, _052605_, _052606_, _052607_, _052608_, _052609_, _052610_, _052611_, _052612_, _052613_, _052614_, _052615_, _052616_, _052617_, _052618_, _052619_, _052620_, _052621_, _052622_, _052623_, _052624_, _052625_, _052626_, _052627_, _052628_, _052629_, _052630_, _052631_, _052632_, _052633_, _052634_, _052635_, _052636_, _052637_, _052638_, _052639_, _052640_, _052641_, _052642_, _052643_, _052644_, _052645_, _052646_, _052647_, _052648_, _052649_, _052650_, _052651_, _052652_, _052653_, _052654_, _052655_, _052656_, _052657_, _052658_, _052659_, _052660_, _052661_, _052662_, _052663_, _052664_, _052665_, _052666_, _052667_, _052668_, _052669_, _052670_, _052671_, _052672_, _052673_, _052674_, _052675_, _052676_, _052677_, _052678_, _052679_, _052680_, _052681_, _052682_, _052683_, _052684_, _052685_, _052686_, _052687_, _052688_, _052689_, _052690_, _052691_, _052692_, _052693_, _052694_, _052695_, _052696_, _052697_, _052698_, _052699_, _052700_, _052701_, _052702_, _052703_, _052704_, _052705_, _052706_, _052707_, _052708_, _052709_, _052710_, _052711_, _052712_, _052713_, _052714_, _052715_, _052716_, _052717_, _052718_, _052719_, _052720_, _052721_, _052722_, _052723_, _052724_, _052725_, _052726_, _052727_, _052728_, _052729_, _052730_, _052731_, _052732_, _052733_, _052734_, _052735_, _052736_, _052737_, _052738_, _052739_, _052740_, _052741_, _052742_, _052743_, _052744_, _052745_, _052746_, _052747_, _052748_, _052749_, _052750_, _052751_, _052752_, _052753_, _052754_, _052755_, _052756_, _052757_, _052758_, _052759_, _052760_, _052761_, _052762_, _052763_, _052764_, _052765_, _052766_, _052767_, _052768_, _052769_, _052770_, _052771_, _052772_, _052773_, _052774_, _052775_, _052776_, _052777_, _052778_, _052779_, _052780_, _052781_, _052782_, _052783_, _052784_, _052785_, _052786_, _052787_, _052788_, _052789_, _052790_, _052791_, _052792_, _052793_, _052794_, _052795_, _052796_, _052797_, _052798_, _052799_, _052800_, _052801_, _052802_, _052803_, _052804_, _052805_, _052806_, _052807_, _052808_, _052809_, _052810_, _052811_, _052812_, _052813_, _052814_, _052815_, _052816_, _052817_, _052818_, _052819_, _052820_, _052821_, _052822_, _052823_, _052824_, _052825_, _052826_, _052827_, _052828_, _052829_, _052830_, _052831_, _052832_, _052833_, _052834_, _052835_, _052836_, _052837_, _052838_, _052839_, _052840_, _052841_, _052842_, _052843_, _052844_, _052845_, _052846_, _052847_, _052848_, _052849_, _052850_, _052851_, _052852_, _052853_, _052854_, _052855_, _052856_, _052857_, _052858_, _052859_, _052860_, _052861_, _052862_, _052863_, _052864_, _052865_, _052866_, _052867_, _052868_, _052869_, _052870_, _052871_, _052872_, _052873_, _052874_, _052875_, _052876_, _052877_, _052878_, _052879_, _052880_, _052881_, _052882_, _052883_, _052884_, _052885_, _052886_, _052887_, _052888_, _052889_, _052890_, _052891_, _052892_, _052893_, _052894_, _052895_, _052896_, _052897_, _052898_, _052899_, _052900_, _052901_, _052902_, _052903_, _052904_, _052905_, _052906_, _052907_, _052908_, _052909_, _052910_, _052911_, _052912_, _052913_, _052914_, _052915_, _052916_, _052917_, _052918_, _052919_, _052920_, _052921_, _052922_, _052923_, _052924_, _052925_, _052926_, _052927_, _052928_, _052929_, _052930_, _052931_, _052932_, _052933_, _052934_, _052935_, _052936_, _052937_, _052938_, _052939_, _052940_, _052941_, _052942_, _052943_, _052944_, _052945_, _052946_, _052947_, _052948_, _052949_, _052950_, _052951_, _052952_, _052953_, _052954_, _052955_, _052956_, _052957_, _052958_, _052959_, _052960_, _052961_, _052962_, _052963_, _052964_, _052965_, _052966_, _052967_, _052968_, _052969_, _052970_, _052971_, _052972_, _052973_, _052974_, _052975_, _052976_, _052977_, _052978_, _052979_, _052980_, _052981_, _052982_, _052983_, _052984_, _052985_, _052986_, _052987_, _052988_, _052989_, _052990_, _052991_, _052992_, _052993_, _052994_, _052995_, _052996_, _052997_, _052998_, _052999_, _053000_, _053001_, _053002_, _053003_, _053004_, _053005_, _053006_, _053007_, _053008_, _053009_, _053010_, _053011_, _053012_, _053013_, _053014_, _053015_, _053016_, _053017_, _053018_, _053019_, _053020_, _053021_, _053022_, _053023_, _053024_, _053025_, _053026_, _053027_, _053028_, _053029_, _053030_, _053031_, _053032_, _053033_, _053034_, _053035_, _053036_, _053037_, _053038_, _053039_, _053040_, _053041_, _053042_, _053043_, _053044_, _053045_, _053046_, _053047_, _053048_, _053049_, _053050_, _053051_, _053052_, _053053_, _053054_, _053055_, _053056_, _053057_, _053058_, _053059_, _053060_, _053061_, _053062_, _053063_, _053064_, _053065_, _053066_, _053067_, _053068_, _053069_, _053070_, _053071_, _053072_, _053073_, _053074_, _053075_, _053076_, _053077_, _053078_, _053079_, _053080_, _053081_, _053082_, _053083_, _053084_, _053085_, _053086_, _053087_, _053088_, _053089_, _053090_, _053091_, _053092_, _053093_, _053094_, _053095_, _053096_, _053097_, _053098_, _053099_, _053100_, _053101_, _053102_, _053103_, _053104_, _053105_, _053106_, _053107_, _053108_, _053109_, _053110_, _053111_, _053112_, _053113_, _053114_, _053115_, _053116_, _053117_, _053118_, _053119_, _053120_, _053121_, _053122_, _053123_, _053124_, _053125_, _053126_, _053127_, _053128_, _053129_, _053130_, _053131_, _053132_, _053133_, _053134_, _053135_, _053136_, _053137_, _053138_, _053139_, _053140_, _053141_, _053142_, _053143_, _053144_, _053145_, _053146_, _053147_, _053148_, _053149_, _053150_, _053151_, _053152_, _053153_, _053154_, _053155_, _053156_, _053157_, _053158_, _053159_, _053160_, _053161_, _053162_, _053163_, _053164_, _053165_, _053166_, _053167_, _053168_, _053169_, _053170_, _053171_, _053172_, _053173_, _053174_, _053175_, _053176_, _053177_, _053178_, _053179_, _053180_, _053181_, _053182_, _053183_, _053184_, _053185_, _053186_, _053187_, _053188_, _053189_, _053190_, _053191_, _053192_, _053193_, _053194_, _053195_, _053196_, _053197_, _053198_, _053199_, _053200_, _053201_, _053202_, _053203_, _053204_, _053205_, _053206_, _053207_, _053208_, _053209_, _053210_, _053211_, _053212_, _053213_, _053214_, _053215_, _053216_, _053217_, _053218_, _053219_, _053220_, _053221_, _053222_, _053223_, _053224_, _053225_, _053226_, _053227_, _053228_, _053229_, _053230_, _053231_, _053232_, _053233_, _053234_, _053235_, _053236_, _053237_, _053238_, _053239_, _053240_, _053241_, _053242_, _053243_, _053244_, _053245_, _053246_, _053247_, _053248_, _053249_, _053250_, _053251_, _053252_, _053253_, _053254_, _053255_, _053256_, _053257_, _053258_, _053259_, _053260_, _053261_, _053262_, _053263_, _053264_, _053265_, _053266_, _053267_, _053268_, _053269_, _053270_, _053271_, _053272_, _053273_, _053274_, _053275_, _053276_, _053277_, _053278_, _053279_, _053280_, _053281_, _053282_, _053283_, _053284_, _053285_, _053286_, _053287_, _053288_, _053289_, _053290_, _053291_, _053292_, _053293_, _053294_, _053295_, _053296_, _053297_, _053298_, _053299_, _053300_, _053301_, _053302_, _053303_, _053304_, _053305_, _053306_, _053307_, _053308_, _053309_, _053310_, _053311_, _053312_, _053313_, _053314_, _053315_, _053316_, _053317_, _053318_, _053319_, _053320_, _053321_, _053322_, _053323_, _053324_, _053325_, _053326_, _053327_, _053328_, _053329_, _053330_, _053331_, _053332_, _053333_, _053334_, _053335_, _053336_, _053337_, _053338_, _053339_, _053340_, _053341_, _053342_, _053343_, _053344_, _053345_, _053346_, _053347_, _053348_, _053349_, _053350_, _053351_, _053352_, _053353_, _053354_, _053355_, _053356_, _053357_, _053358_, _053359_, _053360_, _053361_, _053362_, _053363_, _053364_, _053365_, _053366_, _053367_, _053368_, _053369_, _053370_, _053371_, _053372_, _053373_, _053374_, _053375_, _053376_, _053377_, _053378_, _053379_, _053380_, _053381_, _053382_, _053383_, _053384_, _053385_, _053386_, _053387_, _053388_, _053389_, _053390_, _053391_, _053392_, _053393_, _053394_, _053395_, _053396_, _053397_, _053398_, _053399_, _053400_, _053401_, _053402_, _053403_, _053404_, _053405_, _053406_, _053407_, _053408_, _053409_, _053410_, _053411_, _053412_, _053413_, _053414_, _053415_, _053416_, _053417_, _053418_, _053419_, _053420_, _053421_, _053422_, _053423_, _053424_, _053425_, _053426_, _053427_, _053428_, _053429_, _053430_, _053431_, _053432_, _053433_, _053434_, _053435_, _053436_, _053437_, _053438_, _053439_, _053440_, _053441_, _053442_, _053443_, _053444_, _053445_, _053446_, _053447_, _053448_, _053449_, _053450_, _053451_, _053452_, _053453_, _053454_, _053455_, _053456_, _053457_, _053458_, _053459_, _053460_, _053461_, _053462_, _053463_, _053464_, _053465_, _053466_, _053467_, _053468_, _053469_, _053470_, _053471_, _053472_, _053473_, _053474_, _053475_, _053476_, _053477_, _053478_, _053479_, _053480_, _053481_, _053482_, _053483_, _053484_, _053485_, _053486_, _053487_, _053488_, _053489_, _053490_, _053491_, _053492_, _053493_, _053494_, _053495_, _053496_, _053497_, _053498_, _053499_, _053500_, _053501_, _053502_, _053503_, _053504_, _053505_, _053506_, _053507_, _053508_, _053509_, _053510_, _053511_, _053512_, _053513_, _053514_, _053515_, _053516_, _053517_, _053518_, _053519_, _053520_, _053521_, _053522_, _053523_, _053524_, _053525_, _053526_, _053527_, _053528_, _053529_, _053530_, _053531_, _053532_, _053533_, _053534_, _053535_, _053536_, _053537_, _053538_, _053539_, _053540_, _053541_, _053542_, _053543_, _053544_, _053545_, _053546_, _053547_, _053548_, _053549_, _053550_, _053551_, _053552_, _053553_, _053554_, _053555_, _053556_, _053557_, _053558_, _053559_, _053560_, _053561_, _053562_, _053563_, _053564_, _053565_, _053566_, _053567_, _053568_, _053569_, _053570_, _053571_, _053572_, _053573_, _053574_, _053575_, _053576_, _053577_, _053578_, _053579_, _053580_, _053581_, _053582_, _053583_, _053584_, _053585_, _053586_, _053587_, _053588_, _053589_, _053590_, _053591_, _053592_, _053593_, _053594_, _053595_, _053596_, _053597_, _053598_, _053599_, _053600_, _053601_, _053602_, _053603_, _053604_, _053605_, _053606_, _053607_, _053608_, _053609_, _053610_, _053611_, _053612_, _053613_, _053614_, _053615_, _053616_, _053617_, _053618_, _053619_, _053620_, _053621_, _053622_, _053623_, _053624_, _053625_, _053626_, _053627_, _053628_, _053629_, _053630_, _053631_, _053632_, _053633_, _053634_, _053635_, _053636_, _053637_, _053638_, _053639_, _053640_, _053641_, _053642_, _053643_, _053644_, _053645_, _053646_, _053647_, _053648_, _053649_, _053650_, _053651_, _053652_, _053653_, _053654_, _053655_, _053656_, _053657_, _053658_, _053659_, _053660_, _053661_, _053662_, _053663_, _053664_, _053665_, _053666_, _053667_, _053668_, _053669_, _053670_, _053671_, _053672_, _053673_, _053674_, _053675_, _053676_, _053677_, _053678_, _053679_, _053680_, _053681_, _053682_, _053683_, _053684_, _053685_, _053686_, _053687_, _053688_, _053689_, _053690_, _053691_, _053692_, _053693_, _053694_, _053695_, _053696_, _053697_, _053698_, _053699_, _053700_, _053701_, _053702_, _053703_, _053704_, _053705_, _053706_, _053707_, _053708_, _053709_, _053710_, _053711_, _053712_, _053713_, _053714_, _053715_, _053716_, _053717_, _053718_, _053719_, _053720_, _053721_, _053722_, _053723_, _053724_, _053725_, _053726_, _053727_, _053728_, _053729_, _053730_, _053731_, _053732_, _053733_, _053734_, _053735_, _053736_, _053737_, _053738_, _053739_, _053740_, _053741_, _053742_, _053743_, _053744_, _053745_, _053746_, _053747_, _053748_, _053749_, _053750_, _053751_, _053752_, _053753_, _053754_, _053755_, _053756_, _053757_, _053758_, _053759_, _053760_, _053761_, _053762_, _053763_, _053764_, _053765_, _053766_, _053767_, _053768_, _053769_, _053770_, _053771_, _053772_, _053773_, _053774_, _053775_, _053776_, _053777_, _053778_, _053779_, _053780_, _053781_, _053782_, _053783_, _053784_, _053785_, _053786_, _053787_, _053788_, _053789_, _053790_, _053791_, _053792_, _053793_, _053794_, _053795_, _053796_, _053797_, _053798_, _053799_, _053800_, _053801_, _053802_, _053803_, _053804_, _053805_, _053806_, _053807_, _053808_, _053809_, _053810_, _053811_, _053812_, _053813_, _053814_, _053815_, _053816_, _053817_, _053818_, _053819_, _053820_, _053821_, _053822_, _053823_, _053824_, _053825_, _053826_, _053827_, _053828_, _053829_, _053830_, _053831_, _053832_, _053833_, _053834_, _053835_, _053836_, _053837_, _053838_, _053839_, _053840_, _053841_, _053842_, _053843_, _053844_, _053845_, _053846_, _053847_, _053848_, _053849_, _053850_, _053851_, _053852_, _053853_, _053854_, _053855_, _053856_, _053857_, _053858_, _053859_, _053860_, _053861_, _053862_, _053863_, _053864_, _053865_, _053866_, _053867_, _053868_, _053869_, _053870_, _053871_, _053872_, _053873_, _053874_, _053875_, _053876_, _053877_, _053878_, _053879_, _053880_, _053881_, _053882_, _053883_, _053884_, _053885_, _053886_, _053887_, _053888_, _053889_, _053890_, _053891_, _053892_, _053893_, _053894_, _053895_, _053896_, _053897_, _053898_, _053899_, _053900_, _053901_, _053902_, _053903_, _053904_, _053905_, _053906_, _053907_, _053908_, _053909_, _053910_, _053911_, _053912_, _053913_, _053914_, _053915_, _053916_, _053917_, _053918_, _053919_, _053920_, _053921_, _053922_, _053923_, _053924_, _053925_, _053926_, _053927_, _053928_, _053929_, _053930_, _053931_, _053932_, _053933_, _053934_, _053935_, _053936_, _053937_, _053938_, _053939_, _053940_, _053941_, _053942_, _053943_, _053944_, _053945_, _053946_, _053947_, _053948_, _053949_, _053950_, _053951_, _053952_, _053953_, _053954_, _053955_, _053956_, _053957_, _053958_, _053959_, _053960_, _053961_, _053962_, _053963_, _053964_, _053965_, _053966_, _053967_, _053968_, _053969_, _053970_, _053971_, _053972_, _053973_, _053974_, _053975_, _053976_, _053977_, _053978_, _053979_, _053980_, _053981_, _053982_, _053983_, _053984_, _053985_, _053986_, _053987_, _053988_, _053989_, _053990_, _053991_, _053992_, _053993_, _053994_, _053995_, _053996_, _053997_, _053998_, _053999_, _054000_, _054001_, _054002_, _054003_, _054004_, _054005_, _054006_, _054007_, _054008_, _054009_, _054010_, _054011_, _054012_, _054013_, _054014_, _054015_, _054016_, _054017_, _054018_, _054019_, _054020_, _054021_, _054022_, _054023_, _054024_, _054025_, _054026_, _054027_, _054028_, _054029_, _054030_, _054031_, _054032_, _054033_, _054034_, _054035_, _054036_, _054037_, _054038_, _054039_, _054040_, _054041_, _054042_, _054043_, _054044_, _054045_, _054046_, _054047_, _054048_, _054049_, _054050_, _054051_, _054052_, _054053_, _054054_, _054055_, _054056_, _054057_, _054058_, _054059_, _054060_, _054061_, _054062_, _054063_, _054064_, _054065_, _054066_, _054067_, _054068_, _054069_, _054070_, _054071_, _054072_, _054073_, _054074_, _054075_, _054076_, _054077_, _054078_, _054079_, _054080_, _054081_, _054082_, _054083_, _054084_, _054085_, _054086_, _054087_, _054088_, _054089_, _054090_, _054091_, _054092_, _054093_, _054094_, _054095_, _054096_, _054097_, _054098_, _054099_, _054100_, _054101_, _054102_, _054103_, _054104_, _054105_, _054106_, _054107_, _054108_, _054109_, _054110_, _054111_, _054112_, _054113_, _054114_, _054115_, _054116_, _054117_, _054118_, _054119_, _054120_, _054121_, _054122_, _054123_, _054124_, _054125_, _054126_, _054127_, _054128_, _054129_, _054130_, _054131_, _054132_, _054133_, _054134_, _054135_, _054136_, _054137_, _054138_, _054139_, _054140_, _054141_, _054142_, _054143_, _054144_, _054145_, _054146_, _054147_, _054148_, _054149_, _054150_, _054151_, _054152_, _054153_, _054154_, _054155_, _054156_, _054157_, _054158_, _054159_, _054160_, _054161_, _054162_, _054163_, _054164_, _054165_, _054166_, _054167_, _054168_, _054169_, _054170_, _054171_, _054172_, _054173_, _054174_, _054175_, _054176_, _054177_, _054178_, _054179_, _054180_, _054181_, _054182_, _054183_, _054184_, _054185_, _054186_, _054187_, _054188_, _054189_, _054190_, _054191_, _054192_, _054193_, _054194_, _054195_, _054196_, _054197_, _054198_, _054199_, _054200_, _054201_, _054202_, _054203_, _054204_, _054205_, _054206_, _054207_, _054208_, _054209_, _054210_, _054211_, _054212_, _054213_, _054214_, _054215_, _054216_, _054217_, _054218_, _054219_, _054220_, _054221_, _054222_, _054223_, _054224_, _054225_, _054226_, _054227_, _054228_, _054229_, _054230_, _054231_, _054232_, _054233_, _054234_, _054235_, _054236_, _054237_, _054238_, _054239_, _054240_, _054241_, _054242_, _054243_, _054244_, _054245_, _054246_, _054247_, _054248_, _054249_, _054250_, _054251_, _054252_, _054253_, _054254_, _054255_, _054256_, _054257_, _054258_, _054259_, _054260_, _054261_, _054262_, _054263_, _054264_, _054265_, _054266_, _054267_, _054268_, _054269_, _054270_, _054271_, _054272_, _054273_, _054274_, _054275_, _054276_, _054277_, _054278_, _054279_, _054280_, _054281_, _054282_, _054283_, _054284_, _054285_, _054286_, _054287_, _054288_, _054289_, _054290_, _054291_, _054292_, _054293_, _054294_, _054295_, _054296_, _054297_, _054298_, _054299_, _054300_, _054301_, _054302_, _054303_, _054304_, _054305_, _054306_, _054307_, _054308_, _054309_, _054310_, _054311_, _054312_, _054313_, _054314_, _054315_, _054316_, _054317_, _054318_, _054319_, _054320_, _054321_, _054322_, _054323_, _054324_, _054325_, _054326_, _054327_, _054328_, _054329_, _054330_, _054331_, _054332_, _054333_, _054334_, _054335_, _054336_, _054337_, _054338_, _054339_, _054340_, _054341_, _054342_, _054343_, _054344_, _054345_, _054346_, _054347_, _054348_, _054349_, _054350_, _054351_, _054352_, _054353_, _054354_, _054355_, _054356_, _054357_, _054358_, _054359_, _054360_, _054361_, _054362_, _054363_, _054364_, _054365_, _054366_, _054367_, _054368_, _054369_, _054370_, _054371_, _054372_, _054373_, _054374_, _054375_, _054376_, _054377_, _054378_, _054379_, _054380_, _054381_, _054382_, _054383_, _054384_, _054385_, _054386_, _054387_, _054388_, _054389_, _054390_, _054391_, _054392_, _054393_, _054394_, _054395_, _054396_, _054397_, _054398_, _054399_, _054400_, _054401_, _054402_, _054403_, _054404_, _054405_, _054406_, _054407_, _054408_, _054409_, _054410_, _054411_, _054412_, _054413_, _054414_, _054415_, _054416_, _054417_, _054418_, _054419_, _054420_, _054421_, _054422_, _054423_, _054424_, _054425_, _054426_, _054427_, _054428_, _054429_, _054430_, _054431_, _054432_, _054433_, _054434_, _054435_, _054436_, _054437_, _054438_, _054439_, _054440_, _054441_, _054442_, _054443_, _054444_, _054445_, _054446_, _054447_, _054448_, _054449_, _054450_, _054451_, _054452_, _054453_, _054454_, _054455_, _054456_, _054457_, _054458_, _054459_, _054460_, _054461_, _054462_, _054463_, _054464_, _054465_, _054466_, _054467_, _054468_, _054469_, _054470_, _054471_, _054472_, _054473_, _054474_, _054475_, _054476_, _054477_, _054478_, _054479_, _054480_, _054481_, _054482_, _054483_, _054484_, _054485_, _054486_, _054487_, _054488_, _054489_, _054490_, _054491_, _054492_, _054493_, _054494_, _054495_, _054496_, _054497_, _054498_, _054499_, _054500_, _054501_, _054502_, _054503_, _054504_, _054505_, _054506_, _054507_, _054508_, _054509_, _054510_, _054511_, _054512_, _054513_, _054514_, _054515_, _054516_, _054517_, _054518_, _054519_, _054520_, _054521_, _054522_, _054523_, _054524_, _054525_, _054526_, _054527_, _054528_, _054529_, _054530_, _054531_, _054532_, _054533_, _054534_, _054535_, _054536_, _054537_, _054538_, _054539_, _054540_, _054541_, _054542_, _054543_, _054544_, _054545_, _054546_, _054547_, _054548_, _054549_, _054550_, _054551_, _054552_, _054553_, _054554_, _054555_, _054556_, _054557_, _054558_, _054559_, _054560_, _054561_, _054562_, _054563_, _054564_, _054565_, _054566_, _054567_, _054568_, _054569_, _054570_, _054571_, _054572_, _054573_, _054574_, _054575_, _054576_, _054577_, _054578_, _054579_, _054580_, _054581_, _054582_, _054583_, _054584_, _054585_, _054586_, _054587_, _054588_, _054589_, _054590_, _054591_, _054592_, _054593_, _054594_, _054595_, _054596_, _054597_, _054598_, _054599_, _054600_, _054601_, _054602_, _054603_, _054604_, _054605_, _054606_, _054607_, _054608_, _054609_, _054610_, _054611_, _054612_, _054613_, _054614_, _054615_, _054616_, _054617_, _054618_, _054619_, _054620_, _054621_, _054622_, _054623_, _054624_, _054625_, _054626_, _054627_, _054628_, _054629_, _054630_, _054631_, _054632_, _054633_, _054634_, _054635_, _054636_, _054637_, _054638_, _054639_, _054640_, _054641_, _054642_, _054643_, _054644_, _054645_, _054646_, _054647_, _054648_, _054649_, _054650_, _054651_, _054652_, _054653_, _054654_, _054655_, _054656_, _054657_, _054658_, _054659_, _054660_, _054661_, _054662_, _054663_, _054664_, _054665_, _054666_, _054667_, _054668_, _054669_, _054670_, _054671_, _054672_, _054673_, _054674_, _054675_, _054676_, _054677_, _054678_, _054679_, _054680_, _054681_, _054682_, _054683_, _054684_, _054685_, _054686_, _054687_, _054688_, _054689_, _054690_, _054691_, _054692_, _054693_, _054694_, _054695_, _054696_, _054697_, _054698_, _054699_, _054700_, _054701_, _054702_, _054703_, _054704_, _054705_, _054706_, _054707_, _054708_, _054709_, _054710_, _054711_, _054712_, _054713_, _054714_, _054715_, _054716_, _054717_, _054718_, _054719_, _054720_, _054721_, _054722_, _054723_, _054724_, _054725_, _054726_, _054727_, _054728_, _054729_, _054730_, _054731_, _054732_, _054733_, _054734_, _054735_, _054736_, _054737_, _054738_, _054739_, _054740_, _054741_, _054742_, _054743_, _054744_, _054745_, _054746_, _054747_, _054748_, _054749_, _054750_, _054751_, _054752_, _054753_, _054754_, _054755_, _054756_, _054757_, _054758_, _054759_, _054760_, _054761_, _054762_, _054763_, _054764_, _054765_, _054766_, _054767_, _054768_, _054769_, _054770_, _054771_, _054772_, _054773_, _054774_, _054775_, _054776_, _054777_, _054778_, _054779_, _054780_, _054781_, _054782_, _054783_, _054784_, _054785_, _054786_, _054787_, _054788_, _054789_, _054790_, _054791_, _054792_, _054793_, _054794_, _054795_, _054796_, _054797_, _054798_, _054799_, _054800_, _054801_, _054802_, _054803_, _054804_, _054805_, _054806_, _054807_, _054808_, _054809_, _054810_, _054811_, _054812_, _054813_, _054814_, _054815_, _054816_, _054817_, _054818_, _054819_, _054820_, _054821_, _054822_, _054823_, _054824_, _054825_, _054826_, _054827_, _054828_, _054829_, _054830_, _054831_, _054832_, _054833_, _054834_, _054835_, _054836_, _054837_, _054838_, _054839_, _054840_, _054841_, _054842_, _054843_, _054844_, _054845_, _054846_, _054847_, _054848_, _054849_, _054850_, _054851_, _054852_, _054853_, _054854_, _054855_, _054856_, _054857_, _054858_, _054859_, _054860_, _054861_, _054862_, _054863_, _054864_, _054865_, _054866_, _054867_, _054868_, _054869_, _054870_, _054871_, _054872_, _054873_, _054874_, _054875_, _054876_, _054877_, _054878_, _054879_, _054880_, _054881_, _054882_, _054883_, _054884_, _054885_, _054886_, _054887_, _054888_, _054889_, _054890_, _054891_, _054892_, _054893_, _054894_, _054895_, _054896_, _054897_, _054898_, _054899_, _054900_, _054901_, _054902_, _054903_, _054904_, _054905_, _054906_, _054907_, _054908_, _054909_, _054910_, _054911_, _054912_, _054913_, _054914_, _054915_, _054916_, _054917_, _054918_, _054919_, _054920_, _054921_, _054922_, _054923_, _054924_, _054925_, _054926_, _054927_, _054928_, _054929_, _054930_, _054931_, _054932_, _054933_, _054934_, _054935_, _054936_, _054937_, _054938_, _054939_, _054940_, _054941_, _054942_, _054943_, _054944_, _054945_, _054946_, _054947_, _054948_, _054949_, _054950_, _054951_, _054952_, _054953_, _054954_, _054955_, _054956_, _054957_, _054958_, _054959_, _054960_, _054961_, _054962_, _054963_, _054964_, _054965_, _054966_, _054967_, _054968_, _054969_, _054970_, _054971_, _054972_, _054973_, _054974_, _054975_, _054976_, _054977_, _054978_, _054979_, _054980_, _054981_, _054982_, _054983_, _054984_, _054985_, _054986_, _054987_, _054988_, _054989_, _054990_, _054991_, _054992_, _054993_, _054994_, _054995_, _054996_, _054997_, _054998_, _054999_, _055000_, _055001_, _055002_, _055003_, _055004_, _055005_, _055006_, _055007_, _055008_, _055009_, _055010_, _055011_, _055012_, _055013_, _055014_, _055015_, _055016_, _055017_, _055018_, _055019_, _055020_, _055021_, _055022_, _055023_, _055024_, _055025_, _055026_, _055027_, _055028_, _055029_, _055030_, _055031_, _055032_, _055033_, _055034_, _055035_, _055036_, _055037_, _055038_, _055039_, _055040_, _055041_, _055042_, _055043_, _055044_, _055045_, _055046_, _055047_, _055048_, _055049_, _055050_, _055051_, _055052_, _055053_, _055054_, _055055_, _055056_, _055057_, _055058_, _055059_, _055060_, _055061_, _055062_, _055063_, _055064_, _055065_, _055066_, _055067_, _055068_, _055069_, _055070_, _055071_, _055072_, _055073_, _055074_, _055075_, _055076_, _055077_, _055078_, _055079_, _055080_, _055081_, _055082_, _055083_, _055084_, _055085_, _055086_, _055087_, _055088_, _055089_, _055090_, _055091_, _055092_, _055093_, _055094_, _055095_, _055096_, _055097_, _055098_, _055099_, _055100_, _055101_, _055102_, _055103_, _055104_, _055105_, _055106_, _055107_, _055108_, _055109_, _055110_, _055111_, _055112_, _055113_, _055114_, _055115_, _055116_, _055117_, _055118_, _055119_, _055120_, _055121_, _055122_, _055123_, _055124_, _055125_, _055126_, _055127_, _055128_, _055129_, _055130_, _055131_, _055132_, _055133_, _055134_, _055135_, _055136_, _055137_, _055138_, _055139_, _055140_, _055141_, _055142_, _055143_, _055144_, _055145_, _055146_, _055147_, _055148_, _055149_, _055150_, _055151_, _055152_, _055153_, _055154_, _055155_, _055156_, _055157_, _055158_, _055159_, _055160_, _055161_, _055162_, _055163_, _055164_, _055165_, _055166_, _055167_, _055168_, _055169_, _055170_, _055171_, _055172_, _055173_, _055174_, _055175_, _055176_, _055177_, _055178_, _055179_, _055180_, _055181_, _055182_, _055183_, _055184_, _055185_, _055186_, _055187_, _055188_, _055189_, _055190_, _055191_, _055192_, _055193_, _055194_, _055195_, _055196_, _055197_, _055198_, _055199_, _055200_, _055201_, _055202_, _055203_, _055204_, _055205_, _055206_, _055207_, _055208_, _055209_, _055210_, _055211_, _055212_, _055213_, _055214_, _055215_, _055216_, _055217_, _055218_, _055219_, _055220_, _055221_, _055222_, _055223_, _055224_, _055225_, _055226_, _055227_, _055228_, _055229_, _055230_, _055231_, _055232_, _055233_, _055234_, _055235_, _055236_, _055237_, _055238_, _055239_, _055240_, _055241_, _055242_, _055243_, _055244_, _055245_, _055246_, _055247_, _055248_, _055249_, _055250_, _055251_, _055252_, _055253_, _055254_, _055255_, _055256_, _055257_, _055258_, _055259_, _055260_, _055261_, _055262_, _055263_, _055264_, _055265_, _055266_, _055267_, _055268_, _055269_, _055270_, _055271_, _055272_, _055273_, _055274_, _055275_, _055276_, _055277_, _055278_, _055279_, _055280_, _055281_, _055282_, _055283_, _055284_, _055285_, _055286_, _055287_, _055288_, _055289_, _055290_, _055291_, _055292_, _055293_, _055294_, _055295_, _055296_, _055297_, _055298_, _055299_, _055300_, _055301_, _055302_, _055303_, _055304_, _055305_, _055306_, _055307_, _055308_, _055309_, _055310_, _055311_, _055312_, _055313_, _055314_, _055315_, _055316_, _055317_, _055318_, _055319_, _055320_, _055321_, _055322_, _055323_, _055324_, _055325_, _055326_, _055327_, _055328_, _055329_, _055330_, _055331_, _055332_, _055333_, _055334_, _055335_, _055336_, _055337_, _055338_, _055339_, _055340_, _055341_, _055342_, _055343_, _055344_, _055345_, _055346_, _055347_, _055348_, _055349_, _055350_, _055351_, _055352_, _055353_, _055354_, _055355_, _055356_, _055357_, _055358_, _055359_, _055360_, _055361_, _055362_, _055363_, _055364_, _055365_, _055366_, _055367_, _055368_, _055369_, _055370_, _055371_, _055372_, _055373_, _055374_, _055375_, _055376_, _055377_, _055378_, _055379_, _055380_, _055381_, _055382_, _055383_, _055384_, _055385_, _055386_, _055387_, _055388_, _055389_, _055390_, _055391_, _055392_, _055393_, _055394_, _055395_, _055396_, _055397_, _055398_, _055399_, _055400_, _055401_, _055402_, _055403_, _055404_, _055405_, _055406_, _055407_, _055408_, _055409_, _055410_, _055411_, _055412_, _055413_, _055414_, _055415_, _055416_, _055417_, _055418_, _055419_, _055420_, _055421_, _055422_, _055423_, _055424_, _055425_, _055426_, _055427_, _055428_, _055429_, _055430_, _055431_, _055432_, _055433_, _055434_, _055435_, _055436_, _055437_, _055438_, _055439_, _055440_, _055441_, _055442_, _055443_, _055444_, _055445_, _055446_, _055447_, _055448_, _055449_, _055450_, _055451_, _055452_, _055453_, _055454_, _055455_, _055456_, _055457_, _055458_, _055459_, _055460_, _055461_, _055462_, _055463_, _055464_, _055465_, _055466_, _055467_, _055468_, _055469_, _055470_, _055471_, _055472_, _055473_, _055474_, _055475_, _055476_, _055477_, _055478_, _055479_, _055480_, _055481_, _055482_, _055483_, _055484_, _055485_, _055486_, _055487_, _055488_, _055489_, _055490_, _055491_, _055492_, _055493_, _055494_, _055495_, _055496_, _055497_, _055498_, _055499_, _055500_, _055501_, _055502_, _055503_, _055504_, _055505_, _055506_, _055507_, _055508_, _055509_, _055510_, _055511_, _055512_, _055513_, _055514_, _055515_, _055516_, _055517_, _055518_, _055519_, _055520_, _055521_, _055522_, _055523_, _055524_, _055525_, _055526_, _055527_, _055528_, _055529_, _055530_, _055531_, _055532_, _055533_, _055534_, _055535_, _055536_, _055537_, _055538_, _055539_, _055540_, _055541_, _055542_, _055543_, _055544_, _055545_, _055546_, _055547_, _055548_, _055549_, _055550_, _055551_, _055552_, _055553_, _055554_, _055555_, _055556_, _055557_, _055558_, _055559_, _055560_, _055561_, _055562_, _055563_, _055564_, _055565_, _055566_, _055567_, _055568_, _055569_, _055570_, _055571_, _055572_, _055573_, _055574_, _055575_, _055576_, _055577_, _055578_, _055579_, _055580_, _055581_, _055582_, _055583_, _055584_, _055585_, _055586_, _055587_, _055588_, _055589_, _055590_, _055591_, _055592_, _055593_, _055594_, _055595_, _055596_, _055597_, _055598_, _055599_, _055600_, _055601_, _055602_, _055603_, _055604_, _055605_, _055606_, _055607_, _055608_, _055609_, _055610_, _055611_, _055612_, _055613_, _055614_, _055615_, _055616_, _055617_, _055618_, _055619_, _055620_, _055621_, _055622_, _055623_, _055624_, _055625_, _055626_, _055627_, _055628_, _055629_, _055630_, _055631_, _055632_, _055633_, _055634_, _055635_, _055636_, _055637_, _055638_, _055639_, _055640_, _055641_, _055642_, _055643_, _055644_, _055645_, _055646_, _055647_, _055648_, _055649_, _055650_, _055651_, _055652_, _055653_, _055654_, _055655_, _055656_, _055657_, _055658_, _055659_, _055660_, _055661_, _055662_, _055663_, _055664_, _055665_, _055666_, _055667_, _055668_, _055669_, _055670_, _055671_, _055672_, _055673_, _055674_, _055675_, _055676_, _055677_, _055678_, _055679_, _055680_, _055681_, _055682_, _055683_, _055684_, _055685_, _055686_, _055687_, _055688_, _055689_, _055690_, _055691_, _055692_, _055693_, _055694_, _055695_, _055696_, _055697_, _055698_, _055699_, _055700_, _055701_, _055702_, _055703_, _055704_, _055705_, _055706_, _055707_, _055708_, _055709_, _055710_, _055711_, _055712_, _055713_, _055714_, _055715_, _055716_, _055717_, _055718_, _055719_, _055720_, _055721_, _055722_, _055723_, _055724_, _055725_, _055726_, _055727_, _055728_, _055729_, _055730_, _055731_, _055732_, _055733_, _055734_, _055735_, _055736_, _055737_, _055738_, _055739_, _055740_, _055741_, _055742_, _055743_, _055744_, _055745_, _055746_, _055747_, _055748_, _055749_, _055750_, _055751_, _055752_, _055753_, _055754_, _055755_, _055756_, _055757_, _055758_, _055759_, _055760_, _055761_, _055762_, _055763_, _055764_, _055765_, _055766_, _055767_, _055768_, _055769_, _055770_, _055771_, _055772_, _055773_, _055774_, _055775_, _055776_, _055777_, _055778_, _055779_, _055780_, _055781_, _055782_, _055783_, _055784_, _055785_, _055786_, _055787_, _055788_, _055789_, _055790_, _055791_, _055792_, _055793_, _055794_, _055795_, _055796_, _055797_, _055798_, _055799_, _055800_, _055801_, _055802_, _055803_, _055804_, _055805_, _055806_, _055807_, _055808_, _055809_, _055810_, _055811_, _055812_, _055813_, _055814_, _055815_, _055816_, _055817_, _055818_, _055819_, _055820_, _055821_, _055822_, _055823_, _055824_, _055825_, _055826_, _055827_, _055828_, _055829_, _055830_, _055831_, _055832_, _055833_, _055834_, _055835_, _055836_, _055837_, _055838_, _055839_, _055840_, _055841_, _055842_, _055843_, _055844_, _055845_, _055846_, _055847_, _055848_, _055849_, _055850_, _055851_, _055852_, _055853_, _055854_, _055855_, _055856_, _055857_, _055858_, _055859_, _055860_, _055861_, _055862_, _055863_, _055864_, _055865_, _055866_, _055867_, _055868_, _055869_, _055870_, _055871_, _055872_, _055873_, _055874_, _055875_, _055876_, _055877_, _055878_, _055879_, _055880_, _055881_, _055882_, _055883_, _055884_, _055885_, _055886_, _055887_, _055888_, _055889_, _055890_, _055891_, _055892_, _055893_, _055894_, _055895_, _055896_, _055897_, _055898_, _055899_, _055900_, _055901_, _055902_, _055903_, _055904_, _055905_, _055906_, _055907_, _055908_, _055909_, _055910_, _055911_, _055912_, _055913_, _055914_, _055915_, _055916_, _055917_, _055918_, _055919_, _055920_, _055921_, _055922_, _055923_, _055924_, _055925_, _055926_, _055927_, _055928_, _055929_, _055930_, _055931_, _055932_, _055933_, _055934_, _055935_, _055936_, _055937_, _055938_, _055939_, _055940_, _055941_, _055942_, _055943_, _055944_, _055945_, _055946_, _055947_, _055948_, _055949_, _055950_, _055951_, _055952_, _055953_, _055954_, _055955_, _055956_, _055957_, _055958_, _055959_, _055960_, _055961_, _055962_, _055963_, _055964_, _055965_, _055966_, _055967_, _055968_, _055969_, _055970_, _055971_, _055972_, _055973_, _055974_, _055975_, _055976_, _055977_, _055978_, _055979_, _055980_, _055981_, _055982_, _055983_, _055984_, _055985_, _055986_, _055987_, _055988_, _055989_, _055990_, _055991_, _055992_, _055993_, _055994_, _055995_, _055996_, _055997_, _055998_, _055999_, _056000_, _056001_, _056002_, _056003_, _056004_, _056005_, _056006_, _056007_, _056008_, _056009_, _056010_, _056011_, _056012_, _056013_, _056014_, _056015_, _056016_, _056017_, _056018_, _056019_, _056020_, _056021_, _056022_, _056023_, _056024_, _056025_, _056026_, _056027_, _056028_, _056029_, _056030_, _056031_, _056032_, _056033_, _056034_, _056035_, _056036_, _056037_, _056038_, _056039_, _056040_, _056041_, _056042_, _056043_, _056044_, _056045_, _056046_, _056047_, _056048_, _056049_, _056050_, _056051_, _056052_, _056053_, _056054_, _056055_, _056056_, _056057_, _056058_, _056059_, _056060_, _056061_, _056062_, _056063_, _056064_, _056065_, _056066_, _056067_, _056068_, _056069_, _056070_, _056071_, _056072_, _056073_, _056074_, _056075_, _056076_, _056077_, _056078_, _056079_, _056080_, _056081_, _056082_, _056083_, _056084_, _056085_, _056086_, _056087_, _056088_, _056089_, _056090_, _056091_, _056092_, _056093_, _056094_, _056095_, _056096_, _056097_, _056098_, _056099_, _056100_, _056101_, _056102_, _056103_, _056104_, _056105_, _056106_, _056107_, _056108_, _056109_, _056110_, _056111_, _056112_, _056113_, _056114_, _056115_, _056116_, _056117_, _056118_, _056119_, _056120_, _056121_, _056122_, _056123_, _056124_, _056125_, _056126_, _056127_, _056128_, _056129_, _056130_, _056131_, _056132_, _056133_, _056134_, _056135_, _056136_, _056137_, _056138_, _056139_, _056140_, _056141_, _056142_, _056143_, _056144_, _056145_, _056146_, _056147_, _056148_, _056149_, _056150_, _056151_, _056152_, _056153_, _056154_, _056155_, _056156_, _056157_, _056158_, _056159_, _056160_, _056161_, _056162_, _056163_, _056164_, _056165_, _056166_, _056167_, _056168_, _056169_, _056170_, _056171_, _056172_, _056173_, _056174_, _056175_, _056176_, _056177_, _056178_, _056179_, _056180_, _056181_, _056182_, _056183_, _056184_, _056185_, _056186_, _056187_, _056188_, _056189_, _056190_, _056191_, _056192_, _056193_, _056194_, _056195_, _056196_, _056197_, _056198_, _056199_, _056200_, _056201_, _056202_, _056203_, _056204_, _056205_, _056206_, _056207_, _056208_, _056209_, _056210_, _056211_, _056212_, _056213_, _056214_, _056215_, _056216_, _056217_, _056218_, _056219_, _056220_, _056221_, _056222_, _056223_, _056224_, _056225_, _056226_, _056227_, _056228_, _056229_, _056230_, _056231_, _056232_, _056233_, _056234_, _056235_, _056236_, _056237_, _056238_, _056239_, _056240_, _056241_, _056242_, _056243_, _056244_, _056245_, _056246_, _056247_, _056248_, _056249_, _056250_, _056251_, _056252_, _056253_, _056254_, _056255_, _056256_, _056257_, _056258_, _056259_, _056260_, _056261_, _056262_, _056263_, _056264_, _056265_, _056266_, _056267_, _056268_, _056269_, _056270_, _056271_, _056272_, _056273_, _056274_, _056275_, _056276_, _056277_, _056278_, _056279_, _056280_, _056281_, _056282_, _056283_, _056284_, _056285_, _056286_, _056287_, _056288_, _056289_, _056290_, _056291_, _056292_, _056293_, _056294_, _056295_, _056296_, _056297_, _056298_, _056299_, _056300_, _056301_, _056302_, _056303_, _056304_, _056305_, _056306_, _056307_, _056308_, _056309_, _056310_, _056311_, _056312_, _056313_, _056314_, _056315_, _056316_, _056317_, _056318_, _056319_, _056320_, _056321_, _056322_, _056323_, _056324_, _056325_, _056326_, _056327_, _056328_, _056329_, _056330_, _056331_, _056332_, _056333_, _056334_, _056335_, _056336_, _056337_, _056338_, _056339_, _056340_, _056341_, _056342_, _056343_, _056344_, _056345_, _056346_, _056347_, _056348_, _056349_, _056350_, _056351_, _056352_, _056353_, _056354_, _056355_, _056356_, _056357_, _056358_, _056359_, _056360_, _056361_, _056362_, _056363_, _056364_, _056365_, _056366_, _056367_, _056368_, _056369_, _056370_, _056371_, _056372_, _056373_, _056374_, _056375_, _056376_, _056377_, _056378_, _056379_, _056380_, _056381_, _056382_, _056383_, _056384_, _056385_, _056386_, _056387_, _056388_, _056389_, _056390_, _056391_, _056392_, _056393_, _056394_, _056395_, _056396_, _056397_, _056398_, _056399_, _056400_, _056401_, _056402_, _056403_, _056404_, _056405_, _056406_, _056407_, _056408_, _056409_, _056410_, _056411_, _056412_, _056413_, _056414_, _056415_, _056416_, _056417_, _056418_, _056419_, _056420_, _056421_, _056422_, _056423_, _056424_, _056425_, _056426_, _056427_, _056428_, _056429_, _056430_, _056431_, _056432_, _056433_, _056434_, _056435_, _056436_, _056437_, _056438_, _056439_, _056440_, _056441_, _056442_, _056443_, _056444_, _056445_, _056446_, _056447_, _056448_, _056449_, _056450_, _056451_, _056452_, _056453_, _056454_, _056455_, _056456_, _056457_, _056458_, _056459_, _056460_, _056461_, _056462_, _056463_, _056464_, _056465_, _056466_, _056467_, _056468_, _056469_, _056470_, _056471_, _056472_, _056473_, _056474_, _056475_, _056476_, _056477_, _056478_, _056479_, _056480_, _056481_, _056482_, _056483_, _056484_, _056485_, _056486_, _056487_, _056488_, _056489_, _056490_, _056491_, _056492_, _056493_, _056494_, _056495_, _056496_, _056497_, _056498_, _056499_, _056500_, _056501_, _056502_, _056503_, _056504_, _056505_, _056506_, _056507_, _056508_, _056509_, _056510_, _056511_, _056512_, _056513_, _056514_, _056515_, _056516_, _056517_, _056518_, _056519_, _056520_, _056521_, _056522_, _056523_, _056524_, _056525_, _056526_, _056527_, _056528_, _056529_, _056530_, _056531_, _056532_, _056533_, _056534_, _056535_, _056536_, _056537_, _056538_, _056539_, _056540_, _056541_, _056542_, _056543_, _056544_, _056545_, _056546_, _056547_, _056548_, _056549_, _056550_, _056551_, _056552_, _056553_, _056554_, _056555_, _056556_, _056557_, _056558_, _056559_, _056560_, _056561_, _056562_, _056563_, _056564_, _056565_, _056566_, _056567_, _056568_, _056569_, _056570_, _056571_, _056572_, _056573_, _056574_, _056575_, _056576_, _056577_, _056578_, _056579_, _056580_, _056581_, _056582_, _056583_, _056584_, _056585_, _056586_, _056587_, _056588_, _056589_, _056590_, _056591_, _056592_, _056593_, _056594_, _056595_, _056596_, _056597_, _056598_, _056599_, _056600_, _056601_, _056602_, _056603_, _056604_, _056605_, _056606_, _056607_, _056608_, _056609_, _056610_, _056611_, _056612_, _056613_, _056614_, _056615_, _056616_, _056617_, _056618_, _056619_, _056620_, _056621_, _056622_, _056623_, _056624_, _056625_, _056626_, _056627_, _056628_, _056629_, _056630_, _056631_, _056632_, _056633_, _056634_, _056635_, _056636_, _056637_, _056638_, _056639_, _056640_, _056641_, _056642_, _056643_, _056644_, _056645_, _056646_, _056647_, _056648_, _056649_, _056650_, _056651_, _056652_, _056653_, _056654_, _056655_, _056656_, _056657_, _056658_, _056659_, _056660_, _056661_, _056662_, _056663_, _056664_, _056665_, _056666_, _056667_, _056668_, _056669_, _056670_, _056671_, _056672_, _056673_, _056674_, _056675_, _056676_, _056677_, _056678_, _056679_, _056680_, _056681_, _056682_, _056683_, _056684_, _056685_, _056686_, _056687_, _056688_, _056689_, _056690_, _056691_, _056692_, _056693_, _056694_, _056695_, _056696_, _056697_, _056698_, _056699_, _056700_, _056701_, _056702_, _056703_, _056704_, _056705_, _056706_, _056707_, _056708_, _056709_, _056710_, _056711_, _056712_, _056713_, _056714_, _056715_, _056716_, _056717_, _056718_, _056719_, _056720_, _056721_, _056722_, _056723_, _056724_, _056725_, _056726_, _056727_, _056728_, _056729_, _056730_, _056731_, _056732_, _056733_, _056734_, _056735_, _056736_, _056737_, _056738_, _056739_, _056740_, _056741_, _056742_, _056743_, _056744_, _056745_, _056746_, _056747_, _056748_, _056749_, _056750_, _056751_, _056752_, _056753_, _056754_, _056755_, _056756_, _056757_, _056758_, _056759_, _056760_, _056761_, _056762_, _056763_, _056764_, _056765_, _056766_, _056767_, _056768_, _056769_, _056770_, _056771_, _056772_, _056773_, _056774_, _056775_, _056776_, _056777_, _056778_, _056779_, _056780_, _056781_, _056782_, _056783_, _056784_, _056785_, _056786_, _056787_, _056788_, _056789_, _056790_, _056791_, _056792_, _056793_, _056794_, _056795_, _056796_, _056797_, _056798_, _056799_, _056800_, _056801_, _056802_, _056803_, _056804_, _056805_, _056806_, _056807_, _056808_, _056809_, _056810_, _056811_, _056812_, _056813_, _056814_, _056815_, _056816_, _056817_, _056818_, _056819_, _056820_, _056821_, _056822_, _056823_, _056824_, _056825_, _056826_, _056827_, _056828_, _056829_, _056830_, _056831_, _056832_, _056833_, _056834_, _056835_, _056836_, _056837_, _056838_, _056839_, _056840_, _056841_, _056842_, _056843_, _056844_, _056845_, _056846_, _056847_, _056848_, _056849_, _056850_, _056851_, _056852_, _056853_, _056854_, _056855_, _056856_, _056857_, _056858_, _056859_, _056860_, _056861_, _056862_, _056863_, _056864_, _056865_, _056866_, _056867_, _056868_, _056869_, _056870_, _056871_, _056872_, _056873_, _056874_, _056875_, _056876_, _056877_, _056878_, _056879_, _056880_, _056881_, _056882_, _056883_, _056884_, _056885_, _056886_, _056887_, _056888_, _056889_, _056890_, _056891_, _056892_, _056893_, _056894_, _056895_, _056896_, _056897_, _056898_, _056899_, _056900_, _056901_, _056902_, _056903_, _056904_, _056905_, _056906_, _056907_, _056908_, _056909_, _056910_, _056911_, _056912_, _056913_, _056914_, _056915_, _056916_, _056917_, _056918_, _056919_, _056920_, _056921_, _056922_, _056923_, _056924_, _056925_, _056926_, _056927_, _056928_, _056929_, _056930_, _056931_, _056932_, _056933_, _056934_, _056935_, _056936_, _056937_, _056938_, _056939_, _056940_, _056941_, _056942_, _056943_, _056944_, _056945_, _056946_, _056947_, _056948_, _056949_, _056950_, _056951_, _056952_, _056953_, _056954_, _056955_, _056956_, _056957_, _056958_, _056959_, _056960_, _056961_, _056962_, _056963_, _056964_, _056965_, _056966_, _056967_, _056968_, _056969_, _056970_, _056971_, _056972_, _056973_, _056974_, _056975_, _056976_, _056977_, _056978_, _056979_, _056980_, _056981_, _056982_, _056983_, _056984_, _056985_, _056986_, _056987_, _056988_, _056989_, _056990_, _056991_, _056992_, _056993_, _056994_, _056995_, _056996_, _056997_, _056998_, _056999_, _057000_, _057001_, _057002_, _057003_, _057004_, _057005_, _057006_, _057007_, _057008_, _057009_, _057010_, _057011_, _057012_, _057013_, _057014_, _057015_, _057016_, _057017_, _057018_, _057019_, _057020_, _057021_, _057022_, _057023_, _057024_, _057025_, _057026_, _057027_, _057028_, _057029_, _057030_, _057031_, _057032_, _057033_, _057034_, _057035_, _057036_, _057037_, _057038_, _057039_, _057040_, _057041_, _057042_, _057043_, _057044_, _057045_, _057046_, _057047_, _057048_, _057049_, _057050_, _057051_, _057052_, _057053_, _057054_, _057055_, _057056_, _057057_, _057058_, _057059_, _057060_, _057061_, _057062_, _057063_, _057064_, _057065_, _057066_, _057067_, _057068_, _057069_, _057070_, _057071_, _057072_, _057073_, _057074_, _057075_, _057076_, _057077_, _057078_, _057079_, _057080_, _057081_, _057082_, _057083_, _057084_, _057085_, _057086_, _057087_, _057088_, _057089_, _057090_, _057091_, _057092_, _057093_, _057094_, _057095_, _057096_, _057097_, _057098_, _057099_, _057100_, _057101_, _057102_, _057103_, _057104_, _057105_, _057106_, _057107_, _057108_, _057109_, _057110_, _057111_, _057112_, _057113_, _057114_, _057115_, _057116_, _057117_, _057118_, _057119_, _057120_, _057121_, _057122_, _057123_, _057124_, _057125_, _057126_, _057127_, _057128_, _057129_, _057130_, _057131_, _057132_, _057133_, _057134_, _057135_, _057136_, _057137_, _057138_, _057139_, _057140_, _057141_, _057142_, _057143_, _057144_, _057145_, _057146_, _057147_, _057148_, _057149_, _057150_, _057151_, _057152_, _057153_, _057154_, _057155_, _057156_, _057157_, _057158_, _057159_, _057160_, _057161_, _057162_, _057163_, _057164_, _057165_, _057166_, _057167_, _057168_, _057169_, _057170_, _057171_, _057172_, _057173_, _057174_, _057175_, _057176_, _057177_, _057178_, _057179_, _057180_, _057181_, _057182_, _057183_, _057184_, _057185_, _057186_, _057187_, _057188_, _057189_, _057190_, _057191_, _057192_, _057193_, _057194_, _057195_, _057196_, _057197_, _057198_, _057199_, _057200_, _057201_, _057202_, _057203_, _057204_, _057205_, _057206_, _057207_, _057208_, _057209_, _057210_, _057211_, _057212_, _057213_, _057214_, _057215_, _057216_, _057217_, _057218_, _057219_, _057220_, _057221_, _057222_, _057223_, _057224_, _057225_, _057226_, _057227_, _057228_, _057229_, _057230_, _057231_, _057232_, _057233_, _057234_, _057235_, _057236_, _057237_, _057238_, _057239_, _057240_, _057241_, _057242_, _057243_, _057244_, _057245_, _057246_, _057247_, _057248_, _057249_, _057250_, _057251_, _057252_, _057253_, _057254_, _057255_, _057256_, _057257_, _057258_, _057259_, _057260_, _057261_, _057262_, _057263_, _057264_, _057265_, _057266_, _057267_, _057268_, _057269_, _057270_, _057271_, _057272_, _057273_, _057274_, _057275_, _057276_, _057277_, _057278_, _057279_, _057280_, _057281_, _057282_, _057283_, _057284_, _057285_, _057286_, _057287_, _057288_, _057289_, _057290_, _057291_, _057292_, _057293_, _057294_, _057295_, _057296_, _057297_, _057298_, _057299_, _057300_, _057301_, _057302_, _057303_, _057304_, _057305_, _057306_, _057307_, _057308_, _057309_, _057310_, _057311_, _057312_, _057313_, _057314_, _057315_, _057316_, _057317_, _057318_, _057319_, _057320_, _057321_, _057322_, _057323_, _057324_, _057325_, _057326_, _057327_, _057328_, _057329_, _057330_, _057331_, _057332_, _057333_, _057334_, _057335_, _057336_, _057337_, _057338_, _057339_, _057340_, _057341_, _057342_, _057343_, _057344_, _057345_, _057346_, _057347_, _057348_, _057349_, _057350_, _057351_, _057352_, _057353_, _057354_, _057355_, _057356_, _057357_, _057358_, _057359_, _057360_, _057361_, _057362_, _057363_, _057364_, _057365_, _057366_, _057367_, _057368_, _057369_, _057370_, _057371_, _057372_, _057373_, _057374_, _057375_, _057376_, _057377_, _057378_, _057379_, _057380_, _057381_, _057382_, _057383_, _057384_, _057385_, _057386_, _057387_, _057388_, _057389_, _057390_, _057391_, _057392_, _057393_, _057394_, _057395_, _057396_, _057397_, _057398_, _057399_, _057400_, _057401_, _057402_, _057403_, _057404_, _057405_, _057406_, _057407_, _057408_, _057409_, _057410_, _057411_, _057412_, _057413_, _057414_, _057415_, _057416_, _057417_, _057418_, _057419_, _057420_, _057421_, _057422_, _057423_, _057424_, _057425_, _057426_, _057427_, _057428_, _057429_, _057430_, _057431_, _057432_, _057433_, _057434_, _057435_, _057436_, _057437_, _057438_, _057439_, _057440_, _057441_, _057442_, _057443_, _057444_, _057445_, _057446_, _057447_, _057448_, _057449_, _057450_, _057451_, _057452_, _057453_, _057454_, _057455_, _057456_, _057457_, _057458_, _057459_, _057460_, _057461_, _057462_, _057463_, _057464_, _057465_, _057466_, _057467_, _057468_, _057469_, _057470_, _057471_, _057472_, _057473_, _057474_, _057475_, _057476_, _057477_, _057478_, _057479_, _057480_, _057481_, _057482_, _057483_, _057484_, _057485_, _057486_, _057487_, _057488_, _057489_, _057490_, _057491_, _057492_, _057493_, _057494_, _057495_, _057496_, _057497_, _057498_, _057499_, _057500_, _057501_, _057502_, _057503_, _057504_, _057505_, _057506_, _057507_, _057508_, _057509_, _057510_, _057511_, _057512_, _057513_, _057514_, _057515_, _057516_, _057517_, _057518_, _057519_, _057520_, _057521_, _057522_, _057523_, _057524_, _057525_, _057526_, _057527_, _057528_, _057529_, _057530_, _057531_, _057532_, _057533_, _057534_, _057535_, _057536_, _057537_, _057538_, _057539_, _057540_, _057541_, _057542_, _057543_, _057544_, _057545_, _057546_, _057547_, _057548_, _057549_, _057550_, _057551_, _057552_, _057553_, _057554_, _057555_, _057556_, _057557_, _057558_, _057559_, _057560_, _057561_, _057562_, _057563_, _057564_, _057565_, _057566_, _057567_, _057568_, _057569_, _057570_, _057571_, _057572_, _057573_, _057574_, _057575_, _057576_, _057577_, _057578_, _057579_, _057580_, _057581_, _057582_, _057583_, _057584_, _057585_, _057586_, _057587_, _057588_, _057589_, _057590_, _057591_, _057592_, _057593_, _057594_, _057595_, _057596_, _057597_, _057598_, _057599_, _057600_, _057601_, _057602_, _057603_, _057604_, _057605_, _057606_, _057607_, _057608_, _057609_, _057610_, _057611_, _057612_, _057613_, _057614_, _057615_, _057616_, _057617_, _057618_, _057619_, _057620_, _057621_, _057622_, _057623_, _057624_, _057625_, _057626_, _057627_, _057628_, _057629_, _057630_, _057631_, _057632_, _057633_, _057634_, _057635_, _057636_, _057637_, _057638_, _057639_, _057640_, _057641_, _057642_, _057643_, _057644_, _057645_, _057646_, _057647_, _057648_, _057649_, _057650_, _057651_, _057652_, _057653_, _057654_, _057655_, _057656_, _057657_, _057658_, _057659_, _057660_, _057661_, _057662_, _057663_, _057664_, _057665_, _057666_, _057667_, _057668_, _057669_, _057670_, _057671_, _057672_, _057673_, _057674_, _057675_, _057676_, _057677_, _057678_, _057679_, _057680_, _057681_, _057682_, _057683_, _057684_, _057685_, _057686_, _057687_, _057688_, _057689_, _057690_, _057691_, _057692_, _057693_, _057694_, _057695_, _057696_, _057697_, _057698_, _057699_, _057700_, _057701_, _057702_, _057703_, _057704_, _057705_, _057706_, _057707_, _057708_, _057709_, _057710_, _057711_, _057712_, _057713_, _057714_, _057715_, _057716_, _057717_, _057718_, _057719_, _057720_, _057721_, _057722_, _057723_, _057724_, _057725_, _057726_, _057727_, _057728_, _057729_, _057730_, _057731_, _057732_, _057733_, _057734_, _057735_, _057736_, _057737_, _057738_, _057739_, _057740_, _057741_, _057742_, _057743_, _057744_, _057745_, _057746_, _057747_, _057748_, _057749_, _057750_, _057751_, _057752_, _057753_, _057754_, _057755_, _057756_, _057757_, _057758_, _057759_, _057760_, _057761_, _057762_, _057763_, _057764_, _057765_, _057766_, _057767_, _057768_, _057769_, _057770_, _057771_, _057772_, _057773_, _057774_, _057775_, _057776_, _057777_, _057778_, _057779_, _057780_, _057781_, _057782_, _057783_, _057784_, _057785_, _057786_, _057787_, _057788_, _057789_, _057790_, _057791_, _057792_, _057793_, _057794_, _057795_, _057796_, _057797_, _057798_, _057799_, _057800_, _057801_, _057802_, _057803_, _057804_, _057805_, _057806_, _057807_, _057808_, _057809_, _057810_, _057811_, _057812_, _057813_, _057814_, _057815_, _057816_, _057817_, _057818_, _057819_, _057820_, _057821_, _057822_, _057823_, _057824_, _057825_, _057826_, _057827_, _057828_, _057829_, _057830_, _057831_, _057832_, _057833_, _057834_, _057835_, _057836_, _057837_, _057838_, _057839_, _057840_, _057841_, _057842_, _057843_, _057844_, _057845_, _057846_, _057847_, _057848_, _057849_, _057850_, _057851_, _057852_, _057853_, _057854_, _057855_, _057856_, _057857_, _057858_, _057859_, _057860_, _057861_, _057862_, _057863_, _057864_, _057865_, _057866_, _057867_, _057868_, _057869_, _057870_, _057871_, _057872_, _057873_, _057874_, _057875_, _057876_, _057877_, _057878_, _057879_, _057880_, _057881_, _057882_, _057883_, _057884_, _057885_, _057886_, _057887_, _057888_, _057889_, _057890_, _057891_, _057892_, _057893_, _057894_, _057895_, _057896_, _057897_, _057898_, _057899_, _057900_, _057901_, _057902_, _057903_, _057904_, _057905_, _057906_, _057907_, _057908_, _057909_, _057910_, _057911_, _057912_, _057913_, _057914_, _057915_, _057916_, _057917_, _057918_, _057919_, _057920_, _057921_, _057922_, _057923_, _057924_, _057925_, _057926_, _057927_, _057928_, _057929_, _057930_, _057931_, _057932_, _057933_, _057934_, _057935_, _057936_, _057937_, _057938_, _057939_, _057940_, _057941_, _057942_, _057943_, _057944_, _057945_, _057946_, _057947_, _057948_, _057949_, _057950_, _057951_, _057952_, _057953_, _057954_, _057955_, _057956_, _057957_, _057958_, _057959_, _057960_, _057961_, _057962_, _057963_, _057964_, _057965_, _057966_, _057967_, _057968_, _057969_, _057970_, _057971_, _057972_, _057973_, _057974_, _057975_, _057976_, _057977_, _057978_, _057979_, _057980_, _057981_, _057982_, _057983_, _057984_, _057985_, _057986_, _057987_, _057988_, _057989_, _057990_, _057991_, _057992_, _057993_, _057994_, _057995_, _057996_, _057997_, _057998_, _057999_, _058000_, _058001_, _058002_, _058003_, _058004_, _058005_, _058006_, _058007_, _058008_, _058009_, _058010_, _058011_, _058012_, _058013_, _058014_, _058015_, _058016_, _058017_, _058018_, _058019_, _058020_, _058021_, _058022_, _058023_, _058024_, _058025_, _058026_, _058027_, _058028_, _058029_, _058030_, _058031_, _058032_, _058033_, _058034_, _058035_, _058036_, _058037_, _058038_, _058039_, _058040_, _058041_, _058042_, _058043_, _058044_, _058045_, _058046_, _058047_, _058048_, _058049_, _058050_, _058051_, _058052_, _058053_, _058054_, _058055_, _058056_, _058057_, _058058_, _058059_, _058060_, _058061_, _058062_, _058063_, _058064_, _058065_, _058066_, _058067_, _058068_, _058069_, _058070_, _058071_, _058072_, _058073_, _058074_, _058075_, _058076_, _058077_, _058078_, _058079_, _058080_, _058081_, _058082_, _058083_, _058084_, _058085_, _058086_, _058087_, _058088_, _058089_, _058090_, _058091_, _058092_, _058093_, _058094_, _058095_, _058096_, _058097_, _058098_, _058099_, _058100_, _058101_, _058102_, _058103_, _058104_, _058105_, _058106_, _058107_, _058108_, _058109_, _058110_, _058111_, _058112_, _058113_, _058114_, _058115_, _058116_, _058117_, _058118_, _058119_, _058120_, _058121_, _058122_, _058123_, _058124_, _058125_, _058126_, _058127_, _058128_, _058129_, _058130_, _058131_, _058132_, _058133_, _058134_, _058135_, _058136_, _058137_, _058138_, _058139_, _058140_, _058141_, _058142_, _058143_, _058144_, _058145_, _058146_, _058147_, _058148_, _058149_, _058150_, _058151_, _058152_, _058153_, _058154_, _058155_, _058156_, _058157_, _058158_, _058159_, _058160_, _058161_, _058162_, _058163_, _058164_, _058165_, _058166_, _058167_, _058168_, _058169_, _058170_, _058171_, _058172_, _058173_, _058174_, _058175_, _058176_, _058177_, _058178_, _058179_, _058180_, _058181_, _058182_, _058183_, _058184_, _058185_, _058186_, _058187_, _058188_, _058189_, _058190_, _058191_, _058192_, _058193_, _058194_, _058195_, _058196_, _058197_, _058198_, _058199_, _058200_, _058201_, _058202_, _058203_, _058204_, _058205_, _058206_, _058207_, _058208_, _058209_, _058210_, _058211_, _058212_, _058213_, _058214_, _058215_, _058216_, _058217_, _058218_, _058219_, _058220_, _058221_, _058222_, _058223_, _058224_, _058225_, _058226_, _058227_, _058228_, _058229_, _058230_, _058231_, _058232_, _058233_, _058234_, _058235_, _058236_, _058237_, _058238_, _058239_, _058240_, _058241_, _058242_, _058243_, _058244_, _058245_, _058246_, _058247_, _058248_, _058249_, _058250_, _058251_, _058252_, _058253_, _058254_, _058255_, _058256_, _058257_, _058258_, _058259_, _058260_, _058261_, _058262_, _058263_, _058264_, _058265_, _058266_, _058267_, _058268_, _058269_, _058270_, _058271_, _058272_, _058273_, _058274_, _058275_, _058276_, _058277_, _058278_, _058279_, _058280_, _058281_, _058282_, _058283_, _058284_, _058285_, _058286_, _058287_, _058288_, _058289_, _058290_, _058291_, _058292_, _058293_, _058294_, _058295_, _058296_, _058297_, _058298_, _058299_, _058300_, _058301_, _058302_, _058303_, _058304_, _058305_, _058306_, _058307_, _058308_, _058309_, _058310_, _058311_, _058312_, _058313_, _058314_, _058315_, _058316_, _058317_, _058318_, _058319_, _058320_, _058321_, _058322_, _058323_, _058324_, _058325_, _058326_, _058327_, _058328_, _058329_, _058330_, _058331_, _058332_, _058333_, _058334_, _058335_, _058336_, _058337_, _058338_, _058339_, _058340_, _058341_, _058342_, _058343_, _058344_, _058345_, _058346_, _058347_, _058348_, _058349_, _058350_, _058351_, _058352_, _058353_, _058354_, _058355_, _058356_, _058357_, _058358_, _058359_, _058360_, _058361_, _058362_, _058363_, _058364_, _058365_, _058366_, _058367_, _058368_, _058369_, _058370_, _058371_, _058372_, _058373_, _058374_, _058375_, _058376_, _058377_, _058378_, _058379_, _058380_, _058381_, _058382_, _058383_, _058384_, _058385_, _058386_, _058387_, _058388_, _058389_, _058390_, _058391_, _058392_, _058393_, _058394_, _058395_, _058396_, _058397_, _058398_, _058399_, _058400_, _058401_, _058402_, _058403_, _058404_, _058405_, _058406_, _058407_, _058408_, _058409_, _058410_, _058411_, _058412_, _058413_, _058414_, _058415_, _058416_, _058417_, _058418_, _058419_, _058420_, _058421_, _058422_, _058423_, _058424_, _058425_, _058426_, _058427_, _058428_, _058429_, _058430_, _058431_, _058432_, _058433_, _058434_, _058435_, _058436_, _058437_, _058438_, _058439_, _058440_, _058441_, _058442_, _058443_, _058444_, _058445_, _058446_, _058447_, _058448_, _058449_, _058450_, _058451_, _058452_, _058453_, _058454_, _058455_, _058456_, _058457_, _058458_, _058459_, _058460_, _058461_, _058462_, _058463_, _058464_, _058465_, _058466_, _058467_, _058468_, _058469_, _058470_, _058471_, _058472_, _058473_, _058474_, _058475_, _058476_, _058477_, _058478_, _058479_, _058480_, _058481_, _058482_, _058483_, _058484_, _058485_, _058486_, _058487_, _058488_, _058489_, _058490_, _058491_, _058492_, _058493_, _058494_, _058495_, _058496_, _058497_, _058498_, _058499_, _058500_, _058501_, _058502_, _058503_, _058504_, _058505_, _058506_, _058507_, _058508_, _058509_, _058510_, _058511_, _058512_, _058513_, _058514_, _058515_, _058516_, _058517_, _058518_, _058519_, _058520_, _058521_, _058522_, _058523_, _058524_, _058525_, _058526_, _058527_, _058528_, _058529_, _058530_, _058531_, _058532_, _058533_, _058534_, _058535_, _058536_, _058537_, _058538_, _058539_, _058540_, _058541_, _058542_, _058543_, _058544_, _058545_, _058546_, _058547_, _058548_, _058549_, _058550_, _058551_, _058552_, _058553_, _058554_, _058555_, _058556_, _058557_, _058558_, _058559_, _058560_, _058561_, _058562_, _058563_, _058564_, _058565_, _058566_, _058567_, _058568_, _058569_, _058570_, _058571_, _058572_, _058573_, _058574_, _058575_, _058576_, _058577_, _058578_, _058579_, _058580_, _058581_, _058582_, _058583_, _058584_, _058585_, _058586_, _058587_, _058588_, _058589_, _058590_, _058591_, _058592_, _058593_, _058594_, _058595_, _058596_, _058597_, _058598_, _058599_, _058600_, _058601_, _058602_, _058603_, _058604_, _058605_, _058606_, _058607_, _058608_, _058609_, _058610_, _058611_, _058612_, _058613_, _058614_, _058615_, _058616_, _058617_, _058618_, _058619_, _058620_, _058621_, _058622_, _058623_, _058624_, _058625_, _058626_, _058627_, _058628_, _058629_, _058630_, _058631_, _058632_, _058633_, _058634_, _058635_, _058636_, _058637_, _058638_, _058639_, _058640_, _058641_, _058642_, _058643_, _058644_, _058645_, _058646_, _058647_, _058648_, _058649_, _058650_, _058651_, _058652_, _058653_, _058654_, _058655_, _058656_, _058657_, _058658_, _058659_, _058660_, _058661_, _058662_, _058663_, _058664_, _058665_, _058666_, _058667_, _058668_, _058669_, _058670_, _058671_, _058672_, _058673_, _058674_, _058675_, _058676_, _058677_, _058678_, _058679_, _058680_, _058681_, _058682_, _058683_, _058684_, _058685_, _058686_, _058687_, _058688_, _058689_, _058690_, _058691_, _058692_, _058693_, _058694_, _058695_, _058696_, _058697_, _058698_, _058699_, _058700_, _058701_, _058702_, _058703_, _058704_, _058705_, _058706_, _058707_, _058708_, _058709_, _058710_, _058711_, _058712_, _058713_, _058714_, _058715_, _058716_, _058717_, _058718_, _058719_, _058720_, _058721_, _058722_, _058723_, _058724_, _058725_, _058726_, _058727_, _058728_, _058729_, _058730_, _058731_, _058732_, _058733_, _058734_, _058735_, _058736_, _058737_, _058738_, _058739_, _058740_, _058741_, _058742_, _058743_, _058744_, _058745_, _058746_, _058747_, _058748_, _058749_, _058750_, _058751_, _058752_, _058753_, _058754_, _058755_, _058756_, _058757_, _058758_, _058759_, _058760_, _058761_, _058762_, _058763_, _058764_, _058765_, _058766_, _058767_, _058768_, _058769_, _058770_, _058771_, _058772_, _058773_, _058774_, _058775_, _058776_, _058777_, _058778_, _058779_, _058780_, _058781_, _058782_, _058783_, _058784_, _058785_, _058786_, _058787_, _058788_, _058789_, _058790_, _058791_, _058792_, _058793_, _058794_, _058795_, _058796_, _058797_, _058798_, _058799_, _058800_, _058801_, _058802_, _058803_, _058804_, _058805_, _058806_, _058807_, _058808_, _058809_, _058810_, _058811_, _058812_, _058813_, _058814_, _058815_, _058816_, _058817_, _058818_, _058819_, _058820_, _058821_, _058822_, _058823_, _058824_, _058825_, _058826_, _058827_, _058828_, _058829_, _058830_, _058831_, _058832_, _058833_, _058834_, _058835_, _058836_, _058837_, _058838_, _058839_, _058840_, _058841_, _058842_, _058843_, _058844_, _058845_, _058846_, _058847_, _058848_, _058849_, _058850_, _058851_, _058852_, _058853_, _058854_, _058855_, _058856_, _058857_, _058858_, _058859_, _058860_, _058861_, _058862_, _058863_, _058864_, _058865_, _058866_, _058867_, _058868_, _058869_, _058870_, _058871_, _058872_, _058873_, _058874_, _058875_, _058876_, _058877_, _058878_, _058879_, _058880_, _058881_, _058882_, _058883_, _058884_, _058885_, _058886_, _058887_, _058888_, _058889_, _058890_, _058891_, _058892_, _058893_, _058894_, _058895_, _058896_, _058897_, _058898_, _058899_, _058900_, _058901_, _058902_, _058903_, _058904_, _058905_, _058906_, _058907_, _058908_, _058909_, _058910_, _058911_, _058912_, _058913_, _058914_, _058915_, _058916_, _058917_, _058918_, _058919_, _058920_, _058921_, _058922_, _058923_, _058924_, _058925_, _058926_, _058927_, _058928_, _058929_, _058930_, _058931_, _058932_, _058933_, _058934_, _058935_, _058936_, _058937_, _058938_, _058939_, _058940_, _058941_, _058942_, _058943_, _058944_, _058945_, _058946_, _058947_, _058948_, _058949_, _058950_, _058951_, _058952_, _058953_, _058954_, _058955_, _058956_, _058957_, _058958_, _058959_, _058960_, _058961_, _058962_, _058963_, _058964_, _058965_, _058966_, _058967_, _058968_, _058969_, _058970_, _058971_, _058972_, _058973_, _058974_, _058975_, _058976_, _058977_, _058978_, _058979_, _058980_, _058981_, _058982_, _058983_, _058984_, _058985_, _058986_, _058987_, _058988_, _058989_, _058990_, _058991_, _058992_, _058993_, _058994_, _058995_, _058996_, _058997_, _058998_, _058999_, _059000_, _059001_, _059002_, _059003_, _059004_, _059005_, _059006_, _059007_, _059008_, _059009_, _059010_, _059011_, _059012_, _059013_, _059014_, _059015_, _059016_, _059017_, _059018_, _059019_, _059020_, _059021_, _059022_, _059023_, _059024_, _059025_, _059026_, _059027_, _059028_, _059029_, _059030_, _059031_, _059032_, _059033_, _059034_, _059035_, _059036_, _059037_, _059038_, _059039_, _059040_, _059041_, _059042_, _059043_, _059044_, _059045_, _059046_, _059047_, _059048_, _059049_, _059050_, _059051_, _059052_, _059053_, _059054_, _059055_, _059056_, _059057_, _059058_, _059059_, _059060_, _059061_, _059062_, _059063_, _059064_, _059065_, _059066_, _059067_, _059068_, _059069_, _059070_, _059071_, _059072_, _059073_, _059074_, _059075_, _059076_, _059077_, _059078_, _059079_, _059080_, _059081_, _059082_, _059083_, _059084_, _059085_, _059086_, _059087_, _059088_, _059089_, _059090_, _059091_, _059092_, _059093_, _059094_, _059095_, _059096_, _059097_, _059098_, _059099_, _059100_, _059101_, _059102_, _059103_, _059104_, _059105_, _059106_, _059107_, _059108_, _059109_, _059110_, _059111_, _059112_, _059113_, _059114_, _059115_, _059116_, _059117_, _059118_, _059119_, _059120_, _059121_, _059122_, _059123_, _059124_, _059125_, _059126_, _059127_, _059128_, _059129_, _059130_, _059131_, _059132_, _059133_, _059134_, _059135_, _059136_, _059137_, _059138_, _059139_, _059140_, _059141_, _059142_, _059143_, _059144_, _059145_, _059146_, _059147_, _059148_, _059149_, _059150_, _059151_, _059152_, _059153_, _059154_, _059155_, _059156_, _059157_, _059158_, _059159_, _059160_, _059161_, _059162_, _059163_, _059164_, _059165_, _059166_, _059167_, _059168_, _059169_, _059170_, _059171_, _059172_, _059173_, _059174_, _059175_, _059176_, _059177_, _059178_, _059179_, _059180_, _059181_, _059182_, _059183_, _059184_, _059185_, _059186_, _059187_, _059188_, _059189_, _059190_, _059191_, _059192_, _059193_, _059194_, _059195_, _059196_, _059197_, _059198_, _059199_, _059200_, _059201_, _059202_, _059203_, _059204_, _059205_, _059206_, _059207_, _059208_, _059209_, _059210_, _059211_, _059212_, _059213_, _059214_, _059215_, _059216_, _059217_, _059218_, _059219_, _059220_, _059221_, _059222_, _059223_, _059224_, _059225_, _059226_, _059227_, _059228_, _059229_, _059230_, _059231_, _059232_, _059233_, _059234_, _059235_, _059236_, _059237_, _059238_, _059239_, _059240_, _059241_, _059242_, _059243_, _059244_, _059245_, _059246_, _059247_, _059248_, _059249_, _059250_, _059251_, _059252_, _059253_, _059254_, _059255_, _059256_, _059257_, _059258_, _059259_, _059260_, _059261_, _059262_, _059263_, _059264_, _059265_, _059266_, _059267_, _059268_, _059269_, _059270_, _059271_, _059272_, _059273_, _059274_, _059275_, _059276_, _059277_, _059278_, _059279_, _059280_, _059281_, _059282_, _059283_, _059284_, _059285_, _059286_, _059287_, _059288_, _059289_, _059290_, _059291_, _059292_, _059293_, _059294_, _059295_, _059296_, _059297_, _059298_, _059299_, _059300_, _059301_, _059302_, _059303_, _059304_, _059305_, _059306_, _059307_, _059308_, _059309_, _059310_, _059311_, _059312_, _059313_, _059314_, _059315_, _059316_, _059317_, _059318_, _059319_, _059320_, _059321_, _059322_, _059323_, _059324_, _059325_, _059326_, _059327_, _059328_, _059329_, _059330_, _059331_, _059332_, _059333_, _059334_, _059335_, _059336_, _059337_, _059338_, _059339_, _059340_, _059341_, _059342_, _059343_, _059344_, _059345_, _059346_, _059347_, _059348_, _059349_, _059350_, _059351_, _059352_, _059353_, _059354_, _059355_, _059356_, _059357_, _059358_, _059359_, _059360_, _059361_, _059362_, _059363_, _059364_, _059365_, _059366_, _059367_, _059368_, _059369_, _059370_, _059371_, _059372_, _059373_, _059374_, _059375_, _059376_, _059377_, _059378_, _059379_, _059380_, _059381_, _059382_, _059383_, _059384_, _059385_, _059386_, _059387_, _059388_, _059389_, _059390_, _059391_, _059392_, _059393_, _059394_, _059395_, _059396_, _059397_, _059398_, _059399_, _059400_, _059401_, _059402_, _059403_, _059404_, _059405_, _059406_, _059407_, _059408_, _059409_, _059410_, _059411_, _059412_, _059413_, _059414_, _059415_, _059416_, _059417_, _059418_, _059419_, _059420_, _059421_, _059422_, _059423_, _059424_, _059425_, _059426_, _059427_, _059428_, _059429_, _059430_, _059431_, _059432_, _059433_, _059434_, _059435_, _059436_, _059437_, _059438_, _059439_, _059440_, _059441_, _059442_, _059443_, _059444_, _059445_, _059446_, _059447_, _059448_, _059449_, _059450_, _059451_, _059452_, _059453_, _059454_, _059455_, _059456_, _059457_, _059458_, _059459_, _059460_, _059461_, _059462_, _059463_, _059464_, _059465_, _059466_, _059467_, _059468_, _059469_, _059470_, _059471_, _059472_, _059473_, _059474_, _059475_, _059476_, _059477_, _059478_, _059479_, _059480_, _059481_, _059482_, _059483_, _059484_, _059485_, _059486_, _059487_, _059488_, _059489_, _059490_, _059491_, _059492_, _059493_, _059494_, _059495_, _059496_, _059497_, _059498_, _059499_, _059500_, _059501_, _059502_, _059503_, _059504_, _059505_, _059506_, _059507_, _059508_, _059509_, _059510_, _059511_, _059512_, _059513_, _059514_, _059515_, _059516_, _059517_, _059518_, _059519_, _059520_, _059521_, _059522_, _059523_, _059524_, _059525_, _059526_, _059527_, _059528_, _059529_, _059530_, _059531_, _059532_, _059533_, _059534_, _059535_, _059536_, _059537_, _059538_, _059539_, _059540_, _059541_, _059542_, _059543_, _059544_, _059545_, _059546_, _059547_, _059548_, _059549_, _059550_, _059551_, _059552_, _059553_, _059554_, _059555_, _059556_, _059557_, _059558_, _059559_, _059560_, _059561_, _059562_, _059563_, _059564_, _059565_, _059566_, _059567_, _059568_, _059569_, _059570_, _059571_, _059572_, _059573_, _059574_, _059575_, _059576_, _059577_, _059578_, _059579_, _059580_, _059581_, _059582_, _059583_, _059584_, _059585_, _059586_, _059587_, _059588_, _059589_, _059590_, _059591_, _059592_, _059593_, _059594_, _059595_, _059596_, _059597_, _059598_, _059599_, _059600_, _059601_, _059602_, _059603_, _059604_, _059605_, _059606_, _059607_, _059608_, _059609_, _059610_, _059611_, _059612_, _059613_, _059614_, _059615_, _059616_, _059617_, _059618_, _059619_, _059620_, _059621_, _059622_, _059623_, _059624_, _059625_, _059626_, _059627_, _059628_, _059629_, _059630_, _059631_, _059632_, _059633_, _059634_, _059635_, _059636_, _059637_, _059638_, _059639_, _059640_, _059641_, _059642_, _059643_, _059644_, _059645_, _059646_, _059647_, _059648_, _059649_, _059650_, _059651_, _059652_, _059653_, _059654_, _059655_, _059656_, _059657_, _059658_, _059659_, _059660_, _059661_, _059662_, _059663_, _059664_, _059665_, _059666_, _059667_, _059668_, _059669_, _059670_, _059671_, _059672_, _059673_, _059674_, _059675_, _059676_, _059677_, _059678_, _059679_, _059680_, _059681_, _059682_, _059683_, _059684_, _059685_, _059686_, _059687_, _059688_, _059689_, _059690_, _059691_, _059692_, _059693_, _059694_, _059695_, _059696_, _059697_, _059698_, _059699_, _059700_, _059701_, _059702_, _059703_, _059704_, _059705_, _059706_, _059707_, _059708_, _059709_, _059710_, _059711_, _059712_, _059713_, _059714_, _059715_, _059716_, _059717_, _059718_, _059719_, _059720_, _059721_, _059722_, _059723_, _059724_, _059725_, _059726_, _059727_, _059728_, _059729_, _059730_, _059731_, _059732_, _059733_, _059734_, _059735_, _059736_, _059737_, _059738_, _059739_, _059740_, _059741_, _059742_, _059743_, _059744_, _059745_, _059746_, _059747_, _059748_, _059749_, _059750_, _059751_, _059752_, _059753_, _059754_, _059755_, _059756_, _059757_, _059758_, _059759_, _059760_, _059761_, _059762_, _059763_, _059764_, _059765_, _059766_, _059767_, _059768_, _059769_, _059770_, _059771_, _059772_, _059773_, _059774_, _059775_, _059776_, _059777_, _059778_, _059779_, _059780_, _059781_, _059782_, _059783_, _059784_, _059785_, _059786_, _059787_, _059788_, _059789_, _059790_, _059791_, _059792_, _059793_, _059794_, _059795_, _059796_, _059797_, _059798_, _059799_, _059800_, _059801_, _059802_, _059803_, _059804_, _059805_, _059806_, _059807_, _059808_, _059809_, _059810_, _059811_, _059812_, _059813_, _059814_, _059815_, _059816_, _059817_, _059818_, _059819_, _059820_, _059821_, _059822_, _059823_, _059824_, _059825_, _059826_, _059827_, _059828_, _059829_, _059830_, _059831_, _059832_, _059833_, _059834_, _059835_, _059836_, _059837_, _059838_, _059839_, _059840_, _059841_, _059842_, _059843_, _059844_, _059845_, _059846_, _059847_, _059848_, _059849_, _059850_, _059851_, _059852_, _059853_, _059854_, _059855_, _059856_, _059857_, _059858_, _059859_, _059860_, _059861_, _059862_, _059863_, _059864_, _059865_, _059866_, _059867_, _059868_, _059869_, _059870_, _059871_, _059872_, _059873_, _059874_, _059875_, _059876_, _059877_, _059878_, _059879_, _059880_, _059881_, _059882_, _059883_, _059884_, _059885_, _059886_, _059887_, _059888_, _059889_, _059890_, _059891_, _059892_, _059893_, _059894_, _059895_, _059896_, _059897_, _059898_, _059899_, _059900_, _059901_, _059902_, _059903_, _059904_, _059905_, _059906_, _059907_, _059908_, _059909_, _059910_, _059911_, _059912_, _059913_, _059914_, _059915_, _059916_, _059917_, _059918_, _059919_, _059920_, _059921_, _059922_, _059923_, _059924_, _059925_, _059926_, _059927_, _059928_, _059929_, _059930_, _059931_, _059932_, _059933_, _059934_, _059935_, _059936_, _059937_, _059938_, _059939_, _059940_, _059941_, _059942_, _059943_, _059944_, _059945_, _059946_, _059947_, _059948_, _059949_, _059950_, _059951_, _059952_, _059953_, _059954_, _059955_, _059956_, _059957_, _059958_, _059959_, _059960_, _059961_, _059962_, _059963_, _059964_, _059965_, _059966_, _059967_, _059968_, _059969_, _059970_, _059971_, _059972_, _059973_, _059974_, _059975_, _059976_, _059977_, _059978_, _059979_, _059980_, _059981_, _059982_, _059983_, _059984_, _059985_, _059986_, _059987_, _059988_, _059989_, _059990_, _059991_, _059992_, _059993_, _059994_, _059995_, _059996_, _059997_, _059998_, _059999_, _060000_, _060001_, _060002_, _060003_, _060004_, _060005_, _060006_, _060007_, _060008_, _060009_, _060010_, _060011_, _060012_, _060013_, _060014_, _060015_, _060016_, _060017_, _060018_, _060019_, _060020_, _060021_, _060022_, _060023_, _060024_, _060025_, _060026_, _060027_, _060028_, _060029_, _060030_, _060031_, _060032_, _060033_, _060034_, _060035_, _060036_, _060037_, _060038_, _060039_, _060040_, _060041_, _060042_, _060043_, _060044_, _060045_, _060046_, _060047_, _060048_, _060049_, _060050_, _060051_, _060052_, _060053_, _060054_, _060055_, _060056_, _060057_, _060058_, _060059_, _060060_, _060061_, _060062_, _060063_, _060064_, _060065_, _060066_, _060067_, _060068_, _060069_, _060070_, _060071_, _060072_, _060073_, _060074_, _060075_, _060076_, _060077_, _060078_, _060079_, _060080_, _060081_, _060082_, _060083_, _060084_, _060085_, _060086_, _060087_, _060088_, _060089_, _060090_, _060091_, _060092_, _060093_, _060094_, _060095_, _060096_, _060097_, _060098_, _060099_, _060100_, _060101_, _060102_, _060103_, _060104_, _060105_, _060106_, _060107_, _060108_, _060109_, _060110_, _060111_, _060112_, _060113_, _060114_, _060115_, _060116_, _060117_, _060118_, _060119_, _060120_, _060121_, _060122_, _060123_, _060124_, _060125_, _060126_, _060127_, _060128_, _060129_, _060130_, _060131_, _060132_, _060133_, _060134_, _060135_, _060136_, _060137_, _060138_, _060139_, _060140_, _060141_, _060142_, _060143_, _060144_, _060145_, _060146_, _060147_, _060148_, _060149_, _060150_, _060151_, _060152_, _060153_, _060154_, _060155_, _060156_, _060157_, _060158_, _060159_, _060160_, _060161_, _060162_, _060163_, _060164_, _060165_, _060166_, _060167_, _060168_, _060169_, _060170_, _060171_, _060172_, _060173_, _060174_, _060175_, _060176_, _060177_, _060178_, _060179_, _060180_, _060181_, _060182_, _060183_, _060184_, _060185_, _060186_, _060187_, _060188_, _060189_, _060190_, _060191_, _060192_, _060193_, _060194_, _060195_, _060196_, _060197_, _060198_, _060199_, _060200_, _060201_, _060202_, _060203_, _060204_, _060205_, _060206_, _060207_, _060208_, _060209_, _060210_, _060211_, _060212_, _060213_, _060214_, _060215_, _060216_, _060217_, _060218_, _060219_, _060220_, _060221_, _060222_, _060223_, _060224_, _060225_, _060226_, _060227_, _060228_, _060229_, _060230_, _060231_, _060232_, _060233_, _060234_, _060235_, _060236_, _060237_, _060238_, _060239_, _060240_, _060241_, _060242_, _060243_, _060244_, _060245_, _060246_, _060247_, _060248_, _060249_, _060250_, _060251_, _060252_, _060253_, _060254_, _060255_, _060256_, _060257_, _060258_, _060259_, _060260_, _060261_, _060262_, _060263_, _060264_, _060265_, _060266_, _060267_, _060268_, _060269_, _060270_, _060271_, _060272_, _060273_, _060274_, _060275_, _060276_, _060277_, _060278_, _060279_, _060280_, _060281_, _060282_, _060283_, _060284_, _060285_, _060286_, _060287_, _060288_, _060289_, _060290_, _060291_, _060292_, _060293_, _060294_, _060295_, _060296_, _060297_, _060298_, _060299_, _060300_, _060301_, _060302_, _060303_, _060304_, _060305_, _060306_, _060307_, _060308_, _060309_, _060310_, _060311_, _060312_, _060313_, _060314_, _060315_, _060316_, _060317_, _060318_, _060319_, _060320_, _060321_, _060322_, _060323_, _060324_, _060325_, _060326_, _060327_, _060328_, _060329_, _060330_, _060331_, _060332_, _060333_, _060334_, _060335_, _060336_, _060337_, _060338_, _060339_, _060340_, _060341_, _060342_, _060343_, _060344_, _060345_, _060346_, _060347_, _060348_, _060349_, _060350_, _060351_, _060352_, _060353_, _060354_, _060355_, _060356_, _060357_, _060358_, _060359_, _060360_, _060361_, _060362_, _060363_, _060364_, _060365_, _060366_, _060367_, _060368_, _060369_, _060370_, _060371_, _060372_, _060373_, _060374_, _060375_, _060376_, _060377_, _060378_, _060379_, _060380_, _060381_, _060382_, _060383_, _060384_, _060385_, _060386_, _060387_, _060388_, _060389_, _060390_, _060391_, _060392_, _060393_, _060394_, _060395_, _060396_, _060397_, _060398_, _060399_, _060400_, _060401_, _060402_, _060403_, _060404_, _060405_, _060406_, _060407_, _060408_, _060409_, _060410_, _060411_, _060412_, _060413_, _060414_, _060415_, _060416_, _060417_, _060418_, _060419_, _060420_, _060421_, _060422_, _060423_, _060424_, _060425_, _060426_, _060427_, _060428_, _060429_, _060430_, _060431_, _060432_, _060433_, _060434_, _060435_, _060436_, _060437_, _060438_, _060439_, _060440_, _060441_, _060442_, _060443_, _060444_, _060445_, _060446_, _060447_, _060448_, _060449_, _060450_, _060451_, _060452_, _060453_, _060454_, _060455_, _060456_, _060457_, _060458_, _060459_, _060460_, _060461_, _060462_, _060463_, _060464_, _060465_, _060466_, _060467_, _060468_, _060469_, _060470_, _060471_, _060472_, _060473_, _060474_, _060475_, _060476_, _060477_, _060478_, _060479_, _060480_, _060481_, _060482_, _060483_, _060484_, _060485_, _060486_, _060487_, _060488_, _060489_, _060490_, _060491_, _060492_, _060493_, _060494_, _060495_, _060496_, _060497_, _060498_, _060499_, _060500_, _060501_, _060502_, _060503_, _060504_, _060505_, _060506_, _060507_, _060508_, _060509_, _060510_, _060511_, _060512_, _060513_, _060514_, _060515_, _060516_, _060517_, _060518_, _060519_, _060520_, _060521_, _060522_, _060523_, _060524_, _060525_, _060526_, _060527_, _060528_, _060529_, _060530_, _060531_, _060532_, _060533_, _060534_, _060535_, _060536_, _060537_, _060538_, _060539_, _060540_, _060541_, _060542_, _060543_, _060544_, _060545_, _060546_, _060547_, _060548_, _060549_, _060550_, _060551_, _060552_, _060553_, _060554_, _060555_, _060556_, _060557_, _060558_, _060559_, _060560_, _060561_, _060562_, _060563_, _060564_, _060565_, _060566_, _060567_, _060568_, _060569_, _060570_, _060571_, _060572_, _060573_, _060574_, _060575_, _060576_, _060577_, _060578_, _060579_, _060580_, _060581_, _060582_, _060583_, _060584_, _060585_, _060586_, _060587_, _060588_, _060589_, _060590_, _060591_, _060592_, _060593_, _060594_, _060595_, _060596_, _060597_, _060598_, _060599_, _060600_, _060601_, _060602_, _060603_, _060604_, _060605_, _060606_, _060607_, _060608_, _060609_, _060610_, _060611_, _060612_, _060613_, _060614_, _060615_, _060616_, _060617_, _060618_, _060619_, _060620_, _060621_, _060622_, _060623_, _060624_, _060625_, _060626_, _060627_, _060628_, _060629_, _060630_, _060631_, _060632_, _060633_, _060634_, _060635_, _060636_, _060637_, _060638_, _060639_, _060640_, _060641_, _060642_, _060643_, _060644_, _060645_, _060646_, _060647_, _060648_, _060649_, _060650_, _060651_, _060652_, _060653_, _060654_, _060655_, _060656_, _060657_, _060658_, _060659_, _060660_, _060661_, _060662_, _060663_, _060664_, _060665_, _060666_, _060667_, _060668_, _060669_, _060670_, _060671_, _060672_, _060673_, _060674_, _060675_, _060676_, _060677_, _060678_, _060679_, _060680_, _060681_, _060682_, _060683_, _060684_, _060685_, _060686_, _060687_, _060688_, _060689_, _060690_, _060691_, _060692_, _060693_, _060694_, _060695_, _060696_, _060697_, _060698_, _060699_, _060700_, _060701_, _060702_, _060703_, _060704_, _060705_, _060706_, _060707_, _060708_, _060709_, _060710_, _060711_, _060712_, _060713_, _060714_, _060715_, _060716_, _060717_, _060718_, _060719_, _060720_, _060721_, _060722_, _060723_, _060724_, _060725_, _060726_, _060727_, _060728_, _060729_, _060730_, _060731_, _060732_, _060733_, _060734_, _060735_, _060736_, _060737_, _060738_, _060739_, _060740_, _060741_, _060742_, _060743_, _060744_, _060745_, _060746_, _060747_, _060748_, _060749_, _060750_, _060751_, _060752_, _060753_, _060754_, _060755_, _060756_, _060757_, _060758_, _060759_, _060760_, _060761_, _060762_, _060763_, _060764_, _060765_, _060766_, _060767_, _060768_, _060769_, _060770_, _060771_, _060772_, _060773_, _060774_, _060775_, _060776_, _060777_, _060778_, _060779_, _060780_, _060781_, _060782_, _060783_, _060784_, _060785_, _060786_, _060787_, _060788_, _060789_, _060790_, _060791_, _060792_, _060793_, _060794_, _060795_, _060796_, _060797_, _060798_, _060799_, _060800_, _060801_, _060802_, _060803_, _060804_, _060805_, _060806_, _060807_, _060808_, _060809_, _060810_, _060811_, _060812_, _060813_, _060814_, _060815_, _060816_, _060817_, _060818_, _060819_, _060820_, _060821_, _060822_, _060823_, _060824_, _060825_, _060826_, _060827_, _060828_, _060829_, _060830_, _060831_, _060832_, _060833_, _060834_, _060835_, _060836_, _060837_, _060838_, _060839_, _060840_, _060841_, _060842_, _060843_, _060844_, _060845_, _060846_, _060847_, _060848_, _060849_, _060850_, _060851_, _060852_, _060853_, _060854_, _060855_, _060856_, _060857_, _060858_, _060859_, _060860_, _060861_, _060862_, _060863_, _060864_, _060865_, _060866_, _060867_, _060868_, _060869_, _060870_, _060871_, _060872_, _060873_, _060874_, _060875_, _060876_, _060877_, _060878_, _060879_, _060880_, _060881_, _060882_, _060883_, _060884_, _060885_, _060886_, _060887_, _060888_, _060889_, _060890_, _060891_, _060892_, _060893_, _060894_, _060895_, _060896_, _060897_, _060898_, _060899_, _060900_, _060901_, _060902_, _060903_, _060904_, _060905_, _060906_, _060907_, _060908_, _060909_, _060910_, _060911_, _060912_, _060913_, _060914_, _060915_, _060916_, _060917_, _060918_, _060919_, _060920_, _060921_, _060922_, _060923_, _060924_, _060925_, _060926_, _060927_, _060928_, _060929_, _060930_, _060931_, _060932_, _060933_, _060934_, _060935_, _060936_, _060937_, _060938_, _060939_, _060940_, _060941_, _060942_, _060943_, _060944_, _060945_, _060946_, _060947_, _060948_, _060949_, _060950_, _060951_, _060952_, _060953_, _060954_, _060955_, _060956_, _060957_, _060958_, _060959_, _060960_, _060961_, _060962_, _060963_, _060964_, _060965_, _060966_, _060967_, _060968_, _060969_, _060970_, _060971_, _060972_, _060973_, _060974_, _060975_, _060976_, _060977_, _060978_, _060979_, _060980_, _060981_, _060982_, _060983_, _060984_, _060985_, _060986_, _060987_, _060988_, _060989_, _060990_, _060991_, _060992_, _060993_, _060994_, _060995_, _060996_, _060997_, _060998_, _060999_, _061000_, _061001_, _061002_, _061003_, _061004_, _061005_, _061006_, _061007_, _061008_, _061009_, _061010_, _061011_, _061012_, _061013_, _061014_, _061015_, _061016_, _061017_, _061018_, _061019_, _061020_, _061021_, _061022_, _061023_, _061024_, _061025_, _061026_, _061027_, _061028_, _061029_, _061030_, _061031_, _061032_, _061033_, _061034_, _061035_, _061036_, _061037_, _061038_, _061039_, _061040_, _061041_, _061042_, _061043_, _061044_, _061045_, _061046_, _061047_, _061048_, _061049_, _061050_, _061051_, _061052_, _061053_, _061054_, _061055_, _061056_, _061057_, _061058_, _061059_, _061060_, _061061_, _061062_, _061063_, _061064_, _061065_, _061066_, _061067_, _061068_, _061069_, _061070_, _061071_, _061072_, _061073_, _061074_, _061075_, _061076_, _061077_, _061078_, _061079_, _061080_, _061081_, _061082_, _061083_, _061084_, _061085_, _061086_, _061087_, _061088_, _061089_, _061090_, _061091_, _061092_, _061093_, _061094_, _061095_, _061096_, _061097_, _061098_, _061099_, _061100_, _061101_, _061102_, _061103_, _061104_, _061105_, _061106_, _061107_, _061108_, _061109_, _061110_, _061111_, _061112_, _061113_, _061114_, _061115_, _061116_, _061117_, _061118_, _061119_, _061120_, _061121_, _061122_, _061123_, _061124_, _061125_, _061126_, _061127_, _061128_, _061129_, _061130_, _061131_, _061132_, _061133_, _061134_, _061135_, _061136_, _061137_, _061138_, _061139_, _061140_, _061141_, _061142_, _061143_, _061144_, _061145_, _061146_, _061147_, _061148_, _061149_, _061150_, _061151_, _061152_, _061153_, _061154_, _061155_, _061156_, _061157_, _061158_, _061159_, _061160_, _061161_, _061162_, _061163_, _061164_, _061165_, _061166_, _061167_, _061168_, _061169_, _061170_, _061171_, _061172_, _061173_, _061174_, _061175_, _061176_, _061177_, _061178_, _061179_, _061180_, _061181_, _061182_, _061183_, _061184_, _061185_, _061186_, _061187_, _061188_, _061189_, _061190_, _061191_, _061192_, _061193_, _061194_, _061195_, _061196_, _061197_, _061198_, _061199_, _061200_, _061201_, _061202_, _061203_, _061204_, _061205_, _061206_, _061207_, _061208_, _061209_, _061210_, _061211_, _061212_, _061213_, _061214_, _061215_, _061216_, _061217_, _061218_, _061219_, _061220_, _061221_, _061222_, _061223_, _061224_, _061225_, _061226_, _061227_, _061228_, _061229_, _061230_, _061231_, _061232_, _061233_, _061234_, _061235_, _061236_, _061237_, _061238_, _061239_, _061240_, _061241_, _061242_, _061243_, _061244_, _061245_, _061246_, _061247_, _061248_, _061249_, _061250_, _061251_, _061252_, _061253_, _061254_, _061255_, _061256_, _061257_, _061258_, _061259_, _061260_, _061261_, _061262_, _061263_, _061264_, _061265_, _061266_, _061267_, _061268_, _061269_, _061270_, _061271_, _061272_, _061273_, _061274_, _061275_, _061276_, _061277_, _061278_, _061279_, _061280_, _061281_, _061282_, _061283_, _061284_, _061285_, _061286_, _061287_, _061288_, _061289_, _061290_, _061291_, _061292_, _061293_, _061294_, _061295_, _061296_, _061297_, _061298_, _061299_, _061300_, _061301_, _061302_, _061303_, _061304_, _061305_, _061306_, _061307_, _061308_, _061309_, _061310_, _061311_, _061312_, _061313_, _061314_, _061315_, _061316_, _061317_, _061318_, _061319_, _061320_, _061321_, _061322_, _061323_, _061324_, _061325_, _061326_, _061327_, _061328_, _061329_, _061330_, _061331_, _061332_, _061333_, _061334_, _061335_, _061336_, _061337_, _061338_, _061339_, _061340_, _061341_, _061342_, _061343_, _061344_, _061345_, _061346_, _061347_, _061348_, _061349_, _061350_, _061351_, _061352_, _061353_, _061354_, _061355_, _061356_, _061357_, _061358_, _061359_, _061360_, _061361_, _061362_, _061363_, _061364_, _061365_, _061366_, _061367_, _061368_, _061369_, _061370_, _061371_, _061372_, _061373_, _061374_, _061375_, _061376_, _061377_, _061378_, _061379_, _061380_, _061381_, _061382_, _061383_, _061384_, _061385_, _061386_, _061387_, _061388_, _061389_, _061390_, _061391_, _061392_, _061393_, _061394_, _061395_, _061396_, _061397_, _061398_, _061399_, _061400_, _061401_, _061402_, _061403_, _061404_, _061405_, _061406_, _061407_, _061408_, _061409_, _061410_, _061411_, _061412_, _061413_, _061414_, _061415_, _061416_, _061417_, _061418_, _061419_, _061420_, _061421_, _061422_, _061423_, _061424_, _061425_, _061426_, _061427_, _061428_, _061429_, _061430_, _061431_, _061432_, _061433_, _061434_, _061435_, _061436_, _061437_, _061438_, _061439_, _061440_, _061441_, _061442_, _061443_, _061444_, _061445_, _061446_, _061447_, _061448_, _061449_, _061450_, _061451_, _061452_, _061453_, _061454_, _061455_, _061456_, _061457_, _061458_, _061459_, _061460_, _061461_, _061462_, _061463_, _061464_, _061465_, _061466_, _061467_, _061468_, _061469_, _061470_, _061471_, _061472_, _061473_, _061474_, _061475_, _061476_, _061477_, _061478_, _061479_, _061480_, _061481_, _061482_, _061483_, _061484_, _061485_, _061486_, _061487_, _061488_, _061489_, _061490_, _061491_, _061492_, _061493_, _061494_, _061495_, _061496_, _061497_, _061498_, _061499_, _061500_, _061501_, _061502_, _061503_, _061504_, _061505_, _061506_, _061507_, _061508_, _061509_, _061510_, _061511_, _061512_, _061513_, _061514_, _061515_, _061516_, _061517_, _061518_, _061519_, _061520_, _061521_, _061522_, _061523_, _061524_, _061525_, _061526_, _061527_, _061528_, _061529_, _061530_, _061531_, _061532_, _061533_, _061534_, _061535_, _061536_, _061537_, _061538_, _061539_, _061540_, _061541_, _061542_, _061543_, _061544_, _061545_, _061546_, _061547_, _061548_, _061549_, _061550_, _061551_, _061552_, _061553_, _061554_, _061555_, _061556_, _061557_, _061558_, _061559_, _061560_, _061561_, _061562_, _061563_, _061564_, _061565_, _061566_, _061567_, _061568_, _061569_, _061570_, _061571_, _061572_, _061573_, _061574_, _061575_, _061576_, _061577_, _061578_, _061579_, _061580_, _061581_, _061582_, _061583_, _061584_, _061585_, _061586_, _061587_, _061588_, _061589_, _061590_, _061591_, _061592_, _061593_, _061594_, _061595_, _061596_, _061597_, _061598_, _061599_, _061600_, _061601_, _061602_, _061603_, _061604_, _061605_, _061606_, _061607_, _061608_, _061609_, _061610_, _061611_, _061612_, _061613_, _061614_, _061615_, _061616_, _061617_, _061618_, _061619_, _061620_, _061621_, _061622_, _061623_, _061624_, _061625_, _061626_, _061627_, _061628_, _061629_, _061630_, _061631_, _061632_, _061633_, _061634_, _061635_, _061636_, _061637_, _061638_, _061639_, _061640_, _061641_, _061642_, _061643_, _061644_, _061645_, _061646_, _061647_, _061648_, _061649_, _061650_, _061651_, _061652_, _061653_, _061654_, _061655_, _061656_, _061657_, _061658_, _061659_, _061660_, _061661_, _061662_, _061663_, _061664_, _061665_, _061666_, _061667_, _061668_, _061669_, _061670_, _061671_, _061672_, _061673_, _061674_, _061675_, _061676_, _061677_, _061678_, _061679_, _061680_, _061681_, _061682_, _061683_, _061684_, _061685_, _061686_, _061687_, _061688_, _061689_, _061690_, _061691_, _061692_, _061693_, _061694_, _061695_, _061696_, _061697_, _061698_, _061699_, _061700_, _061701_, _061702_, _061703_, _061704_, _061705_, _061706_, _061707_, _061708_, _061709_, _061710_, _061711_, _061712_, _061713_, _061714_, _061715_, _061716_, _061717_, _061718_, _061719_, _061720_, _061721_, _061722_, _061723_, _061724_, _061725_, _061726_, _061727_, _061728_, _061729_, _061730_, _061731_, _061732_, _061733_, _061734_, _061735_, _061736_, _061737_, _061738_, _061739_, _061740_, _061741_, _061742_, _061743_, _061744_, _061745_, _061746_, _061747_, _061748_, _061749_, _061750_, _061751_, _061752_, _061753_, _061754_, _061755_, _061756_, _061757_, _061758_, _061759_, _061760_, _061761_, _061762_, _061763_, _061764_, _061765_, _061766_, _061767_, _061768_, _061769_, _061770_, _061771_, _061772_, _061773_, _061774_, _061775_, _061776_, _061777_, _061778_, _061779_, _061780_, _061781_, _061782_, _061783_, _061784_, _061785_, _061786_, _061787_, _061788_, _061789_, _061790_, _061791_, _061792_, _061793_, _061794_, _061795_, _061796_, _061797_, _061798_, _061799_, _061800_, _061801_, _061802_, _061803_, _061804_, _061805_, _061806_, _061807_, _061808_, _061809_, _061810_, _061811_, _061812_, _061813_, _061814_, _061815_, _061816_, _061817_, _061818_, _061819_, _061820_, _061821_, _061822_, _061823_, _061824_, _061825_, _061826_, _061827_, _061828_, _061829_, _061830_, _061831_, _061832_, _061833_, _061834_, _061835_, _061836_, _061837_, _061838_, _061839_, _061840_, _061841_, _061842_, _061843_, _061844_, _061845_, _061846_, _061847_, _061848_, _061849_, _061850_, _061851_, _061852_, _061853_, _061854_, _061855_, _061856_, _061857_, _061858_, _061859_, _061860_, _061861_, _061862_, _061863_, _061864_, _061865_, _061866_, _061867_, _061868_, _061869_, _061870_, _061871_, _061872_, _061873_, _061874_, _061875_, _061876_, _061877_, _061878_, _061879_, _061880_, _061881_, _061882_, _061883_, _061884_, _061885_, _061886_, _061887_, _061888_, _061889_, _061890_, _061891_, _061892_, _061893_, _061894_, _061895_, _061896_, _061897_, _061898_, _061899_, _061900_, _061901_, _061902_, _061903_, _061904_, _061905_, _061906_, _061907_, _061908_, _061909_, _061910_, _061911_, _061912_, _061913_, _061914_, _061915_, _061916_, _061917_, _061918_, _061919_, _061920_, _061921_, _061922_, _061923_, _061924_, _061925_, _061926_, _061927_, _061928_, _061929_, _061930_, _061931_, _061932_, _061933_, _061934_, _061935_, _061936_, _061937_, _061938_, _061939_, _061940_, _061941_, _061942_, _061943_, _061944_, _061945_, _061946_, _061947_, _061948_, _061949_, _061950_, _061951_, _061952_, _061953_, _061954_, _061955_, _061956_, _061957_, _061958_, _061959_, _061960_, _061961_, _061962_, _061963_, _061964_, _061965_, _061966_, _061967_, _061968_, _061969_, _061970_, _061971_, _061972_, _061973_, _061974_, _061975_, _061976_, _061977_, _061978_, _061979_, _061980_, _061981_, _061982_, _061983_, _061984_, _061985_, _061986_, _061987_, _061988_, _061989_, _061990_, _061991_, _061992_, _061993_, _061994_, _061995_, _061996_, _061997_, _061998_, _061999_, _062000_, _062001_, _062002_, _062003_, _062004_, _062005_, _062006_, _062007_, _062008_, _062009_, _062010_, _062011_, _062012_, _062013_, _062014_, _062015_, _062016_, _062017_, _062018_, _062019_, _062020_, _062021_, _062022_, _062023_, _062024_, _062025_, _062026_, _062027_, _062028_, _062029_, _062030_, _062031_, _062032_, _062033_, _062034_, _062035_, _062036_, _062037_, _062038_, _062039_, _062040_, _062041_, _062042_, _062043_, _062044_, _062045_, _062046_, _062047_, _062048_, _062049_, _062050_, _062051_, _062052_, _062053_, _062054_, _062055_, _062056_, _062057_, _062058_, _062059_, _062060_, _062061_, _062062_, _062063_, _062064_, _062065_, _062066_, _062067_, _062068_, _062069_, _062070_, _062071_, _062072_, _062073_, _062074_, _062075_, _062076_, _062077_, _062078_, _062079_, _062080_, _062081_, _062082_, _062083_, _062084_, _062085_, _062086_, _062087_, _062088_, _062089_, _062090_, _062091_, _062092_, _062093_, _062094_, _062095_, _062096_, _062097_, _062098_, _062099_, _062100_, _062101_, _062102_, _062103_, _062104_, _062105_, _062106_, _062107_, _062108_, _062109_, _062110_, _062111_, _062112_, _062113_, _062114_, _062115_, _062116_, _062117_, _062118_, _062119_, _062120_, _062121_, _062122_, _062123_, _062124_, _062125_, _062126_, _062127_, _062128_, _062129_, _062130_, _062131_, _062132_, _062133_, _062134_, _062135_, _062136_, _062137_, _062138_, _062139_, _062140_, _062141_, _062142_, _062143_, _062144_, _062145_, _062146_, _062147_, _062148_, _062149_, _062150_, _062151_, _062152_, _062153_, _062154_, _062155_, _062156_, _062157_, _062158_, _062159_, _062160_, _062161_, _062162_, _062163_, _062164_, _062165_, _062166_, _062167_, _062168_, _062169_, _062170_, _062171_, _062172_, _062173_, _062174_, _062175_, _062176_, _062177_, _062178_, _062179_, _062180_, _062181_, _062182_, _062183_, _062184_, _062185_, _062186_, _062187_, _062188_, _062189_, _062190_, _062191_, _062192_, _062193_, _062194_, _062195_, _062196_, _062197_, _062198_, _062199_, _062200_, _062201_, _062202_, _062203_, _062204_, _062205_, _062206_, _062207_, _062208_, _062209_, _062210_, _062211_, _062212_, _062213_, _062214_, _062215_, _062216_, _062217_, _062218_, _062219_, _062220_, _062221_, _062222_, _062223_, _062224_, _062225_, _062226_, _062227_, _062228_, _062229_, _062230_, _062231_, _062232_, _062233_, _062234_, _062235_, _062236_, _062237_, _062238_, _062239_, _062240_, _062241_, _062242_, _062243_, _062244_, _062245_, _062246_, _062247_, _062248_, _062249_, _062250_, _062251_, _062252_, _062253_, _062254_, _062255_, _062256_, _062257_, _062258_, _062259_, _062260_, _062261_, _062262_, _062263_, _062264_, _062265_, _062266_, _062267_, _062268_, _062269_, _062270_, _062271_, _062272_, _062273_, _062274_, _062275_, _062276_, _062277_, _062278_, _062279_, _062280_, _062281_, _062282_, _062283_, _062284_, _062285_, _062286_, _062287_, _062288_, _062289_, _062290_, _062291_, _062292_, _062293_, _062294_, _062295_, _062296_, _062297_, _062298_, _062299_, _062300_, _062301_, _062302_, _062303_, _062304_, _062305_, _062306_, _062307_, _062308_, _062309_, _062310_, _062311_, _062312_, _062313_, _062314_, _062315_, _062316_, _062317_, _062318_, _062319_, _062320_, _062321_, _062322_, _062323_, _062324_, _062325_, _062326_, _062327_, _062328_, _062329_, _062330_, _062331_, _062332_, _062333_, _062334_, _062335_, _062336_, _062337_, _062338_, _062339_, _062340_, _062341_, _062342_, _062343_, _062344_, _062345_, _062346_, _062347_, _062348_, _062349_, _062350_, _062351_, _062352_, _062353_, _062354_, _062355_, _062356_, _062357_, _062358_, _062359_, _062360_, _062361_, _062362_, _062363_, _062364_, _062365_, _062366_, _062367_, _062368_, _062369_, _062370_, _062371_, _062372_, _062373_, _062374_, _062375_, _062376_, _062377_, _062378_, _062379_, _062380_, _062381_, _062382_, _062383_, _062384_, _062385_, _062386_, _062387_, _062388_, _062389_, _062390_, _062391_, _062392_, _062393_, _062394_, _062395_, _062396_, _062397_, _062398_, _062399_, _062400_, _062401_, _062402_, _062403_, _062404_, _062405_, _062406_, _062407_, _062408_, _062409_, _062410_, _062411_, _062412_, _062413_, _062414_, _062415_, _062416_, _062417_, _062418_, _062419_, _062420_, _062421_, _062422_, _062423_, _062424_, _062425_, _062426_, _062427_, _062428_, _062429_, _062430_, _062431_, _062432_, _062433_, _062434_, _062435_, _062436_, _062437_, _062438_, _062439_, _062440_, _062441_, _062442_, _062443_, _062444_, _062445_, _062446_, _062447_, _062448_, _062449_, _062450_, _062451_, _062452_, _062453_, _062454_, _062455_, _062456_, _062457_, _062458_, _062459_, _062460_, _062461_, _062462_, _062463_, _062464_, _062465_, _062466_, _062467_, _062468_, _062469_, _062470_, _062471_, _062472_, _062473_, _062474_, _062475_, _062476_, _062477_, _062478_, _062479_, _062480_, _062481_, _062482_, _062483_, _062484_, _062485_, _062486_, _062487_, _062488_, _062489_, _062490_, _062491_, _062492_, _062493_, _062494_, _062495_, _062496_, _062497_, _062498_, _062499_, _062500_, _062501_, _062502_, _062503_, _062504_, _062505_, _062506_, _062507_, _062508_, _062509_, _062510_, _062511_, _062512_, _062513_, _062514_, _062515_, _062516_, _062517_, _062518_, _062519_, _062520_, _062521_, _062522_, _062523_, _062524_, _062525_, _062526_, _062527_, _062528_, _062529_, _062530_, _062531_, _062532_, _062533_, _062534_, _062535_, _062536_, _062537_, _062538_, _062539_, _062540_, _062541_, _062542_, _062543_, _062544_, _062545_, _062546_, _062547_, _062548_, _062549_, _062550_, _062551_, _062552_, _062553_, _062554_, _062555_, _062556_, _062557_, _062558_, _062559_, _062560_, _062561_, _062562_, _062563_, _062564_, _062565_, _062566_, _062567_, _062568_, _062569_, _062570_, _062571_, _062572_, _062573_, _062574_, _062575_, _062576_, _062577_, _062578_, _062579_, _062580_, _062581_, _062582_, _062583_, _062584_, _062585_, _062586_, _062587_, _062588_, _062589_, _062590_, _062591_, _062592_, _062593_, _062594_, _062595_, _062596_, _062597_, _062598_, _062599_, _062600_, _062601_, _062602_, _062603_, _062604_, _062605_, _062606_, _062607_, _062608_, _062609_, _062610_, _062611_, _062612_, _062613_, _062614_, _062615_, _062616_, _062617_, _062618_, _062619_, _062620_, _062621_, _062622_, _062623_, _062624_, _062625_, _062626_, _062627_, _062628_, _062629_, _062630_, _062631_, _062632_, _062633_, _062634_, _062635_, _062636_, _062637_, _062638_, _062639_, _062640_, _062641_, _062642_, _062643_, _062644_, _062645_, _062646_, _062647_, _062648_, _062649_, _062650_, _062651_, _062652_, _062653_, _062654_, _062655_, _062656_, _062657_, _062658_, _062659_, _062660_, _062661_, _062662_, _062663_, _062664_, _062665_, _062666_, _062667_, _062668_, _062669_, _062670_, _062671_, _062672_, _062673_, _062674_, _062675_, _062676_, _062677_, _062678_, _062679_, _062680_, _062681_, _062682_, _062683_, _062684_, _062685_, _062686_, _062687_, _062688_, _062689_, _062690_, _062691_, _062692_, _062693_, _062694_, _062695_, _062696_, _062697_, _062698_, _062699_, _062700_, _062701_, _062702_, _062703_, _062704_, _062705_, _062706_, _062707_, _062708_, _062709_, _062710_, _062711_, _062712_, _062713_, _062714_, _062715_, _062716_, _062717_, _062718_, _062719_, _062720_, _062721_, _062722_, _062723_, _062724_, _062725_, _062726_, _062727_, _062728_, _062729_, _062730_, _062731_, _062732_, _062733_, _062734_, _062735_, _062736_, _062737_, _062738_, _062739_, _062740_, _062741_, _062742_, _062743_, _062744_, _062745_, _062746_, _062747_, _062748_, _062749_, _062750_, _062751_, _062752_, _062753_, _062754_, _062755_, _062756_, _062757_, _062758_, _062759_, _062760_, _062761_, _062762_, _062763_, _062764_, _062765_, _062766_, _062767_, _062768_, _062769_, _062770_, _062771_, _062772_, _062773_, _062774_, _062775_, _062776_, _062777_, _062778_, _062779_, _062780_, _062781_, _062782_, _062783_, _062784_, _062785_, _062786_, _062787_, _062788_, _062789_, _062790_, _062791_, _062792_, _062793_, _062794_, _062795_, _062796_, _062797_, _062798_, _062799_, _062800_, _062801_, _062802_, _062803_, _062804_, _062805_, _062806_, _062807_, _062808_, _062809_, _062810_, _062811_, _062812_, _062813_, _062814_, _062815_, _062816_, _062817_, _062818_, _062819_, _062820_, _062821_, _062822_, _062823_, _062824_, _062825_, _062826_, _062827_, _062828_, _062829_, _062830_, _062831_, _062832_, _062833_, _062834_, _062835_, _062836_, _062837_, _062838_, _062839_, _062840_, _062841_, _062842_, _062843_, _062844_, _062845_, _062846_, _062847_, _062848_, _062849_, _062850_, _062851_, _062852_, _062853_, _062854_, _062855_, _062856_, _062857_, _062858_, _062859_, _062860_, _062861_, _062862_, _062863_, _062864_, _062865_, _062866_, _062867_, _062868_, _062869_, _062870_, _062871_, _062872_, _062873_, _062874_, _062875_, _062876_, _062877_, _062878_, _062879_, _062880_, _062881_, _062882_, _062883_, _062884_, _062885_, _062886_, _062887_, _062888_, _062889_, _062890_, _062891_, _062892_, _062893_, _062894_, _062895_, _062896_, _062897_, _062898_, _062899_, _062900_, _062901_, _062902_, _062903_, _062904_, _062905_, _062906_, _062907_, _062908_, _062909_, _062910_, _062911_, _062912_, _062913_, _062914_, _062915_, _062916_, _062917_, _062918_, _062919_, _062920_, _062921_, _062922_, _062923_, _062924_, _062925_, _062926_, _062927_, _062928_, _062929_, _062930_, _062931_, _062932_, _062933_, _062934_, _062935_, _062936_, _062937_, _062938_, _062939_, _062940_, _062941_, _062942_, _062943_, _062944_, _062945_, _062946_, _062947_, _062948_, _062949_, _062950_, _062951_, _062952_, _062953_, _062954_, _062955_, _062956_, _062957_, _062958_, _062959_, _062960_, _062961_, _062962_, _062963_, _062964_, _062965_, _062966_, _062967_, _062968_, _062969_, _062970_, _062971_, _062972_, _062973_, _062974_, _062975_, _062976_, _062977_, _062978_, _062979_, _062980_, _062981_, _062982_, _062983_, _062984_, _062985_, _062986_, _062987_, _062988_, _062989_, _062990_, _062991_, _062992_, _062993_, _062994_, _062995_, _062996_, _062997_, _062998_, _062999_, _063000_, _063001_, _063002_, _063003_, _063004_, _063005_, _063006_, _063007_, _063008_, _063009_, _063010_, _063011_, _063012_, _063013_, _063014_, _063015_, _063016_, _063017_, _063018_, _063019_, _063020_, _063021_, _063022_, _063023_, _063024_, _063025_, _063026_, _063027_, _063028_, _063029_, _063030_, _063031_, _063032_, _063033_, _063034_, _063035_, _063036_, _063037_, _063038_, _063039_, _063040_, _063041_, _063042_, _063043_, _063044_, _063045_, _063046_, _063047_, _063048_, _063049_, _063050_, _063051_, _063052_, _063053_, _063054_, _063055_, _063056_, _063057_, _063058_, _063059_, _063060_, _063061_, _063062_, _063063_, _063064_, _063065_, _063066_, _063067_, _063068_, _063069_, _063070_, _063071_, _063072_, _063073_, _063074_, _063075_, _063076_, _063077_, _063078_, _063079_, _063080_, _063081_, _063082_, _063083_, _063084_, _063085_, _063086_, _063087_, _063088_, _063089_, _063090_, _063091_, _063092_, _063093_, _063094_, _063095_, _063096_, _063097_, _063098_, _063099_, _063100_, _063101_, _063102_, _063103_, _063104_, _063105_, _063106_, _063107_, _063108_, _063109_, _063110_, _063111_, _063112_, _063113_, _063114_, _063115_, _063116_, _063117_, _063118_, _063119_, _063120_, _063121_, _063122_, _063123_, _063124_, _063125_, _063126_, _063127_, _063128_, _063129_, _063130_, _063131_, _063132_, _063133_, _063134_, _063135_, _063136_, _063137_, _063138_, _063139_, _063140_, _063141_, _063142_, _063143_, _063144_, _063145_, _063146_, _063147_, _063148_, _063149_, _063150_, _063151_, _063152_, _063153_, _063154_, _063155_, _063156_, _063157_, _063158_, _063159_, _063160_, _063161_, _063162_, _063163_, _063164_, _063165_, _063166_, _063167_, _063168_, _063169_, _063170_, _063171_, _063172_, _063173_, _063174_, _063175_, _063176_, _063177_, _063178_, _063179_, _063180_, _063181_, _063182_, _063183_, _063184_, _063185_, _063186_, _063187_, _063188_, _063189_, _063190_, _063191_, _063192_, _063193_, _063194_, _063195_, _063196_, _063197_, _063198_, _063199_, _063200_, _063201_, _063202_, _063203_, _063204_, _063205_, _063206_, _063207_, _063208_, _063209_, _063210_, _063211_, _063212_, _063213_, _063214_, _063215_, _063216_, _063217_, _063218_, _063219_, _063220_, _063221_, _063222_, _063223_, _063224_, _063225_, _063226_, _063227_, _063228_, _063229_, _063230_, _063231_, _063232_, _063233_, _063234_, _063235_, _063236_, _063237_, _063238_, _063239_, _063240_, _063241_, _063242_, _063243_, _063244_, _063245_, _063246_, _063247_, _063248_, _063249_, _063250_, _063251_, _063252_, _063253_, _063254_, _063255_, _063256_, _063257_, _063258_, _063259_, _063260_, _063261_, _063262_, _063263_, _063264_, _063265_, _063266_, _063267_, _063268_, _063269_, _063270_, _063271_, _063272_, _063273_, _063274_, _063275_, _063276_, _063277_, _063278_, _063279_, _063280_, _063281_, _063282_, _063283_, _063284_, _063285_, _063286_, _063287_, _063288_, _063289_, _063290_, _063291_, _063292_, _063293_, _063294_, _063295_, _063296_, _063297_, _063298_, _063299_, _063300_, _063301_, _063302_, _063303_, _063304_, _063305_, _063306_, _063307_, _063308_, _063309_, _063310_, _063311_, _063312_, _063313_, _063314_, _063315_, _063316_, _063317_, _063318_, _063319_, _063320_, _063321_, _063322_, _063323_, _063324_, _063325_, _063326_, _063327_, _063328_, _063329_, _063330_, _063331_, _063332_, _063333_, _063334_, _063335_, _063336_, _063337_, _063338_, _063339_, _063340_, _063341_, _063342_, _063343_, _063344_, _063345_, _063346_, _063347_, _063348_, _063349_, _063350_, _063351_, _063352_, _063353_, _063354_, _063355_, _063356_, _063357_, _063358_, _063359_, _063360_, _063361_, _063362_, _063363_, _063364_, _063365_, _063366_, _063367_, _063368_, _063369_, _063370_, _063371_, _063372_, _063373_, _063374_, _063375_, _063376_, _063377_, _063378_, _063379_, _063380_, _063381_, _063382_, _063383_, _063384_, _063385_, _063386_, _063387_, _063388_, _063389_, _063390_, _063391_, _063392_, _063393_, _063394_, _063395_, _063396_, _063397_, _063398_, _063399_, _063400_, _063401_, _063402_, _063403_, _063404_, _063405_, _063406_, _063407_, _063408_, _063409_, _063410_, _063411_, _063412_, _063413_, _063414_, _063415_, _063416_, _063417_, _063418_, _063419_, _063420_, _063421_, _063422_, _063423_, _063424_, _063425_, _063426_, _063427_, _063428_, _063429_, _063430_, _063431_, _063432_, _063433_, _063434_, _063435_, _063436_, _063437_, _063438_, _063439_, _063440_, _063441_, _063442_, _063443_, _063444_, _063445_, _063446_, _063447_, _063448_, _063449_, _063450_, _063451_, _063452_, _063453_, _063454_, _063455_, _063456_, _063457_, _063458_, _063459_, _063460_, _063461_, _063462_, _063463_, _063464_, _063465_, _063466_, _063467_, _063468_, _063469_, _063470_, _063471_, _063472_, _063473_, _063474_, _063475_, _063476_, _063477_, _063478_, _063479_, _063480_, _063481_, _063482_, _063483_, _063484_, _063485_, _063486_, _063487_, _063488_, _063489_, _063490_, _063491_, _063492_, _063493_, _063494_, _063495_, _063496_, _063497_, _063498_, _063499_, _063500_, _063501_, _063502_, _063503_, _063504_, _063505_, _063506_, _063507_, _063508_, _063509_, _063510_, _063511_, _063512_, _063513_, _063514_, _063515_, _063516_, _063517_, _063518_, _063519_, _063520_, _063521_, _063522_, _063523_, _063524_, _063525_, _063526_, _063527_, _063528_, _063529_, _063530_, _063531_, _063532_, _063533_, _063534_, _063535_, _063536_, _063537_, _063538_, _063539_, _063540_, _063541_, _063542_, _063543_, _063544_, _063545_, _063546_, _063547_, _063548_, _063549_, _063550_, _063551_, _063552_, _063553_, _063554_, _063555_, _063556_, _063557_, _063558_, _063559_, _063560_, _063561_, _063562_, _063563_, _063564_, _063565_, _063566_, _063567_, _063568_, _063569_, _063570_, _063571_, _063572_, _063573_, _063574_, _063575_, _063576_, _063577_, _063578_, _063579_, _063580_, _063581_, _063582_, _063583_, _063584_, _063585_, _063586_, _063587_, _063588_, _063589_, _063590_, _063591_, _063592_, _063593_, _063594_, _063595_, _063596_, _063597_, _063598_, _063599_, _063600_, _063601_, _063602_, _063603_, _063604_, _063605_, _063606_, _063607_, _063608_, _063609_, _063610_, _063611_, _063612_, _063613_, _063614_, _063615_, _063616_, _063617_, _063618_, _063619_, _063620_, _063621_, _063622_, _063623_, _063624_, _063625_, _063626_, _063627_, _063628_, _063629_, _063630_, _063631_, _063632_, _063633_, _063634_, _063635_, _063636_, _063637_, _063638_, _063639_, _063640_, _063641_, _063642_, _063643_, _063644_, _063645_, _063646_, _063647_, _063648_, _063649_, _063650_, _063651_, _063652_, _063653_, _063654_, _063655_, _063656_, _063657_, _063658_, _063659_, _063660_, _063661_, _063662_, _063663_, _063664_, _063665_, _063666_, _063667_, _063668_, _063669_, _063670_, _063671_, _063672_, _063673_, _063674_, _063675_, _063676_, _063677_, _063678_, _063679_, _063680_, _063681_, _063682_, _063683_, _063684_, _063685_, _063686_, _063687_, _063688_, _063689_, _063690_, _063691_, _063692_, _063693_, _063694_, _063695_, _063696_, _063697_, _063698_, _063699_, _063700_, _063701_, _063702_, _063703_, _063704_, _063705_, _063706_, _063707_, _063708_, _063709_, _063710_, _063711_, _063712_, _063713_, _063714_, _063715_, _063716_, _063717_, _063718_, _063719_, _063720_, _063721_, _063722_, _063723_, _063724_, _063725_, _063726_, _063727_, _063728_, _063729_, _063730_, _063731_, _063732_, _063733_, _063734_, _063735_, _063736_, _063737_, _063738_, _063739_, _063740_, _063741_, _063742_, _063743_, _063744_, _063745_, _063746_, _063747_, _063748_, _063749_, _063750_, _063751_, _063752_, _063753_, _063754_, _063755_, _063756_, _063757_, _063758_, _063759_, _063760_, _063761_, _063762_, _063763_, _063764_, _063765_, _063766_, _063767_, _063768_, _063769_, _063770_, _063771_, _063772_, _063773_, _063774_, _063775_, _063776_, _063777_, _063778_, _063779_, _063780_, _063781_, _063782_, _063783_, _063784_, _063785_, _063786_, _063787_, _063788_, _063789_, _063790_, _063791_, _063792_, _063793_, _063794_, _063795_, _063796_, _063797_, _063798_, _063799_, _063800_, _063801_, _063802_, _063803_, _063804_, _063805_, _063806_, _063807_, _063808_, _063809_, _063810_, _063811_, _063812_, _063813_, _063814_, _063815_, _063816_, _063817_, _063818_, _063819_, _063820_, _063821_, _063822_, _063823_, _063824_, _063825_, _063826_, _063827_, _063828_, _063829_, _063830_, _063831_, _063832_, _063833_, _063834_, _063835_, _063836_, _063837_, _063838_, _063839_, _063840_, _063841_, _063842_, _063843_, _063844_, _063845_, _063846_, _063847_, _063848_, _063849_, _063850_, _063851_, _063852_, _063853_, _063854_, _063855_, _063856_, _063857_, _063858_, _063859_, _063860_, _063861_, _063862_, _063863_, _063864_, _063865_, _063866_, _063867_, _063868_, _063869_, _063870_, _063871_, _063872_, _063873_, _063874_, _063875_, _063876_, _063877_, _063878_, _063879_, _063880_, _063881_, _063882_, _063883_, _063884_, _063885_, _063886_, _063887_, _063888_, _063889_, _063890_, _063891_, _063892_, _063893_, _063894_, _063895_, _063896_, _063897_, _063898_, _063899_, _063900_, _063901_, _063902_, _063903_, _063904_, _063905_, _063906_, _063907_, _063908_, _063909_, _063910_, _063911_, _063912_, _063913_, _063914_, _063915_, _063916_, _063917_, _063918_, _063919_, _063920_, _063921_, _063922_, _063923_, _063924_, _063925_, _063926_, _063927_, _063928_, _063929_, _063930_, _063931_, _063932_, _063933_, _063934_, _063935_, _063936_, _063937_, _063938_, _063939_, _063940_, _063941_, _063942_, _063943_, _063944_, _063945_, _063946_, _063947_, _063948_, _063949_, _063950_, _063951_, _063952_, _063953_, _063954_, _063955_, _063956_, _063957_, _063958_, _063959_, _063960_, _063961_, _063962_, _063963_, _063964_, _063965_, _063966_, _063967_, _063968_, _063969_, _063970_, _063971_, _063972_, _063973_, _063974_, _063975_, _063976_, _063977_, _063978_, _063979_, _063980_, _063981_, _063982_, _063983_, _063984_, _063985_, _063986_, _063987_, _063988_, _063989_, _063990_, _063991_, _063992_, _063993_, _063994_, _063995_, _063996_, _063997_, _063998_, _063999_, _064000_, _064001_, _064002_, _064003_, _064004_, _064005_, _064006_, _064007_, _064008_, _064009_, _064010_, _064011_, _064012_, _064013_, _064014_, _064015_, _064016_, _064017_, _064018_, _064019_, _064020_, _064021_, _064022_, _064023_, _064024_, _064025_, _064026_, _064027_, _064028_, _064029_, _064030_, _064031_, _064032_, _064033_, _064034_, _064035_, _064036_, _064037_, _064038_, _064039_, _064040_, _064041_, _064042_, _064043_, _064044_, _064045_, _064046_, _064047_, _064048_, _064049_, _064050_, _064051_, _064052_, _064053_, _064054_, _064055_, _064056_, _064057_, _064058_, _064059_, _064060_, _064061_, _064062_, _064063_, _064064_, _064065_, _064066_, _064067_, _064068_, _064069_, _064070_, _064071_, _064072_, _064073_, _064074_, _064075_, _064076_, _064077_, _064078_, _064079_, _064080_, _064081_, _064082_, _064083_, _064084_, _064085_, _064086_, _064087_, _064088_, _064089_, _064090_, _064091_, _064092_, _064093_, _064094_, _064095_, _064096_, _064097_, _064098_, _064099_, _064100_, _064101_, _064102_, _064103_, _064104_, _064105_, _064106_, _064107_, _064108_, _064109_, _064110_, _064111_, _064112_, _064113_, _064114_, _064115_, _064116_, _064117_, _064118_, _064119_, _064120_, _064121_, _064122_, _064123_, _064124_, _064125_, _064126_, _064127_, _064128_, _064129_, _064130_, _064131_, _064132_, _064133_, _064134_, _064135_, _064136_, _064137_, _064138_, _064139_, _064140_, _064141_, _064142_, _064143_, _064144_, _064145_, _064146_, _064147_, _064148_, _064149_, _064150_, _064151_, _064152_, _064153_, _064154_, _064155_, _064156_, _064157_, _064158_, _064159_, _064160_, _064161_, _064162_, _064163_, _064164_, _064165_, _064166_, _064167_, _064168_, _064169_, _064170_, _064171_, _064172_, _064173_, _064174_, _064175_, _064176_, _064177_, _064178_, _064179_, _064180_, _064181_, _064182_, _064183_, _064184_, _064185_, _064186_, _064187_, _064188_, _064189_, _064190_, _064191_, _064192_, _064193_, _064194_, _064195_, _064196_, _064197_, _064198_, _064199_, _064200_, _064201_, _064202_, _064203_, _064204_, _064205_, _064206_, _064207_, _064208_, _064209_, _064210_, _064211_, _064212_, _064213_, _064214_, _064215_, _064216_, _064217_, _064218_, _064219_, _064220_, _064221_, _064222_, _064223_, _064224_, _064225_, _064226_, _064227_, _064228_, _064229_, _064230_, _064231_, _064232_, _064233_, _064234_, _064235_, _064236_, _064237_, _064238_, _064239_, _064240_, _064241_, _064242_, _064243_, _064244_, _064245_, _064246_, _064247_, _064248_, _064249_, _064250_, _064251_, _064252_, _064253_, _064254_, _064255_, _064256_, _064257_, _064258_, _064259_, _064260_, _064261_, _064262_, _064263_, _064264_, _064265_, _064266_, _064267_, _064268_, _064269_, _064270_, _064271_, _064272_, _064273_, _064274_, _064275_, _064276_, _064277_, _064278_, _064279_, _064280_, _064281_, _064282_, _064283_, _064284_, _064285_, _064286_, _064287_, _064288_, _064289_, _064290_, _064291_, _064292_, _064293_, _064294_, _064295_, _064296_, _064297_, _064298_, _064299_, _064300_, _064301_, _064302_, _064303_, _064304_, _064305_, _064306_, _064307_, _064308_, _064309_, _064310_, _064311_, _064312_, _064313_, _064314_, _064315_, _064316_, _064317_, _064318_, _064319_, _064320_, _064321_, _064322_, _064323_, _064324_, _064325_, _064326_, _064327_, _064328_, _064329_, _064330_, _064331_, _064332_, _064333_, _064334_, _064335_, _064336_, _064337_, _064338_, _064339_, _064340_, _064341_, _064342_, _064343_, _064344_, _064345_, _064346_, _064347_, _064348_, _064349_, _064350_, _064351_, _064352_, _064353_, _064354_, _064355_, _064356_, _064357_, _064358_, _064359_, _064360_, _064361_, _064362_, _064363_, _064364_, _064365_, _064366_, _064367_, _064368_, _064369_, _064370_, _064371_, _064372_, _064373_, _064374_, _064375_, _064376_, _064377_, _064378_, _064379_, _064380_, _064381_, _064382_, _064383_, _064384_, _064385_, _064386_, _064387_, _064388_, _064389_, _064390_, _064391_, _064392_, _064393_, _064394_, _064395_, _064396_, _064397_, _064398_, _064399_, _064400_, _064401_, _064402_, _064403_, _064404_, _064405_, _064406_, _064407_, _064408_, _064409_, _064410_, _064411_, _064412_, _064413_, _064414_, _064415_, _064416_, _064417_, _064418_, _064419_, _064420_, _064421_, _064422_, _064423_, _064424_, _064425_, _064426_, _064427_, _064428_, _064429_, _064430_, _064431_, _064432_, _064433_, _064434_, _064435_, _064436_, _064437_, _064438_, _064439_, _064440_, _064441_, _064442_, _064443_, _064444_, _064445_, _064446_, _064447_, _064448_, _064449_, _064450_, _064451_, _064452_, _064453_, _064454_, _064455_, _064456_, _064457_, _064458_, _064459_, _064460_, _064461_, _064462_, _064463_, _064464_, _064465_, _064466_, _064467_, _064468_, _064469_, _064470_, _064471_, _064472_, _064473_, _064474_, _064475_, _064476_, _064477_, _064478_, _064479_, _064480_, _064481_, _064482_, _064483_, _064484_, _064485_, _064486_, _064487_, _064488_, _064489_, _064490_, _064491_, _064492_, _064493_, _064494_, _064495_, _064496_, _064497_, _064498_, _064499_, _064500_, _064501_, _064502_, _064503_, _064504_, _064505_, _064506_, _064507_, _064508_, _064509_, _064510_, _064511_, _064512_, _064513_, _064514_, _064515_, _064516_, _064517_, _064518_, _064519_, _064520_, _064521_, _064522_, _064523_, _064524_, _064525_, _064526_, _064527_, _064528_, _064529_, _064530_, _064531_, _064532_, _064533_, _064534_, _064535_, _064536_, _064537_, _064538_, _064539_, _064540_, _064541_, _064542_, _064543_, _064544_, _064545_, _064546_, _064547_, _064548_, _064549_, _064550_, _064551_, _064552_, _064553_, _064554_, _064555_, _064556_, _064557_, _064558_, _064559_, _064560_, _064561_, _064562_, _064563_, _064564_, _064565_, _064566_, _064567_, _064568_, _064569_, _064570_, _064571_, _064572_, _064573_, _064574_, _064575_, _064576_, _064577_, _064578_, _064579_, _064580_, _064581_, _064582_, _064583_, _064584_, _064585_, _064586_, _064587_, _064588_, _064589_, _064590_, _064591_, _064592_, _064593_, _064594_, _064595_, _064596_, _064597_, _064598_, _064599_, _064600_, _064601_, _064602_, _064603_, _064604_, _064605_, _064606_, _064607_, _064608_, _064609_, _064610_, _064611_, _064612_, _064613_, _064614_, _064615_, _064616_, _064617_, _064618_, _064619_, _064620_, _064621_, _064622_, _064623_, _064624_, _064625_, _064626_, _064627_, _064628_, _064629_, _064630_, _064631_, _064632_, _064633_, _064634_, _064635_, _064636_, _064637_, _064638_, _064639_, _064640_, _064641_, _064642_, _064643_, _064644_, _064645_, _064646_, _064647_, _064648_, _064649_, _064650_, _064651_, _064652_, _064653_, _064654_, _064655_, _064656_, _064657_, _064658_, _064659_, _064660_, _064661_, _064662_, _064663_, _064664_, _064665_, _064666_, _064667_, _064668_, _064669_, _064670_, _064671_, _064672_, _064673_, _064674_, _064675_, _064676_, _064677_, _064678_, _064679_, _064680_, _064681_, _064682_, _064683_, _064684_, _064685_, _064686_, _064687_, _064688_, _064689_, _064690_, _064691_, _064692_, _064693_, _064694_, _064695_, _064696_, _064697_, _064698_, _064699_, _064700_, _064701_, _064702_, _064703_, _064704_, _064705_, _064706_, _064707_, _064708_, _064709_, _064710_, _064711_, _064712_, _064713_, _064714_, _064715_, _064716_, _064717_, _064718_, _064719_, _064720_, _064721_, _064722_, _064723_, _064724_, _064725_, _064726_, _064727_, _064728_, _064729_, _064730_, _064731_, _064732_, _064733_, _064734_, _064735_, _064736_, _064737_, _064738_, _064739_, _064740_, _064741_, _064742_, _064743_, _064744_, _064745_, _064746_, _064747_, _064748_, _064749_, _064750_, _064751_, _064752_, _064753_, _064754_, _064755_, _064756_, _064757_, _064758_, _064759_, _064760_, _064761_, _064762_, _064763_, _064764_, _064765_, _064766_, _064767_, _064768_, _064769_, _064770_, _064771_, _064772_, _064773_, _064774_, _064775_, _064776_, _064777_, _064778_, _064779_, _064780_, _064781_, _064782_, _064783_, _064784_, _064785_, _064786_, _064787_, _064788_, _064789_, _064790_, _064791_, _064792_, _064793_, _064794_, _064795_, _064796_, _064797_, _064798_, _064799_, _064800_, _064801_, _064802_, _064803_, _064804_, _064805_, _064806_, _064807_, _064808_, _064809_, _064810_, _064811_, _064812_, _064813_, _064814_, _064815_, _064816_, _064817_, _064818_, _064819_, _064820_, _064821_, _064822_, _064823_, _064824_, _064825_, _064826_, _064827_, _064828_, _064829_, _064830_, _064831_, _064832_, _064833_, _064834_, _064835_, _064836_, _064837_, _064838_, _064839_, _064840_, _064841_, _064842_, _064843_, _064844_, _064845_, _064846_, _064847_, _064848_, _064849_, _064850_, _064851_, _064852_, _064853_, _064854_, _064855_, _064856_, _064857_, _064858_, _064859_, _064860_, _064861_, _064862_, _064863_, _064864_, _064865_, _064866_, _064867_, _064868_, _064869_, _064870_, _064871_, _064872_, _064873_, _064874_, _064875_, _064876_, _064877_, _064878_, _064879_, _064880_, _064881_, _064882_, _064883_, _064884_, _064885_, _064886_, _064887_, _064888_, _064889_, _064890_, _064891_, _064892_, _064893_, _064894_, _064895_, _064896_, _064897_, _064898_, _064899_, _064900_, _064901_, _064902_, _064903_, _064904_, _064905_, _064906_, _064907_, _064908_, _064909_, _064910_, _064911_, _064912_, _064913_, _064914_, _064915_, _064916_, _064917_, _064918_, _064919_, _064920_, _064921_, _064922_, _064923_, _064924_, _064925_, _064926_, _064927_, _064928_, _064929_, _064930_, _064931_, _064932_, _064933_, _064934_, _064935_, _064936_, _064937_, _064938_, _064939_, _064940_, _064941_, _064942_, _064943_, _064944_, _064945_, _064946_, _064947_, _064948_, _064949_, _064950_, _064951_, _064952_, _064953_, _064954_, _064955_, _064956_, _064957_, _064958_, _064959_, _064960_, _064961_, _064962_, _064963_, _064964_, _064965_, _064966_, _064967_, _064968_, _064969_, _064970_, _064971_, _064972_, _064973_, _064974_, _064975_, _064976_, _064977_, _064978_, _064979_, _064980_, _064981_, _064982_, _064983_, _064984_, _064985_, _064986_, _064987_, _064988_, _064989_, _064990_, _064991_, _064992_, _064993_, _064994_, _064995_, _064996_, _064997_, _064998_, _064999_, _065000_, _065001_, _065002_, _065003_, _065004_, _065005_, _065006_, _065007_, _065008_, _065009_, _065010_, _065011_, _065012_, _065013_, _065014_, _065015_, _065016_, _065017_, _065018_, _065019_, _065020_, _065021_, _065022_, _065023_, _065024_, _065025_, _065026_, _065027_, _065028_, _065029_, _065030_, _065031_, _065032_, _065033_, _065034_, _065035_, _065036_, _065037_, _065038_, _065039_, _065040_, _065041_, _065042_, _065043_, _065044_, _065045_, _065046_, _065047_, _065048_, _065049_, _065050_, _065051_, _065052_, _065053_, _065054_, _065055_, _065056_, _065057_, _065058_, _065059_, _065060_, _065061_, _065062_, _065063_, _065064_, _065065_, _065066_, _065067_, _065068_, _065069_, _065070_, _065071_, _065072_, _065073_, _065074_, _065075_, _065076_, _065077_, _065078_, _065079_, _065080_, _065081_, _065082_, _065083_, _065084_, _065085_, _065086_, _065087_, _065088_, _065089_, _065090_, _065091_, _065092_, _065093_, _065094_, _065095_, _065096_, _065097_, _065098_, _065099_, _065100_, _065101_, _065102_, _065103_, _065104_, _065105_, _065106_, _065107_, _065108_, _065109_, _065110_, _065111_, _065112_, _065113_, _065114_, _065115_, _065116_, _065117_, _065118_, _065119_, _065120_, _065121_, _065122_, _065123_, _065124_, _065125_, _065126_, _065127_, _065128_, _065129_, _065130_, _065131_, _065132_, _065133_, _065134_, _065135_, _065136_, _065137_, _065138_, _065139_, _065140_, _065141_, _065142_, _065143_, _065144_, _065145_, _065146_, _065147_, _065148_, _065149_, _065150_, _065151_, _065152_, _065153_, _065154_, _065155_, _065156_, _065157_, _065158_, _065159_, _065160_, _065161_, _065162_, _065163_, _065164_, _065165_, _065166_, _065167_, _065168_, _065169_, _065170_, _065171_, _065172_, _065173_, _065174_, _065175_, _065176_, _065177_, _065178_, _065179_, _065180_, _065181_, _065182_, _065183_, _065184_, _065185_, _065186_, _065187_, _065188_, _065189_, _065190_, _065191_, _065192_, _065193_, _065194_, _065195_, _065196_, _065197_, _065198_, _065199_, _065200_, _065201_, _065202_, _065203_, _065204_, _065205_, _065206_, _065207_, _065208_, _065209_, _065210_, _065211_, _065212_, _065213_, _065214_, _065215_, _065216_, _065217_, _065218_, _065219_, _065220_, _065221_, _065222_, _065223_, _065224_, _065225_, _065226_, _065227_, _065228_, _065229_, _065230_, _065231_, _065232_, _065233_, _065234_, _065235_, _065236_, _065237_, _065238_, _065239_, _065240_, _065241_, _065242_, _065243_, _065244_, _065245_, _065246_, _065247_, _065248_, _065249_, _065250_, _065251_, _065252_, _065253_, _065254_, _065255_, _065256_, _065257_, _065258_, _065259_, _065260_, _065261_, _065262_, _065263_, _065264_, _065265_, _065266_, _065267_, _065268_, _065269_, _065270_, _065271_, _065272_, _065273_, _065274_, _065275_, _065276_, _065277_, _065278_, _065279_, _065280_, _065281_, _065282_, _065283_, _065284_, _065285_, _065286_, _065287_, _065288_, _065289_, _065290_, _065291_, _065292_, _065293_, _065294_, _065295_, _065296_, _065297_, _065298_, _065299_, _065300_, _065301_, _065302_, _065303_, _065304_, _065305_, _065306_, _065307_, _065308_, _065309_, _065310_, _065311_, _065312_, _065313_, _065314_, _065315_, _065316_, _065317_, _065318_, _065319_, _065320_, _065321_, _065322_, _065323_, _065324_, _065325_, _065326_, _065327_, _065328_, _065329_, _065330_, _065331_, _065332_, _065333_, _065334_, _065335_, _065336_, _065337_, _065338_, _065339_, _065340_, _065341_, _065342_, _065343_, _065344_, _065345_, _065346_, _065347_, _065348_, _065349_, _065350_, _065351_, _065352_, _065353_, _065354_, _065355_, _065356_, _065357_, _065358_, _065359_, _065360_, _065361_, _065362_, _065363_, _065364_, _065365_, _065366_, _065367_, _065368_, _065369_, _065370_, _065371_, _065372_, _065373_, _065374_, _065375_, _065376_, _065377_, _065378_, _065379_, _065380_, _065381_, _065382_, _065383_, _065384_, _065385_, _065386_, _065387_, _065388_, _065389_, _065390_, _065391_, _065392_, _065393_, _065394_, _065395_, _065396_, _065397_, _065398_, _065399_, _065400_, _065401_, _065402_, _065403_, _065404_, _065405_, _065406_, _065407_, _065408_, _065409_, _065410_, _065411_, _065412_, _065413_, _065414_, _065415_, _065416_, _065417_, _065418_, _065419_, _065420_, _065421_, _065422_, _065423_, _065424_, _065425_, _065426_, _065427_, _065428_, _065429_, _065430_, _065431_, _065432_, _065433_, _065434_, _065435_, _065436_, _065437_, _065438_, _065439_, _065440_, _065441_, _065442_, _065443_, _065444_, _065445_, _065446_, _065447_, _065448_, _065449_, _065450_, _065451_, _065452_, _065453_, _065454_, _065455_, _065456_, _065457_, _065458_, _065459_, _065460_, _065461_, _065462_, _065463_, _065464_, _065465_, _065466_, _065467_, _065468_, _065469_, _065470_, _065471_, _065472_, _065473_, _065474_, _065475_, _065476_, _065477_, _065478_, _065479_, _065480_, _065481_, _065482_, _065483_, _065484_, _065485_, _065486_, _065487_, _065488_, _065489_, _065490_, _065491_, _065492_, _065493_, _065494_, _065495_, _065496_, _065497_, _065498_, _065499_, _065500_, _065501_, _065502_, _065503_, _065504_, _065505_, _065506_, _065507_, _065508_, _065509_, _065510_, _065511_, _065512_, _065513_, _065514_, _065515_, _065516_, _065517_, _065518_, _065519_, _065520_, _065521_, _065522_, _065523_, _065524_, _065525_, _065526_, _065527_, _065528_, _065529_, _065530_, _065531_, _065532_, _065533_, _065534_, _065535_, _065536_, _065537_, _065538_, _065539_, _065540_, _065541_, _065542_, _065543_, _065544_, _065545_, _065546_, _065547_, _065548_, _065549_, _065550_, _065551_, _065552_, _065553_, _065554_, _065555_, _065556_, _065557_, _065558_, _065559_, _065560_, _065561_, _065562_, _065563_, _065564_, _065565_, _065566_, _065567_, _065568_, _065569_, _065570_, _065571_, _065572_, _065573_, _065574_, _065575_, _065576_, _065577_, _065578_, _065579_, _065580_, _065581_, _065582_, _065583_, _065584_, _065585_, _065586_, _065587_, _065588_, _065589_, _065590_, _065591_, _065592_, _065593_, _065594_, _065595_, _065596_, _065597_, _065598_, _065599_, _065600_, _065601_, _065602_, _065603_, _065604_, _065605_, _065606_, _065607_, _065608_, _065609_, _065610_, _065611_, _065612_, _065613_, _065614_, _065615_, _065616_, _065617_, _065618_, _065619_, _065620_, _065621_, _065622_, _065623_, _065624_, _065625_, _065626_, _065627_, _065628_, _065629_, _065630_, _065631_, _065632_, _065633_, _065634_, _065635_, _065636_, _065637_, _065638_, _065639_, _065640_, _065641_, _065642_, _065643_, _065644_, _065645_, _065646_, _065647_, _065648_, _065649_, _065650_, _065651_, _065652_, _065653_, _065654_, _065655_, _065656_, _065657_, _065658_, _065659_, _065660_, _065661_, _065662_, _065663_, _065664_, _065665_, _065666_, _065667_, _065668_, _065669_, _065670_, _065671_, _065672_, _065673_, _065674_, _065675_, _065676_, _065677_, _065678_, _065679_, _065680_, _065681_, _065682_, _065683_, _065684_, _065685_, _065686_, _065687_, _065688_, _065689_, _065690_, _065691_, _065692_, _065693_, _065694_, _065695_, _065696_, _065697_, _065698_, _065699_, _065700_, _065701_, _065702_, _065703_, _065704_, _065705_, _065706_, _065707_, _065708_, _065709_, _065710_, _065711_, _065712_, _065713_, _065714_, _065715_, _065716_, _065717_, _065718_, _065719_, _065720_, _065721_, _065722_, _065723_, _065724_, _065725_, _065726_, _065727_, _065728_, _065729_, _065730_, _065731_, _065732_, _065733_, _065734_, _065735_, _065736_, _065737_, _065738_, _065739_, _065740_, _065741_, _065742_, _065743_, _065744_, _065745_, _065746_, _065747_, _065748_, _065749_, _065750_, _065751_, _065752_, _065753_, _065754_, _065755_, _065756_, _065757_, _065758_, _065759_, _065760_, _065761_, _065762_, _065763_, _065764_, _065765_, _065766_, _065767_, _065768_, _065769_, _065770_, _065771_, _065772_, _065773_, _065774_, _065775_, _065776_, _065777_, _065778_, _065779_, _065780_, _065781_, _065782_, _065783_, _065784_, _065785_, _065786_, _065787_, _065788_, _065789_, _065790_, _065791_, _065792_, _065793_, _065794_, _065795_, _065796_, _065797_, _065798_, _065799_, _065800_, _065801_, _065802_, _065803_, _065804_, _065805_, _065806_, _065807_, _065808_, _065809_, _065810_, _065811_, _065812_, _065813_, _065814_, _065815_, _065816_, _065817_, _065818_, _065819_, _065820_, _065821_, _065822_, _065823_, _065824_, _065825_, _065826_, _065827_, _065828_, _065829_, _065830_, _065831_, _065832_, _065833_, _065834_, _065835_, _065836_, _065837_, _065838_, _065839_, _065840_, _065841_, _065842_, _065843_, _065844_, _065845_, _065846_, _065847_, _065848_, _065849_, _065850_, _065851_, _065852_, _065853_, _065854_, _065855_, _065856_, _065857_, _065858_, _065859_, _065860_, _065861_, _065862_, _065863_, _065864_, _065865_, _065866_, _065867_, _065868_, _065869_, _065870_, _065871_, _065872_, _065873_, _065874_, _065875_, _065876_, _065877_, _065878_, _065879_, _065880_, _065881_, _065882_, _065883_, _065884_, _065885_, _065886_, _065887_, _065888_, _065889_, _065890_, _065891_, _065892_, _065893_, _065894_, _065895_, _065896_, _065897_, _065898_, _065899_, _065900_, _065901_, _065902_, _065903_, _065904_, _065905_, _065906_, _065907_, _065908_, _065909_, _065910_, _065911_, _065912_, _065913_, _065914_, _065915_, _065916_, _065917_, _065918_, _065919_, _065920_, _065921_, _065922_, _065923_, _065924_, _065925_, _065926_, _065927_, _065928_, _065929_, _065930_, _065931_, _065932_, _065933_, _065934_, _065935_, _065936_, _065937_, _065938_, _065939_, _065940_, _065941_, _065942_, _065943_, _065944_, _065945_, _065946_, _065947_, _065948_, _065949_, _065950_, _065951_, _065952_, _065953_, _065954_, _065955_, _065956_, _065957_, _065958_, _065959_, _065960_, _065961_, _065962_, _065963_, _065964_, _065965_, _065966_, _065967_, _065968_, _065969_, _065970_, _065971_, _065972_, _065973_, _065974_, _065975_, _065976_, _065977_, _065978_, _065979_, _065980_, _065981_, _065982_, _065983_, _065984_, _065985_, _065986_, _065987_, _065988_, _065989_, _065990_, _065991_, _065992_, _065993_, _065994_, _065995_, _065996_, _065997_, _065998_, _065999_, _066000_, _066001_, _066002_, _066003_, _066004_, _066005_, _066006_, _066007_, _066008_, _066009_, _066010_, _066011_, _066012_, _066013_, _066014_, _066015_, _066016_, _066017_, _066018_, _066019_, _066020_, _066021_, _066022_, _066023_, _066024_, _066025_, _066026_, _066027_, _066028_, _066029_, _066030_, _066031_, _066032_, _066033_, _066034_, _066035_, _066036_, _066037_, _066038_, _066039_, _066040_, _066041_, _066042_, _066043_, _066044_, _066045_, _066046_, _066047_, _066048_, _066049_, _066050_, _066051_, _066052_, _066053_, _066054_, _066055_, _066056_, _066057_, _066058_, _066059_, _066060_, _066061_, _066062_, _066063_, _066064_, _066065_, _066066_, _066067_, _066068_, _066069_, _066070_, _066071_, _066072_, _066073_, _066074_, _066075_, _066076_, _066077_, _066078_, _066079_, _066080_, _066081_, _066082_, _066083_, _066084_, _066085_, _066086_, _066087_, _066088_, _066089_, _066090_, _066091_, _066092_, _066093_, _066094_, _066095_, _066096_, _066097_, _066098_, _066099_, _066100_, _066101_, _066102_, _066103_, _066104_, _066105_, _066106_, _066107_, _066108_, _066109_, _066110_, _066111_, _066112_, _066113_, _066114_, _066115_, _066116_, _066117_, _066118_, _066119_, _066120_, _066121_, _066122_, _066123_, _066124_, _066125_, _066126_, _066127_, _066128_, _066129_, _066130_, _066131_, _066132_, _066133_, _066134_, _066135_, _066136_, _066137_, _066138_, _066139_, _066140_, _066141_, _066142_, _066143_, _066144_, _066145_, _066146_, _066147_, _066148_, _066149_, _066150_, _066151_, _066152_, _066153_, _066154_, _066155_, _066156_, _066157_, _066158_, _066159_, _066160_, _066161_, _066162_, _066163_, _066164_, _066165_, _066166_, _066167_, _066168_, _066169_, _066170_, _066171_, _066172_, _066173_, _066174_, _066175_, _066176_, _066177_, _066178_, _066179_, _066180_, _066181_, _066182_, _066183_, _066184_, _066185_, _066186_, _066187_, _066188_, _066189_, _066190_, _066191_, _066192_, _066193_, _066194_, _066195_, _066196_, _066197_, _066198_, _066199_, _066200_, _066201_, _066202_, _066203_, _066204_, _066205_, _066206_, _066207_, _066208_, _066209_, _066210_, _066211_, _066212_, _066213_, _066214_, _066215_, _066216_, _066217_, _066218_, _066219_, _066220_, _066221_, _066222_, _066223_, _066224_, _066225_, _066226_, _066227_, _066228_, _066229_, _066230_, _066231_, _066232_, _066233_, _066234_, _066235_, _066236_, _066237_, _066238_, _066239_, _066240_, _066241_, _066242_, _066243_, _066244_, _066245_, _066246_, _066247_, _066248_, _066249_, _066250_, _066251_, _066252_, _066253_, _066254_, _066255_, _066256_, _066257_, _066258_, _066259_, _066260_, _066261_, _066262_, _066263_, _066264_, _066265_, _066266_, _066267_, _066268_, _066269_, _066270_, _066271_, _066272_, _066273_, _066274_, _066275_, _066276_, _066277_, _066278_, _066279_, _066280_, _066281_, _066282_, _066283_, _066284_, _066285_, _066286_, _066287_, _066288_, _066289_, _066290_, _066291_, _066292_, _066293_, _066294_, _066295_, _066296_, _066297_, _066298_, _066299_, _066300_, _066301_, _066302_, _066303_, _066304_, _066305_, _066306_, _066307_, _066308_, _066309_, _066310_, _066311_, _066312_, _066313_, _066314_, _066315_, _066316_, _066317_, _066318_, _066319_, _066320_, _066321_, _066322_, _066323_, _066324_, _066325_, _066326_, _066327_, _066328_, _066329_, _066330_, _066331_, _066332_, _066333_, _066334_, _066335_, _066336_, _066337_, _066338_, _066339_, _066340_, _066341_, _066342_, _066343_, _066344_, _066345_, _066346_, _066347_, _066348_, _066349_, _066350_, _066351_, _066352_, _066353_, _066354_, _066355_, _066356_, _066357_, _066358_, _066359_, _066360_, _066361_, _066362_, _066363_, _066364_, _066365_, _066366_, _066367_, _066368_, _066369_, _066370_, _066371_, _066372_, _066373_, _066374_, _066375_, _066376_, _066377_, _066378_, _066379_, _066380_, _066381_, _066382_, _066383_, _066384_, _066385_, _066386_, _066387_, _066388_, _066389_, _066390_, _066391_, _066392_, _066393_, _066394_, _066395_, _066396_, _066397_, _066398_, _066399_, _066400_, _066401_, _066402_, _066403_, _066404_, _066405_, _066406_, _066407_, _066408_, _066409_, _066410_, _066411_, _066412_, _066413_, _066414_, _066415_, _066416_, _066417_, _066418_, _066419_, _066420_, _066421_, _066422_, _066423_, _066424_, _066425_, _066426_, _066427_, _066428_, _066429_, _066430_, _066431_, _066432_, _066433_, _066434_, _066435_, _066436_, _066437_, _066438_, _066439_, _066440_, _066441_, _066442_, _066443_, _066444_, _066445_, _066446_, _066447_, _066448_, _066449_, _066450_, _066451_, _066452_, _066453_, _066454_, _066455_, _066456_, _066457_, _066458_, _066459_, _066460_, _066461_, _066462_, _066463_, _066464_, _066465_, _066466_, _066467_, _066468_, _066469_, _066470_, _066471_, _066472_, _066473_, _066474_, _066475_, _066476_, _066477_, _066478_, _066479_, _066480_, _066481_, _066482_, _066483_, _066484_, _066485_, _066486_, _066487_, _066488_, _066489_, _066490_, _066491_, _066492_, _066493_, _066494_, _066495_, _066496_, _066497_, _066498_, _066499_, _066500_, _066501_, _066502_, _066503_, _066504_, _066505_, _066506_, _066507_, _066508_, _066509_, _066510_, _066511_, _066512_, _066513_, _066514_, _066515_, _066516_, _066517_, _066518_, _066519_, _066520_, _066521_, _066522_, _066523_, _066524_, _066525_, _066526_, _066527_, _066528_, _066529_, _066530_, _066531_, _066532_, _066533_, _066534_, _066535_, _066536_, _066537_, _066538_, _066539_, _066540_, _066541_, _066542_, _066543_, _066544_, _066545_, _066546_, _066547_, _066548_, _066549_, _066550_, _066551_, _066552_, _066553_, _066554_, _066555_, _066556_, _066557_, _066558_, _066559_, _066560_, _066561_, _066562_, _066563_, _066564_, _066565_, _066566_, _066567_, _066568_, _066569_, _066570_, _066571_, _066572_, _066573_, _066574_, _066575_, _066576_, _066577_, _066578_, _066579_, _066580_, _066581_, _066582_, _066583_, _066584_, _066585_, _066586_, _066587_, _066588_, _066589_, _066590_, _066591_, _066592_, _066593_, _066594_, _066595_, _066596_, _066597_, _066598_, _066599_, _066600_, _066601_, _066602_, _066603_, _066604_, _066605_, _066606_, _066607_, _066608_, _066609_, _066610_, _066611_, _066612_, _066613_, _066614_, _066615_, _066616_, _066617_, _066618_, _066619_, _066620_, _066621_, _066622_, _066623_, _066624_, _066625_, _066626_, _066627_, _066628_, _066629_, _066630_, _066631_, _066632_, _066633_, _066634_, _066635_, _066636_, _066637_, _066638_, _066639_, _066640_, _066641_, _066642_, _066643_, _066644_, _066645_, _066646_, _066647_, _066648_, _066649_, _066650_, _066651_, _066652_, _066653_, _066654_, _066655_, _066656_, _066657_, _066658_, _066659_, _066660_, _066661_, _066662_, _066663_, _066664_, _066665_, _066666_, _066667_, _066668_, _066669_, _066670_, _066671_, _066672_, _066673_, _066674_, _066675_, _066676_, _066677_, _066678_, _066679_, _066680_, _066681_, _066682_, _066683_, _066684_, _066685_, _066686_, _066687_, _066688_, _066689_, _066690_, _066691_, _066692_, _066693_, _066694_, _066695_, _066696_, _066697_, _066698_, _066699_, _066700_, _066701_, _066702_, _066703_, _066704_, _066705_, _066706_, _066707_, _066708_, _066709_, _066710_, _066711_, _066712_, _066713_, _066714_, _066715_, _066716_, _066717_, _066718_, _066719_, _066720_, _066721_, _066722_, _066723_, _066724_, _066725_, _066726_, _066727_, _066728_, _066729_, _066730_, _066731_, _066732_, _066733_, _066734_, _066735_, _066736_, _066737_, _066738_, _066739_, _066740_, _066741_, _066742_, _066743_, _066744_, _066745_, _066746_, _066747_, _066748_, _066749_, _066750_, _066751_, _066752_, _066753_, _066754_, _066755_, _066756_, _066757_, _066758_, _066759_, _066760_, _066761_, _066762_, _066763_, _066764_, _066765_, _066766_, _066767_, _066768_, _066769_, _066770_, _066771_, _066772_, _066773_, _066774_, _066775_, _066776_, _066777_, _066778_, _066779_, _066780_, _066781_, _066782_, _066783_, _066784_, _066785_, _066786_, _066787_, _066788_, _066789_, _066790_, _066791_, _066792_, _066793_, _066794_, _066795_, _066796_, _066797_, _066798_, _066799_, _066800_, _066801_, _066802_, _066803_, _066804_, _066805_, _066806_, _066807_, _066808_, _066809_, _066810_, _066811_, _066812_, _066813_, _066814_, _066815_, _066816_, _066817_, _066818_, _066819_, _066820_, _066821_, _066822_, _066823_, _066824_, _066825_, _066826_, _066827_, _066828_, _066829_, _066830_, _066831_, _066832_, _066833_, _066834_, _066835_, _066836_, _066837_, _066838_, _066839_, _066840_, _066841_, _066842_, _066843_, _066844_, _066845_, _066846_, _066847_, _066848_, _066849_, _066850_, _066851_, _066852_, _066853_, _066854_, _066855_, _066856_, _066857_, _066858_, _066859_, _066860_, _066861_, _066862_, _066863_, _066864_, _066865_, _066866_, _066867_, _066868_, _066869_, _066870_, _066871_, _066872_, _066873_, _066874_, _066875_, _066876_, _066877_, _066878_, _066879_, _066880_, _066881_, _066882_, _066883_, _066884_, _066885_, _066886_, _066887_, _066888_, _066889_, _066890_, _066891_, _066892_, _066893_, _066894_, _066895_, _066896_, _066897_, _066898_, _066899_, _066900_, _066901_, _066902_, _066903_, _066904_, _066905_, _066906_, _066907_, _066908_, _066909_, _066910_, _066911_, _066912_, _066913_, _066914_, _066915_, _066916_, _066917_, _066918_, _066919_, _066920_, _066921_, _066922_, _066923_, _066924_, _066925_, _066926_, _066927_, _066928_, _066929_, _066930_, _066931_, _066932_, _066933_, _066934_, _066935_, _066936_, _066937_, _066938_, _066939_, _066940_, _066941_, _066942_, _066943_, _066944_, _066945_, _066946_, _066947_, _066948_, _066949_, _066950_, _066951_, _066952_, _066953_, _066954_, _066955_, _066956_, _066957_, _066958_, _066959_, _066960_, _066961_, _066962_, _066963_, _066964_, _066965_, _066966_, _066967_, _066968_, _066969_, _066970_, _066971_, _066972_, _066973_, _066974_, _066975_, _066976_, _066977_, _066978_, _066979_, _066980_, _066981_, _066982_, _066983_, _066984_, _066985_, _066986_, _066987_, _066988_, _066989_, _066990_, _066991_, _066992_, _066993_, _066994_, _066995_, _066996_, _066997_, _066998_, _066999_, _067000_, _067001_, _067002_, _067003_, _067004_, _067005_, _067006_, _067007_, _067008_, _067009_, _067010_, _067011_, _067012_, _067013_, _067014_, _067015_, _067016_, _067017_, _067018_, _067019_, _067020_, _067021_, _067022_, _067023_, _067024_, _067025_, _067026_, _067027_, _067028_, _067029_, _067030_, _067031_, _067032_, _067033_, _067034_, _067035_, _067036_, _067037_, _067038_, _067039_, _067040_, _067041_, _067042_, _067043_, _067044_, _067045_, _067046_, _067047_, _067048_, _067049_, _067050_, _067051_, _067052_, _067053_, _067054_, _067055_, _067056_, _067057_, _067058_, _067059_, _067060_, _067061_, _067062_, _067063_, _067064_, _067065_, _067066_, _067067_, _067068_, _067069_, _067070_, _067071_, _067072_, _067073_, _067074_, _067075_, _067076_, _067077_, _067078_, _067079_, _067080_, _067081_, _067082_, _067083_, _067084_, _067085_, _067086_, _067087_, _067088_, _067089_, _067090_, _067091_, _067092_, _067093_, _067094_, _067095_, _067096_, _067097_, _067098_, _067099_, _067100_, _067101_, _067102_, _067103_, _067104_, _067105_, _067106_, _067107_, _067108_, _067109_, _067110_, _067111_, _067112_, _067113_, _067114_, _067115_, _067116_, _067117_, _067118_, _067119_, _067120_, _067121_, _067122_, _067123_, _067124_, _067125_, _067126_, _067127_, _067128_, _067129_, _067130_, _067131_, _067132_, _067133_, _067134_, _067135_, _067136_, _067137_, _067138_, _067139_, _067140_, _067141_, _067142_, _067143_, _067144_, _067145_, _067146_, _067147_, _067148_, _067149_, _067150_, _067151_, _067152_, _067153_, _067154_, _067155_, _067156_, _067157_, _067158_, _067159_, _067160_, _067161_, _067162_, _067163_, _067164_, _067165_, _067166_, _067167_, _067168_, _067169_, _067170_, _067171_, _067172_, _067173_, _067174_, _067175_, _067176_, _067177_, _067178_, _067179_, _067180_, _067181_, _067182_, _067183_, _067184_, _067185_, _067186_, _067187_, _067188_, _067189_, _067190_, _067191_, _067192_, _067193_, _067194_, _067195_, _067196_, _067197_, _067198_, _067199_, _067200_, _067201_, _067202_, _067203_, _067204_, _067205_, _067206_, _067207_, _067208_, _067209_, _067210_, _067211_, _067212_, _067213_, _067214_, _067215_, _067216_, _067217_, _067218_, _067219_, _067220_, _067221_, _067222_, _067223_, _067224_, _067225_, _067226_, _067227_, _067228_, _067229_, _067230_, _067231_, _067232_, _067233_, _067234_, _067235_, _067236_, _067237_, _067238_, _067239_, _067240_, _067241_, _067242_, _067243_, _067244_, _067245_, _067246_, _067247_, _067248_, _067249_, _067250_, _067251_, _067252_, _067253_, _067254_, _067255_, _067256_, _067257_, _067258_, _067259_, _067260_, _067261_, _067262_, _067263_, _067264_, _067265_, _067266_, _067267_, _067268_, _067269_, _067270_, _067271_, _067272_, _067273_, _067274_, _067275_, _067276_, _067277_, _067278_, _067279_, _067280_, _067281_, _067282_, _067283_, _067284_, _067285_, _067286_, _067287_, _067288_, _067289_, _067290_, _067291_, _067292_, _067293_, _067294_, _067295_, _067296_, _067297_, _067298_, _067299_, _067300_, _067301_, _067302_, _067303_, _067304_, _067305_, _067306_, _067307_, _067308_, _067309_, _067310_, _067311_, _067312_, _067313_, _067314_, _067315_, _067316_, _067317_, _067318_, _067319_, _067320_, _067321_, _067322_, _067323_, _067324_, _067325_, _067326_, _067327_, _067328_, _067329_, _067330_, _067331_, _067332_, _067333_, _067334_, _067335_, _067336_, _067337_, _067338_, _067339_, _067340_, _067341_, _067342_, _067343_, _067344_, _067345_, _067346_, _067347_, _067348_, _067349_, _067350_, _067351_, _067352_, _067353_, _067354_, _067355_, _067356_, _067357_, _067358_, _067359_, _067360_, _067361_, _067362_, _067363_, _067364_, _067365_, _067366_, _067367_, _067368_, _067369_, _067370_, _067371_, _067372_, _067373_, _067374_, _067375_, _067376_, _067377_, _067378_, _067379_, _067380_, _067381_, _067382_, _067383_, _067384_, _067385_, _067386_, _067387_, _067388_, _067389_, _067390_, _067391_, _067392_, _067393_, _067394_, _067395_, _067396_, _067397_, _067398_, _067399_, _067400_, _067401_, _067402_, _067403_, _067404_, _067405_, _067406_, _067407_, _067408_, _067409_, _067410_, _067411_, _067412_, _067413_, _067414_, _067415_, _067416_, _067417_, _067418_, _067419_, _067420_, _067421_, _067422_, _067423_, _067424_, _067425_, _067426_, _067427_, _067428_, _067429_, _067430_, _067431_, _067432_, _067433_, _067434_, _067435_, _067436_, _067437_, _067438_, _067439_, _067440_, _067441_, _067442_, _067443_, _067444_, _067445_, _067446_, _067447_, _067448_, _067449_, _067450_, _067451_, _067452_, _067453_, _067454_, _067455_, _067456_, _067457_, _067458_, _067459_, _067460_, _067461_, _067462_, _067463_, _067464_, _067465_, _067466_, _067467_, _067468_, _067469_, _067470_, _067471_, _067472_, _067473_, _067474_, _067475_, _067476_, _067477_, _067478_, _067479_, _067480_, _067481_, _067482_, _067483_, _067484_, _067485_, _067486_, _067487_, _067488_, _067489_, _067490_, _067491_, _067492_, _067493_, _067494_, _067495_, _067496_, _067497_, _067498_, _067499_, _067500_, _067501_, _067502_, _067503_, _067504_, _067505_, _067506_, _067507_, _067508_, _067509_, _067510_, _067511_, _067512_, _067513_, _067514_, _067515_, _067516_, _067517_, _067518_, _067519_, _067520_, _067521_, _067522_, _067523_, _067524_, _067525_, _067526_, _067527_, _067528_, _067529_, _067530_, _067531_, _067532_, _067533_, _067534_, _067535_, _067536_, _067537_, _067538_, _067539_, _067540_, _067541_, _067542_, _067543_, _067544_, _067545_, _067546_, _067547_, _067548_, _067549_, _067550_, _067551_, _067552_, _067553_, _067554_, _067555_, _067556_, _067557_, _067558_, _067559_, _067560_, _067561_, _067562_, _067563_, _067564_, _067565_, _067566_, _067567_, _067568_, _067569_, _067570_, _067571_, _067572_, _067573_, _067574_, _067575_, _067576_, _067577_, _067578_, _067579_, _067580_, _067581_, _067582_, _067583_, _067584_, _067585_, _067586_, _067587_, _067588_, _067589_, _067590_, _067591_, _067592_, _067593_, _067594_, _067595_, _067596_, _067597_, _067598_, _067599_, _067600_, _067601_, _067602_, _067603_, _067604_, _067605_, _067606_, _067607_, _067608_, _067609_, _067610_, _067611_, _067612_, _067613_, _067614_, _067615_, _067616_, _067617_, _067618_, _067619_, _067620_, _067621_, _067622_, _067623_, _067624_, _067625_, _067626_, _067627_, _067628_, _067629_, _067630_, _067631_, _067632_, _067633_, _067634_, _067635_, _067636_, _067637_, _067638_, _067639_, _067640_, _067641_, _067642_, _067643_, _067644_, _067645_, _067646_, _067647_, _067648_, _067649_, _067650_, _067651_, _067652_, _067653_, _067654_, _067655_, _067656_, _067657_, _067658_, _067659_, _067660_, _067661_, _067662_, _067663_, _067664_, _067665_, _067666_, _067667_, _067668_, _067669_, _067670_, _067671_, _067672_, _067673_, _067674_, _067675_, _067676_, _067677_, _067678_, _067679_, _067680_, _067681_, _067682_, _067683_, _067684_, _067685_, _067686_, _067687_, _067688_, _067689_, _067690_, _067691_, _067692_, _067693_, _067694_, _067695_, _067696_, _067697_, _067698_, _067699_, _067700_, _067701_, _067702_, _067703_, _067704_, _067705_, _067706_, _067707_, _067708_, _067709_, _067710_, _067711_, _067712_, _067713_, _067714_, _067715_, _067716_, _067717_, _067718_, _067719_, _067720_, _067721_, _067722_, _067723_, _067724_, _067725_, _067726_, _067727_, _067728_, _067729_, _067730_, _067731_, _067732_, _067733_, _067734_, _067735_, _067736_, _067737_, _067738_, _067739_, _067740_, _067741_, _067742_, _067743_, _067744_, _067745_, _067746_, _067747_, _067748_, _067749_, _067750_, _067751_, _067752_, _067753_, _067754_, _067755_, _067756_, _067757_, _067758_, _067759_, _067760_, _067761_, _067762_, _067763_, _067764_, _067765_, _067766_, _067767_, _067768_, _067769_, _067770_, _067771_, _067772_, _067773_, _067774_, _067775_, _067776_, _067777_, _067778_, _067779_, _067780_, _067781_, _067782_, _067783_, _067784_, _067785_, _067786_, _067787_, _067788_, _067789_, _067790_, _067791_, _067792_, _067793_, _067794_, _067795_, _067796_, _067797_, _067798_, _067799_, _067800_, _067801_, _067802_, _067803_, _067804_, _067805_, _067806_, _067807_, _067808_, _067809_, _067810_, _067811_, _067812_, _067813_, _067814_, _067815_, _067816_, _067817_, _067818_, _067819_, _067820_, _067821_, _067822_, _067823_, _067824_, _067825_, _067826_, _067827_, _067828_, _067829_, _067830_, _067831_, _067832_, _067833_, _067834_, _067835_, _067836_, _067837_, _067838_, _067839_, _067840_, _067841_, _067842_, _067843_, _067844_, _067845_, _067846_, _067847_, _067848_, _067849_, _067850_, _067851_, _067852_, _067853_, _067854_, _067855_, _067856_, _067857_, _067858_, _067859_, _067860_, _067861_, _067862_, _067863_, _067864_, _067865_, _067866_, _067867_, _067868_, _067869_, _067870_, _067871_, _067872_, _067873_, _067874_, _067875_, _067876_, _067877_, _067878_, _067879_, _067880_, _067881_, _067882_, _067883_, _067884_, _067885_, _067886_, _067887_, _067888_, _067889_, _067890_, _067891_, _067892_, _067893_, _067894_, _067895_, _067896_, _067897_, _067898_, _067899_, _067900_, _067901_, _067902_, _067903_, _067904_, _067905_, _067906_, _067907_, _067908_, _067909_, _067910_, _067911_, _067912_, _067913_, _067914_, _067915_, _067916_, _067917_, _067918_, _067919_, _067920_, _067921_, _067922_, _067923_, _067924_, _067925_, _067926_, _067927_, _067928_, _067929_, _067930_, _067931_, _067932_, _067933_, _067934_, _067935_, _067936_, _067937_, _067938_, _067939_, _067940_, _067941_, _067942_, _067943_, _067944_, _067945_, _067946_, _067947_, _067948_, _067949_, _067950_, _067951_, _067952_, _067953_, _067954_, _067955_, _067956_, _067957_, _067958_, _067959_, _067960_, _067961_, _067962_, _067963_, _067964_, _067965_, _067966_, _067967_, _067968_, _067969_, _067970_, _067971_, _067972_, _067973_, _067974_, _067975_, _067976_, _067977_, _067978_, _067979_, _067980_, _067981_, _067982_, _067983_, _067984_, _067985_, _067986_, _067987_, _067988_, _067989_, _067990_, _067991_, _067992_, _067993_, _067994_, _067995_, _067996_, _067997_, _067998_, _067999_, _068000_, _068001_, _068002_, _068003_, _068004_, _068005_, _068006_, _068007_, _068008_, _068009_, _068010_, _068011_, _068012_, _068013_, _068014_, _068015_, _068016_, _068017_, _068018_, _068019_, _068020_, _068021_, _068022_, _068023_, _068024_, _068025_, _068026_, _068027_, _068028_, _068029_, _068030_, _068031_, _068032_, _068033_, _068034_, _068035_, _068036_, _068037_, _068038_, _068039_, _068040_, _068041_, _068042_, _068043_, _068044_, _068045_, _068046_, _068047_, _068048_, _068049_, _068050_, _068051_, _068052_, _068053_, _068054_, _068055_, _068056_, _068057_, _068058_, _068059_, _068060_, _068061_, _068062_, _068063_, _068064_, _068065_, _068066_, _068067_, _068068_, _068069_, _068070_, _068071_, _068072_, _068073_, _068074_, _068075_, _068076_, _068077_, _068078_, _068079_, _068080_, _068081_, _068082_, _068083_, _068084_, _068085_, _068086_, _068087_, _068088_, _068089_, _068090_, _068091_, _068092_, _068093_, _068094_, _068095_, _068096_, _068097_, _068098_, _068099_, _068100_, _068101_, _068102_, _068103_, _068104_, _068105_, _068106_, _068107_, _068108_, _068109_, _068110_, _068111_, _068112_, _068113_, _068114_, _068115_, _068116_, _068117_, _068118_, _068119_, _068120_, _068121_, _068122_, _068123_, _068124_, _068125_, _068126_, _068127_, _068128_, _068129_, _068130_, _068131_, _068132_, _068133_, _068134_, _068135_, _068136_, _068137_, _068138_, _068139_, _068140_, _068141_, _068142_, _068143_, _068144_, _068145_, _068146_, _068147_, _068148_, _068149_, _068150_, _068151_, _068152_, _068153_, _068154_, _068155_, _068156_, _068157_, _068158_, _068159_, _068160_, _068161_, _068162_, _068163_, _068164_, _068165_, _068166_, _068167_, _068168_, _068169_, _068170_, _068171_, _068172_, _068173_, _068174_, _068175_, _068176_, _068177_, _068178_, _068179_, _068180_, _068181_, _068182_, _068183_, _068184_, _068185_, _068186_, _068187_, _068188_, _068189_, _068190_, _068191_, _068192_, _068193_, _068194_, _068195_, _068196_, _068197_, _068198_, _068199_, _068200_, _068201_, _068202_, _068203_, _068204_, _068205_, _068206_, _068207_, _068208_, _068209_, _068210_, _068211_, _068212_, _068213_, _068214_, _068215_, _068216_, _068217_, _068218_, _068219_, _068220_, _068221_, _068222_, _068223_, _068224_, _068225_, _068226_, _068227_, _068228_, _068229_, _068230_, _068231_, _068232_, _068233_, _068234_, _068235_, _068236_, _068237_, _068238_, _068239_, _068240_, _068241_, _068242_, _068243_, _068244_, _068245_, _068246_, _068247_, _068248_, _068249_, _068250_, _068251_, _068252_, _068253_, _068254_, _068255_, _068256_, _068257_, _068258_, _068259_, _068260_, _068261_, _068262_, _068263_, _068264_, _068265_, _068266_, _068267_, _068268_, _068269_, _068270_, _068271_, _068272_, _068273_, _068274_, _068275_, _068276_, _068277_, _068278_, _068279_, _068280_, _068281_, _068282_, _068283_, _068284_, _068285_, _068286_, _068287_, _068288_, _068289_, _068290_, _068291_, _068292_, _068293_, _068294_, _068295_, _068296_, _068297_, _068298_, _068299_, _068300_, _068301_, _068302_, _068303_, _068304_, _068305_, _068306_, _068307_, _068308_, _068309_, _068310_, _068311_, _068312_, _068313_, _068314_, _068315_, _068316_, _068317_, _068318_, _068319_, _068320_, _068321_, _068322_, _068323_, _068324_, _068325_, _068326_, _068327_, _068328_, _068329_, _068330_, _068331_, _068332_, _068333_, _068334_, _068335_, _068336_, _068337_, _068338_, _068339_, _068340_, _068341_, _068342_, _068343_, _068344_, _068345_, _068346_, _068347_, _068348_, _068349_, _068350_, _068351_, _068352_, _068353_, _068354_, _068355_, _068356_, _068357_, _068358_, _068359_, _068360_, _068361_, _068362_, _068363_, _068364_, _068365_, _068366_, _068367_, _068368_, _068369_, _068370_, _068371_, _068372_, _068373_, _068374_, _068375_, _068376_, _068377_, _068378_, _068379_, _068380_, _068381_, _068382_, _068383_, _068384_, _068385_, _068386_, _068387_, _068388_, _068389_, _068390_, _068391_, _068392_, _068393_, _068394_, _068395_, _068396_, _068397_, _068398_, _068399_, _068400_, _068401_, _068402_, _068403_, _068404_, _068405_, _068406_, _068407_, _068408_, _068409_, _068410_, _068411_, _068412_, _068413_, _068414_, _068415_, _068416_, _068417_, _068418_, _068419_, _068420_, _068421_, _068422_, _068423_, _068424_, _068425_, _068426_, _068427_, _068428_, _068429_, _068430_, _068431_, _068432_, _068433_, _068434_, _068435_, _068436_, _068437_, _068438_, _068439_, _068440_, _068441_, _068442_, _068443_, _068444_, _068445_, _068446_, _068447_, _068448_, _068449_, _068450_, _068451_, _068452_, _068453_, _068454_, _068455_, _068456_, _068457_, _068458_, _068459_, _068460_, _068461_, _068462_, _068463_, _068464_, _068465_, _068466_, _068467_, _068468_, _068469_, _068470_, _068471_, _068472_, _068473_, _068474_, _068475_, _068476_, _068477_, _068478_, _068479_, _068480_, _068481_, _068482_, _068483_, _068484_, _068485_, _068486_, _068487_, _068488_, _068489_, _068490_, _068491_, _068492_, _068493_, _068494_, _068495_, _068496_, _068497_, _068498_, _068499_, _068500_, _068501_, _068502_, _068503_, _068504_, _068505_, _068506_, _068507_, _068508_, _068509_, _068510_, _068511_, _068512_, _068513_, _068514_, _068515_, _068516_, _068517_, _068518_, _068519_, _068520_, _068521_, _068522_, _068523_, _068524_, _068525_, _068526_, _068527_, _068528_, _068529_, _068530_, _068531_, _068532_, _068533_, _068534_, _068535_, _068536_, _068537_, _068538_, _068539_, _068540_, _068541_, _068542_, _068543_, _068544_, _068545_, _068546_, _068547_, _068548_, _068549_, _068550_, _068551_, _068552_, _068553_, _068554_, _068555_, _068556_, _068557_, _068558_, _068559_, _068560_, _068561_, _068562_, _068563_, _068564_, _068565_, _068566_, _068567_, _068568_, _068569_, _068570_, _068571_, _068572_, _068573_, _068574_, _068575_, _068576_, _068577_, _068578_, _068579_, _068580_, _068581_, _068582_, _068583_, _068584_, _068585_, _068586_, _068587_, _068588_, _068589_, _068590_, _068591_, _068592_, _068593_, _068594_, _068595_, _068596_, _068597_, _068598_, _068599_, _068600_, _068601_, _068602_, _068603_, _068604_, _068605_, _068606_, _068607_, _068608_, _068609_, _068610_, _068611_, _068612_, _068613_, _068614_, _068615_, _068616_, _068617_, _068618_, _068619_, _068620_, _068621_, _068622_, _068623_, _068624_, _068625_, _068626_, _068627_, _068628_, _068629_, _068630_, _068631_, _068632_, _068633_, _068634_, _068635_, _068636_, _068637_, _068638_, _068639_, _068640_, _068641_, _068642_, _068643_, _068644_, _068645_, _068646_, _068647_, _068648_, _068649_, _068650_, _068651_, _068652_, _068653_, _068654_, _068655_, _068656_, _068657_, _068658_, _068659_, _068660_, _068661_, _068662_, _068663_, _068664_, _068665_, _068666_, _068667_, _068668_, _068669_, _068670_, _068671_, _068672_, _068673_, _068674_, _068675_, _068676_, _068677_, _068678_, _068679_, _068680_, _068681_, _068682_, _068683_, _068684_, _068685_, _068686_, _068687_, _068688_, _068689_, _068690_, _068691_, _068692_, _068693_, _068694_, _068695_, _068696_, _068697_, _068698_, _068699_, _068700_, _068701_, _068702_, _068703_, _068704_, _068705_, _068706_, _068707_, _068708_, _068709_, _068710_, _068711_, _068712_, _068713_, _068714_, _068715_, _068716_, _068717_, _068718_, _068719_, _068720_, _068721_, _068722_, _068723_, _068724_, _068725_, _068726_, _068727_, _068728_, _068729_, _068730_, _068731_, _068732_, _068733_, _068734_, _068735_, _068736_, _068737_, _068738_, _068739_, _068740_, _068741_, _068742_, _068743_, _068744_, _068745_, _068746_, _068747_, _068748_, _068749_, _068750_, _068751_, _068752_, _068753_, _068754_, _068755_, _068756_, _068757_, _068758_, _068759_, _068760_, _068761_, _068762_, _068763_, _068764_, _068765_, _068766_, _068767_, _068768_, _068769_, _068770_, _068771_, _068772_, _068773_, _068774_, _068775_, _068776_, _068777_, _068778_, _068779_, _068780_, _068781_, _068782_, _068783_, _068784_, _068785_, _068786_, _068787_, _068788_, _068789_, _068790_, _068791_, _068792_, _068793_, _068794_, _068795_, _068796_, _068797_, _068798_, _068799_, _068800_, _068801_, _068802_, _068803_, _068804_, _068805_, _068806_, _068807_, _068808_, _068809_, _068810_, _068811_, _068812_, _068813_, _068814_, _068815_, _068816_, _068817_, _068818_, _068819_, _068820_, _068821_, _068822_, _068823_, _068824_, _068825_, _068826_, _068827_, _068828_, _068829_, _068830_, _068831_, _068832_, _068833_, _068834_, _068835_, _068836_, _068837_, _068838_, _068839_, _068840_, _068841_, _068842_, _068843_, _068844_, _068845_, _068846_, _068847_, _068848_, _068849_, _068850_, _068851_, _068852_, _068853_, _068854_, _068855_, _068856_, _068857_, _068858_, _068859_, _068860_, _068861_, _068862_, _068863_, _068864_, _068865_, _068866_, _068867_, _068868_, _068869_, _068870_, _068871_, _068872_, _068873_, _068874_, _068875_, _068876_, _068877_, _068878_, _068879_, _068880_, _068881_, _068882_, _068883_, _068884_, _068885_, _068886_, _068887_, _068888_, _068889_, _068890_, _068891_, _068892_, _068893_, _068894_, _068895_, _068896_, _068897_, _068898_, _068899_, _068900_, _068901_, _068902_, _068903_, _068904_, _068905_, _068906_, _068907_, _068908_, _068909_, _068910_, _068911_, _068912_, _068913_, _068914_, _068915_, _068916_, _068917_, _068918_, _068919_, _068920_, _068921_, _068922_, _068923_, _068924_, _068925_, _068926_, _068927_, _068928_, _068929_, _068930_, _068931_, _068932_, _068933_, _068934_, _068935_, _068936_, _068937_, _068938_, _068939_, _068940_, _068941_, _068942_, _068943_, _068944_, _068945_, _068946_, _068947_, _068948_, _068949_, _068950_, _068951_, _068952_, _068953_, _068954_, _068955_, _068956_, _068957_, _068958_, _068959_, _068960_, _068961_, _068962_, _068963_, _068964_, _068965_, _068966_, _068967_, _068968_, _068969_, _068970_, _068971_, _068972_, _068973_, _068974_, _068975_, _068976_, _068977_, _068978_, _068979_, _068980_, _068981_, _068982_, _068983_, _068984_, _068985_, _068986_, _068987_, _068988_, _068989_, _068990_, _068991_, _068992_, _068993_, _068994_, _068995_, _068996_, _068997_, _068998_, _068999_, _069000_, _069001_, _069002_, _069003_, _069004_, _069005_, _069006_, _069007_, _069008_, _069009_, _069010_, _069011_, _069012_, _069013_, _069014_, _069015_, _069016_, _069017_, _069018_, _069019_, _069020_, _069021_, _069022_, _069023_, _069024_, _069025_, _069026_, _069027_, _069028_, _069029_, _069030_, _069031_, _069032_, _069033_, _069034_, _069035_, _069036_, _069037_, _069038_, _069039_, _069040_, _069041_, _069042_, _069043_, _069044_, _069045_, _069046_, _069047_, _069048_, _069049_, _069050_, _069051_, _069052_, _069053_, _069054_, _069055_, _069056_, _069057_, _069058_, _069059_, _069060_, _069061_, _069062_, _069063_, _069064_, _069065_, _069066_, _069067_, _069068_, _069069_, _069070_, _069071_, _069072_, _069073_, _069074_, _069075_, _069076_, _069077_, _069078_, _069079_, _069080_, _069081_, _069082_, _069083_, _069084_, _069085_, _069086_, _069087_, _069088_, _069089_, _069090_, _069091_, _069092_, _069093_, _069094_, _069095_, _069096_, _069097_, _069098_, _069099_, _069100_, _069101_, _069102_, _069103_, _069104_, _069105_, _069106_, _069107_, _069108_, _069109_, _069110_, _069111_, _069112_, _069113_, _069114_, _069115_, _069116_, _069117_, _069118_, _069119_, _069120_, _069121_, _069122_, _069123_, _069124_, _069125_, _069126_, _069127_, _069128_, _069129_, _069130_, _069131_, _069132_, _069133_, _069134_, _069135_, _069136_, _069137_, _069138_, _069139_, _069140_, _069141_, _069142_, _069143_, _069144_, _069145_, _069146_, _069147_, _069148_, _069149_, _069150_, _069151_, _069152_, _069153_, _069154_, _069155_, _069156_, _069157_, _069158_, _069159_, _069160_, _069161_, _069162_, _069163_, _069164_, _069165_, _069166_, _069167_, _069168_, _069169_, _069170_, _069171_, _069172_, _069173_, _069174_, _069175_, _069176_, _069177_, _069178_, _069179_, _069180_, _069181_, _069182_, _069183_, _069184_, _069185_, _069186_, _069187_, _069188_, _069189_, _069190_, _069191_, _069192_, _069193_, _069194_, _069195_, _069196_, _069197_, _069198_, _069199_, _069200_, _069201_, _069202_, _069203_, _069204_, _069205_, _069206_, _069207_, _069208_, _069209_, _069210_, _069211_, _069212_, _069213_, _069214_, _069215_, _069216_, _069217_, _069218_, _069219_, _069220_, _069221_, _069222_, _069223_, _069224_, _069225_, _069226_, _069227_, _069228_, _069229_, _069230_, _069231_, _069232_, _069233_, _069234_, _069235_, _069236_, _069237_, _069238_, _069239_, _069240_, _069241_, _069242_, _069243_, _069244_, _069245_, _069246_, _069247_, _069248_, _069249_, _069250_, _069251_, _069252_, _069253_, _069254_, _069255_, _069256_, _069257_, _069258_, _069259_, _069260_, _069261_, _069262_, _069263_, _069264_, _069265_, _069266_, _069267_, _069268_, _069269_, _069270_, _069271_, _069272_, _069273_, _069274_, _069275_, _069276_, _069277_, _069278_, _069279_, _069280_, _069281_, _069282_, _069283_, _069284_, _069285_, _069286_, _069287_, _069288_, _069289_, _069290_, _069291_, _069292_, _069293_, _069294_, _069295_, _069296_, _069297_, _069298_, _069299_, _069300_, _069301_, _069302_, _069303_, _069304_, _069305_, _069306_, _069307_, _069308_, _069309_, _069310_, _069311_, _069312_, _069313_, _069314_, _069315_, _069316_, _069317_, _069318_, _069319_, _069320_, _069321_, _069322_, _069323_, _069324_, _069325_, _069326_, _069327_, _069328_, _069329_, _069330_, _069331_, _069332_, _069333_, _069334_, _069335_, _069336_, _069337_, _069338_, _069339_, _069340_, _069341_, _069342_, _069343_, _069344_, _069345_, _069346_, _069347_, _069348_, _069349_, _069350_, _069351_, _069352_, _069353_, _069354_, _069355_, _069356_, _069357_, _069358_, _069359_, _069360_, _069361_, _069362_, _069363_, _069364_, _069365_, _069366_, _069367_, _069368_, _069369_, _069370_, _069371_, _069372_, _069373_, _069374_, _069375_, _069376_, _069377_, _069378_, _069379_, _069380_, _069381_, _069382_, _069383_, _069384_, _069385_, _069386_, _069387_, _069388_, _069389_, _069390_, _069391_, _069392_, _069393_, _069394_, _069395_, _069396_, _069397_, _069398_, _069399_, _069400_, _069401_, _069402_, _069403_, _069404_, _069405_, _069406_, _069407_, _069408_, _069409_, _069410_, _069411_, _069412_, _069413_, _069414_, _069415_, _069416_, _069417_, _069418_, _069419_, _069420_, _069421_, _069422_, _069423_, _069424_, _069425_, _069426_, _069427_, _069428_, _069429_, _069430_, _069431_, _069432_, _069433_, _069434_, _069435_, _069436_, _069437_, _069438_, _069439_, _069440_, _069441_, _069442_, _069443_, _069444_, _069445_, _069446_, _069447_, _069448_, _069449_, _069450_, _069451_, _069452_, _069453_, _069454_, _069455_, _069456_, _069457_, _069458_, _069459_, _069460_, _069461_, _069462_, _069463_, _069464_, _069465_, _069466_, _069467_, _069468_, _069469_, _069470_, _069471_, _069472_, _069473_, _069474_, _069475_, _069476_, _069477_, _069478_, _069479_, _069480_, _069481_, _069482_, _069483_, _069484_, _069485_, _069486_, _069487_, _069488_, _069489_, _069490_, _069491_, _069492_, _069493_, _069494_, _069495_, _069496_, _069497_, _069498_, _069499_, _069500_, _069501_, _069502_, _069503_, _069504_, _069505_, _069506_, _069507_, _069508_, _069509_, _069510_, _069511_, _069512_, _069513_, _069514_, _069515_, _069516_, _069517_, _069518_, _069519_, _069520_, _069521_, _069522_, _069523_, _069524_, _069525_, _069526_, _069527_, _069528_, _069529_, _069530_, _069531_, _069532_, _069533_, _069534_, _069535_, _069536_, _069537_, _069538_, _069539_, _069540_, _069541_, _069542_, _069543_, _069544_, _069545_, _069546_, _069547_, _069548_, _069549_, _069550_, _069551_, _069552_, _069553_, _069554_, _069555_, _069556_, _069557_, _069558_, _069559_, _069560_, _069561_, _069562_, _069563_, _069564_, _069565_, _069566_, _069567_, _069568_, _069569_, _069570_, _069571_, _069572_, _069573_, _069574_, _069575_, _069576_, _069577_, _069578_, _069579_, _069580_, _069581_, _069582_, _069583_, _069584_, _069585_, _069586_, _069587_, _069588_, _069589_, _069590_, _069591_, _069592_, _069593_, _069594_, _069595_, _069596_, _069597_, _069598_, _069599_, _069600_, _069601_, _069602_, _069603_, _069604_, _069605_, _069606_, _069607_, _069608_, _069609_, _069610_, _069611_, _069612_, _069613_, _069614_, _069615_, _069616_, _069617_, _069618_, _069619_, _069620_, _069621_, _069622_, _069623_, _069624_, _069625_, _069626_, _069627_, _069628_, _069629_, _069630_, _069631_, _069632_, _069633_, _069634_, _069635_, _069636_, _069637_, _069638_, _069639_, _069640_, _069641_, _069642_, _069643_, _069644_, _069645_, _069646_, _069647_, _069648_, _069649_, _069650_, _069651_, _069652_, _069653_, _069654_, _069655_, _069656_, _069657_, _069658_, _069659_, _069660_, _069661_, _069662_, _069663_, _069664_, _069665_, _069666_, _069667_, _069668_, _069669_, _069670_, _069671_, _069672_, _069673_, _069674_, _069675_, _069676_, _069677_, _069678_, _069679_, _069680_, _069681_, _069682_, _069683_, _069684_, _069685_, _069686_, _069687_, _069688_, _069689_, _069690_, _069691_, _069692_, _069693_, _069694_, _069695_, _069696_, _069697_, _069698_, _069699_, _069700_, _069701_, _069702_, _069703_, _069704_, _069705_, _069706_, _069707_, _069708_, _069709_, _069710_, _069711_, _069712_, _069713_, _069714_, _069715_, _069716_, _069717_, _069718_, _069719_, _069720_, _069721_, _069722_, _069723_, _069724_, _069725_, _069726_, _069727_, _069728_, _069729_, _069730_, _069731_, _069732_, _069733_, _069734_, _069735_, _069736_, _069737_, _069738_, _069739_, _069740_, _069741_, _069742_, _069743_, _069744_, _069745_, _069746_, _069747_, _069748_, _069749_, _069750_, _069751_, _069752_, _069753_, _069754_, _069755_, _069756_, _069757_, _069758_, _069759_, _069760_, _069761_, _069762_, _069763_, _069764_, _069765_, _069766_, _069767_, _069768_, _069769_, _069770_, _069771_, _069772_, _069773_, _069774_, _069775_, _069776_, _069777_, _069778_, _069779_, _069780_, _069781_, _069782_, _069783_, _069784_, _069785_, _069786_, _069787_, _069788_, _069789_, _069790_, _069791_, _069792_, _069793_, _069794_, _069795_, _069796_, _069797_, _069798_, _069799_, _069800_, _069801_, _069802_, _069803_, _069804_, _069805_, _069806_, _069807_, _069808_, _069809_, _069810_, _069811_, _069812_, _069813_, _069814_, _069815_, _069816_, _069817_, _069818_, _069819_, _069820_, _069821_, _069822_, _069823_, _069824_, _069825_, _069826_, _069827_, _069828_, _069829_, _069830_, _069831_, _069832_, _069833_, _069834_, _069835_, _069836_, _069837_, _069838_, _069839_, _069840_, _069841_, _069842_, _069843_, _069844_, _069845_, _069846_, _069847_, _069848_, _069849_, _069850_, _069851_, _069852_, _069853_, _069854_, _069855_, _069856_, _069857_, _069858_, _069859_, _069860_, _069861_, _069862_, _069863_, _069864_, _069865_, _069866_, _069867_, _069868_, _069869_, _069870_, _069871_, _069872_, _069873_, _069874_, _069875_, _069876_, _069877_, _069878_, _069879_, _069880_, _069881_, _069882_, _069883_, _069884_, _069885_, _069886_, _069887_, _069888_, _069889_, _069890_, _069891_, _069892_, _069893_, _069894_, _069895_, _069896_, _069897_, _069898_, _069899_, _069900_, _069901_, _069902_, _069903_, _069904_, _069905_, _069906_, _069907_, _069908_, _069909_, _069910_, _069911_, _069912_, _069913_, _069914_, _069915_, _069916_, _069917_, _069918_, _069919_, _069920_, _069921_, _069922_, _069923_, _069924_, _069925_, _069926_, _069927_, _069928_, _069929_, _069930_, _069931_, _069932_, _069933_, _069934_, _069935_, _069936_, _069937_, _069938_, _069939_, _069940_, _069941_, _069942_, _069943_, _069944_, _069945_, _069946_, _069947_, _069948_, _069949_, _069950_, _069951_, _069952_, _069953_, _069954_, _069955_, _069956_, _069957_, _069958_, _069959_, _069960_, _069961_, _069962_, _069963_, _069964_, _069965_, _069966_, _069967_, _069968_, _069969_, _069970_, _069971_, _069972_, _069973_, _069974_, _069975_, _069976_, _069977_, _069978_, _069979_, _069980_, _069981_, _069982_, _069983_, _069984_, _069985_, _069986_, _069987_, _069988_, _069989_, _069990_, _069991_, _069992_, _069993_, _069994_, _069995_, _069996_, _069997_, _069998_, _069999_, _070000_, _070001_, _070002_, _070003_, _070004_, _070005_, _070006_, _070007_, _070008_, _070009_, _070010_, _070011_, _070012_, _070013_, _070014_, _070015_, _070016_, _070017_, _070018_, _070019_, _070020_, _070021_, _070022_, _070023_, _070024_, _070025_, _070026_, _070027_, _070028_, _070029_, _070030_, _070031_, _070032_, _070033_, _070034_, _070035_, _070036_, _070037_, _070038_, _070039_, _070040_, _070041_, _070042_, _070043_, _070044_, _070045_, _070046_, _070047_, _070048_, _070049_, _070050_, _070051_, _070052_, _070053_, _070054_, _070055_, _070056_, _070057_, _070058_, _070059_, _070060_, _070061_, _070062_, _070063_, _070064_, _070065_, _070066_, _070067_, _070068_, _070069_, _070070_, _070071_, _070072_, _070073_, _070074_, _070075_, _070076_, _070077_, _070078_, _070079_, _070080_, _070081_, _070082_, _070083_, _070084_, _070085_, _070086_, _070087_, _070088_, _070089_, _070090_, _070091_, _070092_, _070093_, _070094_, _070095_, _070096_, _070097_, _070098_, _070099_, _070100_, _070101_, _070102_, _070103_, _070104_, _070105_, _070106_, _070107_, _070108_, _070109_, _070110_, _070111_, _070112_, _070113_, _070114_, _070115_, _070116_, _070117_, _070118_, _070119_, _070120_, _070121_, _070122_, _070123_, _070124_, _070125_, _070126_, _070127_, _070128_, _070129_, _070130_, _070131_, _070132_, _070133_, _070134_, _070135_, _070136_, _070137_, _070138_, _070139_, _070140_, _070141_, _070142_, _070143_, _070144_, _070145_, _070146_, _070147_, _070148_, _070149_, _070150_, _070151_, _070152_, _070153_, _070154_, _070155_, _070156_, _070157_, _070158_, _070159_, _070160_, _070161_, _070162_, _070163_, _070164_, _070165_, _070166_, _070167_, _070168_, _070169_, _070170_, _070171_, _070172_, _070173_, _070174_, _070175_, _070176_, _070177_, _070178_, _070179_, _070180_, _070181_, _070182_, _070183_, _070184_, _070185_, _070186_, _070187_, _070188_, _070189_, _070190_, _070191_, _070192_, _070193_, _070194_, _070195_, _070196_, _070197_, _070198_, _070199_, _070200_, _070201_, _070202_, _070203_, _070204_, _070205_, _070206_, _070207_, _070208_, _070209_, _070210_, _070211_, _070212_, _070213_, _070214_, _070215_, _070216_, _070217_, _070218_, _070219_, _070220_, _070221_, _070222_, _070223_, _070224_, _070225_, _070226_, _070227_, _070228_, _070229_, _070230_, _070231_, _070232_, _070233_, _070234_, _070235_, _070236_, _070237_, _070238_, _070239_, _070240_, _070241_, _070242_, _070243_, _070244_, _070245_, _070246_, _070247_, _070248_, _070249_, _070250_, _070251_, _070252_, _070253_, _070254_, _070255_, _070256_, _070257_, _070258_, _070259_, _070260_, _070261_, _070262_, _070263_, _070264_, _070265_, _070266_, _070267_, _070268_, _070269_, _070270_, _070271_, _070272_, _070273_, _070274_, _070275_, _070276_, _070277_, _070278_, _070279_, _070280_, _070281_, _070282_, _070283_, _070284_, _070285_, _070286_, _070287_, _070288_, _070289_, _070290_, _070291_, _070292_, _070293_, _070294_, _070295_, _070296_, _070297_, _070298_, _070299_, _070300_, _070301_, _070302_, _070303_, _070304_, _070305_, _070306_, _070307_, _070308_, _070309_, _070310_, _070311_, _070312_, _070313_, _070314_, _070315_, _070316_, _070317_, _070318_, _070319_, _070320_, _070321_, _070322_, _070323_, _070324_, _070325_, _070326_, _070327_, _070328_, _070329_, _070330_, _070331_, _070332_, _070333_, _070334_, _070335_, _070336_, _070337_, _070338_, _070339_, _070340_, _070341_, _070342_, _070343_, _070344_, _070345_, _070346_, _070347_, _070348_, _070349_, _070350_, _070351_, _070352_, _070353_, _070354_, _070355_, _070356_, _070357_, _070358_, _070359_, _070360_, _070361_, _070362_, _070363_, _070364_, _070365_, _070366_, _070367_, _070368_, _070369_, _070370_, _070371_, _070372_, _070373_, _070374_, _070375_, _070376_, _070377_, _070378_, _070379_, _070380_, _070381_, _070382_, _070383_, _070384_, _070385_, _070386_, _070387_, _070388_, _070389_, _070390_, _070391_, _070392_, _070393_, _070394_, _070395_, _070396_, _070397_, _070398_, _070399_, _070400_, _070401_, _070402_, _070403_, _070404_, _070405_, _070406_, _070407_, _070408_, _070409_, _070410_, _070411_, _070412_, _070413_, _070414_, _070415_, _070416_, _070417_, _070418_, _070419_, _070420_, _070421_, _070422_, _070423_, _070424_, _070425_, _070426_, _070427_, _070428_, _070429_, _070430_, _070431_, _070432_, _070433_, _070434_, _070435_, _070436_, _070437_, _070438_, _070439_, _070440_, _070441_, _070442_, _070443_, _070444_, _070445_, _070446_, _070447_, _070448_, _070449_, _070450_, _070451_, _070452_, _070453_, _070454_, _070455_, _070456_, _070457_, _070458_, _070459_, _070460_, _070461_, _070462_, _070463_, _070464_, _070465_, _070466_, _070467_, _070468_, _070469_, _070470_, _070471_, _070472_, _070473_, _070474_, _070475_, _070476_, _070477_, _070478_, _070479_, _070480_, _070481_, _070482_, _070483_, _070484_, _070485_, _070486_, _070487_, _070488_, _070489_, _070490_, _070491_, _070492_, _070493_, _070494_, _070495_, _070496_, _070497_, _070498_, _070499_, _070500_, _070501_, _070502_, _070503_, _070504_, _070505_, _070506_, _070507_, _070508_, _070509_, _070510_, _070511_, _070512_, _070513_, _070514_, _070515_, _070516_, _070517_, _070518_, _070519_, _070520_, _070521_, _070522_, _070523_, _070524_, _070525_, _070526_, _070527_, _070528_, _070529_, _070530_, _070531_, _070532_, _070533_, _070534_, _070535_, _070536_, _070537_, _070538_, _070539_, _070540_, _070541_, _070542_, _070543_, _070544_, _070545_, _070546_, _070547_, _070548_, _070549_, _070550_, _070551_, _070552_, _070553_, _070554_, _070555_, _070556_, _070557_, _070558_, _070559_, _070560_, _070561_, _070562_, _070563_, _070564_, _070565_, _070566_, _070567_, _070568_, _070569_, _070570_, _070571_, _070572_, _070573_, _070574_, _070575_, _070576_, _070577_, _070578_, _070579_, _070580_, _070581_, _070582_, _070583_, _070584_, _070585_, _070586_, _070587_, _070588_, _070589_, _070590_, _070591_, _070592_, _070593_, _070594_, _070595_, _070596_, _070597_, _070598_, _070599_, _070600_, _070601_, _070602_, _070603_, _070604_, _070605_, _070606_, _070607_, _070608_, _070609_, _070610_, _070611_, _070612_, _070613_, _070614_, _070615_, _070616_, _070617_, _070618_, _070619_, _070620_, _070621_, _070622_, _070623_, _070624_, _070625_, _070626_, _070627_, _070628_, _070629_, _070630_, _070631_, _070632_, _070633_, _070634_, _070635_, _070636_, _070637_, _070638_, _070639_, _070640_, _070641_, _070642_, _070643_, _070644_, _070645_, _070646_, _070647_, _070648_, _070649_, _070650_, _070651_, _070652_, _070653_, _070654_, _070655_, _070656_, _070657_, _070658_, _070659_, _070660_, _070661_, _070662_, _070663_, _070664_, _070665_, _070666_, _070667_, _070668_, _070669_, _070670_, _070671_, _070672_, _070673_, _070674_, _070675_, _070676_, _070677_, _070678_, _070679_, _070680_, _070681_, _070682_, _070683_, _070684_, _070685_, _070686_, _070687_, _070688_, _070689_, _070690_, _070691_, _070692_, _070693_, _070694_, _070695_, _070696_, _070697_, _070698_, _070699_, _070700_, _070701_, _070702_, _070703_, _070704_, _070705_, _070706_, _070707_, _070708_, _070709_, _070710_, _070711_, _070712_, _070713_, _070714_, _070715_, _070716_, _070717_, _070718_, _070719_, _070720_, _070721_, _070722_, _070723_, _070724_, _070725_, _070726_, _070727_, _070728_, _070729_, _070730_, _070731_, _070732_, _070733_, _070734_, _070735_, _070736_, _070737_, _070738_, _070739_, _070740_, _070741_, _070742_, _070743_, _070744_, _070745_, _070746_, _070747_, _070748_, _070749_, _070750_, _070751_, _070752_, _070753_, _070754_, _070755_, _070756_, _070757_, _070758_, _070759_, _070760_, _070761_, _070762_, _070763_, _070764_, _070765_, _070766_, _070767_, _070768_, _070769_, _070770_, _070771_, _070772_, _070773_, _070774_, _070775_, _070776_, _070777_, _070778_, _070779_, _070780_, _070781_, _070782_, _070783_, _070784_, _070785_, _070786_, _070787_, _070788_, _070789_, _070790_, _070791_, _070792_, _070793_, _070794_, _070795_, _070796_, _070797_, _070798_, _070799_, _070800_, _070801_, _070802_, _070803_, _070804_, _070805_, _070806_, _070807_, _070808_, _070809_, _070810_, _070811_, _070812_, _070813_, _070814_, _070815_, _070816_, _070817_, _070818_, _070819_, _070820_, _070821_, _070822_, _070823_, _070824_, _070825_, _070826_, _070827_, _070828_, _070829_, _070830_, _070831_, _070832_, _070833_, _070834_, _070835_, _070836_, _070837_, _070838_, _070839_, _070840_, _070841_, _070842_, _070843_, _070844_, _070845_, _070846_, _070847_, _070848_, _070849_, _070850_, _070851_, _070852_, _070853_, _070854_, _070855_, _070856_, _070857_, _070858_, _070859_, _070860_, _070861_, _070862_, _070863_, _070864_, _070865_, _070866_, _070867_, _070868_, _070869_, _070870_, _070871_, _070872_, _070873_, _070874_, _070875_, _070876_, _070877_, _070878_, _070879_, _070880_, _070881_, _070882_, _070883_, _070884_, _070885_, _070886_, _070887_, _070888_, _070889_, _070890_, _070891_, _070892_, _070893_, _070894_, _070895_, _070896_, _070897_, _070898_, _070899_, _070900_, _070901_, _070902_, _070903_, _070904_, _070905_, _070906_, _070907_, _070908_, _070909_, _070910_, _070911_, _070912_, _070913_, _070914_, _070915_, _070916_, _070917_, _070918_, _070919_, _070920_, _070921_, _070922_, _070923_, _070924_, _070925_, _070926_, _070927_, _070928_, _070929_, _070930_, _070931_, _070932_, _070933_, _070934_, _070935_, _070936_, _070937_, _070938_, _070939_, _070940_, _070941_, _070942_, _070943_, _070944_, _070945_, _070946_, _070947_, _070948_, _070949_, _070950_, _070951_, _070952_, _070953_, _070954_, _070955_, _070956_, _070957_, _070958_, _070959_, _070960_, _070961_, _070962_, _070963_, _070964_, _070965_, _070966_, _070967_, _070968_, _070969_, _070970_, _070971_, _070972_, _070973_, _070974_, _070975_, _070976_, _070977_, _070978_, _070979_, _070980_, _070981_, _070982_, _070983_, _070984_, _070985_, _070986_, _070987_, _070988_, _070989_, _070990_, _070991_, _070992_, _070993_, _070994_, _070995_, _070996_, _070997_, _070998_, _070999_, _071000_, _071001_, _071002_, _071003_, _071004_, _071005_, _071006_, _071007_, _071008_, _071009_, _071010_, _071011_, _071012_, _071013_, _071014_, _071015_, _071016_, _071017_, _071018_, _071019_, _071020_, _071021_, _071022_, _071023_, _071024_, _071025_, _071026_, _071027_, _071028_, _071029_, _071030_, _071031_, _071032_, _071033_, _071034_, _071035_, _071036_, _071037_, _071038_, _071039_, _071040_, _071041_, _071042_, _071043_, _071044_, _071045_, _071046_, _071047_, _071048_, _071049_, _071050_, _071051_, _071052_, _071053_, _071054_, _071055_, _071056_, _071057_, _071058_, _071059_, _071060_, _071061_, _071062_, _071063_, _071064_, _071065_, _071066_, _071067_, _071068_, _071069_, _071070_, _071071_, _071072_, _071073_, _071074_, _071075_, _071076_, _071077_, _071078_, _071079_, _071080_, _071081_, _071082_, _071083_, _071084_, _071085_, _071086_, _071087_, _071088_, _071089_, _071090_, _071091_, _071092_, _071093_, _071094_, _071095_, _071096_, _071097_, _071098_, _071099_, _071100_, _071101_, _071102_, _071103_, _071104_, _071105_, _071106_, _071107_, _071108_, _071109_, _071110_, _071111_, _071112_, _071113_, _071114_, _071115_, _071116_, _071117_, _071118_, _071119_, _071120_, _071121_, _071122_, _071123_, _071124_, _071125_, _071126_, _071127_, _071128_, _071129_, _071130_, _071131_, _071132_, _071133_, _071134_, _071135_, _071136_, _071137_, _071138_, _071139_, _071140_, _071141_, _071142_, _071143_, _071144_, _071145_, _071146_, _071147_, _071148_, _071149_, _071150_, _071151_, _071152_, _071153_, _071154_, _071155_, _071156_, _071157_, _071158_, _071159_, _071160_, _071161_, _071162_, _071163_, _071164_, _071165_, _071166_, _071167_, _071168_, _071169_, _071170_, _071171_, _071172_, _071173_, _071174_, _071175_, _071176_, _071177_, _071178_, _071179_, _071180_, _071181_, _071182_, _071183_, _071184_, _071185_, _071186_, _071187_, _071188_, _071189_, _071190_, _071191_, _071192_, _071193_, _071194_, _071195_, _071196_, _071197_, _071198_, _071199_, _071200_, _071201_, _071202_, _071203_, _071204_, _071205_, _071206_, _071207_, _071208_, _071209_, _071210_, _071211_, _071212_, _071213_, _071214_, _071215_, _071216_, _071217_, _071218_, _071219_, _071220_, _071221_, _071222_, _071223_, _071224_, _071225_, _071226_, _071227_, _071228_, _071229_, _071230_, _071231_, _071232_, _071233_, _071234_, _071235_, _071236_, _071237_, _071238_, _071239_, _071240_, _071241_, _071242_, _071243_, _071244_, _071245_, _071246_, _071247_, _071248_, _071249_, _071250_, _071251_, _071252_, _071253_, _071254_, _071255_, _071256_, _071257_, _071258_, _071259_, _071260_, _071261_, _071262_, _071263_, _071264_, _071265_, _071266_, _071267_, _071268_, _071269_, _071270_, _071271_, _071272_, _071273_, _071274_, _071275_, _071276_, _071277_, _071278_, _071279_, _071280_, _071281_, _071282_, _071283_, _071284_, _071285_, _071286_, _071287_, _071288_, _071289_, _071290_, _071291_, _071292_, _071293_, _071294_, _071295_, _071296_, _071297_, _071298_, _071299_, _071300_, _071301_, _071302_, _071303_, _071304_, _071305_, _071306_, _071307_, _071308_, _071309_, _071310_, _071311_, _071312_, _071313_, _071314_, _071315_, _071316_, _071317_, _071318_, _071319_, _071320_, _071321_, _071322_, _071323_, _071324_, _071325_, _071326_, _071327_, _071328_, _071329_, _071330_, _071331_, _071332_, _071333_, _071334_, _071335_, _071336_, _071337_, _071338_, _071339_, _071340_, _071341_, _071342_, _071343_, _071344_, _071345_, _071346_, _071347_, _071348_, _071349_, _071350_, _071351_, _071352_, _071353_, _071354_, _071355_, _071356_, _071357_, _071358_, _071359_, _071360_, _071361_, _071362_, _071363_, _071364_, _071365_, _071366_, _071367_, _071368_, _071369_, _071370_, _071371_, _071372_, _071373_, _071374_, _071375_, _071376_, _071377_, _071378_, _071379_, _071380_, _071381_, _071382_, _071383_, _071384_, _071385_, _071386_, _071387_, _071388_, _071389_, _071390_, _071391_, _071392_, _071393_, _071394_, _071395_, _071396_, _071397_, _071398_, _071399_, _071400_, _071401_, _071402_, _071403_, _071404_, _071405_, _071406_, _071407_, _071408_, _071409_, _071410_, _071411_, _071412_, _071413_, _071414_, _071415_, _071416_, _071417_, _071418_, _071419_, _071420_, _071421_, _071422_, _071423_, _071424_, _071425_, _071426_, _071427_, _071428_, _071429_, _071430_, _071431_, _071432_, _071433_, _071434_, _071435_, _071436_, _071437_, _071438_, _071439_, _071440_, _071441_, _071442_, _071443_, _071444_, _071445_, _071446_, _071447_, _071448_, _071449_, _071450_, _071451_, _071452_, _071453_, _071454_, _071455_, _071456_, _071457_, _071458_, _071459_, _071460_, _071461_, _071462_, _071463_, _071464_, _071465_, _071466_, _071467_, _071468_, _071469_, _071470_, _071471_, _071472_, _071473_, _071474_, _071475_, _071476_, _071477_, _071478_, _071479_, _071480_, _071481_, _071482_, _071483_, _071484_, _071485_, _071486_, _071487_, _071488_, _071489_, _071490_, _071491_, _071492_, _071493_, _071494_, _071495_, _071496_, _071497_, _071498_, _071499_, _071500_, _071501_, _071502_, _071503_, _071504_, _071505_, _071506_, _071507_, _071508_, _071509_, _071510_, _071511_, _071512_, _071513_, _071514_, _071515_, _071516_, _071517_, _071518_, _071519_, _071520_, _071521_, _071522_, _071523_, _071524_, _071525_, _071526_, _071527_, _071528_, _071529_, _071530_, _071531_, _071532_, _071533_, _071534_, _071535_, _071536_, _071537_, _071538_, _071539_, _071540_, _071541_, _071542_, _071543_, _071544_, _071545_, _071546_, _071547_, _071548_, _071549_, _071550_, _071551_, _071552_, _071553_, _071554_, _071555_, _071556_, _071557_, _071558_, _071559_, _071560_, _071561_, _071562_, _071563_, _071564_, _071565_, _071566_, _071567_, _071568_, _071569_, _071570_, _071571_, _071572_, _071573_, _071574_, _071575_, _071576_, _071577_, _071578_, _071579_, _071580_, _071581_, _071582_, _071583_, _071584_, _071585_, _071586_, _071587_, _071588_, _071589_, _071590_, _071591_, _071592_, _071593_, _071594_, _071595_, _071596_, _071597_, _071598_, _071599_, _071600_, _071601_, _071602_, _071603_, _071604_, _071605_, _071606_, _071607_, _071608_, _071609_, _071610_, _071611_, _071612_, _071613_, _071614_, _071615_, _071616_, _071617_, _071618_, _071619_, _071620_, _071621_, _071622_, _071623_, _071624_, _071625_, _071626_, _071627_, _071628_, _071629_, _071630_, _071631_, _071632_, _071633_, _071634_, _071635_, _071636_, _071637_, _071638_, _071639_, _071640_, _071641_, _071642_, _071643_, _071644_, _071645_, _071646_, _071647_, _071648_, _071649_, _071650_, _071651_, _071652_, _071653_, _071654_, _071655_, _071656_, _071657_, _071658_, _071659_, _071660_, _071661_, _071662_, _071663_, _071664_, _071665_, _071666_, _071667_, _071668_, _071669_, _071670_, _071671_, _071672_, _071673_, _071674_, _071675_, _071676_, _071677_, _071678_, _071679_, _071680_, _071681_, _071682_, _071683_, _071684_, _071685_, _071686_, _071687_, _071688_, _071689_, _071690_, _071691_, _071692_, _071693_, _071694_, _071695_, _071696_, _071697_, _071698_, _071699_, _071700_, _071701_, _071702_, _071703_, _071704_, _071705_, _071706_, _071707_, _071708_, _071709_, _071710_, _071711_, _071712_, _071713_, _071714_, _071715_, _071716_, _071717_, _071718_, _071719_, _071720_, _071721_, _071722_, _071723_, _071724_, _071725_, _071726_, _071727_, _071728_, _071729_, _071730_, _071731_, _071732_, _071733_, _071734_, _071735_, _071736_, _071737_, _071738_, _071739_, _071740_, _071741_, _071742_, _071743_, _071744_, _071745_, _071746_, _071747_, _071748_, _071749_, _071750_, _071751_, _071752_, _071753_, _071754_, _071755_, _071756_, _071757_, _071758_, _071759_, _071760_, _071761_, _071762_, _071763_, _071764_, _071765_, _071766_, _071767_, _071768_, _071769_, _071770_, _071771_, _071772_, _071773_, _071774_, _071775_, _071776_, _071777_, _071778_, _071779_, _071780_, _071781_, _071782_, _071783_, _071784_, _071785_, _071786_, _071787_, _071788_, _071789_, _071790_, _071791_, _071792_, _071793_, _071794_, _071795_, _071796_, _071797_, _071798_, _071799_, _071800_, _071801_, _071802_, _071803_, _071804_, _071805_, _071806_, _071807_, _071808_, _071809_, _071810_, _071811_, _071812_, _071813_, _071814_, _071815_, _071816_, _071817_, _071818_, _071819_, _071820_, _071821_, _071822_, _071823_, _071824_, _071825_, _071826_, _071827_, _071828_, _071829_, _071830_, _071831_, _071832_, _071833_, _071834_, _071835_, _071836_, _071837_, _071838_, _071839_, _071840_, _071841_, _071842_, _071843_, _071844_, _071845_, _071846_, _071847_, _071848_, _071849_, _071850_, _071851_, _071852_, _071853_, _071854_, _071855_, _071856_, _071857_, _071858_, _071859_, _071860_, _071861_, _071862_, _071863_, _071864_, _071865_, _071866_, _071867_, _071868_, _071869_, _071870_, _071871_, _071872_, _071873_, _071874_, _071875_, _071876_, _071877_, _071878_, _071879_, _071880_, _071881_, _071882_, _071883_, _071884_, _071885_, _071886_, _071887_, _071888_, _071889_, _071890_, _071891_, _071892_, _071893_, _071894_, _071895_, _071896_, _071897_, _071898_, _071899_, _071900_, _071901_, _071902_, _071903_, _071904_, _071905_, _071906_, _071907_, _071908_, _071909_, _071910_, _071911_, _071912_, _071913_, _071914_, _071915_, _071916_, _071917_, _071918_, _071919_, _071920_, _071921_, _071922_, _071923_, _071924_, _071925_, _071926_, _071927_, _071928_, _071929_, _071930_, _071931_, _071932_, _071933_, _071934_, _071935_, _071936_, _071937_, _071938_, _071939_, _071940_, _071941_, _071942_, _071943_, _071944_, _071945_, _071946_, _071947_, _071948_, _071949_, _071950_, _071951_, _071952_, _071953_, _071954_, _071955_, _071956_, _071957_, _071958_, _071959_, _071960_, _071961_, _071962_, _071963_, _071964_, _071965_, _071966_, _071967_, _071968_, _071969_, _071970_, _071971_, _071972_, _071973_, _071974_, _071975_, _071976_, _071977_, _071978_, _071979_, _071980_, _071981_, _071982_, _071983_, _071984_, _071985_, _071986_, _071987_, _071988_, _071989_, _071990_, _071991_, _071992_, _071993_, _071994_, _071995_, _071996_, _071997_, _071998_, _071999_, _072000_, _072001_, _072002_, _072003_, _072004_, _072005_, _072006_, _072007_, _072008_, _072009_, _072010_, _072011_, _072012_, _072013_, _072014_, _072015_, _072016_, _072017_, _072018_, _072019_, _072020_, _072021_, _072022_, _072023_, _072024_, _072025_, _072026_, _072027_, _072028_, _072029_, _072030_, _072031_, _072032_, _072033_, _072034_, _072035_, _072036_, _072037_, _072038_, _072039_, _072040_, _072041_, _072042_, _072043_, _072044_, _072045_, _072046_, _072047_, _072048_, _072049_, _072050_, _072051_, _072052_, _072053_, _072054_, _072055_, _072056_, _072057_, _072058_, _072059_, _072060_, _072061_, _072062_, _072063_, _072064_, _072065_, _072066_, _072067_, _072068_, _072069_, _072070_, _072071_, _072072_, _072073_, _072074_, _072075_, _072076_, _072077_, _072078_, _072079_, _072080_, _072081_, _072082_, _072083_, _072084_, _072085_, _072086_, _072087_, _072088_, _072089_, _072090_, _072091_, _072092_, _072093_, _072094_, _072095_, _072096_, _072097_, _072098_, _072099_, _072100_, _072101_, _072102_, _072103_, _072104_, _072105_, _072106_, _072107_, _072108_, _072109_, _072110_, _072111_, _072112_, _072113_, _072114_, _072115_, _072116_, _072117_, _072118_, _072119_, _072120_, _072121_, _072122_, _072123_, _072124_, _072125_, _072126_, _072127_, _072128_, _072129_, _072130_, _072131_, _072132_, _072133_, _072134_, _072135_, _072136_, _072137_, _072138_, _072139_, _072140_, _072141_, _072142_, _072143_, _072144_, _072145_, _072146_, _072147_, _072148_, _072149_, _072150_, _072151_, _072152_, _072153_, _072154_, _072155_, _072156_, _072157_, _072158_, _072159_, _072160_, _072161_, _072162_, _072163_, _072164_, _072165_, _072166_, _072167_, _072168_, _072169_, _072170_, _072171_, _072172_, _072173_, _072174_, _072175_, _072176_, _072177_, _072178_, _072179_, _072180_, _072181_, _072182_, _072183_, _072184_, _072185_, _072186_, _072187_, _072188_, _072189_, _072190_, _072191_, _072192_, _072193_, _072194_, _072195_, _072196_, _072197_, _072198_, _072199_, _072200_, _072201_, _072202_, _072203_, _072204_, _072205_, _072206_, _072207_, _072208_, _072209_, _072210_, _072211_, _072212_, _072213_, _072214_, _072215_, _072216_, _072217_, _072218_, _072219_, _072220_, _072221_, _072222_, _072223_, _072224_, _072225_, _072226_, _072227_, _072228_, _072229_, _072230_, _072231_, _072232_, _072233_, _072234_, _072235_, _072236_, _072237_, _072238_, _072239_, _072240_, _072241_, _072242_, _072243_, _072244_, _072245_, _072246_, _072247_, _072248_, _072249_, _072250_, _072251_, _072252_, _072253_, _072254_, _072255_, _072256_, _072257_, _072258_, _072259_, _072260_, _072261_, _072262_, _072263_, _072264_, _072265_, _072266_, _072267_, _072268_, _072269_, _072270_, _072271_, _072272_, _072273_, _072274_, _072275_, _072276_, _072277_, _072278_, _072279_, _072280_, _072281_, _072282_, _072283_, _072284_, _072285_, _072286_, _072287_, _072288_, _072289_, _072290_, _072291_, _072292_, _072293_, _072294_, _072295_, _072296_, _072297_, _072298_, _072299_, _072300_, _072301_, _072302_, _072303_, _072304_, _072305_, _072306_, _072307_, _072308_, _072309_, _072310_, _072311_, _072312_, _072313_, _072314_, _072315_, _072316_, _072317_, _072318_, _072319_, _072320_, _072321_, _072322_, _072323_, _072324_, _072325_, _072326_, _072327_, _072328_, _072329_, _072330_, _072331_, _072332_, _072333_, _072334_, _072335_, _072336_, _072337_, _072338_, _072339_, _072340_, _072341_, _072342_, _072343_, _072344_, _072345_, _072346_, _072347_, _072348_, _072349_, _072350_, _072351_, _072352_, _072353_, _072354_, _072355_, _072356_, _072357_, _072358_, _072359_, _072360_, _072361_, _072362_, _072363_, _072364_, _072365_, _072366_, _072367_, _072368_, _072369_, _072370_, _072371_, _072372_, _072373_, _072374_, _072375_, _072376_, _072377_, _072378_, _072379_, _072380_, _072381_, _072382_, _072383_, _072384_, _072385_, _072386_, _072387_, _072388_, _072389_, _072390_, _072391_, _072392_, _072393_, _072394_, _072395_, _072396_, _072397_, _072398_, _072399_, _072400_, _072401_, _072402_, _072403_, _072404_, _072405_, _072406_, _072407_, _072408_, _072409_, _072410_, _072411_, _072412_, _072413_, _072414_, _072415_, _072416_, _072417_, _072418_, _072419_, _072420_, _072421_, _072422_, _072423_, _072424_, _072425_, _072426_, _072427_, _072428_, _072429_, _072430_, _072431_, _072432_, _072433_, _072434_, _072435_, _072436_, _072437_, _072438_, _072439_, _072440_, _072441_, _072442_, _072443_, _072444_, _072445_, _072446_, _072447_, _072448_, _072449_, _072450_, _072451_, _072452_, _072453_, _072454_, _072455_, _072456_, _072457_, _072458_, _072459_, _072460_, _072461_, _072462_, _072463_, _072464_, _072465_, _072466_, _072467_, _072468_, _072469_, _072470_, _072471_, _072472_, _072473_, _072474_, _072475_, _072476_, _072477_, _072478_, _072479_, _072480_, _072481_, _072482_, _072483_, _072484_, _072485_, _072486_, _072487_, _072488_, _072489_, _072490_, _072491_, _072492_, _072493_, _072494_, _072495_, _072496_, _072497_, _072498_, _072499_, _072500_, _072501_, _072502_, _072503_, _072504_, _072505_, _072506_, _072507_, _072508_, _072509_, _072510_, _072511_, _072512_, _072513_, _072514_, _072515_, _072516_, _072517_, _072518_, _072519_, _072520_, _072521_, _072522_, _072523_, _072524_, _072525_, _072526_, _072527_, _072528_, _072529_, _072530_, _072531_, _072532_, _072533_, _072534_, _072535_, _072536_, _072537_, _072538_, _072539_, _072540_, _072541_, _072542_, _072543_, _072544_, _072545_, _072546_, _072547_, _072548_, _072549_, _072550_, _072551_, _072552_, _072553_, _072554_, _072555_, _072556_, _072557_, _072558_, _072559_, _072560_, _072561_, _072562_, _072563_, _072564_, _072565_, _072566_, _072567_, _072568_, _072569_, _072570_, _072571_, _072572_, _072573_, _072574_, _072575_, _072576_, _072577_, _072578_, _072579_, _072580_, _072581_, _072582_, _072583_, _072584_, _072585_, _072586_, _072587_, _072588_, _072589_, _072590_, _072591_, _072592_, _072593_, _072594_, _072595_, _072596_, _072597_, _072598_, _072599_, _072600_, _072601_, _072602_, _072603_, _072604_, _072605_, _072606_, _072607_, _072608_, _072609_, _072610_, _072611_, _072612_, _072613_, _072614_, _072615_, _072616_, _072617_, _072618_, _072619_, _072620_, _072621_, _072622_, _072623_, _072624_, _072625_, _072626_, _072627_, _072628_, _072629_, _072630_, _072631_, _072632_, _072633_, _072634_, _072635_, _072636_, _072637_, _072638_, _072639_, _072640_, _072641_, _072642_, _072643_, _072644_, _072645_, _072646_, _072647_, _072648_, _072649_, _072650_, _072651_, _072652_, _072653_, _072654_, _072655_, _072656_, _072657_, _072658_, _072659_, _072660_, _072661_, _072662_, _072663_, _072664_, _072665_, _072666_, _072667_, _072668_, _072669_, _072670_, _072671_, _072672_, _072673_, _072674_, _072675_, _072676_, _072677_, _072678_, _072679_, _072680_, _072681_, _072682_, _072683_, _072684_, _072685_, _072686_, _072687_, _072688_, _072689_, _072690_, _072691_, _072692_, _072693_, _072694_, _072695_, _072696_, _072697_, _072698_, _072699_, _072700_, _072701_, _072702_, _072703_, _072704_, _072705_, _072706_, _072707_, _072708_, _072709_, _072710_, _072711_, _072712_, _072713_, _072714_, _072715_, _072716_, _072717_, _072718_, _072719_, _072720_, _072721_, _072722_, _072723_, _072724_, _072725_, _072726_, _072727_, _072728_, _072729_, _072730_, _072731_, _072732_, _072733_, _072734_, _072735_, _072736_, _072737_, _072738_, _072739_, _072740_, _072741_, _072742_, _072743_, _072744_, _072745_, _072746_, _072747_, _072748_, _072749_, _072750_, _072751_, _072752_, _072753_, _072754_, _072755_, _072756_, _072757_, _072758_, _072759_, _072760_, _072761_, _072762_, _072763_, _072764_, _072765_, _072766_, _072767_, _072768_, _072769_, _072770_, _072771_, _072772_, _072773_, _072774_, _072775_, _072776_, _072777_, _072778_, _072779_, _072780_, _072781_, _072782_, _072783_, _072784_, _072785_, _072786_, _072787_, _072788_, _072789_, _072790_, _072791_, _072792_, _072793_, _072794_, _072795_, _072796_, _072797_, _072798_, _072799_, _072800_, _072801_, _072802_, _072803_, _072804_, _072805_, _072806_, _072807_, _072808_, _072809_, _072810_, _072811_, _072812_, _072813_, _072814_, _072815_, _072816_, _072817_, _072818_, _072819_, _072820_, _072821_, _072822_, _072823_, _072824_, _072825_, _072826_, _072827_, _072828_, _072829_, _072830_, _072831_, _072832_, _072833_, _072834_, _072835_, _072836_, _072837_, _072838_, _072839_, _072840_, _072841_, _072842_, _072843_, _072844_, _072845_, _072846_, _072847_, _072848_, _072849_, _072850_, _072851_, _072852_, _072853_, _072854_, _072855_, _072856_, _072857_, _072858_, _072859_, _072860_, _072861_, _072862_, _072863_, _072864_, _072865_, _072866_, _072867_, _072868_, _072869_, _072870_, _072871_, _072872_, _072873_, _072874_, _072875_, _072876_, _072877_, _072878_, _072879_, _072880_, _072881_, _072882_, _072883_, _072884_, _072885_, _072886_, _072887_, _072888_, _072889_, _072890_, _072891_, _072892_, _072893_, _072894_, _072895_, _072896_, _072897_, _072898_, _072899_, _072900_, _072901_, _072902_, _072903_, _072904_, _072905_, _072906_, _072907_, _072908_, _072909_, _072910_, _072911_, _072912_, _072913_, _072914_, _072915_, _072916_, _072917_, _072918_, _072919_, _072920_, _072921_, _072922_, _072923_, _072924_, _072925_, _072926_, _072927_, _072928_, _072929_, _072930_, _072931_, _072932_, _072933_, _072934_, _072935_, _072936_, _072937_, _072938_, _072939_, _072940_, _072941_, _072942_, _072943_, _072944_, _072945_, _072946_, _072947_, _072948_, _072949_, _072950_, _072951_, _072952_, _072953_, _072954_, _072955_, _072956_, _072957_, _072958_, _072959_, _072960_, _072961_, _072962_, _072963_, _072964_, _072965_, _072966_, _072967_, _072968_, _072969_, _072970_, _072971_, _072972_, _072973_, _072974_, _072975_, _072976_, _072977_, _072978_, _072979_, _072980_, _072981_, _072982_, _072983_, _072984_, _072985_, _072986_, _072987_, _072988_, _072989_, _072990_, _072991_, _072992_, _072993_, _072994_, _072995_, _072996_, _072997_, _072998_, _072999_, _073000_, _073001_, _073002_, _073003_, _073004_, _073005_, _073006_, _073007_, _073008_, _073009_, _073010_, _073011_, _073012_, _073013_, _073014_, _073015_, _073016_, _073017_, _073018_, _073019_, _073020_, _073021_, _073022_, _073023_, _073024_, _073025_, _073026_, _073027_, _073028_, _073029_, _073030_, _073031_, _073032_, _073033_, _073034_, _073035_, _073036_, _073037_, _073038_, _073039_, _073040_, _073041_, _073042_, _073043_, _073044_, _073045_, _073046_, _073047_, _073048_, _073049_, _073050_, _073051_, _073052_, _073053_, _073054_, _073055_, _073056_, _073057_, _073058_, _073059_, _073060_, _073061_, _073062_, _073063_, _073064_, _073065_, _073066_, _073067_, _073068_, _073069_, _073070_, _073071_, _073072_, _073073_, _073074_, _073075_, _073076_, _073077_, _073078_, _073079_, _073080_, _073081_, _073082_, _073083_, _073084_, _073085_, _073086_, _073087_, _073088_, _073089_, _073090_, _073091_, _073092_, _073093_, _073094_, _073095_, _073096_, _073097_, _073098_, _073099_, _073100_, _073101_, _073102_, _073103_, _073104_, _073105_, _073106_, _073107_, _073108_, _073109_, _073110_, _073111_, _073112_, _073113_, _073114_, _073115_, _073116_, _073117_, _073118_, _073119_, _073120_, _073121_, _073122_, _073123_, _073124_, _073125_, _073126_, _073127_, _073128_, _073129_, _073130_, _073131_, _073132_, _073133_, _073134_, _073135_, _073136_, _073137_, _073138_, _073139_, _073140_, _073141_, _073142_, _073143_, _073144_, _073145_, _073146_, _073147_, _073148_, _073149_, _073150_, _073151_, _073152_, _073153_, _073154_, _073155_, _073156_, _073157_, _073158_, _073159_, _073160_, _073161_, _073162_, _073163_, _073164_, _073165_, _073166_, _073167_, _073168_, _073169_, _073170_, _073171_, _073172_, _073173_, _073174_, _073175_, _073176_, _073177_, _073178_, _073179_, _073180_, _073181_, _073182_, _073183_, _073184_, _073185_, _073186_, _073187_, _073188_, _073189_, _073190_, _073191_, _073192_, _073193_, _073194_, _073195_, _073196_, _073197_, _073198_, _073199_, _073200_, _073201_, _073202_, _073203_, _073204_, _073205_, _073206_, _073207_, _073208_, _073209_, _073210_, _073211_, _073212_, _073213_, _073214_, _073215_, _073216_, _073217_, _073218_, _073219_, _073220_, _073221_, _073222_, _073223_, _073224_, _073225_, _073226_, _073227_, _073228_, _073229_, _073230_, _073231_, _073232_, _073233_, _073234_, _073235_, _073236_, _073237_, _073238_, _073239_, _073240_, _073241_, _073242_, _073243_, _073244_, _073245_, _073246_, _073247_, _073248_, _073249_, _073250_, _073251_, _073252_, _073253_, _073254_, _073255_, _073256_, _073257_, _073258_, _073259_, _073260_, _073261_, _073262_, _073263_, _073264_, _073265_, _073266_, _073267_, _073268_, _073269_, _073270_, _073271_, _073272_, _073273_, _073274_, _073275_, _073276_, _073277_, _073278_, _073279_, _073280_, _073281_, _073282_, _073283_, _073284_, _073285_, _073286_, _073287_, _073288_, _073289_, _073290_, _073291_, _073292_, _073293_, _073294_, _073295_, _073296_, _073297_, _073298_, _073299_, _073300_, _073301_, _073302_, _073303_, _073304_, _073305_, _073306_, _073307_, _073308_, _073309_, _073310_, _073311_, _073312_, _073313_, _073314_, _073315_, _073316_, _073317_, _073318_, _073319_, _073320_, _073321_, _073322_, _073323_, _073324_, _073325_, _073326_, _073327_, _073328_, _073329_, _073330_, _073331_, _073332_, _073333_, _073334_, _073335_, _073336_, _073337_, _073338_, _073339_, _073340_, _073341_, _073342_, _073343_, _073344_, _073345_, _073346_, _073347_, _073348_, _073349_, _073350_, _073351_, _073352_, _073353_, _073354_, _073355_, _073356_, _073357_, _073358_, _073359_, _073360_, _073361_, _073362_, _073363_, _073364_, _073365_, _073366_, _073367_, _073368_, _073369_, _073370_, _073371_, _073372_, _073373_, _073374_, _073375_, _073376_, _073377_, _073378_, _073379_, _073380_, _073381_, _073382_, _073383_, _073384_, _073385_, _073386_, _073387_, _073388_, _073389_, _073390_, _073391_, _073392_, _073393_, _073394_, _073395_, _073396_, _073397_, _073398_, _073399_, _073400_, _073401_, _073402_, _073403_, _073404_, _073405_, _073406_, _073407_, _073408_, _073409_, _073410_, _073411_, _073412_, _073413_, _073414_, _073415_, _073416_, _073417_, _073418_, _073419_, _073420_, _073421_, _073422_, _073423_, _073424_, _073425_, _073426_, _073427_, _073428_, _073429_, _073430_, _073431_, _073432_, _073433_, _073434_, _073435_, _073436_, _073437_, _073438_, _073439_, _073440_, _073441_, _073442_, _073443_, _073444_, _073445_, _073446_, _073447_, _073448_, _073449_, _073450_, _073451_, _073452_, _073453_, _073454_, _073455_, _073456_, _073457_, _073458_, _073459_, _073460_, _073461_, _073462_, _073463_, _073464_, _073465_, _073466_, _073467_, _073468_, _073469_, _073470_, _073471_, _073472_, _073473_, _073474_, _073475_, _073476_, _073477_, _073478_, _073479_, _073480_, _073481_, _073482_, _073483_, _073484_, _073485_, _073486_, _073487_, _073488_, _073489_, _073490_, _073491_, _073492_, _073493_, _073494_, _073495_, _073496_, _073497_, _073498_, _073499_, _073500_, _073501_, _073502_, _073503_, _073504_, _073505_, _073506_, _073507_, _073508_, _073509_, _073510_, _073511_, _073512_, _073513_, _073514_, _073515_, _073516_, _073517_, _073518_, _073519_, _073520_, _073521_, _073522_, _073523_, _073524_, _073525_, _073526_, _073527_, _073528_, _073529_, _073530_, _073531_, _073532_, _073533_, _073534_, _073535_, _073536_, _073537_, _073538_, _073539_, _073540_, _073541_, _073542_, _073543_, _073544_, _073545_, _073546_, _073547_, _073548_, _073549_, _073550_, _073551_, _073552_, _073553_, _073554_, _073555_, _073556_, _073557_, _073558_, _073559_, _073560_, _073561_, _073562_, _073563_, _073564_, _073565_, _073566_, _073567_, _073568_, _073569_, _073570_, _073571_, _073572_, _073573_, _073574_, _073575_, _073576_, _073577_, _073578_, _073579_, _073580_, _073581_, _073582_, _073583_, _073584_, _073585_, _073586_, _073587_, _073588_, _073589_, _073590_, _073591_, _073592_, _073593_, _073594_, _073595_, _073596_, _073597_, _073598_, _073599_, _073600_, _073601_, _073602_, _073603_, _073604_, _073605_, _073606_, _073607_, _073608_, _073609_, _073610_, _073611_, _073612_, _073613_, _073614_, _073615_, _073616_, _073617_, _073618_, _073619_, _073620_, _073621_, _073622_, _073623_, _073624_, _073625_, _073626_, _073627_, _073628_, _073629_, _073630_, _073631_, _073632_, _073633_, _073634_, _073635_, _073636_, _073637_, _073638_, _073639_, _073640_, _073641_, _073642_, _073643_, _073644_, _073645_, _073646_, _073647_, _073648_, _073649_, _073650_, _073651_, _073652_, _073653_, _073654_, _073655_, _073656_, _073657_, _073658_, _073659_, _073660_, _073661_, _073662_, _073663_, _073664_, _073665_, _073666_, _073667_, _073668_, _073669_, _073670_, _073671_, _073672_, _073673_, _073674_, _073675_, _073676_, _073677_, _073678_, _073679_, _073680_, _073681_, _073682_, _073683_, _073684_, _073685_, _073686_, _073687_, _073688_, _073689_, _073690_, _073691_, _073692_, _073693_, _073694_, _073695_, _073696_, _073697_, _073698_, _073699_, _073700_, _073701_, _073702_, _073703_, _073704_, _073705_, _073706_, _073707_, _073708_, _073709_, _073710_, _073711_, _073712_, _073713_, _073714_, _073715_, _073716_, _073717_, _073718_, _073719_, _073720_, _073721_, _073722_, _073723_, _073724_, _073725_, _073726_, _073727_, _073728_, _073729_, _073730_, _073731_, _073732_, _073733_, _073734_, _073735_, _073736_, _073737_, _073738_, _073739_, _073740_, _073741_, _073742_, _073743_, _073744_, _073745_, _073746_, _073747_, _073748_, _073749_, _073750_, _073751_, _073752_, _073753_, _073754_, _073755_, _073756_, _073757_, _073758_, _073759_, _073760_, _073761_, _073762_, _073763_, _073764_, _073765_, _073766_, _073767_, _073768_, _073769_, _073770_, _073771_, _073772_, _073773_, _073774_, _073775_, _073776_, _073777_, _073778_, _073779_, _073780_, _073781_, _073782_, _073783_, _073784_, _073785_, _073786_, _073787_, _073788_, _073789_, _073790_, _073791_, _073792_, _073793_, _073794_, _073795_, _073796_, _073797_, _073798_, _073799_, _073800_, _073801_, _073802_, _073803_, _073804_, _073805_, _073806_, _073807_, _073808_, _073809_, _073810_, _073811_, _073812_, _073813_, _073814_, _073815_, _073816_, _073817_, _073818_, _073819_, _073820_, _073821_, _073822_, _073823_, _073824_, _073825_, _073826_, _073827_, _073828_, _073829_, _073830_, _073831_, _073832_, _073833_, _073834_, _073835_, _073836_, _073837_, _073838_, _073839_, _073840_, _073841_, _073842_, _073843_, _073844_, _073845_, _073846_, _073847_, _073848_, _073849_, _073850_, _073851_, _073852_, _073853_, _073854_, _073855_, _073856_, _073857_, _073858_, _073859_, _073860_, _073861_, _073862_, _073863_, _073864_, _073865_, _073866_, _073867_, _073868_, _073869_, _073870_, _073871_, _073872_, _073873_, _073874_, _073875_, _073876_, _073877_, _073878_, _073879_, _073880_, _073881_, _073882_, _073883_, _073884_, _073885_, _073886_, _073887_, _073888_, _073889_, _073890_, _073891_, _073892_, _073893_, _073894_, _073895_, _073896_, _073897_, _073898_, _073899_, _073900_, _073901_, _073902_, _073903_, _073904_, _073905_, _073906_, _073907_, _073908_, _073909_, _073910_, _073911_, _073912_, _073913_, _073914_, _073915_, _073916_, _073917_, _073918_, _073919_, _073920_, _073921_, _073922_, _073923_, _073924_, _073925_, _073926_, _073927_, _073928_, _073929_, _073930_, _073931_, _073932_, _073933_, _073934_, _073935_, _073936_, _073937_, _073938_, _073939_, _073940_, _073941_, _073942_, _073943_, _073944_, _073945_, _073946_, _073947_, _073948_, _073949_, _073950_, _073951_, _073952_, _073953_, _073954_, _073955_, _073956_, _073957_, _073958_, _073959_, _073960_, _073961_, _073962_, _073963_, _073964_, _073965_, _073966_, _073967_, _073968_, _073969_, _073970_, _073971_, _073972_, _073973_, _073974_, _073975_, _073976_, _073977_, _073978_, _073979_, _073980_, _073981_, _073982_, _073983_, _073984_, _073985_, _073986_, _073987_, _073988_, _073989_, _073990_, _073991_, _073992_, _073993_, _073994_, _073995_, _073996_, _073997_, _073998_, _073999_, _074000_, _074001_, _074002_, _074003_, _074004_, _074005_, _074006_, _074007_, _074008_, _074009_, _074010_, _074011_, _074012_, _074013_, _074014_, _074015_, _074016_, _074017_, _074018_, _074019_, _074020_, _074021_, _074022_, _074023_, _074024_, _074025_, _074026_, _074027_, _074028_, _074029_, _074030_, _074031_, _074032_, _074033_, _074034_, _074035_, _074036_, _074037_, _074038_, _074039_, _074040_, _074041_, _074042_, _074043_, _074044_, _074045_, _074046_, _074047_, _074048_, _074049_, _074050_, _074051_, _074052_, _074053_, _074054_, _074055_, _074056_, _074057_, _074058_, _074059_, _074060_, _074061_, _074062_, _074063_, _074064_, _074065_, _074066_, _074067_, _074068_, _074069_, _074070_, _074071_, _074072_, _074073_, _074074_, _074075_, _074076_, _074077_, _074078_, _074079_, _074080_, _074081_, _074082_, _074083_, _074084_, _074085_, _074086_, _074087_, _074088_, _074089_, _074090_, _074091_, _074092_, _074093_, _074094_, _074095_, _074096_, _074097_, _074098_, _074099_, _074100_, _074101_, _074102_, _074103_, _074104_, _074105_, _074106_, _074107_, _074108_, _074109_, _074110_, _074111_, _074112_, _074113_, _074114_, _074115_, _074116_, _074117_, _074118_, _074119_, _074120_, _074121_, _074122_, _074123_, _074124_, _074125_, _074126_, _074127_, _074128_, _074129_, _074130_, _074131_, _074132_, _074133_, _074134_, _074135_, _074136_, _074137_, _074138_, _074139_, _074140_, _074141_, _074142_, _074143_, _074144_, _074145_, _074146_, _074147_, _074148_, _074149_, _074150_, _074151_, _074152_, _074153_, _074154_, _074155_, _074156_, _074157_, _074158_, _074159_, _074160_, _074161_, _074162_, _074163_, _074164_, _074165_, _074166_, _074167_, _074168_, _074169_, _074170_, _074171_, _074172_, _074173_, _074174_, _074175_, _074176_, _074177_, _074178_, _074179_, _074180_, _074181_, _074182_, _074183_, _074184_, _074185_, _074186_, _074187_, _074188_, _074189_, _074190_, _074191_, _074192_, _074193_, _074194_, _074195_, _074196_, _074197_, _074198_, _074199_, _074200_, _074201_, _074202_, _074203_, _074204_, _074205_, _074206_, _074207_, _074208_, _074209_, _074210_, _074211_, _074212_, _074213_, _074214_, _074215_, _074216_, _074217_, _074218_, _074219_, _074220_, _074221_, _074222_, _074223_, _074224_, _074225_, _074226_, _074227_, _074228_, _074229_, _074230_, _074231_, _074232_, _074233_, _074234_, _074235_, _074236_, _074237_, _074238_, _074239_, _074240_, _074241_, _074242_, _074243_, _074244_, _074245_, _074246_, _074247_, _074248_, _074249_, _074250_, _074251_, _074252_, _074253_, _074254_, _074255_, _074256_, _074257_, _074258_, _074259_, _074260_, _074261_, _074262_, _074263_, _074264_, _074265_, _074266_, _074267_, _074268_, _074269_, _074270_, _074271_, _074272_, _074273_, _074274_, _074275_, _074276_, _074277_, _074278_, _074279_, _074280_, _074281_, _074282_, _074283_, _074284_, _074285_, _074286_, _074287_, _074288_, _074289_, _074290_, _074291_, _074292_, _074293_, _074294_, _074295_, _074296_, _074297_, _074298_, _074299_, _074300_, _074301_, _074302_, _074303_, _074304_, _074305_, _074306_, _074307_, _074308_, _074309_, _074310_, _074311_, _074312_, _074313_, _074314_, _074315_, _074316_, _074317_, _074318_, _074319_, _074320_, _074321_, _074322_, _074323_, _074324_, _074325_, _074326_, _074327_, _074328_, _074329_, _074330_, _074331_, _074332_, _074333_, _074334_, _074335_, _074336_, _074337_, _074338_, _074339_, _074340_, _074341_, _074342_, _074343_, _074344_, _074345_, _074346_, _074347_, _074348_, _074349_, _074350_, _074351_, _074352_, _074353_, _074354_, _074355_, _074356_, _074357_, _074358_, _074359_, _074360_, _074361_, _074362_, _074363_, _074364_, _074365_, _074366_, _074367_, _074368_, _074369_, _074370_, _074371_, _074372_, _074373_, _074374_, _074375_, _074376_, _074377_, _074378_, _074379_, _074380_, _074381_, _074382_, _074383_, _074384_, _074385_, _074386_, _074387_, _074388_, _074389_, _074390_, _074391_, _074392_, _074393_, _074394_, _074395_, _074396_, _074397_, _074398_, _074399_, _074400_, _074401_, _074402_, _074403_, _074404_, _074405_, _074406_, _074407_, _074408_, _074409_, _074410_, _074411_, _074412_, _074413_, _074414_, _074415_, _074416_, _074417_, _074418_, _074419_, _074420_, _074421_, _074422_, _074423_, _074424_, _074425_, _074426_, _074427_, _074428_, _074429_, _074430_, _074431_, _074432_, _074433_, _074434_, _074435_, _074436_, _074437_, _074438_, _074439_, _074440_, _074441_, _074442_, _074443_, _074444_, _074445_, _074446_, _074447_, _074448_, _074449_, _074450_, _074451_, _074452_, _074453_, _074454_, _074455_, _074456_, _074457_, _074458_, _074459_, _074460_, _074461_, _074462_, _074463_, _074464_, _074465_, _074466_, _074467_, _074468_, _074469_, _074470_, _074471_, _074472_, _074473_, _074474_, _074475_, _074476_, _074477_, _074478_, _074479_, _074480_, _074481_, _074482_, _074483_, _074484_, _074485_, _074486_, _074487_, _074488_, _074489_, _074490_, _074491_, _074492_, _074493_, _074494_, _074495_, _074496_, _074497_, _074498_, _074499_, _074500_, _074501_, _074502_, _074503_, _074504_, _074505_, _074506_, _074507_, _074508_, _074509_, _074510_, _074511_, _074512_, _074513_, _074514_, _074515_, _074516_, _074517_, _074518_, _074519_, _074520_, _074521_, _074522_, _074523_, _074524_, _074525_, _074526_, _074527_, _074528_, _074529_, _074530_, _074531_, _074532_, _074533_, _074534_, _074535_, _074536_, _074537_, _074538_, _074539_, _074540_, _074541_, _074542_, _074543_, _074544_, _074545_, _074546_, _074547_, _074548_, _074549_, _074550_, _074551_, _074552_, _074553_, _074554_, _074555_, _074556_, _074557_, _074558_, _074559_, _074560_, _074561_, _074562_, _074563_, _074564_, _074565_, _074566_, _074567_, _074568_, _074569_, _074570_, _074571_, _074572_, _074573_, _074574_, _074575_, _074576_, _074577_, _074578_, _074579_, _074580_, _074581_, _074582_, _074583_, _074584_, _074585_, _074586_, _074587_, _074588_, _074589_, _074590_, _074591_, _074592_, _074593_, _074594_, _074595_, _074596_, _074597_, _074598_, _074599_, _074600_, _074601_, _074602_, _074603_, _074604_, _074605_, _074606_, _074607_, _074608_, _074609_, _074610_, _074611_, _074612_, _074613_, _074614_, _074615_, _074616_, _074617_, _074618_, _074619_, _074620_, _074621_, _074622_, _074623_, _074624_, _074625_, _074626_, _074627_, _074628_, _074629_, _074630_, _074631_, _074632_, _074633_, _074634_, _074635_, _074636_, _074637_, _074638_, _074639_, _074640_, _074641_, _074642_, _074643_, _074644_, _074645_, _074646_, _074647_, _074648_, _074649_, _074650_, _074651_, _074652_, _074653_, _074654_, _074655_, _074656_, _074657_, _074658_, _074659_, _074660_, _074661_, _074662_, _074663_, _074664_, _074665_, _074666_, _074667_, _074668_, _074669_, _074670_, _074671_, _074672_, _074673_, _074674_, _074675_, _074676_, _074677_, _074678_, _074679_, _074680_, _074681_, _074682_, _074683_, _074684_, _074685_, _074686_, _074687_, _074688_, _074689_, _074690_, _074691_, _074692_, _074693_, _074694_, _074695_, _074696_, _074697_, _074698_, _074699_, _074700_, _074701_, _074702_, _074703_, _074704_, _074705_, _074706_, _074707_, _074708_, _074709_, _074710_, _074711_, _074712_, _074713_, _074714_, _074715_, _074716_, _074717_, _074718_, _074719_, _074720_, _074721_, _074722_, _074723_, _074724_, _074725_, _074726_, _074727_, _074728_, _074729_, _074730_, _074731_, _074732_, _074733_, _074734_, _074735_, _074736_, _074737_, _074738_, _074739_, _074740_, _074741_, _074742_, _074743_, _074744_, _074745_, _074746_, _074747_, _074748_, _074749_, _074750_, _074751_, _074752_, _074753_, _074754_, _074755_, _074756_, _074757_, _074758_, _074759_, _074760_, _074761_, _074762_, _074763_, _074764_, _074765_, _074766_, _074767_, _074768_, _074769_, _074770_, _074771_, _074772_, _074773_, _074774_, _074775_, _074776_, _074777_, _074778_, _074779_, _074780_, _074781_, _074782_, _074783_, _074784_, _074785_, _074786_, _074787_, _074788_, _074789_, _074790_, _074791_, _074792_, _074793_, _074794_, _074795_, _074796_, _074797_, _074798_, _074799_, _074800_, _074801_, _074802_, _074803_, _074804_, _074805_, _074806_, _074807_, _074808_, _074809_, _074810_, _074811_, _074812_, _074813_, _074814_, _074815_, _074816_, _074817_, _074818_, _074819_, _074820_, _074821_, _074822_, _074823_, _074824_, _074825_, _074826_, _074827_, _074828_, _074829_, _074830_, _074831_, _074832_, _074833_, _074834_, _074835_, _074836_, _074837_, _074838_, _074839_, _074840_, _074841_, _074842_, _074843_, _074844_, _074845_, _074846_, _074847_, _074848_, _074849_, _074850_, _074851_, _074852_, _074853_, _074854_, _074855_, _074856_, _074857_, _074858_, _074859_, _074860_, _074861_, _074862_, _074863_, _074864_, _074865_, _074866_, _074867_, _074868_, _074869_, _074870_, _074871_, _074872_, _074873_, _074874_, _074875_, _074876_, _074877_, _074878_, _074879_, _074880_, _074881_, _074882_, _074883_, _074884_, _074885_, _074886_, _074887_, _074888_, _074889_, _074890_, _074891_, _074892_, _074893_, _074894_, _074895_, _074896_, _074897_, _074898_, _074899_, _074900_, _074901_, _074902_, _074903_, _074904_, _074905_, _074906_, _074907_, _074908_, _074909_, _074910_, _074911_, _074912_, _074913_, _074914_, _074915_, _074916_, _074917_, _074918_, _074919_, _074920_, _074921_, _074922_, _074923_, _074924_, _074925_, _074926_, _074927_, _074928_, _074929_, _074930_, _074931_, _074932_, _074933_, _074934_, _074935_, _074936_, _074937_, _074938_, _074939_, _074940_, _074941_, _074942_, _074943_, _074944_, _074945_, _074946_, _074947_, _074948_, _074949_, _074950_, _074951_, _074952_, _074953_, _074954_, _074955_, _074956_, _074957_, _074958_, _074959_, _074960_, _074961_, _074962_, _074963_, _074964_, _074965_, _074966_, _074967_, _074968_, _074969_, _074970_, _074971_, _074972_, _074973_, _074974_, _074975_, _074976_, _074977_, _074978_, _074979_, _074980_, _074981_, _074982_, _074983_, _074984_, _074985_, _074986_, _074987_, _074988_, _074989_, _074990_, _074991_, _074992_, _074993_, _074994_, _074995_, _074996_, _074997_, _074998_, _074999_, _075000_, _075001_, _075002_, _075003_, _075004_, _075005_, _075006_, _075007_, _075008_, _075009_, _075010_, _075011_, _075012_, _075013_, _075014_, _075015_, _075016_, _075017_, _075018_, _075019_, _075020_, _075021_, _075022_, _075023_, _075024_, _075025_, _075026_, _075027_, _075028_, _075029_, _075030_, _075031_, _075032_, _075033_, _075034_, _075035_, _075036_, _075037_, _075038_, _075039_, _075040_, _075041_, _075042_, _075043_, _075044_, _075045_, _075046_, _075047_, _075048_, _075049_, _075050_, _075051_, _075052_, _075053_, _075054_, _075055_, _075056_, _075057_, _075058_, _075059_, _075060_, _075061_, _075062_, _075063_, _075064_, _075065_, _075066_, _075067_, _075068_, _075069_, _075070_, _075071_, _075072_, _075073_, _075074_, _075075_, _075076_, _075077_, _075078_, _075079_, _075080_, _075081_, _075082_, _075083_, _075084_, _075085_, _075086_, _075087_, _075088_, _075089_, _075090_, _075091_, _075092_, _075093_, _075094_, _075095_, _075096_, _075097_, _075098_, _075099_, _075100_, _075101_, _075102_, _075103_, _075104_, _075105_, _075106_, _075107_, _075108_, _075109_, _075110_, _075111_, _075112_, _075113_, _075114_, _075115_, _075116_, _075117_, _075118_, _075119_, _075120_, _075121_, _075122_, _075123_, _075124_, _075125_, _075126_, _075127_, _075128_, _075129_, _075130_, _075131_, _075132_, _075133_, _075134_, _075135_, _075136_, _075137_, _075138_, _075139_, _075140_, _075141_, _075142_, _075143_, _075144_, _075145_, _075146_, _075147_, _075148_, _075149_, _075150_, _075151_, _075152_, _075153_, _075154_, _075155_, _075156_, _075157_, _075158_, _075159_, _075160_, _075161_, _075162_, _075163_, _075164_, _075165_, _075166_, _075167_, _075168_, _075169_, _075170_, _075171_, _075172_, _075173_, _075174_, _075175_, _075176_, _075177_, _075178_, _075179_, _075180_, _075181_, _075182_, _075183_, _075184_, _075185_, _075186_, _075187_, _075188_, _075189_, _075190_, _075191_, _075192_, _075193_, _075194_, _075195_, _075196_, _075197_, _075198_, _075199_, _075200_, _075201_, _075202_, _075203_, _075204_, _075205_, _075206_, _075207_, _075208_, _075209_, _075210_, _075211_, _075212_, _075213_, _075214_, _075215_, _075216_, _075217_, _075218_, _075219_, _075220_, _075221_, _075222_, _075223_, _075224_, _075225_, _075226_, _075227_, _075228_, _075229_, _075230_, _075231_, _075232_, _075233_, _075234_, _075235_, _075236_, _075237_, _075238_, _075239_, _075240_, _075241_, _075242_, _075243_, _075244_, _075245_, _075246_, _075247_, _075248_, _075249_, _075250_, _075251_, _075252_, _075253_, _075254_, _075255_, _075256_, _075257_, _075258_, _075259_, _075260_, _075261_, _075262_, _075263_, _075264_, _075265_, _075266_, _075267_, _075268_, _075269_, _075270_, _075271_, _075272_, _075273_, _075274_, _075275_, _075276_, _075277_, _075278_, _075279_, _075280_, _075281_, _075282_, _075283_, _075284_, _075285_, _075286_, _075287_, _075288_, _075289_, _075290_, _075291_, _075292_, _075293_, _075294_, _075295_, _075296_, _075297_, _075298_, _075299_, _075300_, _075301_, _075302_, _075303_, _075304_, _075305_, _075306_, _075307_, _075308_, _075309_, _075310_, _075311_, _075312_, _075313_, _075314_, _075315_, _075316_, _075317_, _075318_, _075319_, _075320_, _075321_, _075322_, _075323_, _075324_, _075325_, _075326_, _075327_, _075328_, _075329_, _075330_, _075331_, _075332_, _075333_, _075334_, _075335_, _075336_, _075337_, _075338_, _075339_, _075340_, _075341_, _075342_, _075343_, _075344_, _075345_, _075346_, _075347_, _075348_, _075349_, _075350_, _075351_, _075352_, _075353_, _075354_, _075355_, _075356_, _075357_, _075358_, _075359_, _075360_, _075361_, _075362_, _075363_, _075364_, _075365_, _075366_, _075367_, _075368_, _075369_, _075370_, _075371_, _075372_, _075373_, _075374_, _075375_, _075376_, _075377_, _075378_, _075379_, _075380_, _075381_, _075382_, _075383_, _075384_, _075385_, _075386_, _075387_, _075388_, _075389_, _075390_, _075391_, _075392_, _075393_, _075394_, _075395_, _075396_, _075397_, _075398_, _075399_, _075400_, _075401_, _075402_, _075403_, _075404_, _075405_, _075406_, _075407_, _075408_, _075409_, _075410_, _075411_, _075412_, _075413_, _075414_, _075415_, _075416_, _075417_, _075418_, _075419_, _075420_, _075421_, _075422_, _075423_, _075424_, _075425_, _075426_, _075427_, _075428_, _075429_, _075430_, _075431_, _075432_, _075433_, _075434_, _075435_, _075436_, _075437_, _075438_, _075439_, _075440_, _075441_, _075442_, _075443_, _075444_, _075445_, _075446_, _075447_, _075448_, _075449_, _075450_, _075451_, _075452_, _075453_, _075454_, _075455_, _075456_, _075457_, _075458_, _075459_, _075460_, _075461_, _075462_, _075463_, _075464_, _075465_, _075466_, _075467_, _075468_, _075469_, _075470_, _075471_, _075472_, _075473_, _075474_, _075475_, _075476_, _075477_, _075478_, _075479_, _075480_, _075481_, _075482_, _075483_, _075484_, _075485_, _075486_, _075487_, _075488_, _075489_, _075490_, _075491_, _075492_, _075493_, _075494_, _075495_, _075496_, _075497_, _075498_, _075499_, _075500_, _075501_, _075502_, _075503_, _075504_, _075505_, _075506_, _075507_, _075508_, _075509_, _075510_, _075511_, _075512_, _075513_, _075514_, _075515_, _075516_, _075517_, _075518_, _075519_, _075520_, _075521_, _075522_, _075523_, _075524_, _075525_, _075526_, _075527_, _075528_, _075529_, _075530_, _075531_, _075532_, _075533_, _075534_, _075535_, _075536_, _075537_, _075538_, _075539_, _075540_, _075541_, _075542_, _075543_, _075544_, _075545_, _075546_, _075547_, _075548_, _075549_, _075550_, _075551_, _075552_, _075553_, _075554_, _075555_, _075556_, _075557_, _075558_, _075559_, _075560_, _075561_, _075562_, _075563_, _075564_, _075565_, _075566_, _075567_, _075568_, _075569_, _075570_, _075571_, _075572_, _075573_, _075574_, _075575_, _075576_, _075577_, _075578_, _075579_, _075580_, _075581_, _075582_, _075583_, _075584_, _075585_, _075586_, _075587_, _075588_, _075589_, _075590_, _075591_, _075592_, _075593_, _075594_, _075595_, _075596_, _075597_, _075598_, _075599_, _075600_, _075601_, _075602_, _075603_, _075604_, _075605_, _075606_, _075607_, _075608_, _075609_, _075610_, _075611_, _075612_, _075613_, _075614_, _075615_, _075616_, _075617_, _075618_, _075619_, _075620_, _075621_, _075622_, _075623_, _075624_, _075625_, _075626_, _075627_, _075628_, _075629_, _075630_, _075631_, _075632_, _075633_, _075634_, _075635_, _075636_, _075637_, _075638_, _075639_, _075640_, _075641_, _075642_, _075643_, _075644_, _075645_, _075646_, _075647_, _075648_, _075649_, _075650_, _075651_, _075652_, _075653_, _075654_, _075655_, _075656_, _075657_, _075658_, _075659_, _075660_, _075661_, _075662_, _075663_, _075664_, _075665_, _075666_, _075667_, _075668_, _075669_, _075670_, _075671_, _075672_, _075673_, _075674_, _075675_, _075676_, _075677_, _075678_, _075679_, _075680_, _075681_, _075682_, _075683_, _075684_, _075685_, _075686_, _075687_, _075688_, _075689_, _075690_, _075691_, _075692_, _075693_, _075694_, _075695_, _075696_, _075697_, _075698_, _075699_, _075700_, _075701_, _075702_, _075703_, _075704_, _075705_, _075706_, _075707_, _075708_, _075709_, _075710_, _075711_, _075712_, _075713_, _075714_, _075715_, _075716_, _075717_, _075718_, _075719_, _075720_, _075721_, _075722_, _075723_, _075724_, _075725_, _075726_, _075727_, _075728_, _075729_, _075730_, _075731_, _075732_, _075733_, _075734_, _075735_, _075736_, _075737_, _075738_, _075739_, _075740_, _075741_, _075742_, _075743_, _075744_, _075745_, _075746_, _075747_, _075748_, _075749_, _075750_, _075751_, _075752_, _075753_, _075754_, _075755_, _075756_, _075757_, _075758_, _075759_, _075760_, _075761_, _075762_, _075763_, _075764_, _075765_, _075766_, _075767_, _075768_, _075769_, _075770_, _075771_, _075772_, _075773_, _075774_, _075775_, _075776_, _075777_, _075778_, _075779_, _075780_, _075781_, _075782_, _075783_, _075784_, _075785_, _075786_, _075787_, _075788_, _075789_, _075790_, _075791_, _075792_, _075793_, _075794_, _075795_, _075796_, _075797_, _075798_, _075799_, _075800_, _075801_, _075802_, _075803_, _075804_, _075805_, _075806_, _075807_, _075808_, _075809_, _075810_, _075811_, _075812_, _075813_, _075814_, _075815_, _075816_, _075817_, _075818_, _075819_, _075820_, _075821_, _075822_, _075823_, _075824_, _075825_, _075826_, _075827_, _075828_, _075829_, _075830_, _075831_, _075832_, _075833_, _075834_, _075835_, _075836_, _075837_, _075838_, _075839_, _075840_, _075841_, _075842_, _075843_, _075844_, _075845_, _075846_, _075847_, _075848_, _075849_, _075850_, _075851_, _075852_, _075853_, _075854_, _075855_, _075856_, _075857_, _075858_, _075859_, _075860_, _075861_, _075862_, _075863_, _075864_, _075865_, _075866_, _075867_, _075868_, _075869_, _075870_, _075871_, _075872_, _075873_, _075874_, _075875_, _075876_, _075877_, _075878_, _075879_, _075880_, _075881_, _075882_, _075883_, _075884_, _075885_, _075886_, _075887_, _075888_, _075889_, _075890_, _075891_, _075892_, _075893_, _075894_, _075895_, _075896_, _075897_, _075898_, _075899_, _075900_, _075901_, _075902_, _075903_, _075904_, _075905_, _075906_, _075907_, _075908_, _075909_, _075910_, _075911_, _075912_, _075913_, _075914_, _075915_, _075916_, _075917_, _075918_, _075919_, _075920_, _075921_, _075922_, _075923_, _075924_, _075925_, _075926_, _075927_, _075928_, _075929_, _075930_, _075931_, _075932_, _075933_, _075934_, _075935_, _075936_, _075937_, _075938_, _075939_, _075940_, _075941_, _075942_, _075943_, _075944_, _075945_, _075946_, _075947_, _075948_, _075949_, _075950_, _075951_, _075952_, _075953_, _075954_, _075955_, _075956_, _075957_, _075958_, _075959_, _075960_, _075961_, _075962_, _075963_, _075964_, _075965_, _075966_, _075967_, _075968_, _075969_, _075970_, _075971_, _075972_, _075973_, _075974_, _075975_, _075976_, _075977_, _075978_, _075979_, _075980_, _075981_, _075982_, _075983_, _075984_, _075985_, _075986_, _075987_, _075988_, _075989_, _075990_, _075991_, _075992_, _075993_, _075994_, _075995_, _075996_, _075997_, _075998_, _075999_, _076000_, _076001_, _076002_, _076003_, _076004_, _076005_, _076006_, _076007_, _076008_, _076009_, _076010_, _076011_, _076012_, _076013_, _076014_, _076015_, _076016_, _076017_, _076018_, _076019_, _076020_, _076021_, _076022_, _076023_, _076024_, _076025_, _076026_, _076027_, _076028_, _076029_, _076030_, _076031_, _076032_, _076033_, _076034_, _076035_, _076036_, _076037_, _076038_, _076039_, _076040_, _076041_, _076042_, _076043_, _076044_, _076045_, _076046_, _076047_, _076048_, _076049_, _076050_, _076051_, _076052_, _076053_, _076054_, _076055_, _076056_, _076057_, _076058_, _076059_, _076060_, _076061_, _076062_, _076063_, _076064_, _076065_, _076066_, _076067_, _076068_, _076069_, _076070_, _076071_, _076072_, _076073_, _076074_, _076075_, _076076_, _076077_, _076078_, _076079_, _076080_, _076081_, _076082_, _076083_, _076084_, _076085_, _076086_, _076087_, _076088_, _076089_, _076090_, _076091_, _076092_, _076093_, _076094_, _076095_, _076096_, _076097_, _076098_, _076099_, _076100_, _076101_, _076102_, _076103_, _076104_, _076105_, _076106_, _076107_, _076108_, _076109_, _076110_, _076111_, _076112_, _076113_, _076114_, _076115_, _076116_, _076117_, _076118_, _076119_, _076120_, _076121_, _076122_, _076123_, _076124_, _076125_, _076126_, _076127_, _076128_, _076129_, _076130_, _076131_, _076132_, _076133_, _076134_, _076135_, _076136_, _076137_, _076138_, _076139_, _076140_, _076141_, _076142_, _076143_, _076144_, _076145_, _076146_, _076147_, _076148_, _076149_, _076150_, _076151_, _076152_, _076153_, _076154_, _076155_, _076156_, _076157_, _076158_, _076159_, _076160_, _076161_, _076162_, _076163_, _076164_, _076165_, _076166_, _076167_, _076168_, _076169_, _076170_, _076171_, _076172_, _076173_, _076174_, _076175_, _076176_, _076177_, _076178_, _076179_, _076180_, _076181_, _076182_, _076183_, _076184_, _076185_, _076186_, _076187_, _076188_, _076189_, _076190_, _076191_, _076192_, _076193_, _076194_, _076195_, _076196_, _076197_, _076198_, _076199_, _076200_, _076201_, _076202_, _076203_, _076204_, _076205_, _076206_, _076207_, _076208_, _076209_, _076210_, _076211_, _076212_, _076213_, _076214_, _076215_, _076216_, _076217_, _076218_, _076219_, _076220_, _076221_, _076222_, _076223_, _076224_, _076225_, _076226_, _076227_, _076228_, _076229_, _076230_, _076231_, _076232_, _076233_, _076234_, _076235_, _076236_, _076237_, _076238_, _076239_, _076240_, _076241_, _076242_, _076243_, _076244_, _076245_, _076246_, _076247_, _076248_, _076249_, _076250_, _076251_, _076252_, _076253_, _076254_, _076255_, _076256_, _076257_, _076258_, _076259_, _076260_, _076261_, _076262_, _076263_, _076264_, _076265_, _076266_, _076267_, _076268_, _076269_, _076270_, _076271_, _076272_, _076273_, _076274_, _076275_, _076276_, _076277_, _076278_, _076279_, _076280_, _076281_, _076282_, _076283_, _076284_, _076285_, _076286_, _076287_, _076288_, _076289_, _076290_, _076291_, _076292_, _076293_, _076294_, _076295_, _076296_, _076297_, _076298_, _076299_, _076300_, _076301_, _076302_, _076303_, _076304_, _076305_, _076306_, _076307_, _076308_, _076309_, _076310_, _076311_, _076312_, _076313_, _076314_, _076315_, _076316_, _076317_, _076318_, _076319_, _076320_, _076321_, _076322_, _076323_, _076324_, _076325_, _076326_, _076327_, _076328_, _076329_, _076330_, _076331_, _076332_, _076333_, _076334_, _076335_, _076336_, _076337_, _076338_, _076339_, _076340_, _076341_, _076342_, _076343_, _076344_, _076345_, _076346_, _076347_, _076348_, _076349_, _076350_, _076351_, _076352_, _076353_, _076354_, _076355_, _076356_, _076357_, _076358_, _076359_, _076360_, _076361_, _076362_, _076363_, _076364_, _076365_, _076366_, _076367_, _076368_, _076369_, _076370_, _076371_, _076372_, _076373_, _076374_, _076375_, _076376_, _076377_, _076378_, _076379_, _076380_, _076381_, _076382_, _076383_, _076384_, _076385_, _076386_, _076387_, _076388_, _076389_, _076390_, _076391_, _076392_, _076393_, _076394_, _076395_, _076396_, _076397_, _076398_, _076399_, _076400_, _076401_, _076402_, _076403_, _076404_, _076405_, _076406_, _076407_, _076408_, _076409_, _076410_, _076411_, _076412_, _076413_, _076414_, _076415_, _076416_, _076417_, _076418_, _076419_, _076420_, _076421_, _076422_, _076423_, _076424_, _076425_, _076426_, _076427_, _076428_, _076429_, _076430_, _076431_, _076432_, _076433_, _076434_, _076435_, _076436_, _076437_, _076438_, _076439_, _076440_, _076441_, _076442_, _076443_, _076444_, _076445_, _076446_, _076447_, _076448_, _076449_, _076450_, _076451_, _076452_, _076453_, _076454_, _076455_, _076456_, _076457_, _076458_, _076459_, _076460_, _076461_, _076462_, _076463_, _076464_, _076465_, _076466_, _076467_, _076468_, _076469_, _076470_, _076471_, _076472_, _076473_, _076474_, _076475_, _076476_, _076477_, _076478_, _076479_, _076480_, _076481_, _076482_, _076483_, _076484_, _076485_, _076486_, _076487_, _076488_, _076489_, _076490_, _076491_, _076492_, _076493_, _076494_, _076495_, _076496_, _076497_, _076498_, _076499_, _076500_, _076501_, _076502_, _076503_, _076504_, _076505_, _076506_, _076507_, _076508_, _076509_, _076510_, _076511_, _076512_, _076513_, _076514_, _076515_, _076516_, _076517_, _076518_, _076519_, _076520_, _076521_, _076522_, _076523_, _076524_, _076525_, _076526_, _076527_, _076528_, _076529_, _076530_, _076531_, _076532_, _076533_, _076534_, _076535_, _076536_, _076537_, _076538_, _076539_, _076540_, _076541_, _076542_, _076543_, _076544_, _076545_, _076546_, _076547_, _076548_, _076549_, _076550_, _076551_, _076552_, _076553_, _076554_, _076555_, _076556_, _076557_, _076558_, _076559_, _076560_, _076561_, _076562_, _076563_, _076564_, _076565_, _076566_, _076567_, _076568_, _076569_, _076570_, _076571_, _076572_, _076573_, _076574_, _076575_, _076576_, _076577_, _076578_, _076579_, _076580_, _076581_, _076582_, _076583_, _076584_, _076585_, _076586_, _076587_, _076588_, _076589_, _076590_, _076591_, _076592_, _076593_, _076594_, _076595_, _076596_, _076597_, _076598_, _076599_, _076600_, _076601_, _076602_, _076603_, _076604_, _076605_, _076606_, _076607_, _076608_, _076609_, _076610_, _076611_, _076612_, _076613_, _076614_, _076615_, _076616_, _076617_, _076618_, _076619_, _076620_, _076621_, _076622_, _076623_, _076624_, _076625_, _076626_, _076627_, _076628_, _076629_, _076630_, _076631_, _076632_, _076633_, _076634_, _076635_, _076636_, _076637_, _076638_, _076639_, _076640_, _076641_, _076642_, _076643_, _076644_, _076645_, _076646_, _076647_, _076648_, _076649_, _076650_, _076651_, _076652_, _076653_, _076654_, _076655_, _076656_, _076657_, _076658_, _076659_, _076660_, _076661_, _076662_, _076663_, _076664_, _076665_, _076666_, _076667_, _076668_, _076669_, _076670_, _076671_, _076672_, _076673_, _076674_, _076675_, _076676_, _076677_, _076678_, _076679_, _076680_, _076681_, _076682_, _076683_, _076684_, _076685_, _076686_, _076687_, _076688_, _076689_, _076690_, _076691_, _076692_, _076693_, _076694_, _076695_, _076696_, _076697_, _076698_, _076699_, _076700_, _076701_, _076702_, _076703_, _076704_, _076705_, _076706_, _076707_, _076708_, _076709_, _076710_, _076711_, _076712_, _076713_, _076714_, _076715_, _076716_, _076717_, _076718_, _076719_, _076720_, _076721_, _076722_, _076723_, _076724_, _076725_, _076726_, _076727_, _076728_, _076729_, _076730_, _076731_, _076732_, _076733_, _076734_, _076735_, _076736_, _076737_, _076738_, _076739_, _076740_, _076741_, _076742_, _076743_, _076744_, _076745_, _076746_, _076747_, _076748_, _076749_, _076750_, _076751_, _076752_, _076753_, _076754_, _076755_, _076756_, _076757_, _076758_, _076759_, _076760_, _076761_, _076762_, _076763_, _076764_, _076765_, _076766_, _076767_, _076768_, _076769_, _076770_, _076771_, _076772_, _076773_, _076774_, _076775_, _076776_, _076777_, _076778_, _076779_, _076780_, _076781_, _076782_, _076783_, _076784_, _076785_, _076786_, _076787_, _076788_, _076789_, _076790_, _076791_, _076792_, _076793_, _076794_, _076795_, _076796_, _076797_, _076798_, _076799_, _076800_, _076801_, _076802_, _076803_, _076804_, _076805_, _076806_, _076807_, _076808_, _076809_, _076810_, _076811_, _076812_, _076813_, _076814_, _076815_, _076816_, _076817_, _076818_, _076819_, _076820_, _076821_, _076822_, _076823_, _076824_, _076825_, _076826_, _076827_, _076828_, _076829_, _076830_, _076831_, _076832_, _076833_, _076834_, _076835_, _076836_, _076837_, _076838_, _076839_, _076840_, _076841_, _076842_, _076843_, _076844_, _076845_, _076846_, _076847_, _076848_, _076849_, _076850_, _076851_, _076852_, _076853_, _076854_, _076855_, _076856_, _076857_, _076858_, _076859_, _076860_, _076861_, _076862_, _076863_, _076864_, _076865_, _076866_, _076867_, _076868_, _076869_, _076870_, _076871_, _076872_, _076873_, _076874_, _076875_, _076876_, _076877_, _076878_, _076879_, _076880_, _076881_, _076882_, _076883_, _076884_, _076885_, _076886_, _076887_, _076888_, _076889_, _076890_, _076891_, _076892_, _076893_, _076894_, _076895_, _076896_, _076897_, _076898_, _076899_, _076900_, _076901_, _076902_, _076903_, _076904_, _076905_, _076906_, _076907_, _076908_, _076909_, _076910_, _076911_, _076912_, _076913_, _076914_, _076915_, _076916_, _076917_, _076918_, _076919_, _076920_, _076921_, _076922_, _076923_, _076924_, _076925_, _076926_, _076927_, _076928_, _076929_, _076930_, _076931_, _076932_, _076933_, _076934_, _076935_, _076936_, _076937_, _076938_, _076939_, _076940_, _076941_, _076942_, _076943_, _076944_, _076945_, _076946_, _076947_, _076948_, _076949_, _076950_, _076951_, _076952_, _076953_, _076954_, _076955_, _076956_, _076957_, _076958_, _076959_, _076960_, _076961_, _076962_, _076963_, _076964_, _076965_, _076966_, _076967_, _076968_, _076969_, _076970_, _076971_, _076972_, _076973_, _076974_, _076975_, _076976_, _076977_, _076978_, _076979_, _076980_, _076981_, _076982_, _076983_, _076984_, _076985_, _076986_, _076987_, _076988_, _076989_, _076990_, _076991_, _076992_, _076993_, _076994_, _076995_, _076996_, _076997_, _076998_, _076999_, _077000_, _077001_, _077002_, _077003_, _077004_, _077005_, _077006_, _077007_, _077008_, _077009_, _077010_, _077011_, _077012_, _077013_, _077014_, _077015_, _077016_, _077017_, _077018_, _077019_, _077020_, _077021_, _077022_, _077023_, _077024_, _077025_, _077026_, _077027_, _077028_, _077029_, _077030_, _077031_, _077032_, _077033_, _077034_, _077035_, _077036_, _077037_, _077038_, _077039_, _077040_, _077041_, _077042_, _077043_, _077044_, _077045_, _077046_, _077047_, _077048_, _077049_, _077050_, _077051_, _077052_, _077053_, _077054_, _077055_, _077056_, _077057_, _077058_, _077059_, _077060_, _077061_, _077062_, _077063_, _077064_, _077065_, _077066_, _077067_, _077068_, _077069_, _077070_, _077071_, _077072_, _077073_, _077074_, _077075_, _077076_, _077077_, _077078_, _077079_, _077080_, _077081_, _077082_, _077083_, _077084_, _077085_, _077086_, _077087_, _077088_, _077089_, _077090_, _077091_, _077092_, _077093_, _077094_, _077095_, _077096_, _077097_, _077098_, _077099_, _077100_, _077101_, _077102_, _077103_, _077104_, _077105_, _077106_, _077107_, _077108_, _077109_, _077110_, _077111_, _077112_, _077113_, _077114_, _077115_, _077116_, _077117_, _077118_, _077119_, _077120_, _077121_, _077122_, _077123_, _077124_, _077125_, _077126_, _077127_, _077128_, _077129_, _077130_, _077131_, _077132_, _077133_, _077134_, _077135_, _077136_, _077137_, _077138_, _077139_, _077140_, _077141_, _077142_, _077143_, _077144_, _077145_, _077146_, _077147_, _077148_, _077149_, _077150_, _077151_, _077152_, _077153_, _077154_, _077155_, _077156_, _077157_, _077158_, _077159_, _077160_, _077161_, _077162_, _077163_, _077164_, _077165_, _077166_, _077167_, _077168_, _077169_, _077170_, _077171_, _077172_, _077173_, _077174_, _077175_, _077176_, _077177_, _077178_, _077179_, _077180_, _077181_, _077182_, _077183_, _077184_, _077185_, _077186_, _077187_, _077188_, _077189_, _077190_, _077191_, _077192_, _077193_, _077194_, _077195_, _077196_, _077197_, _077198_, _077199_, _077200_, _077201_, _077202_, _077203_, _077204_, _077205_, _077206_, _077207_, _077208_, _077209_, _077210_, _077211_, _077212_, _077213_, _077214_, _077215_, _077216_, _077217_, _077218_, _077219_, _077220_, _077221_, _077222_, _077223_, _077224_, _077225_, _077226_, _077227_, _077228_, _077229_, _077230_, _077231_, _077232_, _077233_, _077234_, _077235_, _077236_, _077237_, _077238_, _077239_, _077240_, _077241_, _077242_, _077243_, _077244_, _077245_, _077246_, _077247_, _077248_, _077249_, _077250_, _077251_, _077252_, _077253_, _077254_, _077255_, _077256_, _077257_, _077258_, _077259_, _077260_, _077261_, _077262_, _077263_, _077264_, _077265_, _077266_, _077267_, _077268_, _077269_, _077270_, _077271_, _077272_, _077273_, _077274_, _077275_, _077276_, _077277_, _077278_, _077279_, _077280_, _077281_, _077282_, _077283_, _077284_, _077285_, _077286_, _077287_, _077288_, _077289_, _077290_, _077291_, _077292_, _077293_, _077294_, _077295_, _077296_, _077297_, _077298_, _077299_, _077300_, _077301_, _077302_, _077303_, _077304_, _077305_, _077306_, _077307_, _077308_, _077309_, _077310_, _077311_, _077312_, _077313_, _077314_, _077315_, _077316_, _077317_, _077318_, _077319_, _077320_, _077321_, _077322_, _077323_, _077324_, _077325_, _077326_, _077327_, _077328_, _077329_, _077330_, _077331_, _077332_, _077333_, _077334_, _077335_, _077336_, _077337_, _077338_, _077339_, _077340_, _077341_, _077342_, _077343_, _077344_, _077345_, _077346_, _077347_, _077348_, _077349_, _077350_, _077351_, _077352_, _077353_, _077354_, _077355_, _077356_, _077357_, _077358_, _077359_, _077360_, _077361_, _077362_, _077363_, _077364_, _077365_, _077366_, _077367_, _077368_, _077369_, _077370_, _077371_, _077372_, _077373_, _077374_, _077375_, _077376_, _077377_, _077378_, _077379_, _077380_, _077381_, _077382_, _077383_, _077384_, _077385_, _077386_, _077387_, _077388_, _077389_, _077390_, _077391_, _077392_, _077393_, _077394_, _077395_, _077396_, _077397_, _077398_, _077399_, _077400_, _077401_, _077402_, _077403_, _077404_, _077405_, _077406_, _077407_, _077408_, _077409_, _077410_, _077411_, _077412_, _077413_, _077414_, _077415_, _077416_, _077417_, _077418_, _077419_, _077420_, _077421_, _077422_, _077423_, _077424_, _077425_, _077426_, _077427_, _077428_, _077429_, _077430_, _077431_, _077432_, _077433_, _077434_, _077435_, _077436_, _077437_, _077438_, _077439_, _077440_, _077441_, _077442_, _077443_, _077444_, _077445_, _077446_, _077447_, _077448_, _077449_, _077450_, _077451_, _077452_, _077453_, _077454_, _077455_, _077456_, _077457_, _077458_, _077459_, _077460_, _077461_, _077462_, _077463_, _077464_, _077465_, _077466_, _077467_, _077468_, _077469_, _077470_, _077471_, _077472_, _077473_, _077474_, _077475_, _077476_, _077477_, _077478_, _077479_, _077480_, _077481_, _077482_, _077483_, _077484_, _077485_, _077486_, _077487_, _077488_, _077489_, _077490_, _077491_, _077492_, _077493_, _077494_, _077495_, _077496_, _077497_, _077498_, _077499_, _077500_, _077501_, _077502_, _077503_, _077504_, _077505_, _077506_, _077507_, _077508_, _077509_, _077510_, _077511_, _077512_, _077513_, _077514_, _077515_, _077516_, _077517_, _077518_, _077519_, _077520_, _077521_, _077522_, _077523_, _077524_, _077525_, _077526_, _077527_, _077528_, _077529_, _077530_, _077531_, _077532_, _077533_, _077534_, _077535_, _077536_, _077537_, _077538_, _077539_, _077540_, _077541_, _077542_, _077543_, _077544_, _077545_, _077546_, _077547_, _077548_, _077549_, _077550_, _077551_, _077552_, _077553_, _077554_, _077555_, _077556_, _077557_, _077558_, _077559_, _077560_, _077561_, _077562_, _077563_, _077564_, _077565_, _077566_, _077567_, _077568_, _077569_, _077570_, _077571_, _077572_, _077573_, _077574_, _077575_, _077576_, _077577_, _077578_, _077579_, _077580_, _077581_, _077582_, _077583_, _077584_, _077585_, _077586_, _077587_, _077588_, _077589_, _077590_, _077591_, _077592_, _077593_, _077594_, _077595_, _077596_, _077597_, _077598_, _077599_, _077600_, _077601_, _077602_, _077603_, _077604_, _077605_, _077606_, _077607_, _077608_, _077609_, _077610_, _077611_, _077612_, _077613_, _077614_, _077615_, _077616_, _077617_, _077618_, _077619_, _077620_, _077621_, _077622_, _077623_, _077624_, _077625_, _077626_, _077627_, _077628_, _077629_, _077630_, _077631_, _077632_, _077633_, _077634_, _077635_, _077636_, _077637_, _077638_, _077639_, _077640_, _077641_, _077642_, _077643_, _077644_, _077645_, _077646_, _077647_, _077648_, _077649_, _077650_, _077651_, _077652_, _077653_, _077654_, _077655_, _077656_, _077657_, _077658_, _077659_, _077660_, _077661_, _077662_, _077663_, _077664_, _077665_, _077666_, _077667_, _077668_, _077669_, _077670_, _077671_, _077672_, _077673_, _077674_, _077675_, _077676_, _077677_, _077678_, _077679_, _077680_, _077681_, _077682_, _077683_, _077684_, _077685_, _077686_, _077687_, _077688_, _077689_, _077690_, _077691_, _077692_, _077693_, _077694_, _077695_, _077696_, _077697_, _077698_, _077699_, _077700_, _077701_, _077702_, _077703_, _077704_, _077705_, _077706_, _077707_, _077708_, _077709_, _077710_, _077711_, _077712_, _077713_, _077714_, _077715_, _077716_, _077717_, _077718_, _077719_, _077720_, _077721_, _077722_, _077723_, _077724_, _077725_, _077726_, _077727_, _077728_, _077729_, _077730_, _077731_, _077732_, _077733_, _077734_, _077735_, _077736_, _077737_, _077738_, _077739_, _077740_, _077741_, _077742_, _077743_, _077744_, _077745_, _077746_, _077747_, _077748_, _077749_, _077750_, _077751_, _077752_, _077753_, _077754_, _077755_, _077756_, _077757_, _077758_, _077759_, _077760_, _077761_, _077762_, _077763_, _077764_, _077765_, _077766_, _077767_, _077768_, _077769_, _077770_, _077771_, _077772_, _077773_, _077774_, _077775_, _077776_, _077777_, _077778_, _077779_, _077780_, _077781_, _077782_, _077783_, _077784_, _077785_, _077786_, _077787_, _077788_, _077789_, _077790_, _077791_, _077792_, _077793_, _077794_, _077795_, _077796_, _077797_, _077798_, _077799_, _077800_, _077801_, _077802_, _077803_, _077804_, _077805_, _077806_, _077807_, _077808_, _077809_, _077810_, _077811_, _077812_, _077813_, _077814_, _077815_, _077816_, _077817_, _077818_, _077819_, _077820_, _077821_, _077822_, _077823_, _077824_, _077825_, _077826_, _077827_, _077828_, _077829_, _077830_, _077831_, _077832_, _077833_, _077834_, _077835_, _077836_, _077837_, _077838_, _077839_, _077840_, _077841_, _077842_, _077843_, _077844_, _077845_, _077846_, _077847_, _077848_, _077849_, _077850_, _077851_, _077852_, _077853_, _077854_, _077855_, _077856_, _077857_, _077858_, _077859_, _077860_, _077861_, _077862_, _077863_, _077864_, _077865_, _077866_, _077867_, _077868_, _077869_, _077870_, _077871_, _077872_, _077873_, _077874_, _077875_, _077876_, _077877_, _077878_, _077879_, _077880_, _077881_, _077882_, _077883_, _077884_, _077885_, _077886_, _077887_, _077888_, _077889_, _077890_, _077891_, _077892_, _077893_, _077894_, _077895_, _077896_, _077897_, _077898_, _077899_, _077900_, _077901_, _077902_, _077903_, _077904_, _077905_, _077906_, _077907_, _077908_, _077909_, _077910_, _077911_, _077912_, _077913_, _077914_, _077915_, _077916_, _077917_, _077918_, _077919_, _077920_, _077921_, _077922_, _077923_, _077924_, _077925_, _077926_, _077927_, _077928_, _077929_, _077930_, _077931_, _077932_, _077933_, _077934_, _077935_, _077936_, _077937_, _077938_, _077939_, _077940_, _077941_, _077942_, _077943_, _077944_, _077945_, _077946_, _077947_, _077948_, _077949_, _077950_, _077951_, _077952_, _077953_, _077954_, _077955_, _077956_, _077957_, _077958_, _077959_, _077960_, _077961_, _077962_, _077963_, _077964_, _077965_, _077966_, _077967_, _077968_, _077969_, _077970_, _077971_, _077972_, _077973_, _077974_, _077975_, _077976_, _077977_, _077978_, _077979_, _077980_, _077981_, _077982_, _077983_, _077984_, _077985_, _077986_, _077987_, _077988_, _077989_, _077990_, _077991_, _077992_, _077993_, _077994_, _077995_, _077996_, _077997_, _077998_, _077999_, _078000_, _078001_, _078002_, _078003_, _078004_, _078005_, _078006_, _078007_, _078008_, _078009_, _078010_, _078011_, _078012_, _078013_, _078014_, _078015_, _078016_, _078017_, _078018_, _078019_, _078020_, _078021_, _078022_, _078023_, _078024_, _078025_, _078026_, _078027_, _078028_, _078029_, _078030_, _078031_, _078032_, _078033_, _078034_, _078035_, _078036_, _078037_, _078038_, _078039_, _078040_, _078041_, _078042_, _078043_, _078044_, _078045_, _078046_, _078047_, _078048_, _078049_, _078050_, _078051_, _078052_, _078053_, _078054_, _078055_, _078056_, _078057_, _078058_, _078059_, _078060_, _078061_, _078062_, _078063_, _078064_, _078065_, _078066_, _078067_, _078068_, _078069_, _078070_, _078071_, _078072_, _078073_, _078074_, _078075_, _078076_, _078077_, _078078_, _078079_, _078080_, _078081_, _078082_, _078083_, _078084_, _078085_, _078086_, _078087_, _078088_, _078089_, _078090_, _078091_, _078092_, _078093_, _078094_, _078095_, _078096_, _078097_, _078098_, _078099_, _078100_, _078101_, _078102_, _078103_, _078104_, _078105_, _078106_, _078107_, _078108_, _078109_, _078110_, _078111_, _078112_, _078113_, _078114_, _078115_, _078116_, _078117_, _078118_, _078119_, _078120_, _078121_, _078122_, _078123_, _078124_, _078125_, _078126_, _078127_, _078128_, _078129_, _078130_, _078131_, _078132_, _078133_, _078134_, _078135_, _078136_, _078137_, _078138_, _078139_, _078140_, _078141_, _078142_, _078143_, _078144_, _078145_, _078146_, _078147_, _078148_, _078149_, _078150_, _078151_, _078152_, _078153_, _078154_, _078155_, _078156_, _078157_, _078158_, _078159_, _078160_, _078161_, _078162_, _078163_, _078164_, _078165_, _078166_, _078167_, _078168_, _078169_, _078170_, _078171_, _078172_, _078173_, _078174_, _078175_, _078176_, _078177_, _078178_, _078179_, _078180_, _078181_, _078182_, _078183_, _078184_, _078185_, _078186_, _078187_, _078188_, _078189_, _078190_, _078191_, _078192_, _078193_, _078194_, _078195_, _078196_, _078197_, _078198_, _078199_, _078200_, _078201_, _078202_, _078203_, _078204_, _078205_, _078206_, _078207_, _078208_, _078209_, _078210_, _078211_, _078212_, _078213_, _078214_, _078215_, _078216_, _078217_, _078218_, _078219_, _078220_, _078221_, _078222_, _078223_, _078224_, _078225_, _078226_, _078227_, _078228_, _078229_, _078230_, _078231_, _078232_, _078233_, _078234_, _078235_, _078236_, _078237_, _078238_, _078239_, _078240_, _078241_, _078242_, _078243_, _078244_, _078245_, _078246_, _078247_, _078248_, _078249_, _078250_, _078251_, _078252_, _078253_, _078254_, _078255_, _078256_, _078257_, _078258_, _078259_, _078260_, _078261_, _078262_, _078263_, _078264_, _078265_, _078266_, _078267_, _078268_, _078269_, _078270_, _078271_, _078272_, _078273_, _078274_, _078275_, _078276_, _078277_, _078278_, _078279_, _078280_, _078281_, _078282_, _078283_, _078284_, _078285_, _078286_, _078287_, _078288_, _078289_, _078290_, _078291_, _078292_, _078293_, _078294_, _078295_, _078296_, _078297_, _078298_, _078299_, _078300_, _078301_, _078302_, _078303_, _078304_, _078305_, _078306_, _078307_, _078308_, _078309_, _078310_, _078311_, _078312_, _078313_, _078314_, _078315_, _078316_, _078317_, _078318_, _078319_, _078320_, _078321_, _078322_, _078323_, _078324_, _078325_, _078326_, _078327_, _078328_, _078329_, _078330_, _078331_, _078332_, _078333_, _078334_, _078335_, _078336_, _078337_, _078338_, _078339_, _078340_, _078341_, _078342_, _078343_, _078344_, _078345_, _078346_, _078347_, _078348_, _078349_, _078350_, _078351_, _078352_, _078353_, _078354_, _078355_, _078356_, _078357_, _078358_, _078359_, _078360_, _078361_, _078362_, _078363_, _078364_, _078365_, _078366_, _078367_, _078368_, _078369_, _078370_, _078371_, _078372_, _078373_, _078374_, _078375_, _078376_, _078377_, _078378_, _078379_, _078380_, _078381_, _078382_, _078383_, _078384_, _078385_, _078386_, _078387_, _078388_, _078389_, _078390_, _078391_, _078392_, _078393_, _078394_, _078395_, _078396_, _078397_, _078398_, _078399_, _078400_, _078401_, _078402_, _078403_, _078404_, _078405_, _078406_, _078407_, _078408_, _078409_, _078410_, _078411_, _078412_, _078413_, _078414_, _078415_, _078416_, _078417_, _078418_, _078419_, _078420_, _078421_, _078422_, _078423_, _078424_, _078425_, _078426_, _078427_, _078428_, _078429_, _078430_, _078431_, _078432_, _078433_, _078434_, _078435_, _078436_, _078437_, _078438_, _078439_, _078440_, _078441_, _078442_, _078443_, _078444_, _078445_, _078446_, _078447_, _078448_, _078449_, _078450_, _078451_, _078452_, _078453_, _078454_, _078455_, _078456_, _078457_, _078458_, _078459_, _078460_, _078461_, _078462_, _078463_, _078464_, _078465_, _078466_, _078467_, _078468_, _078469_, _078470_, _078471_, _078472_, _078473_, _078474_, _078475_, _078476_, _078477_, _078478_, _078479_, _078480_, _078481_, _078482_, _078483_, _078484_, _078485_, _078486_, _078487_, _078488_, _078489_, _078490_, _078491_, _078492_, _078493_, _078494_, _078495_, _078496_, _078497_, _078498_, _078499_, _078500_, _078501_, _078502_, _078503_, _078504_, _078505_, _078506_, _078507_, _078508_, _078509_, _078510_, _078511_, _078512_, _078513_, _078514_, _078515_, _078516_, _078517_, _078518_, _078519_, _078520_, _078521_, _078522_, _078523_, _078524_, _078525_, _078526_, _078527_, _078528_, _078529_, _078530_, _078531_, _078532_, _078533_, _078534_, _078535_, _078536_, _078537_, _078538_, _078539_, _078540_, _078541_, _078542_, _078543_, _078544_, _078545_, _078546_, _078547_, _078548_, _078549_, _078550_, _078551_, _078552_, _078553_, _078554_, _078555_, _078556_, _078557_, _078558_, _078559_, _078560_, _078561_, _078562_, _078563_, _078564_, _078565_, _078566_, _078567_, _078568_, _078569_, _078570_, _078571_, _078572_, _078573_, _078574_, _078575_, _078576_, _078577_, _078578_, _078579_, _078580_, _078581_, _078582_, _078583_, _078584_, _078585_, _078586_, _078587_, _078588_, _078589_, _078590_, _078591_, _078592_, _078593_, _078594_, _078595_, _078596_, _078597_, _078598_, _078599_, _078600_, _078601_, _078602_, _078603_, _078604_, _078605_, _078606_, _078607_, _078608_, _078609_, _078610_, _078611_, _078612_, _078613_, _078614_, _078615_, _078616_, _078617_, _078618_, _078619_, _078620_, _078621_, _078622_, _078623_, _078624_, _078625_, _078626_, _078627_, _078628_, _078629_, _078630_, _078631_, _078632_, _078633_, _078634_, _078635_, _078636_, _078637_, _078638_, _078639_, _078640_, _078641_, _078642_, _078643_, _078644_, _078645_, _078646_, _078647_, _078648_, _078649_, _078650_, _078651_, _078652_, _078653_, _078654_, _078655_, _078656_, _078657_, _078658_, _078659_, _078660_, _078661_, _078662_, _078663_, _078664_, _078665_, _078666_, _078667_, _078668_, _078669_, _078670_, _078671_, _078672_, _078673_, _078674_, _078675_, _078676_, _078677_, _078678_, _078679_, _078680_, _078681_, _078682_, _078683_, _078684_, _078685_, _078686_, _078687_, _078688_, _078689_, _078690_, _078691_, _078692_, _078693_, _078694_, _078695_, _078696_, _078697_, _078698_, _078699_, _078700_, _078701_, _078702_, _078703_, _078704_, _078705_, _078706_, _078707_, _078708_, _078709_, _078710_, _078711_, _078712_, _078713_, _078714_, _078715_, _078716_, _078717_, _078718_, _078719_, _078720_, _078721_, _078722_, _078723_, _078724_, _078725_, _078726_, _078727_, _078728_, _078729_, _078730_, _078731_, _078732_, _078733_, _078734_, _078735_, _078736_, _078737_, _078738_, _078739_, _078740_, _078741_, _078742_, _078743_, _078744_, _078745_, _078746_, _078747_, _078748_, _078749_, _078750_, _078751_, _078752_, _078753_, _078754_, _078755_, _078756_, _078757_, _078758_, _078759_, _078760_, _078761_, _078762_, _078763_, _078764_, _078765_, _078766_, _078767_, _078768_, _078769_, _078770_, _078771_, _078772_, _078773_, _078774_, _078775_, _078776_, _078777_, _078778_, _078779_, _078780_, _078781_, _078782_, _078783_, _078784_, _078785_, _078786_, _078787_, _078788_, _078789_, _078790_, _078791_, _078792_, _078793_, _078794_, _078795_, _078796_, _078797_, _078798_, _078799_, _078800_, _078801_, _078802_, _078803_, _078804_, _078805_, _078806_, _078807_, _078808_, _078809_, _078810_, _078811_, _078812_, _078813_, _078814_, _078815_, _078816_, _078817_, _078818_, _078819_, _078820_, _078821_, _078822_, _078823_, _078824_, _078825_, _078826_, _078827_, _078828_, _078829_, _078830_, _078831_, _078832_, _078833_, _078834_, _078835_, _078836_, _078837_, _078838_, _078839_, _078840_, _078841_, _078842_, _078843_, _078844_, _078845_, _078846_, _078847_, _078848_, _078849_, _078850_, _078851_, _078852_, _078853_, _078854_, _078855_, _078856_, _078857_, _078858_, _078859_, _078860_, _078861_, _078862_, _078863_, _078864_, _078865_, _078866_, _078867_, _078868_, _078869_, _078870_, _078871_, _078872_, _078873_, _078874_, _078875_, _078876_, _078877_, _078878_, _078879_, _078880_, _078881_, _078882_, _078883_, _078884_, _078885_, _078886_, _078887_, _078888_, _078889_, _078890_, _078891_, _078892_, _078893_, _078894_, _078895_, _078896_, _078897_, _078898_, _078899_, _078900_, _078901_, _078902_, _078903_, _078904_, _078905_, _078906_, _078907_, _078908_, _078909_, _078910_, _078911_, _078912_, _078913_, _078914_, _078915_, _078916_, _078917_, _078918_, _078919_, _078920_, _078921_, _078922_, _078923_, _078924_, _078925_, _078926_, _078927_, _078928_, _078929_, _078930_, _078931_, _078932_, _078933_, _078934_, _078935_, _078936_, _078937_, _078938_, _078939_, _078940_, _078941_, _078942_, _078943_, _078944_, _078945_, _078946_, _078947_, _078948_, _078949_, _078950_, _078951_, _078952_, _078953_, _078954_, _078955_, _078956_, _078957_, _078958_, _078959_, _078960_, _078961_, _078962_, _078963_, _078964_, _078965_, _078966_, _078967_, _078968_, _078969_, _078970_, _078971_, _078972_, _078973_, _078974_, _078975_, _078976_, _078977_, _078978_, _078979_, _078980_, _078981_, _078982_, _078983_, _078984_, _078985_, _078986_, _078987_, _078988_, _078989_, _078990_, _078991_, _078992_, _078993_, _078994_, _078995_, _078996_, _078997_, _078998_, _078999_, _079000_, _079001_, _079002_, _079003_, _079004_, _079005_, _079006_, _079007_, _079008_, _079009_, _079010_, _079011_, _079012_, _079013_, _079014_, _079015_, _079016_, _079017_, _079018_, _079019_, _079020_, _079021_, _079022_, _079023_, _079024_, _079025_, _079026_, _079027_, _079028_, _079029_, _079030_, _079031_, _079032_, _079033_, _079034_, _079035_, _079036_, _079037_, _079038_, _079039_, _079040_, _079041_, _079042_, _079043_, _079044_, _079045_, _079046_, _079047_, _079048_, _079049_, _079050_, _079051_, _079052_, _079053_, _079054_, _079055_, _079056_, _079057_, _079058_, _079059_, _079060_, _079061_, _079062_, _079063_, _079064_, _079065_, _079066_, _079067_, _079068_, _079069_, _079070_, _079071_, _079072_, _079073_, _079074_, _079075_, _079076_, _079077_, _079078_, _079079_, _079080_, _079081_, _079082_, _079083_, _079084_, _079085_, _079086_, _079087_, _079088_, _079089_, _079090_, _079091_, _079092_, _079093_, _079094_, _079095_, _079096_, _079097_, _079098_, _079099_, _079100_, _079101_, _079102_, _079103_, _079104_, _079105_, _079106_, _079107_, _079108_, _079109_, _079110_, _079111_, _079112_, _079113_, _079114_, _079115_, _079116_, _079117_, _079118_, _079119_, _079120_, _079121_, _079122_, _079123_, _079124_, _079125_, _079126_, _079127_, _079128_, _079129_, _079130_, _079131_, _079132_, _079133_, _079134_, _079135_, _079136_, _079137_, _079138_, _079139_, _079140_, _079141_, _079142_, _079143_, _079144_, _079145_, _079146_, _079147_, _079148_, _079149_, _079150_, _079151_, _079152_, _079153_, _079154_, _079155_, _079156_, _079157_, _079158_, _079159_, _079160_, _079161_, _079162_, _079163_, _079164_, _079165_, _079166_, _079167_, _079168_, _079169_, _079170_, _079171_, _079172_, _079173_, _079174_, _079175_, _079176_, _079177_, _079178_, _079179_, _079180_, _079181_, _079182_, _079183_, _079184_, _079185_, _079186_, _079187_, _079188_, _079189_, _079190_, _079191_, _079192_, _079193_, _079194_, _079195_, _079196_, _079197_, _079198_, _079199_, _079200_, _079201_, _079202_, _079203_, _079204_, _079205_, _079206_, _079207_, _079208_, _079209_, _079210_, _079211_, _079212_, _079213_, _079214_, _079215_, _079216_, _079217_, _079218_, _079219_, _079220_, _079221_, _079222_, _079223_, _079224_, _079225_, _079226_, _079227_, _079228_, _079229_, _079230_, _079231_, _079232_, _079233_, _079234_, _079235_, _079236_, _079237_, _079238_, _079239_, _079240_, _079241_, _079242_, _079243_, _079244_, _079245_, _079246_, _079247_, _079248_, _079249_, _079250_, _079251_, _079252_, _079253_, _079254_, _079255_, _079256_, _079257_, _079258_, _079259_, _079260_, _079261_, _079262_, _079263_, _079264_, _079265_, _079266_, _079267_, _079268_, _079269_, _079270_, _079271_, _079272_, _079273_, _079274_, _079275_, _079276_, _079277_, _079278_, _079279_, _079280_, _079281_, _079282_, _079283_, _079284_, _079285_, _079286_, _079287_, _079288_, _079289_, _079290_, _079291_, _079292_, _079293_, _079294_, _079295_, _079296_, _079297_, _079298_, _079299_, _079300_, _079301_, _079302_, _079303_, _079304_, _079305_, _079306_, _079307_, _079308_, _079309_, _079310_, _079311_, _079312_, _079313_, _079314_, _079315_, _079316_, _079317_, _079318_, _079319_, _079320_, _079321_, _079322_, _079323_, _079324_, _079325_, _079326_, _079327_, _079328_, _079329_, _079330_, _079331_, _079332_, _079333_, _079334_, _079335_, _079336_, _079337_, _079338_, _079339_, _079340_, _079341_, _079342_, _079343_, _079344_, _079345_, _079346_, _079347_, _079348_, _079349_, _079350_, _079351_, _079352_, _079353_, _079354_, _079355_, _079356_, _079357_, _079358_, _079359_, _079360_, _079361_, _079362_, _079363_, _079364_, _079365_, _079366_, _079367_, _079368_, _079369_, _079370_, _079371_, _079372_, _079373_, _079374_, _079375_, _079376_, _079377_, _079378_, _079379_, _079380_, _079381_, _079382_, _079383_, _079384_, _079385_, _079386_, _079387_, _079388_, _079389_, _079390_, _079391_, _079392_, _079393_, _079394_, _079395_, _079396_, _079397_, _079398_, _079399_, _079400_, _079401_, _079402_, _079403_, _079404_, _079405_, _079406_, _079407_, _079408_, _079409_, _079410_, _079411_, _079412_, _079413_, _079414_, _079415_, _079416_, _079417_, _079418_, _079419_, _079420_, _079421_, _079422_, _079423_, _079424_, _079425_, _079426_, _079427_, _079428_, _079429_, _079430_, _079431_, _079432_, _079433_, _079434_, _079435_, _079436_, _079437_, _079438_, _079439_, _079440_, _079441_, _079442_, _079443_, _079444_, _079445_, _079446_, _079447_, _079448_, _079449_, _079450_, _079451_, _079452_, _079453_, _079454_, _079455_, _079456_, _079457_, _079458_, _079459_, _079460_, _079461_, _079462_, _079463_, _079464_, _079465_, _079466_, _079467_, _079468_, _079469_, _079470_, _079471_, _079472_, _079473_, _079474_, _079475_, _079476_, _079477_, _079478_, _079479_, _079480_, _079481_, _079482_, _079483_, _079484_, _079485_, _079486_, _079487_, _079488_, _079489_, _079490_, _079491_, _079492_, _079493_, _079494_, _079495_, _079496_, _079497_, _079498_, _079499_, _079500_, _079501_, _079502_, _079503_, _079504_, _079505_, _079506_, _079507_, _079508_, _079509_, _079510_, _079511_, _079512_, _079513_, _079514_, _079515_, _079516_, _079517_, _079518_, _079519_, _079520_, _079521_, _079522_, _079523_, _079524_, _079525_, _079526_, _079527_, _079528_, _079529_, _079530_, _079531_, _079532_, _079533_, _079534_, _079535_, _079536_, _079537_, _079538_, _079539_, _079540_, _079541_, _079542_, _079543_, _079544_, _079545_, _079546_, _079547_, _079548_, _079549_, _079550_, _079551_, _079552_, _079553_, _079554_, _079555_, _079556_, _079557_, _079558_, _079559_, _079560_, _079561_, _079562_, _079563_, _079564_, _079565_, _079566_, _079567_, _079568_, _079569_, _079570_, _079571_, _079572_, _079573_, _079574_, _079575_, _079576_, _079577_, _079578_, _079579_, _079580_, _079581_, _079582_, _079583_, _079584_, _079585_, _079586_, _079587_, _079588_, _079589_, _079590_, _079591_, _079592_, _079593_, _079594_, _079595_, _079596_, _079597_, _079598_, _079599_, _079600_, _079601_, _079602_, _079603_, _079604_, _079605_, _079606_, _079607_, _079608_, _079609_, _079610_, _079611_, _079612_, _079613_, _079614_, _079615_, _079616_, _079617_, _079618_, _079619_, _079620_, _079621_, _079622_, _079623_, _079624_, _079625_, _079626_, _079627_, _079628_, _079629_, _079630_, _079631_, _079632_, _079633_, _079634_, _079635_, _079636_, _079637_, _079638_, _079639_, _079640_, _079641_, _079642_, _079643_, _079644_, _079645_, _079646_, _079647_, _079648_, _079649_, _079650_, _079651_, _079652_, _079653_, _079654_, _079655_, _079656_, _079657_, _079658_, _079659_, _079660_, _079661_, _079662_, _079663_, _079664_, _079665_, _079666_, _079667_, _079668_, _079669_, _079670_, _079671_, _079672_, _079673_, _079674_, _079675_, _079676_, _079677_, _079678_, _079679_, _079680_, _079681_, _079682_, _079683_, _079684_, _079685_, _079686_, _079687_, _079688_, _079689_, _079690_, _079691_, _079692_, _079693_, _079694_, _079695_, _079696_, _079697_, _079698_, _079699_, _079700_, _079701_, _079702_, _079703_, _079704_, _079705_, _079706_, _079707_, _079708_, _079709_, _079710_, _079711_, _079712_, _079713_, _079714_, _079715_, _079716_, _079717_, _079718_, _079719_, _079720_, _079721_, _079722_, _079723_, _079724_, _079725_, _079726_, _079727_, _079728_, _079729_, _079730_, _079731_, _079732_, _079733_, _079734_, _079735_, _079736_, _079737_, _079738_, _079739_, _079740_, _079741_, _079742_, _079743_, _079744_, _079745_, _079746_, _079747_, _079748_, _079749_, _079750_, _079751_, _079752_, _079753_, _079754_, _079755_, _079756_, _079757_, _079758_, _079759_, _079760_, _079761_, _079762_, _079763_, _079764_, _079765_, _079766_, _079767_, _079768_, _079769_, _079770_, _079771_, _079772_, _079773_, _079774_, _079775_, _079776_, _079777_, _079778_, _079779_, _079780_, _079781_, _079782_, _079783_, _079784_, _079785_, _079786_, _079787_, _079788_, _079789_, _079790_, _079791_, _079792_, _079793_, _079794_, _079795_, _079796_, _079797_, _079798_, _079799_, _079800_, _079801_, _079802_, _079803_, _079804_, _079805_, _079806_, _079807_, _079808_, _079809_, _079810_, _079811_, _079812_, _079813_, _079814_, _079815_, _079816_, _079817_, _079818_, _079819_, _079820_, _079821_, _079822_, _079823_, _079824_, _079825_, _079826_, _079827_, _079828_, _079829_, _079830_, _079831_, _079832_, _079833_, _079834_, _079835_, _079836_, _079837_, _079838_, _079839_, _079840_, _079841_, _079842_, _079843_, _079844_, _079845_, _079846_, _079847_, _079848_, _079849_, _079850_, _079851_, _079852_, _079853_, _079854_, _079855_, _079856_, _079857_, _079858_, _079859_, _079860_, _079861_, _079862_, _079863_, _079864_, _079865_, _079866_, _079867_, _079868_, _079869_, _079870_, _079871_, _079872_, _079873_, _079874_, _079875_, _079876_, _079877_, _079878_, _079879_, _079880_, _079881_, _079882_, _079883_, _079884_, _079885_, _079886_, _079887_, _079888_, _079889_, _079890_, _079891_, _079892_, _079893_, _079894_, _079895_, _079896_, _079897_, _079898_, _079899_, _079900_, _079901_, _079902_, _079903_, _079904_, _079905_, _079906_, _079907_, _079908_, _079909_, _079910_, _079911_, _079912_, _079913_, _079914_, _079915_, _079916_, _079917_, _079918_, _079919_, _079920_, _079921_, _079922_, _079923_, _079924_, _079925_, _079926_, _079927_, _079928_, _079929_, _079930_, _079931_, _079932_, _079933_, _079934_, _079935_, _079936_, _079937_, _079938_, _079939_, _079940_, _079941_, _079942_, _079943_, _079944_, _079945_, _079946_, _079947_, _079948_, _079949_, _079950_, _079951_, _079952_, _079953_, _079954_, _079955_, _079956_, _079957_, _079958_, _079959_, _079960_, _079961_, _079962_, _079963_, _079964_, _079965_, _079966_, _079967_, _079968_, _079969_, _079970_, _079971_, _079972_, _079973_, _079974_, _079975_, _079976_, _079977_, _079978_, _079979_, _079980_, _079981_, _079982_, _079983_, _079984_, _079985_, _079986_, _079987_, _079988_, _079989_, _079990_, _079991_, _079992_, _079993_, _079994_, _079995_, _079996_, _079997_, _079998_, _079999_, _080000_, _080001_, _080002_, _080003_, _080004_, _080005_, _080006_, _080007_, _080008_, _080009_, _080010_, _080011_, _080012_, _080013_, _080014_, _080015_, _080016_, _080017_, _080018_, _080019_, _080020_, _080021_, _080022_, _080023_, _080024_, _080025_, _080026_, _080027_, _080028_, _080029_, _080030_, _080031_, _080032_, _080033_, _080034_, _080035_, _080036_, _080037_, _080038_, _080039_, _080040_, _080041_, _080042_, _080043_, _080044_, _080045_, _080046_, _080047_, _080048_, _080049_, _080050_, _080051_, _080052_, _080053_, _080054_, _080055_, _080056_, _080057_, _080058_, _080059_, _080060_, _080061_, _080062_, _080063_, _080064_, _080065_, _080066_, _080067_, _080068_, _080069_, _080070_, _080071_, _080072_, _080073_, _080074_, _080075_, _080076_, _080077_, _080078_, _080079_, _080080_, _080081_, _080082_, _080083_, _080084_, _080085_, _080086_, _080087_, _080088_, _080089_, _080090_, _080091_, _080092_, _080093_, _080094_, _080095_, _080096_, _080097_, _080098_, _080099_, _080100_, _080101_, _080102_, _080103_, _080104_, _080105_, _080106_, _080107_, _080108_, _080109_, _080110_, _080111_, _080112_, _080113_, _080114_, _080115_, _080116_, _080117_, _080118_, _080119_, _080120_, _080121_, _080122_, _080123_, _080124_, _080125_, _080126_, _080127_, _080128_, _080129_, _080130_, _080131_, _080132_, _080133_, _080134_, _080135_, _080136_, _080137_, _080138_, _080139_, _080140_, _080141_, _080142_, _080143_, _080144_, _080145_, _080146_, _080147_, _080148_, _080149_, _080150_, _080151_, _080152_, _080153_, _080154_, _080155_, _080156_, _080157_, _080158_, _080159_, _080160_, _080161_, _080162_, _080163_, _080164_, _080165_, _080166_, _080167_, _080168_, _080169_, _080170_, _080171_, _080172_, _080173_, _080174_, _080175_, _080176_, _080177_, _080178_, _080179_, _080180_, _080181_, _080182_, _080183_, _080184_, _080185_, _080186_, _080187_, _080188_, _080189_, _080190_, _080191_, _080192_, _080193_, _080194_, _080195_, _080196_, _080197_, _080198_, _080199_, _080200_, _080201_, _080202_, _080203_, _080204_, _080205_, _080206_, _080207_, _080208_, _080209_, _080210_, _080211_, _080212_, _080213_, _080214_, _080215_, _080216_, _080217_, _080218_, _080219_, _080220_, _080221_, _080222_, _080223_, _080224_, _080225_, _080226_, _080227_, _080228_, _080229_, _080230_, _080231_, _080232_, _080233_, _080234_, _080235_, _080236_, _080237_, _080238_, _080239_, _080240_, _080241_, _080242_, _080243_, _080244_, _080245_, _080246_, _080247_, _080248_, _080249_, _080250_, _080251_, _080252_, _080253_, _080254_, _080255_, _080256_, _080257_, _080258_, _080259_, _080260_, _080261_, _080262_, _080263_, _080264_, _080265_, _080266_, _080267_, _080268_, _080269_, _080270_, _080271_, _080272_, _080273_, _080274_, _080275_, _080276_, _080277_, _080278_, _080279_, _080280_, _080281_, _080282_, _080283_, _080284_, _080285_, _080286_, _080287_, _080288_, _080289_, _080290_, _080291_, _080292_, _080293_, _080294_, _080295_, _080296_, _080297_, _080298_, _080299_, _080300_, _080301_, _080302_, _080303_, _080304_, _080305_, _080306_, _080307_, _080308_, _080309_, _080310_, _080311_, _080312_, _080313_, _080314_, _080315_, _080316_, _080317_, _080318_, _080319_, _080320_, _080321_, _080322_, _080323_, _080324_, _080325_, _080326_, _080327_, _080328_, _080329_, _080330_, _080331_, _080332_, _080333_, _080334_, _080335_, _080336_, _080337_, _080338_, _080339_, _080340_, _080341_, _080342_, _080343_, _080344_, _080345_, _080346_, _080347_, _080348_, _080349_, _080350_, _080351_, _080352_, _080353_, _080354_, _080355_, _080356_, _080357_, _080358_, _080359_, _080360_, _080361_, _080362_, _080363_, _080364_, _080365_, _080366_, _080367_, _080368_, _080369_, _080370_, _080371_, _080372_, _080373_, _080374_, _080375_, _080376_, _080377_, _080378_, _080379_, _080380_, _080381_, _080382_, _080383_, _080384_, _080385_, _080386_, _080387_, _080388_, _080389_, _080390_, _080391_, _080392_, _080393_, _080394_, _080395_, _080396_, _080397_, _080398_, _080399_, _080400_, _080401_, _080402_, _080403_, _080404_, _080405_, _080406_, _080407_, _080408_, _080409_, _080410_, _080411_, _080412_, _080413_, _080414_, _080415_, _080416_, _080417_, _080418_, _080419_, _080420_, _080421_, _080422_, _080423_, _080424_, _080425_, _080426_, _080427_, _080428_, _080429_, _080430_, _080431_, _080432_, _080433_, _080434_, _080435_, _080436_, _080437_, _080438_, _080439_, _080440_, _080441_, _080442_, _080443_, _080444_, _080445_, _080446_, _080447_, _080448_, _080449_, _080450_, _080451_, _080452_, _080453_, _080454_, _080455_, _080456_, _080457_, _080458_, _080459_, _080460_, _080461_, _080462_, _080463_, _080464_, _080465_, _080466_, _080467_, _080468_, _080469_, _080470_, _080471_, _080472_, _080473_, _080474_, _080475_, _080476_, _080477_, _080478_, _080479_, _080480_, _080481_, _080482_, _080483_, _080484_, _080485_, _080486_, _080487_, _080488_, _080489_, _080490_, _080491_, _080492_, _080493_, _080494_, _080495_, _080496_, _080497_, _080498_, _080499_, _080500_, _080501_, _080502_, _080503_, _080504_, _080505_, _080506_, _080507_, _080508_, _080509_, _080510_, _080511_, _080512_, _080513_, _080514_, _080515_, _080516_, _080517_, _080518_, _080519_, _080520_, _080521_, _080522_, _080523_, _080524_, _080525_, _080526_, _080527_, _080528_, _080529_, _080530_, _080531_, _080532_, _080533_, _080534_, _080535_, _080536_, _080537_, _080538_, _080539_, _080540_, _080541_, _080542_, _080543_, _080544_, _080545_, _080546_, _080547_, _080548_, _080549_, _080550_, _080551_, _080552_, _080553_, _080554_, _080555_, _080556_, _080557_, _080558_, _080559_, _080560_, _080561_, _080562_, _080563_, _080564_, _080565_, _080566_, _080567_, _080568_, _080569_, _080570_, _080571_, _080572_, _080573_, _080574_, _080575_, _080576_, _080577_, _080578_, _080579_, _080580_, _080581_, _080582_, _080583_, _080584_, _080585_, _080586_, _080587_, _080588_, _080589_, _080590_, _080591_, _080592_, _080593_, _080594_, _080595_, _080596_, _080597_, _080598_, _080599_, _080600_, _080601_, _080602_, _080603_, _080604_, _080605_, _080606_, _080607_, _080608_, _080609_, _080610_, _080611_, _080612_, _080613_, _080614_, _080615_, _080616_, _080617_, _080618_, _080619_, _080620_, _080621_, _080622_, _080623_, _080624_, _080625_, _080626_, _080627_, _080628_, _080629_, _080630_, _080631_, _080632_, _080633_, _080634_, _080635_, _080636_, _080637_, _080638_, _080639_, _080640_, _080641_, _080642_, _080643_, _080644_, _080645_, _080646_, _080647_, _080648_, _080649_, _080650_, _080651_, _080652_, _080653_, _080654_, _080655_, _080656_, _080657_, _080658_, _080659_, _080660_, _080661_, _080662_, _080663_, _080664_, _080665_, _080666_, _080667_, _080668_, _080669_, _080670_, _080671_, _080672_, _080673_, _080674_, _080675_, _080676_, _080677_, _080678_, _080679_, _080680_, _080681_, _080682_, _080683_, _080684_, _080685_, _080686_, _080687_, _080688_, _080689_, _080690_, _080691_, _080692_, _080693_, _080694_, _080695_, _080696_, _080697_, _080698_, _080699_, _080700_, _080701_, _080702_, _080703_, _080704_, _080705_, _080706_, _080707_, _080708_, _080709_, _080710_, _080711_, _080712_, _080713_, _080714_, _080715_, _080716_, _080717_, _080718_, _080719_, _080720_, _080721_, _080722_, _080723_, _080724_, _080725_, _080726_, _080727_, _080728_, _080729_, _080730_, _080731_, _080732_, _080733_, _080734_, _080735_, _080736_, _080737_, _080738_, _080739_, _080740_, _080741_, _080742_, _080743_, _080744_, _080745_, _080746_, _080747_, _080748_, _080749_, _080750_, _080751_, _080752_, _080753_, _080754_, _080755_, _080756_, _080757_, _080758_, _080759_, _080760_, _080761_, _080762_, _080763_, _080764_, _080765_, _080766_, _080767_, _080768_, _080769_, _080770_, _080771_, _080772_, _080773_, _080774_, _080775_, _080776_, _080777_, _080778_, _080779_, _080780_, _080781_, _080782_, _080783_, _080784_, _080785_, _080786_, _080787_, _080788_, _080789_, _080790_, _080791_, _080792_, _080793_, _080794_, _080795_, _080796_, _080797_, _080798_, _080799_, _080800_, _080801_, _080802_, _080803_, _080804_, _080805_, _080806_, _080807_, _080808_, _080809_, _080810_, _080811_, _080812_, _080813_, _080814_, _080815_, _080816_, _080817_, _080818_, _080819_, _080820_, _080821_, _080822_, _080823_, _080824_, _080825_, _080826_, _080827_, _080828_, _080829_, _080830_, _080831_, _080832_, _080833_, _080834_, _080835_, _080836_, _080837_, _080838_, _080839_, _080840_, _080841_, _080842_, _080843_, _080844_, _080845_, _080846_, _080847_, _080848_, _080849_, _080850_, _080851_, _080852_, _080853_, _080854_, _080855_, _080856_, _080857_, _080858_, _080859_, _080860_, _080861_, _080862_, _080863_, _080864_, _080865_, _080866_, _080867_, _080868_, _080869_, _080870_, _080871_, _080872_, _080873_, _080874_, _080875_, _080876_, _080877_, _080878_, _080879_, _080880_, _080881_, _080882_, _080883_, _080884_, _080885_, _080886_, _080887_, _080888_, _080889_, _080890_, _080891_, _080892_, _080893_, _080894_, _080895_, _080896_, _080897_, _080898_, _080899_, _080900_, _080901_, _080902_, _080903_, _080904_, _080905_, _080906_, _080907_, _080908_, _080909_, _080910_, _080911_, _080912_, _080913_, _080914_, _080915_, _080916_, _080917_, _080918_, _080919_, _080920_, _080921_, _080922_, _080923_, _080924_, _080925_, _080926_, _080927_, _080928_, _080929_, _080930_, _080931_, _080932_, _080933_, _080934_, _080935_, _080936_, _080937_, _080938_, _080939_, _080940_, _080941_, _080942_, _080943_, _080944_, _080945_, _080946_, _080947_, _080948_, _080949_, _080950_, _080951_, _080952_, _080953_, _080954_, _080955_, _080956_, _080957_, _080958_, _080959_, _080960_, _080961_, _080962_, _080963_, _080964_, _080965_, _080966_, _080967_, _080968_, _080969_, _080970_, _080971_, _080972_, _080973_, _080974_, _080975_, _080976_, _080977_, _080978_, _080979_, _080980_, _080981_, _080982_, _080983_, _080984_, _080985_, _080986_, _080987_, _080988_, _080989_, _080990_, _080991_, _080992_, _080993_, _080994_, _080995_, _080996_, _080997_, _080998_, _080999_, _081000_, _081001_, _081002_, _081003_, _081004_, _081005_, _081006_, _081007_, _081008_, _081009_, _081010_, _081011_, _081012_, _081013_, _081014_, _081015_, _081016_, _081017_, _081018_, _081019_, _081020_, _081021_, _081022_, _081023_, _081024_, _081025_, _081026_, _081027_, _081028_, _081029_, _081030_, _081031_, _081032_, _081033_, _081034_, _081035_, _081036_, _081037_, _081038_, _081039_, _081040_, _081041_, _081042_, _081043_, _081044_, _081045_, _081046_, _081047_, _081048_, _081049_, _081050_, _081051_, _081052_, _081053_, _081054_, _081055_, _081056_, _081057_, _081058_, _081059_, _081060_, _081061_, _081062_, _081063_, _081064_, _081065_, _081066_, _081067_, _081068_, _081069_, _081070_, _081071_, _081072_, _081073_, _081074_, _081075_, _081076_, _081077_, _081078_, _081079_, _081080_, _081081_, _081082_, _081083_, _081084_, _081085_, _081086_, _081087_, _081088_, _081089_, _081090_, _081091_, _081092_, _081093_, _081094_, _081095_, _081096_, _081097_, _081098_, _081099_, _081100_, _081101_, _081102_, _081103_, _081104_, _081105_, _081106_, _081107_, _081108_, _081109_, _081110_, _081111_, _081112_, _081113_, _081114_, _081115_, _081116_, _081117_, _081118_, _081119_, _081120_, _081121_, _081122_, _081123_, _081124_, _081125_, _081126_, _081127_, _081128_, _081129_, _081130_, _081131_, _081132_, _081133_, _081134_, _081135_, _081136_, _081137_, _081138_, _081139_, _081140_, _081141_, _081142_, _081143_, _081144_, _081145_, _081146_, _081147_, _081148_, _081149_, _081150_, _081151_, _081152_, _081153_, _081154_, _081155_, _081156_, _081157_, _081158_, _081159_, _081160_, _081161_, _081162_, _081163_, _081164_, _081165_, _081166_, _081167_, _081168_, _081169_, _081170_, _081171_, _081172_, _081173_, _081174_, _081175_, _081176_, _081177_, _081178_, _081179_, _081180_, _081181_, _081182_, _081183_, _081184_, _081185_, _081186_, _081187_, _081188_, _081189_, _081190_, _081191_, _081192_, _081193_, _081194_, _081195_, _081196_, _081197_, _081198_, _081199_, _081200_, _081201_, _081202_, _081203_, _081204_, _081205_, _081206_, _081207_, _081208_, _081209_, _081210_, _081211_, _081212_, _081213_, _081214_, _081215_, _081216_, _081217_, _081218_, _081219_, _081220_, _081221_, _081222_, _081223_, _081224_, _081225_, _081226_, _081227_, _081228_, _081229_, _081230_, _081231_, _081232_, _081233_, _081234_, _081235_, _081236_, _081237_, _081238_, _081239_, _081240_, _081241_, _081242_, _081243_, _081244_, _081245_, _081246_, _081247_, _081248_, _081249_, _081250_, _081251_, _081252_, _081253_, _081254_, _081255_, _081256_, _081257_, _081258_, _081259_, _081260_, _081261_, _081262_, _081263_, _081264_, _081265_, _081266_, _081267_, _081268_, _081269_, _081270_, _081271_, _081272_, _081273_, _081274_, _081275_, _081276_, _081277_, _081278_, _081279_, _081280_, _081281_, _081282_, _081283_, _081284_, _081285_, _081286_, _081287_, _081288_, _081289_, _081290_, _081291_, _081292_, _081293_, _081294_, _081295_, _081296_, _081297_, _081298_, _081299_, _081300_, _081301_, _081302_, _081303_, _081304_, _081305_, _081306_, _081307_, _081308_, _081309_, _081310_, _081311_, _081312_, _081313_, _081314_, _081315_, _081316_, _081317_, _081318_, _081319_, _081320_, _081321_, _081322_, _081323_, _081324_, _081325_, _081326_, _081327_, _081328_, _081329_, _081330_, _081331_, _081332_, _081333_, _081334_, _081335_, _081336_, _081337_, _081338_, _081339_, _081340_, _081341_, _081342_, _081343_, _081344_, _081345_, _081346_, _081347_, _081348_, _081349_, _081350_, _081351_, _081352_, _081353_, _081354_, _081355_, _081356_, _081357_, _081358_, _081359_, _081360_, _081361_, _081362_, _081363_, _081364_, _081365_, _081366_, _081367_, _081368_, _081369_, _081370_, _081371_, _081372_, _081373_, _081374_, _081375_, _081376_, _081377_, _081378_, _081379_, _081380_, _081381_, _081382_, _081383_, _081384_, _081385_, _081386_, _081387_, _081388_, _081389_, _081390_, _081391_, _081392_, _081393_, _081394_, _081395_, _081396_, _081397_, _081398_, _081399_, _081400_, _081401_, _081402_, _081403_, _081404_, _081405_, _081406_, _081407_, _081408_, _081409_, _081410_, _081411_, _081412_, _081413_, _081414_, _081415_, _081416_, _081417_, _081418_, _081419_, _081420_, _081421_, _081422_, _081423_, _081424_, _081425_, _081426_, _081427_, _081428_, _081429_, _081430_, _081431_, _081432_, _081433_, _081434_, _081435_, _081436_, _081437_, _081438_, _081439_, _081440_, _081441_, _081442_, _081443_, _081444_, _081445_, _081446_, _081447_, _081448_, _081449_, _081450_, _081451_, _081452_, _081453_, _081454_, _081455_, _081456_, _081457_, _081458_, _081459_, _081460_, _081461_, _081462_, _081463_, _081464_, _081465_, _081466_, _081467_, _081468_, _081469_, _081470_, _081471_, _081472_, _081473_, _081474_, _081475_, _081476_, _081477_, _081478_, _081479_, _081480_, _081481_, _081482_, _081483_, _081484_, _081485_, _081486_, _081487_, _081488_, _081489_, _081490_, _081491_, _081492_, _081493_, _081494_, _081495_, _081496_, _081497_, _081498_, _081499_, _081500_, _081501_, _081502_, _081503_, _081504_, _081505_, _081506_, _081507_, _081508_, _081509_, _081510_, _081511_, _081512_, _081513_, _081514_, _081515_, _081516_, _081517_, _081518_, _081519_, _081520_, _081521_, _081522_, _081523_, _081524_, _081525_, _081526_, _081527_, _081528_, _081529_, _081530_, _081531_, _081532_, _081533_, _081534_, _081535_, _081536_, _081537_, _081538_, _081539_, _081540_, _081541_, _081542_, _081543_, _081544_, _081545_, _081546_, _081547_, _081548_, _081549_, _081550_, _081551_, _081552_, _081553_, _081554_, _081555_, _081556_, _081557_, _081558_, _081559_, _081560_, _081561_, _081562_, _081563_, _081564_, _081565_, _081566_, _081567_, _081568_, _081569_, _081570_, _081571_, _081572_, _081573_, _081574_, _081575_, _081576_, _081577_, _081578_, _081579_, _081580_, _081581_, _081582_, _081583_, _081584_, _081585_, _081586_, _081587_, _081588_, _081589_, _081590_, _081591_, _081592_, _081593_, _081594_, _081595_, _081596_, _081597_, _081598_, _081599_, _081600_, _081601_, _081602_, _081603_, _081604_, _081605_, _081606_, _081607_, _081608_, _081609_, _081610_, _081611_, _081612_, _081613_, _081614_, _081615_, _081616_, _081617_, _081618_, _081619_, _081620_, _081621_, _081622_, _081623_, _081624_, _081625_, _081626_, _081627_, _081628_, _081629_, _081630_, _081631_, _081632_, _081633_, _081634_, _081635_, _081636_, _081637_, _081638_, _081639_, _081640_, _081641_, _081642_, _081643_, _081644_, _081645_, _081646_, _081647_, _081648_, _081649_, _081650_, _081651_, _081652_, _081653_, _081654_, _081655_, _081656_, _081657_, _081658_, _081659_, _081660_, _081661_, _081662_, _081663_, _081664_, _081665_, _081666_, _081667_, _081668_, _081669_, _081670_, _081671_, _081672_, _081673_, _081674_, _081675_, _081676_, _081677_, _081678_, _081679_, _081680_, _081681_, _081682_, _081683_, _081684_, _081685_, _081686_, _081687_, _081688_, _081689_, _081690_, _081691_, _081692_, _081693_, _081694_, _081695_, _081696_, _081697_, _081698_, _081699_, _081700_, _081701_, _081702_, _081703_, _081704_, _081705_, _081706_, _081707_, _081708_, _081709_, _081710_, _081711_, _081712_, _081713_, _081714_, _081715_, _081716_, _081717_, _081718_, _081719_, _081720_, _081721_, _081722_, _081723_, _081724_, _081725_, _081726_, _081727_, _081728_, _081729_, _081730_, _081731_, _081732_, _081733_, _081734_, _081735_, _081736_, _081737_, _081738_, _081739_, _081740_, _081741_, _081742_, _081743_, _081744_, _081745_, _081746_, _081747_, _081748_, _081749_, _081750_, _081751_, _081752_, _081753_, _081754_, _081755_, _081756_, _081757_, _081758_, _081759_, _081760_, _081761_, _081762_, _081763_, _081764_, _081765_, _081766_, _081767_, _081768_, _081769_, _081770_, _081771_, _081772_, _081773_, _081774_, _081775_, _081776_, _081777_, _081778_, _081779_, _081780_, _081781_, _081782_, _081783_, _081784_, _081785_, _081786_, _081787_, _081788_, _081789_, _081790_, _081791_, _081792_, _081793_, _081794_, _081795_, _081796_, _081797_, _081798_, _081799_, _081800_, _081801_, _081802_, _081803_, _081804_, _081805_, _081806_, _081807_, _081808_, _081809_, _081810_, _081811_, _081812_, _081813_, _081814_, _081815_, _081816_, _081817_, _081818_, _081819_, _081820_, _081821_, _081822_, _081823_, _081824_, _081825_, _081826_, _081827_, _081828_, _081829_, _081830_, _081831_, _081832_, _081833_, _081834_, _081835_, _081836_, _081837_, _081838_, _081839_, _081840_, _081841_, _081842_, _081843_, _081844_, _081845_, _081846_, _081847_, _081848_, _081849_, _081850_, _081851_, _081852_, _081853_, _081854_, _081855_, _081856_, _081857_, _081858_, _081859_, _081860_, _081861_, _081862_, _081863_, _081864_, _081865_, _081866_, _081867_, _081868_, _081869_, _081870_, _081871_, _081872_, _081873_, _081874_, _081875_, _081876_, _081877_, _081878_, _081879_, _081880_, _081881_, _081882_, _081883_, _081884_, _081885_, _081886_, _081887_, _081888_, _081889_, _081890_, _081891_, _081892_, _081893_, _081894_, _081895_, _081896_, _081897_, _081898_, _081899_, _081900_, _081901_, _081902_, _081903_, _081904_, _081905_, _081906_, _081907_, _081908_, _081909_, _081910_, _081911_, _081912_, _081913_, _081914_, _081915_, _081916_, _081917_, _081918_, _081919_, _081920_, _081921_, _081922_, _081923_, _081924_, _081925_, _081926_, _081927_, _081928_, _081929_, _081930_, _081931_, _081932_, _081933_, _081934_, _081935_, _081936_, _081937_, _081938_, _081939_, _081940_, _081941_, _081942_, _081943_, _081944_, _081945_, _081946_, _081947_, _081948_, _081949_, _081950_, _081951_, _081952_, _081953_, _081954_, _081955_, _081956_, _081957_, _081958_, _081959_, _081960_, _081961_, _081962_, _081963_, _081964_, _081965_, _081966_, _081967_, _081968_, _081969_, _081970_, _081971_, _081972_, _081973_, _081974_, _081975_, _081976_, _081977_, _081978_, _081979_, _081980_, _081981_, _081982_, _081983_, _081984_, _081985_, _081986_, _081987_, _081988_, _081989_, _081990_, _081991_, _081992_, _081993_, _081994_, _081995_, _081996_, _081997_, _081998_, _081999_, _082000_, _082001_, _082002_, _082003_, _082004_, _082005_, _082006_, _082007_, _082008_, _082009_, _082010_, _082011_, _082012_, _082013_, _082014_, _082015_, _082016_, _082017_, _082018_, _082019_, _082020_, _082021_, _082022_, _082023_, _082024_, _082025_, _082026_, _082027_, _082028_, _082029_, _082030_, _082031_, _082032_, _082033_, _082034_, _082035_, _082036_, _082037_, _082038_, _082039_, _082040_, _082041_, _082042_, _082043_, _082044_, _082045_, _082046_, _082047_, _082048_, _082049_, _082050_, _082051_, _082052_, _082053_, _082054_, _082055_, _082056_, _082057_, _082058_, _082059_, _082060_, _082061_, _082062_, _082063_, _082064_, _082065_, _082066_, _082067_, _082068_, _082069_, _082070_, _082071_, _082072_, _082073_, _082074_, _082075_, _082076_, _082077_, _082078_, _082079_, _082080_, _082081_, _082082_, _082083_, _082084_, _082085_, _082086_, _082087_, _082088_, _082089_, _082090_, _082091_, _082092_, _082093_, _082094_, _082095_, _082096_, _082097_, _082098_, _082099_, _082100_, _082101_, _082102_, _082103_, _082104_, _082105_, _082106_, _082107_, _082108_, _082109_, _082110_, _082111_, _082112_, _082113_, _082114_, _082115_, _082116_, _082117_, _082118_, _082119_, _082120_, _082121_, _082122_, _082123_, _082124_, _082125_, _082126_, _082127_, _082128_, _082129_, _082130_, _082131_, _082132_, _082133_, _082134_, _082135_, _082136_, _082137_, _082138_, _082139_, _082140_, _082141_, _082142_, _082143_, _082144_, _082145_, _082146_, _082147_, _082148_, _082149_, _082150_, _082151_, _082152_, _082153_, _082154_, _082155_, _082156_, _082157_, _082158_, _082159_, _082160_, _082161_, _082162_, _082163_, _082164_, _082165_, _082166_, _082167_, _082168_, _082169_, _082170_, _082171_, _082172_, _082173_, _082174_, _082175_, _082176_, _082177_, _082178_, _082179_, _082180_, _082181_, _082182_, _082183_, _082184_, _082185_, _082186_, _082187_, _082188_, _082189_, _082190_, _082191_, _082192_, _082193_, _082194_, _082195_, _082196_, _082197_, _082198_, _082199_, _082200_, _082201_, _082202_, _082203_, _082204_, _082205_, _082206_, _082207_, _082208_, _082209_, _082210_, _082211_, _082212_, _082213_, _082214_, _082215_, _082216_, _082217_, _082218_, _082219_, _082220_, _082221_, _082222_, _082223_, _082224_, _082225_, _082226_, _082227_, _082228_, _082229_, _082230_, _082231_, _082232_, _082233_, _082234_, _082235_, _082236_, _082237_, _082238_, _082239_, _082240_, _082241_, _082242_, _082243_, _082244_, _082245_, _082246_, _082247_, _082248_, _082249_, _082250_, _082251_, _082252_, _082253_, _082254_, _082255_, _082256_, _082257_, _082258_, _082259_, _082260_, _082261_, _082262_, _082263_, _082264_, _082265_, _082266_, _082267_, _082268_, _082269_, _082270_, _082271_, _082272_, _082273_, _082274_, _082275_, _082276_, _082277_, _082278_, _082279_, _082280_, _082281_, _082282_, _082283_, _082284_, _082285_, _082286_, _082287_, _082288_, _082289_, _082290_, _082291_, _082292_, _082293_, _082294_, _082295_, _082296_, _082297_, _082298_, _082299_, _082300_, _082301_, _082302_, _082303_, _082304_, _082305_, _082306_, _082307_, _082308_, _082309_, _082310_, _082311_, _082312_, _082313_, _082314_, _082315_, _082316_, _082317_, _082318_, _082319_, _082320_, _082321_, _082322_, _082323_, _082324_, _082325_, _082326_, _082327_, _082328_, _082329_, _082330_, _082331_, _082332_, _082333_, _082334_, _082335_, _082336_, _082337_, _082338_, _082339_, _082340_, _082341_, _082342_, _082343_, _082344_, _082345_, _082346_, _082347_, _082348_, _082349_, _082350_, _082351_, _082352_, _082353_, _082354_, _082355_, _082356_, _082357_, _082358_, _082359_, _082360_, _082361_, _082362_, _082363_, _082364_, _082365_, _082366_, _082367_, _082368_, _082369_, _082370_, _082371_, _082372_, _082373_, _082374_, _082375_, _082376_, _082377_, _082378_, _082379_, _082380_, _082381_, _082382_, _082383_, _082384_, _082385_, _082386_, _082387_, _082388_, _082389_, _082390_, _082391_, _082392_, _082393_, _082394_, _082395_, _082396_, _082397_, _082398_, _082399_, _082400_, _082401_, _082402_, _082403_, _082404_, _082405_, _082406_, _082407_, _082408_, _082409_, _082410_, _082411_, _082412_, _082413_, _082414_, _082415_, _082416_, _082417_, _082418_, _082419_, _082420_, _082421_, _082422_, _082423_, _082424_, _082425_, _082426_, _082427_, _082428_, _082429_, _082430_, _082431_, _082432_, _082433_, _082434_, _082435_, _082436_, _082437_, _082438_, _082439_, _082440_, _082441_, _082442_, _082443_, _082444_, _082445_, _082446_, _082447_, _082448_, _082449_, _082450_, _082451_, _082452_, _082453_, _082454_, _082455_, _082456_, _082457_, _082458_, _082459_, _082460_, _082461_, _082462_, _082463_, _082464_, _082465_, _082466_, _082467_, _082468_, _082469_, _082470_, _082471_, _082472_, _082473_, _082474_, _082475_, _082476_, _082477_, _082478_, _082479_, _082480_, _082481_, _082482_, _082483_, _082484_, _082485_, _082486_, _082487_, _082488_, _082489_, _082490_, _082491_, _082492_, _082493_, _082494_, _082495_, _082496_, _082497_, _082498_, _082499_, _082500_, _082501_, _082502_, _082503_, _082504_, _082505_, _082506_, _082507_, _082508_, _082509_, _082510_, _082511_, _082512_, _082513_, _082514_, _082515_, _082516_, _082517_, _082518_, _082519_, _082520_, _082521_, _082522_, _082523_, _082524_, _082525_, _082526_, _082527_, _082528_, _082529_, _082530_, _082531_, _082532_, _082533_, _082534_, _082535_, _082536_, _082537_, _082538_, _082539_, _082540_, _082541_, _082542_, _082543_, _082544_, _082545_, _082546_, _082547_, _082548_, _082549_, _082550_, _082551_, _082552_, _082553_, _082554_, _082555_, _082556_, _082557_, _082558_, _082559_, _082560_, _082561_, _082562_, _082563_, _082564_, _082565_, _082566_, _082567_, _082568_, _082569_, _082570_, _082571_, _082572_, _082573_, _082574_, _082575_, _082576_, _082577_, _082578_, _082579_, _082580_, _082581_, _082582_, _082583_, _082584_, _082585_, _082586_, _082587_, _082588_, _082589_, _082590_, _082591_, _082592_, _082593_, _082594_, _082595_, _082596_, _082597_, _082598_, _082599_, _082600_, _082601_, _082602_, _082603_, _082604_, _082605_, _082606_, _082607_, _082608_, _082609_, _082610_, _082611_, _082612_, _082613_, _082614_, _082615_, _082616_, _082617_, _082618_, _082619_, _082620_, _082621_, _082622_, _082623_, _082624_, _082625_, _082626_, _082627_, _082628_, _082629_, _082630_, _082631_, _082632_, _082633_, _082634_, _082635_, _082636_, _082637_, _082638_, _082639_, _082640_, _082641_, _082642_, _082643_, _082644_, _082645_, _082646_, _082647_, _082648_, _082649_, _082650_, _082651_, _082652_, _082653_, _082654_, _082655_, _082656_, _082657_, _082658_, _082659_, _082660_, _082661_, _082662_, _082663_, _082664_, _082665_, _082666_, _082667_, _082668_, _082669_, _082670_, _082671_, _082672_, _082673_, _082674_, _082675_, _082676_, _082677_, _082678_, _082679_, _082680_, _082681_, _082682_, _082683_, _082684_, _082685_, _082686_, _082687_, _082688_, _082689_, _082690_, _082691_, _082692_, _082693_, _082694_, _082695_, _082696_, _082697_, _082698_, _082699_, _082700_, _082701_, _082702_, _082703_, _082704_, _082705_, _082706_, _082707_, _082708_, _082709_, _082710_, _082711_, _082712_, _082713_, _082714_, _082715_, _082716_, _082717_, _082718_, _082719_, _082720_, _082721_, _082722_, _082723_, _082724_, _082725_, _082726_, _082727_, _082728_, _082729_, _082730_, _082731_, _082732_, _082733_, _082734_, _082735_, _082736_, _082737_, _082738_, _082739_, _082740_, _082741_, _082742_, _082743_, _082744_, _082745_, _082746_, _082747_, _082748_, _082749_, _082750_, _082751_, _082752_, _082753_, _082754_, _082755_, _082756_, _082757_, _082758_, _082759_, _082760_, _082761_, _082762_, _082763_, _082764_, _082765_, _082766_, _082767_, _082768_, _082769_, _082770_, _082771_, _082772_, _082773_, _082774_, _082775_, _082776_, _082777_, _082778_, _082779_, _082780_, _082781_, _082782_, _082783_, _082784_, _082785_, _082786_, _082787_, _082788_, _082789_, _082790_, _082791_, _082792_, _082793_, _082794_, _082795_, _082796_, _082797_, _082798_, _082799_, _082800_, _082801_, _082802_, _082803_, _082804_, _082805_, _082806_, _082807_, _082808_, _082809_, _082810_, _082811_, _082812_, _082813_, _082814_, _082815_, _082816_, _082817_, _082818_, _082819_, _082820_, _082821_, _082822_, _082823_, _082824_, _082825_, _082826_, _082827_, _082828_, _082829_, _082830_, _082831_, _082832_, _082833_, _082834_, _082835_, _082836_, _082837_, _082838_, _082839_, _082840_, _082841_, _082842_, _082843_, _082844_, _082845_, _082846_, _082847_, _082848_, _082849_, _082850_, _082851_, _082852_, _082853_, _082854_, _082855_, _082856_, _082857_, _082858_, _082859_, _082860_, _082861_, _082862_, _082863_, _082864_, _082865_, _082866_, _082867_, _082868_, _082869_, _082870_, _082871_, _082872_, _082873_, _082874_, _082875_, _082876_, _082877_, _082878_, _082879_, _082880_, _082881_, _082882_, _082883_, _082884_, _082885_, _082886_, _082887_, _082888_, _082889_, _082890_, _082891_, _082892_, _082893_, _082894_, _082895_, _082896_, _082897_, _082898_, _082899_, _082900_, _082901_, _082902_, _082903_, _082904_, _082905_, _082906_, _082907_, _082908_, _082909_, _082910_, _082911_, _082912_, _082913_, _082914_, _082915_, _082916_, _082917_, _082918_, _082919_, _082920_, _082921_, _082922_, _082923_, _082924_, _082925_, _082926_, _082927_, _082928_, _082929_, _082930_, _082931_, _082932_, _082933_, _082934_, _082935_, _082936_, _082937_, _082938_, _082939_, _082940_, _082941_, _082942_, _082943_, _082944_, _082945_, _082946_, _082947_, _082948_, _082949_, _082950_, _082951_, _082952_, _082953_, _082954_, _082955_, _082956_, _082957_, _082958_, _082959_, _082960_, _082961_, _082962_, _082963_, _082964_, _082965_, _082966_, _082967_, _082968_, _082969_, _082970_, _082971_, _082972_, _082973_, _082974_, _082975_, _082976_, _082977_, _082978_, _082979_, _082980_, _082981_, _082982_, _082983_, _082984_, _082985_, _082986_, _082987_, _082988_, _082989_, _082990_, _082991_, _082992_, _082993_, _082994_, _082995_, _082996_, _082997_, _082998_, _082999_, _083000_, _083001_, _083002_, _083003_, _083004_, _083005_, _083006_, _083007_, _083008_, _083009_, _083010_, _083011_, _083012_, _083013_, _083014_, _083015_, _083016_, _083017_, _083018_, _083019_, _083020_, _083021_, _083022_, _083023_, _083024_, _083025_, _083026_, _083027_, _083028_, _083029_, _083030_, _083031_, _083032_, _083033_, _083034_, _083035_, _083036_, _083037_, _083038_, _083039_, _083040_, _083041_, _083042_, _083043_, _083044_, _083045_, _083046_, _083047_, _083048_, _083049_, _083050_, _083051_, _083052_, _083053_, _083054_, _083055_, _083056_, _083057_, _083058_, _083059_, _083060_, _083061_, _083062_, _083063_, _083064_, _083065_, _083066_, _083067_, _083068_, _083069_, _083070_, _083071_, _083072_, _083073_, _083074_, _083075_, _083076_, _083077_, _083078_, _083079_, _083080_, _083081_, _083082_, _083083_, _083084_, _083085_, _083086_, _083087_, _083088_, _083089_, _083090_, _083091_, _083092_, _083093_, _083094_, _083095_, _083096_, _083097_, _083098_, _083099_, _083100_, _083101_, _083102_, _083103_, _083104_, _083105_, _083106_, _083107_, _083108_, _083109_, _083110_, _083111_, _083112_, _083113_, _083114_, _083115_, _083116_, _083117_, _083118_, _083119_, _083120_, _083121_, _083122_, _083123_, _083124_, _083125_, _083126_, _083127_, _083128_, _083129_, _083130_, _083131_, _083132_, _083133_, _083134_, _083135_, _083136_, _083137_, _083138_, _083139_, _083140_, _083141_, _083142_, _083143_, _083144_, _083145_, _083146_, _083147_, _083148_, _083149_, _083150_, _083151_, _083152_, _083153_, _083154_, _083155_, _083156_, _083157_, _083158_, _083159_, _083160_, _083161_, _083162_, _083163_, _083164_, _083165_, _083166_, _083167_, _083168_, _083169_, _083170_, _083171_, _083172_, _083173_, _083174_, _083175_, _083176_, _083177_, _083178_, _083179_, _083180_, _083181_, _083182_, _083183_, _083184_, _083185_, _083186_, _083187_, _083188_, _083189_, _083190_, _083191_, _083192_, _083193_, _083194_, _083195_, _083196_, _083197_, _083198_, _083199_, _083200_, _083201_, _083202_, _083203_, _083204_, _083205_, _083206_, _083207_, _083208_, _083209_, _083210_, _083211_, _083212_, _083213_, _083214_, _083215_, _083216_, _083217_, _083218_, _083219_, _083220_, _083221_, _083222_, _083223_, _083224_, _083225_, _083226_, _083227_, _083228_, _083229_, _083230_, _083231_, _083232_, _083233_, _083234_, _083235_, _083236_, _083237_, _083238_, _083239_, _083240_, _083241_, _083242_, _083243_, _083244_, _083245_, _083246_, _083247_, _083248_, _083249_, _083250_, _083251_, _083252_, _083253_, _083254_, _083255_, _083256_, _083257_, _083258_, _083259_, _083260_, _083261_, _083262_, _083263_, _083264_, _083265_, _083266_, _083267_, _083268_, _083269_, _083270_, _083271_, _083272_, _083273_, _083274_, _083275_, _083276_, _083277_, _083278_, _083279_, _083280_, _083281_, _083282_, _083283_, _083284_, _083285_, _083286_, _083287_, _083288_, _083289_, _083290_, _083291_, _083292_, _083293_, _083294_, _083295_, _083296_, _083297_, _083298_, _083299_, _083300_, _083301_, _083302_, _083303_, _083304_, _083305_, _083306_, _083307_, _083308_, _083309_, _083310_, _083311_, _083312_, _083313_, _083314_, _083315_, _083316_, _083317_, _083318_, _083319_, _083320_, _083321_, _083322_, _083323_, _083324_, _083325_, _083326_, _083327_, _083328_, _083329_, _083330_, _083331_, _083332_, _083333_, _083334_, _083335_, _083336_, _083337_, _083338_, _083339_, _083340_, _083341_, _083342_, _083343_, _083344_, _083345_, _083346_, _083347_, _083348_, _083349_, _083350_, _083351_, _083352_, _083353_, _083354_, _083355_, _083356_, _083357_, _083358_, _083359_, _083360_, _083361_, _083362_, _083363_, _083364_, _083365_, _083366_, _083367_, _083368_, _083369_, _083370_, _083371_, _083372_, _083373_, _083374_, _083375_, _083376_, _083377_, _083378_, _083379_, _083380_, _083381_, _083382_, _083383_, _083384_, _083385_, _083386_, _083387_, _083388_, _083389_, _083390_, _083391_, _083392_, _083393_, _083394_, _083395_, _083396_, _083397_, _083398_, _083399_, _083400_, _083401_, _083402_, _083403_, _083404_, _083405_, _083406_, _083407_, _083408_, _083409_, _083410_, _083411_, _083412_, _083413_, _083414_, _083415_, _083416_, _083417_, _083418_, _083419_, _083420_, _083421_, _083422_, _083423_, _083424_, _083425_, _083426_, _083427_, _083428_, _083429_, _083430_, _083431_, _083432_, _083433_, _083434_, _083435_, _083436_, _083437_, _083438_, _083439_, _083440_, _083441_, _083442_, _083443_, _083444_, _083445_, _083446_, _083447_, _083448_, _083449_, _083450_, _083451_, _083452_, _083453_, _083454_, _083455_, _083456_, _083457_, _083458_, _083459_, _083460_, _083461_, _083462_, _083463_, _083464_, _083465_, _083466_, _083467_, _083468_, _083469_, _083470_, _083471_, _083472_, _083473_, _083474_, _083475_, _083476_, _083477_, _083478_, _083479_, _083480_, _083481_, _083482_, _083483_, _083484_, _083485_, _083486_, _083487_, _083488_, _083489_, _083490_, _083491_, _083492_, _083493_, _083494_, _083495_, _083496_, _083497_, _083498_, _083499_, _083500_, _083501_, _083502_, _083503_, _083504_, _083505_, _083506_, _083507_, _083508_, _083509_, _083510_, _083511_, _083512_, _083513_, _083514_, _083515_, _083516_, _083517_, _083518_, _083519_, _083520_, _083521_, _083522_, _083523_, _083524_, _083525_, _083526_, _083527_, _083528_, _083529_, _083530_, _083531_, _083532_, _083533_, _083534_, _083535_, _083536_, _083537_, _083538_, _083539_, _083540_, _083541_, _083542_, _083543_, _083544_, _083545_, _083546_, _083547_, _083548_, _083549_, _083550_, _083551_, _083552_, _083553_, _083554_, _083555_, _083556_, _083557_, _083558_, _083559_, _083560_, _083561_, _083562_, _083563_, _083564_, _083565_, _083566_, _083567_, _083568_, _083569_, _083570_, _083571_, _083572_, _083573_, _083574_, _083575_, _083576_, _083577_, _083578_, _083579_, _083580_, _083581_, _083582_, _083583_, _083584_, _083585_, _083586_, _083587_, _083588_, _083589_, _083590_, _083591_, _083592_, _083593_, _083594_, _083595_, _083596_, _083597_, _083598_, _083599_, _083600_, _083601_, _083602_, _083603_, _083604_, _083605_, _083606_, _083607_, _083608_, _083609_, _083610_, _083611_, _083612_, _083613_, _083614_, _083615_, _083616_, _083617_, _083618_, _083619_, _083620_, _083621_, _083622_, _083623_, _083624_, _083625_, _083626_, _083627_, _083628_, _083629_, _083630_, _083631_, _083632_, _083633_, _083634_, _083635_, _083636_, _083637_, _083638_, _083639_, _083640_, _083641_, _083642_, _083643_, _083644_, _083645_, _083646_, _083647_, _083648_, _083649_, _083650_, _083651_, _083652_, _083653_, _083654_, _083655_, _083656_, _083657_, _083658_, _083659_, _083660_, _083661_, _083662_, _083663_, _083664_, _083665_, _083666_, _083667_, _083668_, _083669_, _083670_, _083671_, _083672_, _083673_, _083674_, _083675_, _083676_, _083677_, _083678_, _083679_, _083680_, _083681_, _083682_, _083683_, _083684_, _083685_, _083686_, _083687_, _083688_, _083689_, _083690_, _083691_, _083692_, _083693_, _083694_, _083695_, _083696_, _083697_, _083698_, _083699_, _083700_, _083701_, _083702_, _083703_, _083704_, _083705_, _083706_, _083707_, _083708_, _083709_, _083710_, _083711_, _083712_, _083713_, _083714_, _083715_, _083716_, _083717_, _083718_, _083719_, _083720_, _083721_, _083722_, _083723_, _083724_, _083725_, _083726_, _083727_, _083728_, _083729_, _083730_, _083731_, _083732_, _083733_, _083734_, _083735_, _083736_, _083737_, _083738_, _083739_, _083740_, _083741_, _083742_, _083743_, _083744_, _083745_, _083746_, _083747_, _083748_, _083749_, _083750_, _083751_, _083752_, _083753_, _083754_, _083755_, _083756_, _083757_, _083758_, _083759_, _083760_, _083761_, _083762_, _083763_, _083764_, _083765_, _083766_, _083767_, _083768_, _083769_, _083770_, _083771_, _083772_, _083773_, _083774_, _083775_, _083776_, _083777_, _083778_, _083779_, _083780_, _083781_, _083782_, _083783_, _083784_, _083785_, _083786_, _083787_, _083788_, _083789_, _083790_, _083791_, _083792_, _083793_, _083794_, _083795_, _083796_, _083797_, _083798_, _083799_, _083800_, _083801_, _083802_, _083803_, _083804_, _083805_, _083806_, _083807_, _083808_, _083809_, _083810_, _083811_, _083812_, _083813_, _083814_, _083815_, _083816_, _083817_, _083818_, _083819_, _083820_, _083821_, _083822_, _083823_, _083824_, _083825_, _083826_, _083827_, _083828_, _083829_, _083830_, _083831_, _083832_, _083833_, _083834_, _083835_, _083836_, _083837_, _083838_, _083839_, _083840_, _083841_, _083842_, _083843_, _083844_, _083845_, _083846_, _083847_, _083848_, _083849_, _083850_, _083851_, _083852_, _083853_, _083854_, _083855_, _083856_, _083857_, _083858_, _083859_, _083860_, _083861_, _083862_, _083863_, _083864_, _083865_, _083866_, _083867_, _083868_, _083869_, _083870_, _083871_, _083872_, _083873_, _083874_, _083875_, _083876_, _083877_, _083878_, _083879_, _083880_, _083881_, _083882_, _083883_, _083884_, _083885_, _083886_, _083887_, _083888_, _083889_, _083890_, _083891_, _083892_, _083893_, _083894_, _083895_, _083896_, _083897_, _083898_, _083899_, _083900_, _083901_, _083902_, _083903_, _083904_, _083905_, _083906_, _083907_, _083908_, _083909_, _083910_, _083911_, _083912_, _083913_, _083914_, _083915_, _083916_, _083917_, _083918_, _083919_, _083920_, _083921_, _083922_, _083923_, _083924_, _083925_, _083926_, _083927_, _083928_, _083929_, _083930_, _083931_, _083932_, _083933_, _083934_, _083935_, _083936_, _083937_, _083938_, _083939_, _083940_, _083941_, _083942_, _083943_, _083944_, _083945_, _083946_, _083947_, _083948_, _083949_, _083950_, _083951_, _083952_, _083953_, _083954_, _083955_, _083956_, _083957_, _083958_, _083959_, _083960_, _083961_, _083962_, _083963_, _083964_, _083965_, _083966_, _083967_, _083968_, _083969_, _083970_, _083971_, _083972_, _083973_, _083974_, _083975_, _083976_, _083977_, _083978_, _083979_, _083980_, _083981_, _083982_, _083983_, _083984_, _083985_, _083986_, _083987_, _083988_, _083989_, _083990_, _083991_, _083992_, _083993_, _083994_, _083995_, _083996_, _083997_, _083998_, _083999_, _084000_, _084001_, _084002_, _084003_, _084004_, _084005_, _084006_, _084007_, _084008_, _084009_, _084010_, _084011_, _084012_, _084013_, _084014_, _084015_, _084016_, _084017_, _084018_, _084019_, _084020_, _084021_, _084022_, _084023_, _084024_, _084025_, _084026_, _084027_, _084028_, _084029_, _084030_, _084031_, _084032_, _084033_, _084034_, _084035_, _084036_, _084037_, _084038_, _084039_, _084040_, _084041_, _084042_, _084043_, _084044_, _084045_, _084046_, _084047_, _084048_, _084049_, _084050_, _084051_, _084052_, _084053_, _084054_, _084055_, _084056_, _084057_, _084058_, _084059_, _084060_, _084061_, _084062_, _084063_, _084064_, _084065_, _084066_, _084067_, _084068_, _084069_, _084070_, _084071_, _084072_, _084073_, _084074_, _084075_, _084076_, _084077_, _084078_, _084079_, _084080_, _084081_, _084082_, _084083_, _084084_, _084085_, _084086_, _084087_, _084088_, _084089_, _084090_, _084091_, _084092_, _084093_, _084094_, _084095_, _084096_, _084097_, _084098_, _084099_, _084100_, _084101_, _084102_, _084103_, _084104_, _084105_, _084106_, _084107_, _084108_, _084109_, _084110_, _084111_, _084112_, _084113_, _084114_, _084115_, _084116_, _084117_, _084118_, _084119_, _084120_, _084121_, _084122_, _084123_, _084124_, _084125_, _084126_, _084127_, _084128_, _084129_, _084130_, _084131_, _084132_, _084133_, _084134_, _084135_, _084136_, _084137_, _084138_, _084139_, _084140_, _084141_, _084142_, _084143_, _084144_, _084145_, _084146_, _084147_, _084148_, _084149_, _084150_, _084151_, _084152_, _084153_, _084154_, _084155_, _084156_, _084157_, _084158_, _084159_, _084160_, _084161_, _084162_, _084163_, _084164_, _084165_, _084166_, _084167_, _084168_, _084169_, _084170_, _084171_, _084172_, _084173_, _084174_, _084175_, _084176_, _084177_, _084178_, _084179_, _084180_, _084181_, _084182_, _084183_, _084184_, _084185_, _084186_, _084187_, _084188_, _084189_, _084190_, _084191_, _084192_, _084193_, _084194_, _084195_, _084196_, _084197_, _084198_, _084199_, _084200_, _084201_, _084202_, _084203_, _084204_, _084205_, _084206_, _084207_, _084208_, _084209_, _084210_, _084211_, _084212_, _084213_, _084214_, _084215_, _084216_, _084217_, _084218_, _084219_, _084220_, _084221_, _084222_, _084223_, _084224_, _084225_, _084226_, _084227_, _084228_, _084229_, _084230_, _084231_, _084232_, _084233_, _084234_, _084235_, _084236_, _084237_, _084238_, _084239_, _084240_, _084241_, _084242_, _084243_, _084244_, _084245_, _084246_, _084247_, _084248_, _084249_, _084250_, _084251_, _084252_, _084253_, _084254_, _084255_, _084256_, _084257_, _084258_, _084259_, _084260_, _084261_, _084262_, _084263_, _084264_, _084265_, _084266_, _084267_, _084268_, _084269_, _084270_, _084271_, _084272_, _084273_, _084274_, _084275_, _084276_, _084277_, _084278_, _084279_, _084280_, _084281_, _084282_, _084283_, _084284_, _084285_, _084286_, _084287_, _084288_, _084289_, _084290_, _084291_, _084292_, _084293_, _084294_, _084295_, _084296_, _084297_, _084298_, _084299_, _084300_, _084301_, _084302_, _084303_, _084304_, _084305_, _084306_, _084307_, _084308_, _084309_, _084310_, _084311_, _084312_, _084313_, _084314_, _084315_, _084316_, _084317_, _084318_, _084319_, _084320_, _084321_, _084322_, _084323_, _084324_, _084325_, _084326_, _084327_, _084328_, _084329_, _084330_, _084331_, _084332_, _084333_, _084334_, _084335_, _084336_, _084337_, _084338_, _084339_, _084340_, _084341_, _084342_, _084343_, _084344_, _084345_, _084346_, _084347_, _084348_, _084349_, _084350_, _084351_, _084352_, _084353_, _084354_, _084355_, _084356_, _084357_, _084358_, _084359_, _084360_, _084361_, _084362_, _084363_, _084364_, _084365_, _084366_, _084367_, _084368_, _084369_, _084370_, _084371_, _084372_, _084373_, _084374_, _084375_, _084376_, _084377_, _084378_, _084379_, _084380_, _084381_, _084382_, _084383_, _084384_, _084385_, _084386_, _084387_, _084388_, _084389_, _084390_, _084391_, _084392_, _084393_, _084394_, _084395_, _084396_, _084397_, _084398_, _084399_, _084400_, _084401_, _084402_, _084403_, _084404_, _084405_, _084406_, _084407_, _084408_, _084409_, _084410_, _084411_, _084412_, _084413_, _084414_, _084415_, _084416_, _084417_, _084418_, _084419_, _084420_, _084421_, _084422_, _084423_, _084424_, _084425_, _084426_, _084427_, _084428_, _084429_, _084430_, _084431_, _084432_, _084433_, _084434_, _084435_, _084436_, _084437_, _084438_, _084439_, _084440_, _084441_, _084442_, _084443_, _084444_, _084445_, _084446_, _084447_, _084448_, _084449_, _084450_, _084451_, _084452_, _084453_, _084454_, _084455_, _084456_, _084457_, _084458_, _084459_, _084460_, _084461_, _084462_, _084463_, _084464_, _084465_, _084466_, _084467_, _084468_, _084469_, _084470_, _084471_, _084472_, _084473_, _084474_, _084475_, _084476_, _084477_, _084478_, _084479_, _084480_, _084481_, _084482_, _084483_, _084484_, _084485_, _084486_, _084487_, _084488_, _084489_, _084490_, _084491_, _084492_, _084493_, _084494_, _084495_, _084496_, _084497_, _084498_, _084499_, _084500_, _084501_, _084502_, _084503_, _084504_, _084505_, _084506_, _084507_, _084508_, _084509_, _084510_, _084511_, _084512_, _084513_, _084514_, _084515_, _084516_, _084517_, _084518_, _084519_, _084520_, _084521_, _084522_, _084523_, _084524_, _084525_, _084526_, _084527_, _084528_, _084529_, _084530_, _084531_, _084532_, _084533_, _084534_, _084535_, _084536_, _084537_, _084538_, _084539_, _084540_, _084541_, _084542_, _084543_, _084544_, _084545_, _084546_, _084547_, _084548_, _084549_, _084550_, _084551_, _084552_, _084553_, _084554_, _084555_, _084556_, _084557_, _084558_, _084559_, _084560_, _084561_, _084562_, _084563_, _084564_, _084565_, _084566_, _084567_, _084568_, _084569_, _084570_, _084571_, _084572_, _084573_, _084574_, _084575_, _084576_, _084577_, _084578_, _084579_, _084580_, _084581_, _084582_, _084583_, _084584_, _084585_, _084586_, _084587_, _084588_, _084589_, _084590_, _084591_, _084592_, _084593_, _084594_, _084595_, _084596_, _084597_, _084598_, _084599_, _084600_, _084601_, _084602_, _084603_, _084604_, _084605_, _084606_, _084607_, _084608_, _084609_, _084610_, _084611_, _084612_, _084613_, _084614_, _084615_, _084616_, , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , ;
  input [479:0] set1;
  input [479:0] set2;
  input set1[0], set1[1], set1[2], set1[3], set1[4], set1[5], set1[6], set1[7], set1[8], set1[9], set1[10], set1[11], set1[12], set1[13], set1[14], set1[15], set1[16], set1[17], set1[18], set1[19], set1[20], set1[21], set1[22], set1[23], set1[24], set1[25], set1[26], set1[27], set1[28], set1[29], set1[30], set1[31], set1[32], set1[33], set1[34], set1[35], set1[36], set1[37], set1[38], set1[39], set1[40], set1[41], set1[42], set1[43], set1[44], set1[45], set1[46], set1[47], set1[48], set1[49], set1[50], set1[51], set1[52], set1[53], set1[54], set1[55], set1[56], set1[57], set1[58], set1[59], set1[60], set1[61], set1[62], set1[63], set1[64], set1[65], set1[66], set1[67], set1[68], set1[69], set1[70], set1[71], set1[72], set1[73], set1[74], set1[75], set1[76], set1[77], set1[78], set1[79], set1[80], set1[81], set1[82], set1[83], set1[84], set1[85], set1[86], set1[87], set1[88], set1[89], set1[90], set1[91], set1[92], set1[93], set1[94], set1[95], set1[96], set1[97], set1[98], set1[99], set1[100], set1[101], set1[102], set1[103], set1[104], set1[105], set1[106], set1[107], set1[108], set1[109], set1[110], set1[111], set1[112], set1[113], set1[114], set1[115], set1[116], set1[117], set1[118], set1[119], set1[120], set1[121], set1[122], set1[123], set1[124], set1[125], set1[126], set1[127], set1[128], set1[129], set1[130], set1[131], set1[132], set1[133], set1[134], set1[135], set1[136], set1[137], set1[138], set1[139], set1[140], set1[141], set1[142], set1[143], set1[144], set1[145], set1[146], set1[147], set1[148], set1[149], set1[150], set1[151], set1[152], set1[153], set1[154], set1[155], set1[156], set1[157], set1[158], set1[159], set1[160], set1[161], set1[162], set1[163], set1[164], set1[165], set1[166], set1[167], set1[168], set1[169], set1[170], set1[171], set1[172], set1[173], set1[174], set1[175], set1[176], set1[177], set1[178], set1[179], set1[180], set1[181], set1[182], set1[183], set1[184], set1[185], set1[186], set1[187], set1[188], set1[189], set1[190], set1[191], set1[192], set1[193], set1[194], set1[195], set1[196], set1[197], set1[198], set1[199], set1[200], set1[201], set1[202], set1[203], set1[204], set1[205], set1[206], set1[207], set1[208], set1[209], set1[210], set1[211], set1[212], set1[213], set1[214], set1[215], set1[216], set1[217], set1[218], set1[219], set1[220], set1[221], set1[222], set1[223], set1[224], set1[225], set1[226], set1[227], set1[228], set1[229], set1[230], set1[231], set1[232], set1[233], set1[234], set1[235], set1[236], set1[237], set1[238], set1[239], set1[240], set1[241], set1[242], set1[243], set1[244], set1[245], set1[246], set1[247], set1[248], set1[249], set1[250], set1[251], set1[252], set1[253], set1[254], set1[255], set1[256], set1[257], set1[258], set1[259], set1[260], set1[261], set1[262], set1[263], set1[264], set1[265], set1[266], set1[267], set1[268], set1[269], set1[270], set1[271], set1[272], set1[273], set1[274], set1[275], set1[276], set1[277], set1[278], set1[279], set1[280], set1[281], set1[282], set1[283], set1[284], set1[285], set1[286], set1[287], set1[288], set1[289], set1[290], set1[291], set1[292], set1[293], set1[294], set1[295], set1[296], set1[297], set1[298], set1[299], set1[300], set1[301], set1[302], set1[303], set1[304], set1[305], set1[306], set1[307], set1[308], set1[309], set1[310], set1[311], set1[312], set1[313], set1[314], set1[315], set1[316], set1[317], set1[318], set1[319], set1[320], set1[321], set1[322], set1[323], set1[324], set1[325], set1[326], set1[327], set1[328], set1[329], set1[330], set1[331], set1[332], set1[333], set1[334], set1[335], set1[336], set1[337], set1[338], set1[339], set1[340], set1[341], set1[342], set1[343], set1[344], set1[345], set1[346], set1[347], set1[348], set1[349], set1[350], set1[351], set1[352], set1[353], set1[354], set1[355], set1[356], set1[357], set1[358], set1[359], set1[360], set1[361], set1[362], set1[363], set1[364], set1[365], set1[366], set1[367], set1[368], set1[369], set1[370], set1[371], set1[372], set1[373], set1[374], set1[375], set1[376], set1[377], set1[378], set1[379], set1[380], set1[381], set1[382], set1[383], set1[384], set1[385], set1[386], set1[387], set1[388], set1[389], set1[390], set1[391], set1[392], set1[393], set1[394], set1[395], set1[396], set1[397], set1[398], set1[399], set1[400], set1[401], set1[402], set1[403], set1[404], set1[405], set1[406], set1[407], set1[408], set1[409], set1[410], set1[411], set1[412], set1[413], set1[414], set1[415], set1[416], set1[417], set1[418], set1[419], set1[420], set1[421], set1[422], set1[423], set1[424], set1[425], set1[426], set1[427], set1[428], set1[429], set1[430], set1[431], set1[432], set1[433], set1[434], set1[435], set1[436], set1[437], set1[438], set1[439], set1[440], set1[441], set1[442], set1[443], set1[444], set1[445], set1[446], set1[447], set1[448], set1[449], set1[450], set1[451], set1[452], set1[453], set1[454], set1[455], set1[456], set1[457], set1[458], set1[459], set1[460], set1[461], set1[462], set1[463], set1[464], set1[465], set1[466], set1[467], set1[468], set1[469], set1[470], set1[471], set1[472], set1[473], set1[474], set1[475], set1[476], set1[477], set1[478], set1[479], set2[0], set2[1], set2[2], set2[3], set2[4], set2[5], set2[6], set2[7], set2[8], set2[9], set2[10], set2[11], set2[12], set2[13], set2[14], set2[15], set2[16], set2[17], set2[18], set2[19], set2[20], set2[21], set2[22], set2[23], set2[24], set2[25], set2[26], set2[27], set2[28], set2[29], set2[30], set2[31], set2[32], set2[33], set2[34], set2[35], set2[36], set2[37], set2[38], set2[39], set2[40], set2[41], set2[42], set2[43], set2[44], set2[45], set2[46], set2[47], set2[48], set2[49], set2[50], set2[51], set2[52], set2[53], set2[54], set2[55], set2[56], set2[57], set2[58], set2[59], set2[60], set2[61], set2[62], set2[63], set2[64], set2[65], set2[66], set2[67], set2[68], set2[69], set2[70], set2[71], set2[72], set2[73], set2[74], set2[75], set2[76], set2[77], set2[78], set2[79], set2[80], set2[81], set2[82], set2[83], set2[84], set2[85], set2[86], set2[87], set2[88], set2[89], set2[90], set2[91], set2[92], set2[93], set2[94], set2[95], set2[96], set2[97], set2[98], set2[99], set2[100], set2[101], set2[102], set2[103], set2[104], set2[105], set2[106], set2[107], set2[108], set2[109], set2[110], set2[111], set2[112], set2[113], set2[114], set2[115], set2[116], set2[117], set2[118], set2[119], set2[120], set2[121], set2[122], set2[123], set2[124], set2[125], set2[126], set2[127], set2[128], set2[129], set2[130], set2[131], set2[132], set2[133], set2[134], set2[135], set2[136], set2[137], set2[138], set2[139], set2[140], set2[141], set2[142], set2[143], set2[144], set2[145], set2[146], set2[147], set2[148], set2[149], set2[150], set2[151], set2[152], set2[153], set2[154], set2[155], set2[156], set2[157], set2[158], set2[159], set2[160], set2[161], set2[162], set2[163], set2[164], set2[165], set2[166], set2[167], set2[168], set2[169], set2[170], set2[171], set2[172], set2[173], set2[174], set2[175], set2[176], set2[177], set2[178], set2[179], set2[180], set2[181], set2[182], set2[183], set2[184], set2[185], set2[186], set2[187], set2[188], set2[189], set2[190], set2[191], set2[192], set2[193], set2[194], set2[195], set2[196], set2[197], set2[198], set2[199], set2[200], set2[201], set2[202], set2[203], set2[204], set2[205], set2[206], set2[207], set2[208], set2[209], set2[210], set2[211], set2[212], set2[213], set2[214], set2[215], set2[216], set2[217], set2[218], set2[219], set2[220], set2[221], set2[222], set2[223], set2[224], set2[225], set2[226], set2[227], set2[228], set2[229], set2[230], set2[231], set2[232], set2[233], set2[234], set2[235], set2[236], set2[237], set2[238], set2[239], set2[240], set2[241], set2[242], set2[243], set2[244], set2[245], set2[246], set2[247], set2[248], set2[249], set2[250], set2[251], set2[252], set2[253], set2[254], set2[255], set2[256], set2[257], set2[258], set2[259], set2[260], set2[261], set2[262], set2[263], set2[264], set2[265], set2[266], set2[267], set2[268], set2[269], set2[270], set2[271], set2[272], set2[273], set2[274], set2[275], set2[276], set2[277], set2[278], set2[279], set2[280], set2[281], set2[282], set2[283], set2[284], set2[285], set2[286], set2[287], set2[288], set2[289], set2[290], set2[291], set2[292], set2[293], set2[294], set2[295], set2[296], set2[297], set2[298], set2[299], set2[300], set2[301], set2[302], set2[303], set2[304], set2[305], set2[306], set2[307], set2[308], set2[309], set2[310], set2[311], set2[312], set2[313], set2[314], set2[315], set2[316], set2[317], set2[318], set2[319], set2[320], set2[321], set2[322], set2[323], set2[324], set2[325], set2[326], set2[327], set2[328], set2[329], set2[330], set2[331], set2[332], set2[333], set2[334], set2[335], set2[336], set2[337], set2[338], set2[339], set2[340], set2[341], set2[342], set2[343], set2[344], set2[345], set2[346], set2[347], set2[348], set2[349], set2[350], set2[351], set2[352], set2[353], set2[354], set2[355], set2[356], set2[357], set2[358], set2[359], set2[360], set2[361], set2[362], set2[363], set2[364], set2[365], set2[366], set2[367], set2[368], set2[369], set2[370], set2[371], set2[372], set2[373], set2[374], set2[375], set2[376], set2[377], set2[378], set2[379], set2[380], set2[381], set2[382], set2[383], set2[384], set2[385], set2[386], set2[387], set2[388], set2[389], set2[390], set2[391], set2[392], set2[393], set2[394], set2[395], set2[396], set2[397], set2[398], set2[399], set2[400], set2[401], set2[402], set2[403], set2[404], set2[405], set2[406], set2[407], set2[408], set2[409], set2[410], set2[411], set2[412], set2[413], set2[414], set2[415], set2[416], set2[417], set2[418], set2[419], set2[420], set2[421], set2[422], set2[423], set2[424], set2[425], set2[426], set2[427], set2[428], set2[429], set2[430], set2[431], set2[432], set2[433], set2[434], set2[435], set2[436], set2[437], set2[438], set2[439], set2[440], set2[441], set2[442], set2[443], set2[444], set2[445], set2[446], set2[447], set2[448], set2[449], set2[450], set2[451], set2[452], set2[453], set2[454], set2[455], set2[456], set2[457], set2[458], set2[459], set2[460], set2[461], set2[462], set2[463], set2[464], set2[465], set2[466], set2[467], set2[468], set2[469], set2[470], set2[471], set2[472], set2[473], set2[474], set2[475], set2[476], set2[477], set2[478], set2[479];
  output out[0], out[1], out[2], out[3], out[4], out[5], out[6], out[7], out[8], out[9], out[10], out[11], out[12], out[13], out[14], out[15], out[16], out[17], out[18], out[19], out[20], out[21], out[22], out[23], out[24], out[25], out[26], out[27], out[28], out[29], out[30], out[31], out[32], out[33], out[34], out[35], out[36], out[37], out[38], out[39], out[40], out[41], out[42], out[43], out[44], out[45], out[46], out[47], out[48], out[49], out[50], out[51], out[52], out[53], out[54], out[55], out[56], out[57], out[58], out[59], out[60], out[61], out[62], out[63], out[64], out[65], out[66], out[67], out[68], out[69], out[70], out[71], out[72], out[73], out[74], out[75], out[76], out[77], out[78], out[79], out[80], out[81], out[82], out[83], out[84], out[85], out[86], out[87], out[88], out[89], out[90], out[91], out[92], out[93], out[94], out[95], out[96], out[97], out[98], out[99], out[100], out[101], out[102], out[103], out[104], out[105], out[106], out[107], out[108], out[109], out[110], out[111], out[112], out[113], out[114], out[115], out[116], out[117], out[118], out[119], out[120], out[121], out[122], out[123], out[124], out[125], out[126], out[127], out[128], out[129], out[130], out[131], out[132], out[133], out[134], out[135], out[136], out[137], out[138], out[139], out[140], out[141], out[142], out[143], out[144], out[145], out[146], out[147], out[148], out[149], out[150], out[151], out[152], out[153], out[154], out[155], out[156], out[157], out[158], out[159], out[160], out[161], out[162], out[163], out[164], out[165], out[166], out[167], out[168], out[169], out[170], out[171], out[172], out[173], out[174], out[175], out[176], out[177], out[178], out[179], out[180], out[181], out[182], out[183], out[184], out[185], out[186], out[187], out[188], out[189], out[190], out[191], out[192], out[193], out[194], out[195], out[196], out[197], out[198], out[199], out[200], out[201], out[202], out[203], out[204], out[205], out[206], out[207], out[208], out[209], out[210], out[211], out[212], out[213], out[214], out[215], out[216], out[217], out[218], out[219], out[220], out[221], out[222], out[223], out[224], out[225], out[226], out[227], out[228], out[229], out[230], out[231], out[232], out[233], out[234], out[235], out[236], out[237], out[238], out[239], out[240], out[241], out[242], out[243], out[244], out[245], out[246], out[247], out[248], out[249], out[250], out[251], out[252], out[253], out[254], out[255], out[256], out[257], out[258], out[259], out[260], out[261], out[262], out[263], out[264], out[265], out[266], out[267], out[268], out[269], out[270], out[271], out[272], out[273], out[274], out[275], out[276], out[277], out[278], out[279], out[280], out[281], out[282], out[283], out[284], out[285], out[286], out[287], out[288], out[289], out[290], out[291], out[292], out[293], out[294], out[295], out[296], out[297], out[298], out[299], out[300], out[301], out[302], out[303], out[304], out[305], out[306], out[307], out[308], out[309], out[310], out[311], out[312], out[313], out[314], out[315], out[316], out[317], out[318], out[319], out[320], out[321], out[322], out[323], out[324], out[325], out[326], out[327], out[328], out[329], out[330], out[331], out[332], out[333], out[334], out[335], out[336], out[337], out[338], out[339], out[340], out[341], out[342], out[343], out[344], out[345], out[346], out[347], out[348], out[349], out[350], out[351], out[352], out[353], out[354], out[355], out[356], out[357], out[358], out[359], out[360], out[361], out[362], out[363], out[364], out[365], out[366], out[367], out[368], out[369], out[370], out[371], out[372], out[373], out[374], out[375], out[376], out[377], out[378], out[379], out[380], out[381], out[382], out[383], out[384], out[385], out[386], out[387], out[388], out[389], out[390], out[391], out[392], out[393], out[394], out[395], out[396], out[397], out[398], out[399], out[400], out[401], out[402], out[403], out[404], out[405], out[406], out[407], out[408], out[409], out[410], out[411], out[412], out[413], out[414], out[415], out[416], out[417], out[418], out[419], out[420], out[421], out[422], out[423], out[424], out[425], out[426], out[427], out[428], out[429], out[430], out[431], out[432], out[433], out[434], out[435], out[436], out[437], out[438], out[439], out[440], out[441], out[442], out[443], out[444], out[445], out[446], out[447], out[448], out[449], out[450], out[451], out[452], out[453], out[454], out[455], out[456], out[457], out[458], out[459], out[460], out[461], out[462], out[463], out[464], out[465], out[466], out[467], out[468], out[469], out[470], out[471], out[472], out[473], out[474], out[475], out[476], out[477], out[478], out[479], out[480], out[481], out[482], out[483], out[484], out[485], out[486], out[487], out[488], out[489], out[490], out[491], out[492], out[493], out[494], out[495], out[496], out[497], out[498], out[499], out[500], out[501], out[502], out[503], out[504], out[505], out[506], out[507], out[508], out[509], out[510], out[511], out[512], out[513], out[514], out[515], out[516], out[517], out[518], out[519], out[520], out[521], out[522], out[523], out[524], out[525], out[526], out[527], out[528], out[529], out[530], out[531], out[532], out[533], out[534], out[535], out[536], out[537], out[538], out[539], out[540], out[541], out[542], out[543], out[544], out[545], out[546], out[547], out[548], out[549], out[550], out[551], out[552], out[553], out[554], out[555], out[556], out[557], out[558], out[559], out[560], out[561], out[562], out[563], out[564], out[565], out[566], out[567], out[568], out[569], out[570], out[571], out[572], out[573], out[574], out[575], out[576], out[577], out[578], out[579], out[580], out[581], out[582], out[583], out[584], out[585], out[586], out[587], out[588], out[589], out[590], out[591], out[592], out[593], out[594], out[595], out[596], out[597], out[598], out[599], out[600], out[601], out[602], out[603], out[604], out[605], out[606], out[607], out[608], out[609], out[610], out[611], out[612], out[613], out[614], out[615], out[616], out[617], out[618], out[619], out[620], out[621], out[622], out[623], out[624], out[625], out[626], out[627], out[628], out[629], out[630], out[631], out[632], out[633], out[634], out[635], out[636], out[637], out[638], out[639], out[640], out[641], out[642], out[643], out[644], out[645], out[646], out[647], out[648], out[649], out[650], out[651], out[652], out[653], out[654], out[655], out[656], out[657], out[658], out[659], out[660], out[661], out[662], out[663], out[664], out[665], out[666], out[667], out[668], out[669], out[670], out[671], out[672], out[673], out[674], out[675], out[676], out[677], out[678], out[679], out[680], out[681], out[682], out[683], out[684], out[685], out[686], out[687], out[688], out[689], out[690], out[691], out[692], out[693], out[694], out[695], out[696], out[697], out[698], out[699], out[700], out[701], out[702], out[703], out[704], out[705], out[706], out[707], out[708], out[709], out[710], out[711], out[712], out[713], out[714], out[715], out[716], out[717], out[718], out[719], out[720], out[721], out[722], out[723], out[724], out[725], out[726], out[727], out[728], out[729], out[730], out[731], out[732], out[733], out[734], out[735], out[736], out[737], out[738], out[739], out[740], out[741], out[742], out[743], out[744], out[745], out[746], out[747], out[748], out[749], out[750], out[751], out[752], out[753], out[754], out[755], out[756], out[757], out[758], out[759], out[760], out[761], out[762], out[763], out[764], out[765], out[766], out[767], out[768], out[769], out[770], out[771], out[772], out[773], out[774], out[775], out[776], out[777], out[778], out[779], out[780], out[781], out[782], out[783], out[784], out[785], out[786], out[787], out[788], out[789], out[790], out[791], out[792], out[793], out[794], out[795], out[796], out[797], out[798], out[799], out[800], out[801], out[802], out[803], out[804], out[805], out[806], out[807], out[808], out[809], out[810], out[811], out[812], out[813], out[814], out[815], out[816], out[817], out[818], out[819], out[820], out[821], out[822], out[823], out[824], out[825], out[826], out[827], out[828], out[829], out[830], out[831], out[832], out[833], out[834], out[835], out[836], out[837], out[838], out[839], out[840], out[841], out[842], out[843], out[844], out[845], out[846], out[847], out[848], out[849], out[850], out[851], out[852], out[853], out[854], out[855], out[856], out[857], out[858], out[859], out[860], out[861], out[862], out[863], out[864], out[865], out[866], out[867], out[868], out[869], out[870], out[871], out[872], out[873], out[874], out[875], out[876], out[877], out[878], out[879], out[880], out[881], out[882], out[883], out[884], out[885], out[886], out[887], out[888], out[889], out[890], out[891], out[892], out[893], out[894], out[895], out[896], out[897], out[898], out[899], out[900], out[901], out[902], out[903], out[904], out[905], out[906], out[907], out[908], out[909], out[910], out[911], out[912], out[913], out[914], out[915], out[916], out[917], out[918], out[919], out[920], out[921], out[922], out[923], out[924], out[925], out[926], out[927], out[928], out[929], out[930], out[931], out[932], out[933], out[934], out[935], out[936], out[937], out[938], out[939], out[940], out[941], out[942], out[943], out[944], out[945], out[946], out[947], out[948], out[949], out[950], out[951], out[952], out[953], out[954], out[955], out[956], out[957], out[958], out[959], out[960], out[961], out[962], out[963], out[964], out[965], out[966], out[967], out[968], out[969], out[970], out[971], out[972], out[973], out[974], out[975];
  not g_084617_(out[261], _052972_);
  not g_084618_(out[262], _052983_);
  not g_084619_(out[260], _052994_);
  not g_084620_(out[259], _053005_);
  not g_084621_(out[258], _053016_);
  not g_084622_(out[257], _053027_);
  not g_084623_(out[241], _053038_);
  not g_084624_(out[279], _053049_);
  not g_084625_(out[280], _053060_);
  not g_084626_(out[277], _053071_);
  not g_084627_(out[278], _053082_);
  not g_084628_(out[275], _053093_);
  not g_084629_(out[276], _053104_);
  not g_084630_(out[274], _053115_);
  not g_084631_(out[273], _053126_);
  not g_084632_(out[281], _053137_);
  not g_084633_(out[295], _053148_);
  not g_084634_(out[296], _053159_);
  not g_084635_(out[293], _053170_);
  not g_084636_(out[294], _053181_);
  not g_084637_(out[291], _053192_);
  not g_084638_(out[292], _053203_);
  not g_084639_(out[290], _053214_);
  not g_084640_(out[289], _053225_);
  not g_084641_(out[297], _053236_);
  not g_084642_(out[311], _053247_);
  not g_084643_(out[312], _053258_);
  not g_084644_(out[309], _053269_);
  not g_084645_(out[310], _053280_);
  not g_084646_(out[308], _053291_);
  not g_084647_(out[307], _053302_);
  not g_084648_(out[306], _053313_);
  not g_084649_(out[305], _053324_);
  not g_084650_(out[313], _053335_);
  not g_084651_(out[327], _053346_);
  not g_084652_(out[328], _053357_);
  not g_084653_(out[325], _053368_);
  not g_084654_(out[326], _053379_);
  not g_084655_(out[323], _053390_);
  not g_084656_(out[324], _053401_);
  not g_084657_(out[322], _053412_);
  not g_084658_(out[321], _053423_);
  not g_084659_(out[329], _053434_);
  not g_084660_(out[343], _053445_);
  not g_084661_(out[344], _053456_);
  not g_084662_(out[341], _053467_);
  not g_084663_(out[342], _053478_);
  not g_084664_(out[339], _053489_);
  not g_084665_(out[340], _053500_);
  not g_084666_(out[338], _053511_);
  not g_084667_(out[337], _053522_);
  not g_084668_(out[345], _053533_);
  not g_084669_(out[359], _053544_);
  not g_084670_(out[360], _053555_);
  not g_084671_(out[357], _053566_);
  not g_084672_(out[358], _053577_);
  not g_084673_(out[355], _053588_);
  not g_084674_(out[356], _053599_);
  not g_084675_(out[354], _053610_);
  not g_084676_(out[353], _053621_);
  not g_084677_(out[361], _053632_);
  not g_084678_(out[375], _053643_);
  not g_084679_(out[376], _053654_);
  not g_084680_(out[373], _053665_);
  not g_084681_(out[374], _053676_);
  not g_084682_(out[371], _053687_);
  not g_084683_(out[372], _053698_);
  not g_084684_(out[370], _053709_);
  not g_084685_(out[369], _053720_);
  not g_084686_(out[377], _053731_);
  not g_084687_(out[391], _053742_);
  not g_084688_(out[392], _053753_);
  not g_084689_(out[389], _053764_);
  not g_084690_(out[390], _053775_);
  not g_084691_(out[387], _053786_);
  not g_084692_(out[388], _053797_);
  not g_084693_(out[386], _053808_);
  not g_084694_(out[385], _053819_);
  not g_084695_(out[393], _053830_);
  not g_084696_(out[407], _053841_);
  not g_084697_(out[408], _053852_);
  not g_084698_(out[405], _053863_);
  not g_084699_(out[406], _053874_);
  not g_084700_(out[403], _053885_);
  not g_084701_(out[404], _053896_);
  not g_084702_(out[402], _053907_);
  not g_084703_(out[401], _053918_);
  not g_084704_(out[409], _053929_);
  not g_084705_(out[423], _053940_);
  not g_084706_(out[424], _053951_);
  not g_084707_(out[421], _053962_);
  not g_084708_(out[422], _053973_);
  not g_084709_(out[419], _053984_);
  not g_084710_(out[420], _053995_);
  not g_084711_(out[418], _054006_);
  not g_084712_(out[417], _054017_);
  not g_084713_(out[425], _054028_);
  not g_084714_(out[439], _054039_);
  not g_084715_(out[440], _054050_);
  not g_084716_(out[437], _054061_);
  not g_084717_(out[438], _054072_);
  not g_084718_(out[435], _054083_);
  not g_084719_(out[436], _054094_);
  not g_084720_(out[434], _054105_);
  not g_084721_(out[433], _054116_);
  not g_084722_(out[441], _054127_);
  not g_084723_(out[455], _054138_);
  not g_084724_(out[456], _054149_);
  not g_084725_(out[453], _054160_);
  not g_084726_(out[454], _054171_);
  not g_084727_(out[451], _054182_);
  not g_084728_(out[452], _054193_);
  not g_084729_(out[450], _054204_);
  not g_084730_(out[449], _054215_);
  not g_084731_(out[457], _054226_);
  not g_084732_(out[471], _054237_);
  not g_084733_(out[472], _054248_);
  not g_084734_(out[469], _054259_);
  not g_084735_(out[470], _054270_);
  not g_084736_(out[467], _054281_);
  not g_084737_(out[468], _054292_);
  not g_084738_(out[466], _054303_);
  not g_084739_(out[465], _054314_);
  not g_084740_(out[473], _054325_);
  not g_084741_(out[945], _054336_);
  not g_084742_(out[480], _054347_);
  not g_084743_(out[491], _054358_);
  not g_084744_(out[487], _054369_);
  not g_084745_(out[486], _054380_);
  not g_084746_(out[485], _054391_);
  not g_084747_(out[484], _054402_);
  not g_084748_(out[481], _054413_);
  not g_084749_(out[482], _054424_);
  not g_084750_(out[483], _054435_);
  not g_084751_(out[488], _054446_);
  not g_084752_(out[489], _054457_);
  not g_084753_(out[490], _054468_);
  not g_084754_(out[507], _054479_);
  not g_084755_(out[503], _054490_);
  not g_084756_(out[502], _054501_);
  not g_084757_(out[501], _054512_);
  not g_084758_(out[500], _054523_);
  not g_084759_(out[497], _054534_);
  not g_084760_(out[496], _054545_);
  not g_084761_(out[498], _054556_);
  not g_084762_(out[499], _054567_);
  not g_084763_(out[504], _054578_);
  not g_084764_(out[505], _054589_);
  not g_084765_(out[506], _054600_);
  not g_084766_(out[523], _054611_);
  not g_084767_(out[519], _054622_);
  not g_084768_(out[518], _054633_);
  not g_084769_(out[517], _054644_);
  not g_084770_(out[516], _054655_);
  not g_084771_(out[513], _054666_);
  not g_084772_(out[512], _054677_);
  not g_084773_(out[514], _054688_);
  not g_084774_(out[515], _054699_);
  not g_084775_(out[520], _054710_);
  not g_084776_(out[521], _054721_);
  not g_084777_(out[522], _054732_);
  not g_084778_(out[539], _054743_);
  not g_084779_(out[535], _054754_);
  not g_084780_(out[534], _054765_);
  not g_084781_(out[533], _054776_);
  not g_084782_(out[532], _054787_);
  not g_084783_(out[529], _054798_);
  not g_084784_(out[528], _054809_);
  not g_084785_(out[530], _054820_);
  not g_084786_(out[531], _054831_);
  not g_084787_(out[536], _054842_);
  not g_084788_(out[537], _054853_);
  not g_084789_(out[538], _054864_);
  not g_084790_(out[555], _054875_);
  not g_084791_(out[551], _054886_);
  not g_084792_(out[550], _054897_);
  not g_084793_(out[549], _054908_);
  not g_084794_(out[548], _054919_);
  not g_084795_(out[545], _054930_);
  not g_084796_(out[544], _054941_);
  not g_084797_(out[546], _054952_);
  not g_084798_(out[547], _054963_);
  not g_084799_(out[552], _054974_);
  not g_084800_(out[553], _054985_);
  not g_084801_(out[554], _054996_);
  not g_084802_(out[571], _055007_);
  not g_084803_(out[567], _055018_);
  not g_084804_(out[566], _055029_);
  not g_084805_(out[565], _055040_);
  not g_084806_(out[564], _055051_);
  not g_084807_(out[561], _055062_);
  not g_084808_(out[560], _055073_);
  not g_084809_(out[562], _055084_);
  not g_084810_(out[563], _055095_);
  not g_084811_(out[568], _055106_);
  not g_084812_(out[569], _055117_);
  not g_084813_(out[570], _055128_);
  not g_084814_(out[587], _055139_);
  not g_084815_(out[583], _055150_);
  not g_084816_(out[582], _055161_);
  not g_084817_(out[581], _055172_);
  not g_084818_(out[580], _055183_);
  not g_084819_(out[577], _055194_);
  not g_084820_(out[576], _055205_);
  not g_084821_(out[578], _055216_);
  not g_084822_(out[579], _055227_);
  not g_084823_(out[584], _055238_);
  not g_084824_(out[585], _055249_);
  not g_084825_(out[586], _055260_);
  not g_084826_(out[603], _055271_);
  not g_084827_(out[599], _055282_);
  not g_084828_(out[598], _055293_);
  not g_084829_(out[597], _055304_);
  not g_084830_(out[596], _055315_);
  not g_084831_(out[593], _055326_);
  not g_084832_(out[592], _055337_);
  not g_084833_(out[594], _055348_);
  not g_084834_(out[595], _055359_);
  not g_084835_(out[600], _055370_);
  not g_084836_(out[601], _055381_);
  not g_084837_(out[602], _055392_);
  not g_084838_(out[619], _055403_);
  not g_084839_(out[615], _055414_);
  not g_084840_(out[614], _055425_);
  not g_084841_(out[613], _055436_);
  not g_084842_(out[612], _055447_);
  not g_084843_(out[609], _055458_);
  not g_084844_(out[608], _055469_);
  not g_084845_(out[610], _055480_);
  not g_084846_(out[611], _055491_);
  not g_084847_(out[616], _055502_);
  not g_084848_(out[617], _055513_);
  not g_084849_(out[618], _055524_);
  not g_084850_(out[635], _055535_);
  not g_084851_(out[631], _055546_);
  not g_084852_(out[630], _055557_);
  not g_084853_(out[629], _055568_);
  not g_084854_(out[628], _055579_);
  not g_084855_(out[625], _055590_);
  not g_084856_(out[624], _055601_);
  not g_084857_(out[626], _055612_);
  not g_084858_(out[627], _055623_);
  not g_084859_(out[632], _055634_);
  not g_084860_(out[633], _055645_);
  not g_084861_(out[634], _055656_);
  not g_084862_(out[651], _055667_);
  not g_084863_(out[647], _055678_);
  not g_084864_(out[646], _055689_);
  not g_084865_(out[645], _055700_);
  not g_084866_(out[644], _055711_);
  not g_084867_(out[641], _055722_);
  not g_084868_(out[640], _055733_);
  not g_084869_(out[642], _055744_);
  not g_084870_(out[643], _055755_);
  not g_084871_(out[648], _055766_);
  not g_084872_(out[649], _055777_);
  not g_084873_(out[650], _055788_);
  not g_084874_(out[667], _055799_);
  not g_084875_(out[663], _055810_);
  not g_084876_(out[662], _055821_);
  not g_084877_(out[661], _055832_);
  not g_084878_(out[660], _055843_);
  not g_084879_(out[657], _055854_);
  not g_084880_(out[656], _055865_);
  not g_084881_(out[658], _055876_);
  not g_084882_(out[659], _055887_);
  not g_084883_(out[664], _055898_);
  not g_084884_(out[665], _055909_);
  not g_084885_(out[666], _055920_);
  not g_084886_(out[683], _055931_);
  not g_084887_(out[679], _055942_);
  not g_084888_(out[678], _055953_);
  not g_084889_(out[677], _055964_);
  not g_084890_(out[676], _000010_);
  not g_084891_(out[673], _000021_);
  not g_084892_(out[672], _000032_);
  not g_084893_(out[674], _000043_);
  not g_084894_(out[675], _000054_);
  not g_084895_(out[680], _000065_);
  not g_084896_(out[681], _000076_);
  not g_084897_(out[682], _000087_);
  not g_084898_(out[699], _000098_);
  not g_084899_(out[695], _000109_);
  not g_084900_(out[694], _000120_);
  not g_084901_(out[693], _000131_);
  not g_084902_(out[692], _000142_);
  not g_084903_(out[689], _000153_);
  not g_084904_(out[688], _000164_);
  not g_084905_(out[690], _000175_);
  not g_084906_(out[691], _000186_);
  not g_084907_(out[696], _000197_);
  not g_084908_(out[697], _000208_);
  not g_084909_(out[698], _000219_);
  not g_084910_(out[715], _000230_);
  not g_084911_(out[711], _000241_);
  not g_084912_(out[710], _000252_);
  not g_084913_(out[709], _000263_);
  not g_084914_(out[708], _000274_);
  not g_084915_(out[705], _000285_);
  not g_084916_(out[704], _000296_);
  not g_084917_(out[706], _000307_);
  not g_084918_(out[707], _000318_);
  not g_084919_(out[712], _000329_);
  not g_084920_(out[713], _000340_);
  not g_084921_(out[714], _000351_);
  not g_084922_(out[731], _000362_);
  not g_084923_(out[727], _000373_);
  not g_084924_(out[726], _000384_);
  not g_084925_(out[725], _000395_);
  not g_084926_(out[724], _000406_);
  not g_084927_(out[721], _000417_);
  not g_084928_(out[720], _000428_);
  not g_084929_(out[722], _000439_);
  not g_084930_(out[723], _000450_);
  not g_084931_(out[728], _000461_);
  not g_084932_(out[729], _000472_);
  not g_084933_(out[730], _000483_);
  not g_084934_(out[747], _000494_);
  not g_084935_(out[743], _000505_);
  not g_084936_(out[742], _000516_);
  not g_084937_(out[741], _000527_);
  not g_084938_(out[740], _000538_);
  not g_084939_(out[737], _000549_);
  not g_084940_(out[736], _000560_);
  not g_084941_(out[738], _000571_);
  not g_084942_(out[739], _000582_);
  not g_084943_(out[744], _000593_);
  not g_084944_(out[745], _000604_);
  not g_084945_(out[746], _000615_);
  not g_084946_(out[763], _000626_);
  not g_084947_(out[759], _000637_);
  not g_084948_(out[758], _000648_);
  not g_084949_(out[757], _000659_);
  not g_084950_(out[756], _000670_);
  not g_084951_(out[753], _000681_);
  not g_084952_(out[752], _000692_);
  not g_084953_(out[754], _000703_);
  not g_084954_(out[755], _000714_);
  not g_084955_(out[760], _000725_);
  not g_084956_(out[761], _000736_);
  not g_084957_(out[762], _000747_);
  not g_084958_(out[779], _000758_);
  not g_084959_(out[775], _000769_);
  not g_084960_(out[774], _000780_);
  not g_084961_(out[773], _000791_);
  not g_084962_(out[772], _000802_);
  not g_084963_(out[769], _000813_);
  not g_084964_(out[768], _000824_);
  not g_084965_(out[770], _000835_);
  not g_084966_(out[771], _000846_);
  not g_084967_(out[776], _000857_);
  not g_084968_(out[777], _000868_);
  not g_084969_(out[778], _000879_);
  not g_084970_(out[795], _000890_);
  not g_084971_(out[791], _000901_);
  not g_084972_(out[790], _000912_);
  not g_084973_(out[789], _000923_);
  not g_084974_(out[788], _000934_);
  not g_084975_(out[785], _000945_);
  not g_084976_(out[784], _000956_);
  not g_084977_(out[786], _000967_);
  not g_084978_(out[787], _000978_);
  not g_084979_(out[792], _000989_);
  not g_084980_(out[793], _001000_);
  not g_084981_(out[794], _001011_);
  not g_084982_(out[811], _001022_);
  not g_084983_(out[807], _001033_);
  not g_084984_(out[806], _001044_);
  not g_084985_(out[805], _001055_);
  not g_084986_(out[804], _001066_);
  not g_084987_(out[801], _001077_);
  not g_084988_(out[800], _001088_);
  not g_084989_(out[802], _001099_);
  not g_084990_(out[803], _001110_);
  not g_084991_(out[808], _001121_);
  not g_084992_(out[809], _001132_);
  not g_084993_(out[810], _001143_);
  not g_084994_(out[827], _001154_);
  not g_084995_(out[823], _001165_);
  not g_084996_(out[822], _001176_);
  not g_084997_(out[821], _001187_);
  not g_084998_(out[820], _001198_);
  not g_084999_(out[817], _001209_);
  not g_085000_(out[816], _001220_);
  not g_085001_(out[818], _001231_);
  not g_085002_(out[819], _001242_);
  not g_085003_(out[824], _001253_);
  not g_085004_(out[825], _001264_);
  not g_085005_(out[826], _001275_);
  not g_085006_(out[843], _001286_);
  not g_085007_(out[839], _001297_);
  not g_085008_(out[838], _001308_);
  not g_085009_(out[837], _001319_);
  not g_085010_(out[836], _001330_);
  not g_085011_(out[833], _001341_);
  not g_085012_(out[832], _001352_);
  not g_085013_(out[834], _001363_);
  not g_085014_(out[835], _001374_);
  not g_085015_(out[840], _001385_);
  not g_085016_(out[841], _001396_);
  not g_085017_(out[842], _001407_);
  not g_085018_(out[859], _001418_);
  not g_085019_(out[855], _001429_);
  not g_085020_(out[854], _001440_);
  not g_085021_(out[853], _001451_);
  not g_085022_(out[852], _001462_);
  not g_085023_(out[849], _001473_);
  not g_085024_(out[848], _001484_);
  not g_085025_(out[850], _001495_);
  not g_085026_(out[851], _001506_);
  not g_085027_(out[856], _001517_);
  not g_085028_(out[857], _001528_);
  not g_085029_(out[858], _001539_);
  not g_085030_(out[875], _001550_);
  not g_085031_(out[871], _001561_);
  not g_085032_(out[870], _001572_);
  not g_085033_(out[869], _001583_);
  not g_085034_(out[868], _001594_);
  not g_085035_(out[865], _001605_);
  not g_085036_(out[864], _001616_);
  not g_085037_(out[866], _001627_);
  not g_085038_(out[867], _001638_);
  not g_085039_(out[872], _001649_);
  not g_085040_(out[873], _001660_);
  not g_085041_(out[874], _001671_);
  not g_085042_(out[891], _001682_);
  not g_085043_(out[887], _001693_);
  not g_085044_(out[886], _001704_);
  not g_085045_(out[885], _001715_);
  not g_085046_(out[884], _001726_);
  not g_085047_(out[881], _001737_);
  not g_085048_(out[880], _001748_);
  not g_085049_(out[882], _001759_);
  not g_085050_(out[883], _001770_);
  not g_085051_(out[888], _001781_);
  not g_085052_(out[889], _001792_);
  not g_085053_(out[890], _001803_);
  not g_085054_(out[907], _001814_);
  not g_085055_(out[903], _001825_);
  not g_085056_(out[902], _001836_);
  not g_085057_(out[901], _001847_);
  not g_085058_(out[900], _001858_);
  not g_085059_(out[897], _001869_);
  not g_085060_(out[896], _001880_);
  not g_085061_(out[898], _001891_);
  not g_085062_(out[899], _001902_);
  not g_085063_(out[904], _001913_);
  not g_085064_(out[905], _001924_);
  not g_085065_(out[906], _001935_);
  not g_085066_(out[923], _001946_);
  not g_085067_(out[919], _001957_);
  not g_085068_(out[918], _001968_);
  not g_085069_(out[917], _001979_);
  not g_085070_(out[916], _001990_);
  not g_085071_(out[913], _002001_);
  not g_085072_(out[912], _002012_);
  not g_085073_(out[914], _002023_);
  not g_085074_(out[915], _002034_);
  not g_085075_(out[920], _002045_);
  not g_085076_(out[921], _002056_);
  not g_085077_(out[922], _002067_);
  not g_085078_(out[935], _002078_);
  not g_085079_(out[933], _002089_);
  not g_085080_(out[932], _002100_);
  not g_085081_(out[929], _002111_);
  not g_085082_(out[928], _002122_);
  not g_085083_(out[930], _002133_);
  not g_085084_(out[931], _002144_);
  not g_085085_(out[936], _002155_);
  not g_085086_(out[937], _002166_);
  not g_085087_(out[938], _002177_);
  not g_085088_(out[951], _002188_);
  not g_085089_(out[950], _002199_);
  not g_085090_(out[949], _002210_);
  not g_085091_(out[948], _002221_);
  not g_085092_(out[944], _002232_);
  not g_085093_(out[946], _002243_);
  not g_085094_(out[947], _002254_);
  not g_085095_(out[952], _002265_);
  not g_085096_(out[953], _002276_);
  not g_085097_(out[954], _002287_);
  not g_085098_(out[11], _002298_);
  not g_085099_(out[7], _002309_);
  not g_085100_(out[6], _002320_);
  not g_085101_(out[5], _002331_);
  not g_085102_(out[4], _002342_);
  not g_085103_(out[1], _002353_);
  not g_085104_(out[0], _002364_);
  not g_085105_(out[2], _002375_);
  not g_085106_(out[3], _002386_);
  not g_085107_(out[8], _002397_);
  not g_085108_(out[9], _002408_);
  not g_085109_(out[10], _002419_);
  not g_085110_(out[27], _002430_);
  not g_085111_(out[23], _002441_);
  not g_085112_(out[22], _002452_);
  not g_085113_(out[21], _002463_);
  not g_085114_(out[20], _002474_);
  not g_085115_(out[17], _002485_);
  not g_085116_(out[16], _002496_);
  not g_085117_(out[18], _002507_);
  not g_085118_(out[19], _002518_);
  not g_085119_(out[24], _002529_);
  not g_085120_(out[25], _002540_);
  not g_085121_(out[26], _002551_);
  not g_085122_(out[43], _002562_);
  not g_085123_(out[39], _002573_);
  not g_085124_(out[38], _002584_);
  not g_085125_(out[37], _002595_);
  not g_085126_(out[36], _002606_);
  not g_085127_(out[33], _002617_);
  not g_085128_(out[32], _002628_);
  not g_085129_(out[34], _002639_);
  not g_085130_(out[35], _002650_);
  not g_085131_(out[40], _002661_);
  not g_085132_(out[41], _002672_);
  not g_085133_(out[42], _002683_);
  not g_085134_(out[59], _002694_);
  not g_085135_(out[55], _002705_);
  not g_085136_(out[54], _002716_);
  not g_085137_(out[53], _002727_);
  not g_085138_(out[52], _002738_);
  not g_085139_(out[49], _002749_);
  not g_085140_(out[48], _002760_);
  not g_085141_(out[50], _002771_);
  not g_085142_(out[51], _002782_);
  not g_085143_(out[56], _002793_);
  not g_085144_(out[57], _002804_);
  not g_085145_(out[58], _002815_);
  not g_085146_(out[75], _002826_);
  not g_085147_(out[71], _002837_);
  not g_085148_(out[70], _002848_);
  not g_085149_(out[69], _002859_);
  not g_085150_(out[68], _002870_);
  not g_085151_(out[65], _002881_);
  not g_085152_(out[64], _002892_);
  not g_085153_(out[66], _002903_);
  not g_085154_(out[67], _002914_);
  not g_085155_(out[72], _002925_);
  not g_085156_(out[73], _002936_);
  not g_085157_(out[74], _002947_);
  not g_085158_(out[91], _002958_);
  not g_085159_(out[87], _002969_);
  not g_085160_(out[86], _002980_);
  not g_085161_(out[85], _002991_);
  not g_085162_(out[84], _003002_);
  not g_085163_(out[81], _003013_);
  not g_085164_(out[80], _003024_);
  not g_085165_(out[82], _003035_);
  not g_085166_(out[83], _003046_);
  not g_085167_(out[88], _003057_);
  not g_085168_(out[89], _003068_);
  not g_085169_(out[90], _003079_);
  not g_085170_(out[107], _003090_);
  not g_085171_(out[103], _003101_);
  not g_085172_(out[102], _003112_);
  not g_085173_(out[101], _003123_);
  not g_085174_(out[100], _003134_);
  not g_085175_(out[97], _003145_);
  not g_085176_(out[96], _003156_);
  not g_085177_(out[98], _003167_);
  not g_085178_(out[99], _003178_);
  not g_085179_(out[104], _003189_);
  not g_085180_(out[105], _003200_);
  not g_085181_(out[106], _003211_);
  not g_085182_(out[123], _003222_);
  not g_085183_(out[119], _003233_);
  not g_085184_(out[118], _003244_);
  not g_085185_(out[117], _003255_);
  not g_085186_(out[116], _003266_);
  not g_085187_(out[113], _003277_);
  not g_085188_(out[112], _003288_);
  not g_085189_(out[114], _003299_);
  not g_085190_(out[115], _003310_);
  not g_085191_(out[120], _003321_);
  not g_085192_(out[121], _003332_);
  not g_085193_(out[122], _003343_);
  not g_085194_(out[139], _003354_);
  not g_085195_(out[135], _003365_);
  not g_085196_(out[134], _003376_);
  not g_085197_(out[133], _003387_);
  not g_085198_(out[132], _003398_);
  not g_085199_(out[129], _003409_);
  not g_085200_(out[128], _003420_);
  not g_085201_(out[130], _003431_);
  not g_085202_(out[131], _003442_);
  not g_085203_(out[136], _003453_);
  not g_085204_(out[137], _003464_);
  not g_085205_(out[138], _003475_);
  not g_085206_(out[155], _003486_);
  not g_085207_(out[151], _003497_);
  not g_085208_(out[150], _003508_);
  not g_085209_(out[149], _003519_);
  not g_085210_(out[148], _003530_);
  not g_085211_(out[145], _003541_);
  not g_085212_(out[144], _003552_);
  not g_085213_(out[146], _003563_);
  not g_085214_(out[147], _003574_);
  not g_085215_(out[152], _003585_);
  not g_085216_(out[153], _003596_);
  not g_085217_(out[154], _003607_);
  not g_085218_(out[171], _003618_);
  not g_085219_(out[167], _003629_);
  not g_085220_(out[166], _003640_);
  not g_085221_(out[165], _003651_);
  not g_085222_(out[164], _003662_);
  not g_085223_(out[161], _003673_);
  not g_085224_(out[160], _003684_);
  not g_085225_(out[162], _003695_);
  not g_085226_(out[163], _003706_);
  not g_085227_(out[168], _003717_);
  not g_085228_(out[169], _003728_);
  not g_085229_(out[170], _003739_);
  not g_085230_(out[187], _003750_);
  not g_085231_(out[183], _003761_);
  not g_085232_(out[182], _003772_);
  not g_085233_(out[181], _003783_);
  not g_085234_(out[180], _003794_);
  not g_085235_(out[177], _003805_);
  not g_085236_(out[176], _003816_);
  not g_085237_(out[178], _003827_);
  not g_085238_(out[179], _003838_);
  not g_085239_(out[184], _003849_);
  not g_085240_(out[185], _003860_);
  not g_085241_(out[186], _003871_);
  not g_085242_(out[203], _003882_);
  not g_085243_(out[199], _003893_);
  not g_085244_(out[198], _003904_);
  not g_085245_(out[197], _003915_);
  not g_085246_(out[196], _003926_);
  not g_085247_(out[193], _003937_);
  not g_085248_(out[192], _003948_);
  not g_085249_(out[194], _003959_);
  not g_085250_(out[195], _003970_);
  not g_085251_(out[200], _003981_);
  not g_085252_(out[219], _003992_);
  not g_085253_(out[215], _004003_);
  not g_085254_(out[214], _004014_);
  not g_085255_(out[213], _004025_);
  not g_085256_(out[212], _004036_);
  not g_085257_(out[209], _004047_);
  not g_085258_(out[208], _004058_);
  not g_085259_(out[210], _004069_);
  not g_085260_(out[211], _004080_);
  not g_085261_(out[216], _004091_);
  not g_085262_(out[217], _004102_);
  not g_085263_(out[218], _004113_);
  not g_085264_(out[235], _004124_);
  not g_085265_(out[231], _004135_);
  not g_085266_(out[230], _004146_);
  not g_085267_(out[229], _004157_);
  not g_085268_(out[228], _004168_);
  not g_085269_(out[225], _004179_);
  not g_085270_(out[224], _004190_);
  not g_085271_(out[226], _004201_);
  not g_085272_(out[227], _004212_);
  not g_085273_(out[232], _004223_);
  not g_085274_(out[234], _004234_);
  not g_085275_(out[251], _004245_);
  not g_085276_(out[247], _004256_);
  not g_085277_(out[246], _004267_);
  not g_085278_(out[245], _004278_);
  not g_085279_(out[244], _004289_);
  not g_085280_(out[240], _004300_);
  not g_085281_(out[242], _004311_);
  not g_085282_(out[243], _004322_);
  not g_085283_(out[248], _004333_);
  not g_085284_(out[249], _004344_);
  not g_085285_(out[250], _004355_);
  not g_085286_(out[267], _004366_);
  not g_085287_(out[263], _004377_);
  not g_085288_(out[256], _004388_);
  not g_085289_(out[264], _004399_);
  not g_085290_(out[265], _004410_);
  not g_085291_(out[266], _004421_);
  not g_085292_(out[283], _004432_);
  not g_085293_(out[272], _004443_);
  not g_085294_(out[282], _004454_);
  not g_085295_(out[299], _004465_);
  not g_085296_(out[288], _004476_);
  not g_085297_(out[298], _004487_);
  not g_085298_(out[315], _004498_);
  not g_085299_(out[304], _004509_);
  not g_085300_(out[314], _004520_);
  not g_085301_(out[331], _004531_);
  not g_085302_(out[320], _004542_);
  not g_085303_(out[330], _004553_);
  not g_085304_(out[347], _004564_);
  not g_085305_(out[336], _004575_);
  not g_085306_(out[346], _004586_);
  not g_085307_(out[363], _004597_);
  not g_085308_(out[352], _004608_);
  not g_085309_(out[362], _004619_);
  not g_085310_(out[379], _004630_);
  not g_085311_(out[368], _004641_);
  not g_085312_(out[378], _004652_);
  not g_085313_(out[395], _004663_);
  not g_085314_(out[384], _004674_);
  not g_085315_(out[394], _004685_);
  not g_085316_(out[411], _004696_);
  not g_085317_(out[400], _004707_);
  not g_085318_(out[410], _004718_);
  not g_085319_(out[427], _004729_);
  not g_085320_(out[416], _004740_);
  not g_085321_(out[426], _004751_);
  not g_085322_(out[443], _004762_);
  not g_085323_(out[432], _004773_);
  not g_085324_(out[442], _004784_);
  not g_085325_(out[459], _004795_);
  not g_085326_(out[448], _004806_);
  not g_085327_(out[458], _004817_);
  not g_085328_(out[475], _004828_);
  not g_085329_(out[464], _004839_);
  and g_085330_(out[65], out[66], _004850_);
  or g_085331_(out[68], out[67], _004861_);
  or g_085332_(out[67], _004850_, _004872_);
  or g_085333_(_004850_, _004861_, _004883_);
  or g_085334_(out[69], _004883_, _004894_);
  and g_085335_(out[70], _004894_, _004905_);
  and g_085336_(out[71], _004905_, _004916_);
  or g_085337_(out[72], _004916_, _004927_);
  or g_085338_(out[73], _004927_, _004938_);
  or g_085339_(out[74], _004938_, _004949_);
  xor g_085340_(_002826_, _004949_, _004960_);
  xor g_085341_(out[75], _004949_, _004971_);
  and g_085342_(out[49], out[50], _004982_);
  or g_085343_(out[52], out[51], _004993_);
  or g_085344_(out[51], _004982_, _005004_);
  or g_085345_(_004982_, _004993_, _005015_);
  or g_085346_(out[53], _005015_, _005026_);
  and g_085347_(out[54], _005026_, _005037_);
  and g_085348_(out[55], _005037_, _005048_);
  or g_085349_(out[56], _005048_, _005059_);
  or g_085350_(out[57], _005059_, _005070_);
  or g_085351_(out[58], _005070_, _005081_);
  xor g_085352_(_002694_, _005081_, _005092_);
  xor g_085353_(out[59], _005081_, _005103_);
  xor g_085354_(out[58], _005070_, _005114_);
  xor g_085355_(_002815_, _005070_, _005125_);
  and g_085356_(out[33], out[34], _005136_);
  or g_085357_(out[36], out[35], _005147_);
  or g_085358_(out[35], _005136_, _005158_);
  or g_085359_(_005136_, _005147_, _005169_);
  or g_085360_(out[37], _005169_, _005180_);
  and g_085361_(out[38], _005180_, _005191_);
  and g_085362_(out[39], _005191_, _005202_);
  or g_085363_(out[40], _005202_, _005213_);
  or g_085364_(out[41], _005213_, _005224_);
  or g_085365_(out[42], _005224_, _005235_);
  xor g_085366_(out[42], _005224_, _005246_);
  xor g_085367_(_002683_, _005224_, _005257_);
  xor g_085368_(out[39], _005191_, _005268_);
  xor g_085369_(_002573_, _005191_, _005279_);
  and g_085370_(out[1], out[2], _005290_);
  or g_085371_(out[4], out[3], _005301_);
  not g_085372_(_005301_, _005312_);
  or g_085373_(out[3], _005290_, _005323_);
  or g_085374_(_005290_, _005301_, _005334_);
  or g_085375_(out[5], _005334_, _005345_);
  and g_085376_(out[6], _005345_, _005356_);
  and g_085377_(out[7], _005356_, _005367_);
  xor g_085378_(out[7], _005356_, _005378_);
  xor g_085379_(_002309_, _005356_, _005389_);
  or g_085380_(out[8], _005367_, _005400_);
  or g_085381_(out[9], _005400_, _005411_);
  or g_085382_(out[10], _005411_, _005422_);
  xor g_085383_(_002298_, _005422_, _005433_);
  xor g_085384_(out[11], _005422_, _005444_);
  and g_085385_(out[17], out[18], _005455_);
  or g_085386_(out[20], out[19], _005466_);
  not g_085387_(_005466_, _005477_);
  or g_085388_(out[19], _005455_, _005488_);
  or g_085389_(_005455_, _005466_, _005499_);
  or g_085390_(out[21], _005499_, _005510_);
  and g_085391_(out[22], _005510_, _005521_);
  and g_085392_(out[23], _005521_, _005532_);
  or g_085393_(out[24], _005532_, _005543_);
  or g_085394_(out[25], _005543_, _005554_);
  or g_085395_(out[26], _005554_, _005565_);
  xor g_085396_(_002430_, _005565_, _005576_);
  xor g_085397_(out[27], _005565_, _005587_);
  and g_085398_(_005433_, _005587_, _005598_);
  or g_085399_(_005444_, _005576_, _005609_);
  xor g_085400_(out[23], _005521_, _005620_);
  xor g_085401_(_002441_, _005521_, _005631_);
  and g_085402_(_005389_, _005620_, _005642_);
  or g_085403_(_005378_, _005631_, _005653_);
  xor g_085404_(out[6], _005345_, _005664_);
  xor g_085405_(_002320_, _005345_, _005675_);
  xor g_085406_(out[22], _005510_, _005686_);
  xor g_085407_(_002452_, _005510_, _005697_);
  and g_085408_(_005664_, _005697_, _005708_);
  or g_085409_(_005675_, _005686_, _005719_);
  xor g_085410_(out[3], _005290_, _005730_);
  xor g_085411_(_002386_, _005290_, _005741_);
  xor g_085412_(out[19], _005455_, _005752_);
  xor g_085413_(_002518_, _005455_, _005763_);
  and g_085414_(_005730_, _005763_, _005774_);
  or g_085415_(_005741_, _005752_, _005785_);
  and g_085416_(_005741_, _005752_, _005796_);
  or g_085417_(_005730_, _005763_, _005807_);
  or g_085418_(out[17], out[18], _005818_);
  xor g_085419_(out[17], out[18], _005829_);
  xor g_085420_(_002485_, out[18], _005840_);
  or g_085421_(out[1], out[2], _005851_);
  xor g_085422_(out[1], out[2], _005862_);
  not g_085423_(_005862_, _005873_);
  and g_085424_(_005840_, _005862_, _005884_);
  or g_085425_(_005829_, _005873_, _005895_);
  or g_085426_(_005840_, _005862_, _005906_);
  xor g_085427_(_005829_, _005862_, _005917_);
  or g_085428_(_005796_, _005917_, _005928_);
  and g_085429_(_005785_, _005895_, _005939_);
  and g_085430_(_005807_, _005906_, _005950_);
  and g_085431_(_005939_, _005950_, _005961_);
  or g_085432_(_005774_, _005928_, _005972_);
  or g_085433_(out[1], _002485_, _005983_);
  not g_085434_(_005983_, _005994_);
  and g_085435_(out[1], _002485_, _006005_);
  or g_085436_(_002353_, out[17], _006016_);
  and g_085437_(_002364_, out[16], _006027_);
  or g_085438_(out[0], _002496_, _006038_);
  and g_085439_(_005983_, _006038_, _006049_);
  xor g_085440_(out[1], out[17], _006060_);
  and g_085441_(_006016_, _006049_, _006071_);
  or g_085442_(_006027_, _006060_, _006082_);
  and g_085443_(_005983_, _006082_, _006093_);
  or g_085444_(_005994_, _006071_, _006104_);
  and g_085445_(_005961_, _006104_, _006115_);
  or g_085446_(_005972_, _006093_, _006126_);
  and g_085447_(_005785_, _005884_, _006137_);
  or g_085448_(_005774_, _005895_, _006148_);
  and g_085449_(_005807_, _006148_, _006159_);
  or g_085450_(_005796_, _006137_, _006170_);
  and g_085451_(_006126_, _006159_, _006181_);
  or g_085452_(_006115_, _006170_, _006192_);
  xor g_085453_(out[4], _005323_, _006203_);
  xor g_085454_(_002342_, _005323_, _006214_);
  xor g_085455_(out[20], _005488_, _006225_);
  xor g_085456_(_002474_, _005488_, _006236_);
  and g_085457_(_006203_, _006236_, _006247_);
  or g_085458_(_006214_, _006225_, _006258_);
  and g_085459_(out[0], _002496_, _006269_);
  or g_085460_(_002364_, out[16], _006280_);
  and g_085461_(_006071_, _006280_, _006291_);
  or g_085462_(_006082_, _006269_, _006302_);
  and g_085463_(_005961_, _006291_, _006313_);
  or g_085464_(_005972_, _006302_, _006324_);
  and g_085465_(_006258_, _006324_, _006335_);
  or g_085466_(_006247_, _006313_, _006346_);
  and g_085467_(_006192_, _006335_, _006357_);
  or g_085468_(_006181_, _006346_, _006368_);
  xor g_085469_(out[5], _005334_, _006379_);
  xor g_085470_(_002331_, _005334_, _006390_);
  xor g_085471_(out[21], _005499_, _006401_);
  xor g_085472_(_002463_, _005499_, _006412_);
  and g_085473_(_006390_, _006401_, _006423_);
  or g_085474_(_006379_, _006412_, _006434_);
  and g_085475_(_006214_, _006225_, _006445_);
  or g_085476_(_006203_, _006236_, _006456_);
  and g_085477_(_006434_, _006456_, _006467_);
  or g_085478_(_006423_, _006445_, _006478_);
  and g_085479_(_006368_, _006467_, _006489_);
  or g_085480_(_006357_, _006478_, _006500_);
  and g_085481_(_006379_, _006412_, _006511_);
  or g_085482_(_006390_, _006401_, _006522_);
  and g_085483_(_005675_, _005686_, _006533_);
  or g_085484_(_005664_, _005697_, _006544_);
  and g_085485_(_006522_, _006544_, _006555_);
  or g_085486_(_006511_, _006533_, _006566_);
  and g_085487_(_006500_, _006555_, _006577_);
  or g_085488_(_006489_, _006566_, _006588_);
  and g_085489_(_005719_, _006588_, _006599_);
  or g_085490_(_005708_, _006577_, _006610_);
  and g_085491_(_005653_, _006610_, _006621_);
  or g_085492_(_005642_, _006599_, _006632_);
  and g_085493_(_005378_, _005631_, _006643_);
  or g_085494_(_005389_, _005620_, _006654_);
  xor g_085495_(out[24], _005532_, _006665_);
  xor g_085496_(_002529_, _005532_, _006676_);
  xor g_085497_(out[8], _005367_, _006687_);
  xor g_085498_(_002397_, _005367_, _006698_);
  and g_085499_(_006665_, _006698_, _006709_);
  or g_085500_(_006676_, _006687_, _006720_);
  and g_085501_(_006654_, _006720_, _006731_);
  or g_085502_(_006643_, _006709_, _006742_);
  and g_085503_(_006632_, _006731_, _006753_);
  or g_085504_(_006621_, _006742_, _006764_);
  xor g_085505_(out[25], _005543_, _006775_);
  xor g_085506_(_002540_, _005543_, _006786_);
  xor g_085507_(out[9], _005400_, _006797_);
  xor g_085508_(_002408_, _005400_, _006808_);
  and g_085509_(_006786_, _006797_, _006819_);
  or g_085510_(_006775_, _006808_, _006830_);
  and g_085511_(_006676_, _006687_, _006841_);
  or g_085512_(_006665_, _006698_, _006852_);
  and g_085513_(_006830_, _006852_, _006863_);
  or g_085514_(_006819_, _006841_, _006874_);
  and g_085515_(_006764_, _006863_, _006885_);
  or g_085516_(_006753_, _006874_, _006896_);
  and g_085517_(_006775_, _006808_, _006907_);
  or g_085518_(_006786_, _006797_, _006918_);
  xor g_085519_(out[10], _005411_, _006929_);
  xor g_085520_(_002419_, _005411_, _006940_);
  xor g_085521_(out[26], _005554_, _006951_);
  xor g_085522_(_002551_, _005554_, _006962_);
  and g_085523_(_006940_, _006951_, _006973_);
  or g_085524_(_006929_, _006962_, _006984_);
  and g_085525_(_006918_, _006984_, _006995_);
  or g_085526_(_006907_, _006973_, _007006_);
  and g_085527_(_006896_, _006995_, _007017_);
  or g_085528_(_006885_, _007006_, _007028_);
  and g_085529_(_005444_, _005576_, _007039_);
  or g_085530_(_005433_, _005587_, _007050_);
  and g_085531_(_006929_, _006962_, _007061_);
  or g_085532_(_006940_, _006951_, _007072_);
  and g_085533_(_007050_, _007072_, _007083_);
  or g_085534_(_007039_, _007061_, _007094_);
  and g_085535_(_007028_, _007083_, _007105_);
  or g_085536_(_007017_, _007094_, _007116_);
  and g_085537_(_005609_, _007116_, _007127_);
  or g_085538_(_005598_, _007105_, _007138_);
  and g_085539_(_005389_, _007127_, _007149_);
  or g_085540_(_005378_, _007138_, _007160_);
  and g_085541_(_005631_, _007138_, _007171_);
  or g_085542_(_005620_, _007127_, _007182_);
  and g_085543_(_007160_, _007182_, _007193_);
  or g_085544_(_007149_, _007171_, _007204_);
  and g_085545_(_005279_, _007193_, _007215_);
  or g_085546_(_005268_, _007204_, _007226_);
  xor g_085547_(out[38], _005180_, _007237_);
  xor g_085548_(_002584_, _005180_, _007248_);
  and g_085549_(_005675_, _007127_, _007259_);
  or g_085550_(_005664_, _007138_, _007270_);
  and g_085551_(_005697_, _007138_, _007281_);
  or g_085552_(_005686_, _007127_, _007292_);
  and g_085553_(_007270_, _007292_, _007303_);
  or g_085554_(_007259_, _007281_, _007314_);
  and g_085555_(_007248_, _007303_, _007325_);
  or g_085556_(_007237_, _007314_, _007336_);
  and g_085557_(_007226_, _007336_, _007347_);
  or g_085558_(_007215_, _007325_, _007358_);
  xor g_085559_(out[37], _005169_, _007369_);
  xor g_085560_(_002595_, _005169_, _007380_);
  and g_085561_(_006379_, _007127_, _007391_);
  or g_085562_(_006390_, _007138_, _007402_);
  and g_085563_(_006401_, _007138_, _007413_);
  or g_085564_(_006412_, _007127_, _007424_);
  and g_085565_(_007402_, _007424_, _007435_);
  or g_085566_(_007391_, _007413_, _007446_);
  and g_085567_(_007369_, _007435_, _007457_);
  or g_085568_(_007380_, _007446_, _007468_);
  xor g_085569_(out[36], _005158_, _007479_);
  xor g_085570_(_002606_, _005158_, _007490_);
  and g_085571_(_006203_, _007127_, _007501_);
  or g_085572_(_006214_, _007138_, _007512_);
  and g_085573_(_006225_, _007138_, _007523_);
  or g_085574_(_006236_, _007127_, _007534_);
  and g_085575_(_007512_, _007534_, _007545_);
  or g_085576_(_007501_, _007523_, _007556_);
  and g_085577_(_007479_, _007545_, _007567_);
  or g_085578_(_007490_, _007556_, _007578_);
  and g_085579_(_007468_, _007578_, _007589_);
  or g_085580_(_007457_, _007567_, _007600_);
  and g_085581_(_007380_, _007446_, _007611_);
  or g_085582_(_007369_, _007435_, _007622_);
  and g_085583_(_007490_, _007556_, _007633_);
  or g_085584_(_007479_, _007545_, _007644_);
  and g_085585_(_007622_, _007644_, _007655_);
  or g_085586_(_007611_, _007633_, _007666_);
  and g_085587_(_007589_, _007655_, _007677_);
  or g_085588_(_007600_, _007666_, _007688_);
  xor g_085589_(out[35], _005136_, _007699_);
  xor g_085590_(_002650_, _005136_, _007710_);
  and g_085591_(_005730_, _007127_, _007721_);
  or g_085592_(_005741_, _007138_, _007732_);
  and g_085593_(_005752_, _007138_, _007743_);
  or g_085594_(_005763_, _007127_, _007754_);
  and g_085595_(_007732_, _007754_, _007765_);
  or g_085596_(_007721_, _007743_, _007776_);
  and g_085597_(_007710_, _007776_, _007787_);
  not g_085598_(_007787_, _007798_);
  and g_085599_(_007699_, _007765_, _007809_);
  or g_085600_(_007710_, _007776_, _007820_);
  or g_085601_(out[33], out[34], _007831_);
  xor g_085602_(out[33], out[34], _007842_);
  xor g_085603_(_002617_, out[34], _007853_);
  and g_085604_(_005840_, _007138_, _007864_);
  or g_085605_(_005829_, _007127_, _007875_);
  and g_085606_(_005873_, _007127_, _007886_);
  or g_085607_(_005862_, _007138_, _007897_);
  and g_085608_(_007875_, _007897_, _007908_);
  or g_085609_(_007864_, _007886_, _007919_);
  and g_085610_(_007853_, _007908_, _007930_);
  or g_085611_(_007842_, _007919_, _007941_);
  and g_085612_(_007820_, _007941_, _007952_);
  or g_085613_(_007809_, _007930_, _007963_);
  and g_085614_(_007798_, _007963_, _007974_);
  or g_085615_(_007787_, _007952_, _007985_);
  and g_085616_(_007842_, _007919_, _007996_);
  or g_085617_(_007853_, _007908_, _008007_);
  and g_085618_(_007798_, _008007_, _008018_);
  or g_085619_(_007787_, _007996_, _008029_);
  and g_085620_(_007952_, _008018_, _008040_);
  or g_085621_(_007963_, _008029_, _008051_);
  or g_085622_(_002485_, _007127_, _008062_);
  or g_085623_(_002353_, _007138_, _008073_);
  and g_085624_(_008062_, _008073_, _008084_);
  and g_085625_(out[33], _008084_, _008095_);
  not g_085626_(_008095_, _008106_);
  and g_085627_(_007600_, _007622_, _008117_);
  or g_085628_(_007589_, _007611_, _008128_);
  and g_085629_(_002364_, _007127_, _008139_);
  or g_085630_(out[0], _007138_, _008150_);
  and g_085631_(_002496_, _007138_, _008161_);
  or g_085632_(out[16], _007127_, _008172_);
  and g_085633_(_008150_, _008172_, _008183_);
  or g_085634_(_008139_, _008161_, _008194_);
  and g_085635_(out[32], _008194_, _008205_);
  or g_085636_(_002628_, _008183_, _008216_);
  xor g_085637_(out[33], _008084_, _008227_);
  xor g_085638_(_002617_, _008084_, _008238_);
  and g_085639_(_008216_, _008227_, _008249_);
  or g_085640_(_008205_, _008238_, _008260_);
  and g_085641_(_007677_, _008249_, _008271_);
  or g_085642_(_007688_, _008260_, _008282_);
  and g_085643_(_008040_, _008271_, _008293_);
  or g_085644_(_008051_, _008282_, _008304_);
  and g_085645_(_008106_, _008260_, _008315_);
  or g_085646_(_008095_, _008249_, _008326_);
  and g_085647_(_008040_, _008326_, _008337_);
  or g_085648_(_008051_, _008315_, _008348_);
  and g_085649_(_007985_, _008348_, _008359_);
  or g_085650_(_007974_, _008337_, _008370_);
  and g_085651_(_007677_, _008370_, _008381_);
  or g_085652_(_007688_, _008359_, _008392_);
  and g_085653_(_008128_, _008392_, _008403_);
  or g_085654_(_008117_, _008381_, _008414_);
  and g_085655_(_007237_, _007314_, _008425_);
  or g_085656_(_007248_, _007303_, _008436_);
  and g_085657_(_008414_, _008436_, _008447_);
  or g_085658_(_008403_, _008425_, _008458_);
  and g_085659_(_007347_, _008458_, _008469_);
  or g_085660_(_007358_, _008447_, _008480_);
  and g_085661_(_005433_, _005576_, _008491_);
  or g_085662_(_005444_, _005587_, _008502_);
  xor g_085663_(_002562_, _005235_, _008513_);
  xor g_085664_(out[43], _005235_, _008524_);
  and g_085665_(_008491_, _008524_, _008535_);
  or g_085666_(_008502_, _008513_, _008546_);
  and g_085667_(_006929_, _007127_, _008557_);
  or g_085668_(_006940_, _007138_, _008568_);
  and g_085669_(_006951_, _007138_, _008579_);
  or g_085670_(_006962_, _007127_, _008590_);
  and g_085671_(_008568_, _008590_, _008601_);
  or g_085672_(_008557_, _008579_, _008612_);
  and g_085673_(_005246_, _008601_, _008623_);
  or g_085674_(_005257_, _008612_, _008634_);
  and g_085675_(_008546_, _008634_, _008645_);
  or g_085676_(_008535_, _008623_, _008656_);
  and g_085677_(_008502_, _008513_, _008667_);
  or g_085678_(_008491_, _008524_, _008678_);
  and g_085679_(_005257_, _008612_, _008689_);
  or g_085680_(_005246_, _008601_, _008700_);
  and g_085681_(_008678_, _008700_, _008711_);
  or g_085682_(_008667_, _008689_, _008722_);
  xor g_085683_(out[41], _005213_, _008733_);
  xor g_085684_(_002672_, _005213_, _008744_);
  and g_085685_(_006797_, _007127_, _008755_);
  or g_085686_(_006808_, _007138_, _008766_);
  and g_085687_(_006775_, _007138_, _008777_);
  or g_085688_(_006786_, _007127_, _008788_);
  and g_085689_(_008766_, _008788_, _008799_);
  or g_085690_(_008755_, _008777_, _008810_);
  and g_085691_(_008744_, _008810_, _008821_);
  or g_085692_(_008733_, _008799_, _008832_);
  and g_085693_(_008645_, _008711_, _008843_);
  or g_085694_(_008656_, _008722_, _008854_);
  and g_085695_(_008832_, _008843_, _008865_);
  or g_085696_(_008821_, _008854_, _008876_);
  and g_085697_(_008733_, _008799_, _008887_);
  or g_085698_(_008744_, _008810_, _008898_);
  xor g_085699_(out[40], _005202_, _008909_);
  xor g_085700_(_002661_, _005202_, _008920_);
  and g_085701_(_006665_, _007138_, _008931_);
  or g_085702_(_006676_, _007127_, _008942_);
  and g_085703_(_006687_, _007127_, _008953_);
  or g_085704_(_006698_, _007138_, _008964_);
  and g_085705_(_008942_, _008964_, _008975_);
  or g_085706_(_008931_, _008953_, _008986_);
  and g_085707_(_008909_, _008975_, _008997_);
  or g_085708_(_008920_, _008986_, _009008_);
  and g_085709_(_008898_, _009008_, _009019_);
  or g_085710_(_008887_, _008997_, _009030_);
  and g_085711_(_008920_, _008986_, _009041_);
  or g_085712_(_008909_, _008975_, _009052_);
  and g_085713_(_009019_, _009052_, _009063_);
  or g_085714_(_009030_, _009041_, _009074_);
  and g_085715_(_008865_, _009063_, _009085_);
  or g_085716_(_008876_, _009074_, _009096_);
  and g_085717_(_005268_, _007204_, _009107_);
  or g_085718_(_005279_, _007193_, _009118_);
  and g_085719_(_009085_, _009118_, _009129_);
  or g_085720_(_009096_, _009107_, _009140_);
  and g_085721_(_008480_, _009129_, _009151_);
  or g_085722_(_008469_, _009140_, _009162_);
  and g_085723_(_008656_, _008678_, _009173_);
  or g_085724_(_008645_, _008667_, _009184_);
  and g_085725_(_008865_, _009030_, _009195_);
  or g_085726_(_008876_, _009019_, _009206_);
  and g_085727_(_009184_, _009206_, _009217_);
  or g_085728_(_009173_, _009195_, _009228_);
  and g_085729_(_009162_, _009217_, _009239_);
  or g_085730_(_009151_, _009228_, _009250_);
  and g_085731_(_002628_, _008183_, _009261_);
  or g_085732_(out[32], _008194_, _009272_);
  and g_085733_(_008436_, _009118_, _009283_);
  or g_085734_(_008425_, _009107_, _009294_);
  and g_085735_(_009272_, _009283_, _009305_);
  or g_085736_(_009261_, _009294_, _009316_);
  and g_085737_(_007347_, _009305_, _009327_);
  or g_085738_(_007358_, _009316_, _009338_);
  and g_085739_(_008293_, _009327_, _009349_);
  or g_085740_(_008304_, _009338_, _009360_);
  and g_085741_(_009085_, _009349_, _009371_);
  or g_085742_(_009096_, _009360_, _009382_);
  and g_085743_(_009250_, _009382_, _009393_);
  or g_085744_(_009239_, _009371_, _009404_);
  and g_085745_(_005246_, _009393_, _009415_);
  or g_085746_(_005257_, _009404_, _009426_);
  and g_085747_(_008612_, _009404_, _009437_);
  or g_085748_(_008601_, _009393_, _009448_);
  and g_085749_(_009426_, _009448_, _009459_);
  or g_085750_(_009415_, _009437_, _009470_);
  and g_085751_(_005114_, _009459_, _009481_);
  or g_085752_(_005125_, _009470_, _009492_);
  and g_085753_(_008524_, _009393_, _009503_);
  or g_085754_(_008513_, _009404_, _009514_);
  and g_085755_(_008502_, _009404_, _009525_);
  or g_085756_(_008491_, _009393_, _009536_);
  and g_085757_(_009514_, _009536_, _009547_);
  or g_085758_(_009503_, _009525_, _009558_);
  and g_085759_(_005103_, _009547_, _009569_);
  or g_085760_(_005092_, _009558_, _009580_);
  and g_085761_(_009492_, _009580_, _009591_);
  or g_085762_(_009481_, _009569_, _009602_);
  and g_085763_(_005125_, _009470_, _009613_);
  or g_085764_(_005114_, _009459_, _009624_);
  and g_085765_(_005092_, _009558_, _009635_);
  or g_085766_(_005103_, _009547_, _009646_);
  and g_085767_(_009624_, _009646_, _009657_);
  or g_085768_(_009613_, _009635_, _009668_);
  and g_085769_(_009591_, _009657_, _009679_);
  or g_085770_(_009602_, _009668_, _009690_);
  xor g_085771_(out[56], _005048_, _009701_);
  xor g_085772_(_002793_, _005048_, _009712_);
  and g_085773_(_008986_, _009404_, _009723_);
  or g_085774_(_008975_, _009393_, _009734_);
  and g_085775_(_008909_, _009393_, _009745_);
  or g_085776_(_008920_, _009404_, _009756_);
  and g_085777_(_009734_, _009756_, _009767_);
  or g_085778_(_009723_, _009745_, _009778_);
  and g_085779_(_009701_, _009767_, _009789_);
  or g_085780_(_009712_, _009778_, _009800_);
  xor g_085781_(out[57], _005059_, _009811_);
  xor g_085782_(_002804_, _005059_, _009822_);
  and g_085783_(_008810_, _009404_, _009833_);
  or g_085784_(_008799_, _009393_, _009844_);
  and g_085785_(_008733_, _009393_, _009855_);
  or g_085786_(_008744_, _009404_, _009866_);
  and g_085787_(_009844_, _009866_, _009877_);
  or g_085788_(_009833_, _009855_, _009888_);
  and g_085789_(_009811_, _009877_, _009899_);
  or g_085790_(_009822_, _009888_, _009910_);
  and g_085791_(_009800_, _009910_, _009921_);
  or g_085792_(_009789_, _009899_, _009932_);
  and g_085793_(_009822_, _009888_, _009943_);
  or g_085794_(_009811_, _009877_, _009954_);
  and g_085795_(_009712_, _009778_, _009965_);
  or g_085796_(_009701_, _009767_, _009976_);
  xor g_085797_(out[55], _005037_, _009987_);
  xor g_085798_(_002705_, _005037_, _009998_);
  and g_085799_(_007193_, _009404_, _010009_);
  or g_085800_(_007204_, _009393_, _010020_);
  and g_085801_(_005268_, _009393_, _010031_);
  or g_085802_(_005279_, _009404_, _010042_);
  and g_085803_(_010020_, _010042_, _010053_);
  or g_085804_(_010009_, _010031_, _010064_);
  and g_085805_(_009987_, _010053_, _010075_);
  or g_085806_(_009998_, _010064_, _010086_);
  and g_085807_(_009976_, _010086_, _010097_);
  or g_085808_(_009965_, _010075_, _010108_);
  and g_085809_(_009954_, _010097_, _010119_);
  or g_085810_(_009943_, _010108_, _010130_);
  and g_085811_(_009921_, _010119_, _010141_);
  or g_085812_(_009932_, _010130_, _010152_);
  and g_085813_(_009679_, _010141_, _010163_);
  or g_085814_(_009690_, _010152_, _010174_);
  xor g_085815_(out[54], _005026_, _010185_);
  xor g_085816_(_002716_, _005026_, _010196_);
  and g_085817_(_007314_, _009404_, _010207_);
  or g_085818_(_007303_, _009393_, _010218_);
  and g_085819_(_007248_, _009393_, _010229_);
  or g_085820_(_007237_, _009404_, _010240_);
  and g_085821_(_010218_, _010240_, _010251_);
  or g_085822_(_010207_, _010229_, _010262_);
  and g_085823_(_010196_, _010251_, _010273_);
  or g_085824_(_010185_, _010262_, _010284_);
  and g_085825_(_009998_, _010064_, _010295_);
  or g_085826_(_009987_, _010053_, _010306_);
  and g_085827_(_010284_, _010306_, _010317_);
  or g_085828_(_010273_, _010295_, _010328_);
  and g_085829_(_010185_, _010262_, _010339_);
  or g_085830_(_010196_, _010251_, _010350_);
  and g_085831_(_010317_, _010350_, _010361_);
  or g_085832_(_010328_, _010339_, _010372_);
  xor g_085833_(out[53], _005015_, _010383_);
  xor g_085834_(_002727_, _005015_, _010394_);
  and g_085835_(_007435_, _009404_, _010405_);
  or g_085836_(_007446_, _009393_, _010416_);
  and g_085837_(_007380_, _009393_, _010427_);
  or g_085838_(_007369_, _009404_, _010438_);
  and g_085839_(_010416_, _010438_, _010449_);
  or g_085840_(_010405_, _010427_, _010460_);
  and g_085841_(_010383_, _010460_, _010471_);
  or g_085842_(_010394_, _010449_, _010482_);
  xor g_085843_(out[52], _005004_, _010493_);
  xor g_085844_(_002738_, _005004_, _010504_);
  and g_085845_(_007479_, _009393_, _010515_);
  or g_085846_(_007490_, _009404_, _010526_);
  and g_085847_(_007556_, _009404_, _010537_);
  or g_085848_(_007545_, _009393_, _010548_);
  and g_085849_(_010526_, _010548_, _010559_);
  or g_085850_(_010515_, _010537_, _010570_);
  and g_085851_(_010504_, _010570_, _010581_);
  or g_085852_(_010493_, _010559_, _010592_);
  and g_085853_(_010482_, _010592_, _010603_);
  or g_085854_(_010471_, _010581_, _010614_);
  and g_085855_(_010493_, _010559_, _010625_);
  or g_085856_(_010504_, _010570_, _010636_);
  and g_085857_(_010394_, _010449_, _010647_);
  or g_085858_(_010383_, _010460_, _010658_);
  and g_085859_(_010636_, _010658_, _010669_);
  or g_085860_(_010625_, _010647_, _010680_);
  and g_085861_(_010603_, _010669_, _010691_);
  or g_085862_(_010614_, _010680_, _010702_);
  and g_085863_(_010361_, _010691_, _010713_);
  or g_085864_(_010372_, _010702_, _010724_);
  and g_085865_(_010163_, _010713_, _010735_);
  or g_085866_(_010174_, _010724_, _010746_);
  xor g_085867_(out[51], _004982_, _010757_);
  xor g_085868_(_002782_, _004982_, _010768_);
  or g_085869_(_007776_, _009393_, _010779_);
  or g_085870_(_007699_, _009404_, _010790_);
  and g_085871_(_010779_, _010790_, _010801_);
  or g_085872_(_010768_, _010801_, _010812_);
  or g_085873_(out[49], out[50], _010823_);
  xor g_085874_(out[49], out[50], _010834_);
  xor g_085875_(_002749_, out[50], _010845_);
  or g_085876_(_007908_, _009393_, _010856_);
  or g_085877_(_007842_, _009404_, _010867_);
  and g_085878_(_010856_, _010867_, _010878_);
  not g_085879_(_010878_, _010889_);
  and g_085880_(_010768_, _010801_, _010900_);
  or g_085881_(_010834_, _010889_, _010911_);
  xor g_085882_(_010845_, _010878_, _010922_);
  xor g_085883_(_010834_, _010878_, _010933_);
  xor g_085884_(_010768_, _010801_, _010944_);
  xor g_085885_(_010757_, _010801_, _010955_);
  and g_085886_(_010922_, _010944_, _010966_);
  or g_085887_(_010933_, _010955_, _010977_);
  or g_085888_(_002617_, _009404_, _010988_);
  or g_085889_(_008084_, _009393_, _010999_);
  and g_085890_(_010988_, _010999_, _011010_);
  and g_085891_(out[49], _011010_, _011021_);
  not g_085892_(_011021_, _011032_);
  and g_085893_(_008194_, _009404_, _011043_);
  or g_085894_(_008183_, _009393_, _011054_);
  and g_085895_(_002628_, _009393_, _011065_);
  or g_085896_(out[32], _009404_, _011076_);
  and g_085897_(_011054_, _011076_, _011087_);
  or g_085898_(_011043_, _011065_, _011098_);
  and g_085899_(out[48], _011098_, _011109_);
  or g_085900_(_002760_, _011087_, _011120_);
  xor g_085901_(out[49], _011010_, _011131_);
  xor g_085902_(_002749_, _011010_, _011142_);
  and g_085903_(_011120_, _011131_, _011153_);
  or g_085904_(_011109_, _011142_, _011164_);
  and g_085905_(_011032_, _011164_, _011175_);
  or g_085906_(_011021_, _011153_, _011186_);
  and g_085907_(_010966_, _011186_, _011197_);
  or g_085908_(_010977_, _011175_, _011208_);
  or g_085909_(_010900_, _010911_, _011219_);
  and g_085910_(_010812_, _011219_, _011230_);
  not g_085911_(_011230_, _011241_);
  and g_085912_(_011208_, _011230_, _011252_);
  or g_085913_(_011197_, _011241_, _011263_);
  and g_085914_(_010735_, _011263_, _011274_);
  or g_085915_(_010746_, _011252_, _011285_);
  and g_085916_(_010482_, _010636_, _011296_);
  or g_085917_(_010471_, _010625_, _011307_);
  and g_085918_(_010658_, _011307_, _011318_);
  or g_085919_(_010647_, _011296_, _011329_);
  and g_085920_(_010361_, _011318_, _011340_);
  or g_085921_(_010372_, _011329_, _011351_);
  and g_085922_(_010317_, _011351_, _011362_);
  or g_085923_(_010328_, _011340_, _011373_);
  and g_085924_(_010163_, _011373_, _011384_);
  or g_085925_(_010174_, _011362_, _011395_);
  and g_085926_(_009932_, _009954_, _011406_);
  or g_085927_(_009921_, _009943_, _011417_);
  and g_085928_(_009679_, _011406_, _011428_);
  or g_085929_(_009690_, _011417_, _011439_);
  and g_085930_(_009602_, _009646_, _011450_);
  not g_085931_(_011450_, _011461_);
  and g_085932_(_011439_, _011461_, _011472_);
  or g_085933_(_011428_, _011450_, _011483_);
  and g_085934_(_011395_, _011472_, _011494_);
  or g_085935_(_011384_, _011483_, _011505_);
  and g_085936_(_011285_, _011494_, _011516_);
  or g_085937_(_011274_, _011505_, _011527_);
  and g_085938_(_002760_, _011087_, _011538_);
  or g_085939_(_010977_, _011538_, _011549_);
  not g_085940_(_011549_, _011560_);
  and g_085941_(_011153_, _011560_, _011571_);
  not g_085942_(_011571_, _011582_);
  and g_085943_(_010735_, _011571_, _011593_);
  or g_085944_(_010746_, _011582_, _011604_);
  and g_085945_(_011527_, _011604_, _011615_);
  or g_085946_(_011516_, _011593_, _011626_);
  and g_085947_(_005103_, _011615_, _011637_);
  or g_085948_(_005092_, _011626_, _011648_);
  and g_085949_(_009558_, _011626_, _011659_);
  or g_085950_(_009547_, _011615_, _011670_);
  and g_085951_(_011648_, _011670_, _011681_);
  or g_085952_(_011637_, _011659_, _011692_);
  and g_085953_(_004960_, _011681_, _011703_);
  or g_085954_(_004971_, _011692_, _011714_);
  and g_085955_(out[81], out[82], _011725_);
  or g_085956_(out[84], out[83], _011736_);
  or g_085957_(out[83], _011725_, _011747_);
  or g_085958_(_011725_, _011736_, _011758_);
  or g_085959_(out[85], _011758_, _011769_);
  and g_085960_(out[86], _011769_, _011780_);
  and g_085961_(out[87], _011780_, _011791_);
  or g_085962_(out[88], _011791_, _011802_);
  or g_085963_(out[89], _011802_, _011813_);
  or g_085964_(out[90], _011813_, _011824_);
  xor g_085965_(_002958_, _011824_, _011835_);
  xor g_085966_(out[91], _011824_, _011846_);
  and g_085967_(_011703_, _011835_, _011857_);
  or g_085968_(_011714_, _011846_, _011868_);
  and g_085969_(out[97], out[98], _011879_);
  or g_085970_(out[100], out[99], _011890_);
  or g_085971_(out[99], _011879_, _011901_);
  or g_085972_(_011879_, _011890_, _011912_);
  or g_085973_(out[101], _011912_, _011923_);
  and g_085974_(out[102], _011923_, _011934_);
  and g_085975_(out[103], _011934_, _011945_);
  or g_085976_(out[104], _011945_, _011956_);
  or g_085977_(out[105], _011956_, _011967_);
  or g_085978_(out[106], _011967_, _011978_);
  xor g_085979_(out[107], _011978_, _011989_);
  not g_085980_(_011989_, _012000_);
  and g_085981_(_011857_, _012000_, _012011_);
  or g_085982_(_011868_, _011989_, _012022_);
  and g_085983_(out[113], out[114], _012033_);
  or g_085984_(out[116], out[115], _012044_);
  or g_085985_(out[115], _012033_, _012055_);
  or g_085986_(_012033_, _012044_, _012066_);
  or g_085987_(out[117], _012066_, _012077_);
  and g_085988_(out[118], _012077_, _012088_);
  and g_085989_(out[119], _012088_, _012099_);
  or g_085990_(out[120], _012099_, _012110_);
  or g_085991_(out[121], _012110_, _012121_);
  or g_085992_(out[122], _012121_, _012132_);
  xor g_085993_(_003222_, _012132_, _012143_);
  xor g_085994_(out[123], _012132_, _012154_);
  and g_085995_(_012011_, _012143_, _012165_);
  or g_085996_(_012022_, _012154_, _012176_);
  and g_085997_(out[129], out[130], _012187_);
  or g_085998_(out[132], out[131], _012198_);
  or g_085999_(out[131], _012187_, _012209_);
  or g_086000_(_012187_, _012198_, _012220_);
  or g_086001_(out[133], _012220_, _012231_);
  and g_086002_(out[134], _012231_, _012242_);
  and g_086003_(out[135], _012242_, _012253_);
  or g_086004_(out[136], _012253_, _012264_);
  or g_086005_(out[137], _012264_, _012275_);
  or g_086006_(out[138], _012275_, _012286_);
  xor g_086007_(_003354_, _012286_, _012297_);
  xor g_086008_(out[139], _012286_, _012308_);
  and g_086009_(_012165_, _012297_, _012319_);
  or g_086010_(_012176_, _012308_, _012330_);
  and g_086011_(out[145], out[146], _012341_);
  or g_086012_(out[148], out[147], _012352_);
  or g_086013_(out[147], _012341_, _012363_);
  or g_086014_(_012341_, _012352_, _012374_);
  or g_086015_(out[149], _012374_, _012385_);
  and g_086016_(out[150], _012385_, _012396_);
  and g_086017_(out[151], _012396_, _012407_);
  or g_086018_(out[152], _012407_, _012418_);
  or g_086019_(out[153], _012418_, _012429_);
  or g_086020_(out[154], _012429_, _012440_);
  xor g_086021_(_003486_, _012440_, _012451_);
  xor g_086022_(out[155], _012440_, _012462_);
  and g_086023_(_012319_, _012451_, _012473_);
  or g_086024_(_012330_, _012462_, _012484_);
  and g_086025_(out[161], out[162], _012495_);
  or g_086026_(out[164], out[163], _012506_);
  or g_086027_(out[163], _012495_, _012517_);
  or g_086028_(_012495_, _012506_, _012528_);
  or g_086029_(out[165], _012528_, _012539_);
  and g_086030_(out[166], _012539_, _012550_);
  and g_086031_(out[167], _012550_, _012561_);
  or g_086032_(out[168], _012561_, _012572_);
  or g_086033_(out[169], _012572_, _012583_);
  or g_086034_(out[170], _012583_, _012594_);
  xor g_086035_(out[171], _012594_, _012605_);
  not g_086036_(_012605_, _012616_);
  and g_086037_(_012473_, _012616_, _012627_);
  or g_086038_(_012484_, _012605_, _012638_);
  and g_086039_(out[177], out[178], _012649_);
  or g_086040_(out[180], out[179], _012660_);
  or g_086041_(out[179], _012649_, _012671_);
  or g_086042_(_012649_, _012660_, _012682_);
  or g_086043_(out[181], _012682_, _012693_);
  and g_086044_(out[182], _012693_, _012704_);
  and g_086045_(out[183], _012704_, _012715_);
  or g_086046_(out[184], _012715_, _012726_);
  or g_086047_(out[185], _012726_, _012737_);
  or g_086048_(out[186], _012737_, _012748_);
  xor g_086049_(_003750_, _012748_, _012759_);
  xor g_086050_(out[187], _012748_, _012770_);
  and g_086051_(_012627_, _012759_, _012781_);
  or g_086052_(_012638_, _012770_, _012792_);
  and g_086053_(out[193], out[194], _012803_);
  or g_086054_(out[196], out[195], _012814_);
  or g_086055_(out[195], _012803_, _012825_);
  or g_086056_(_012803_, _012814_, _012836_);
  or g_086057_(out[197], _012836_, _012847_);
  and g_086058_(out[198], _012847_, _012858_);
  and g_086059_(out[199], _012858_, _012869_);
  or g_086060_(out[200], _012869_, _012880_);
  or g_086061_(out[201], _012880_, _012891_);
  not g_086062_(_012891_, _012902_);
  or g_086063_(out[202], _012891_, _012913_);
  xor g_086064_(_003882_, _012913_, _012924_);
  xor g_086065_(out[203], _012913_, _012935_);
  and g_086066_(_012781_, _012924_, _012946_);
  or g_086067_(_012792_, _012935_, _012957_);
  and g_086068_(out[209], out[210], _012968_);
  or g_086069_(out[212], out[211], _012979_);
  or g_086070_(out[211], _012968_, _012990_);
  or g_086071_(_012968_, _012979_, _013001_);
  or g_086072_(out[213], _013001_, _013012_);
  and g_086073_(out[214], _013012_, _013023_);
  and g_086074_(out[215], _013023_, _013034_);
  or g_086075_(out[216], _013034_, _013045_);
  or g_086076_(out[217], _013045_, _013056_);
  or g_086077_(out[218], _013056_, _013067_);
  xor g_086078_(_003992_, _013067_, _013078_);
  xor g_086079_(out[219], _013067_, _013089_);
  and g_086080_(_012946_, _013078_, _013100_);
  or g_086081_(_012957_, _013089_, _013111_);
  and g_086082_(out[225], out[226], _013122_);
  or g_086083_(out[228], out[227], _013133_);
  or g_086084_(out[227], _013122_, _013144_);
  or g_086085_(_013122_, _013133_, _013155_);
  or g_086086_(out[229], _013155_, _013166_);
  and g_086087_(out[230], _013166_, _013177_);
  and g_086088_(out[231], _013177_, _013188_);
  or g_086089_(out[232], _013188_, _013199_);
  or g_086090_(out[233], _013199_, _013210_);
  or g_086091_(out[234], _013210_, _013221_);
  xor g_086092_(_004124_, _013221_, _013232_);
  xor g_086093_(out[235], _013221_, _013243_);
  and g_086094_(_013100_, _013232_, _013254_);
  or g_086095_(_013111_, _013243_, _013265_);
  and g_086096_(out[241], out[242], _013276_);
  or g_086097_(out[243], _013276_, _013287_);
  or g_086098_(out[244], _013287_, _013298_);
  or g_086099_(out[245], _013298_, _013309_);
  and g_086100_(out[246], _013309_, _013320_);
  and g_086101_(out[247], _013320_, _013331_);
  or g_086102_(out[248], _013331_, _013342_);
  or g_086103_(out[249], _013342_, _013353_);
  or g_086104_(out[250], _013353_, _013364_);
  xor g_086105_(_004245_, _013364_, _013375_);
  xor g_086106_(out[251], _013364_, _013386_);
  and g_086107_(_013254_, _013375_, _013397_);
  or g_086108_(_013265_, _013386_, _013408_);
  and g_086109_(out[258], out[257], _013419_);
  not g_086110_(_013419_, _013430_);
  or g_086111_(out[259], _013419_, _013441_);
  or g_086112_(out[260], _013441_, _013452_);
  or g_086113_(out[261], _013452_, _013463_);
  and g_086114_(out[262], _013463_, _013474_);
  and g_086115_(out[263], _013474_, _013485_);
  or g_086116_(out[264], _013485_, _013496_);
  or g_086117_(out[265], _013496_, _013507_);
  or g_086118_(out[266], _013507_, _013518_);
  xor g_086119_(out[267], _013518_, _013529_);
  not g_086120_(_013529_, _013540_);
  and g_086121_(_013397_, _013540_, _013551_);
  or g_086122_(_013408_, _013529_, _013562_);
  and g_086123_(out[274], out[273], _013573_);
  or g_086124_(out[275], out[276], _013584_);
  or g_086125_(out[275], _013573_, _013595_);
  or g_086126_(_013573_, _013584_, _013606_);
  or g_086127_(out[277], _013606_, _013617_);
  and g_086128_(out[278], _013617_, _013628_);
  and g_086129_(out[279], _013628_, _013639_);
  or g_086130_(out[280], _013639_, _013650_);
  or g_086131_(out[281], _013650_, _013661_);
  or g_086132_(out[282], _013661_, _013672_);
  xor g_086133_(_004432_, _013672_, _013683_);
  xor g_086134_(out[283], _013672_, _013694_);
  and g_086135_(_013551_, _013683_, _013705_);
  or g_086136_(_013562_, _013694_, _013716_);
  and g_086137_(out[290], out[289], _013727_);
  or g_086138_(out[291], out[292], _013738_);
  or g_086139_(out[291], _013727_, _013749_);
  or g_086140_(_013727_, _013738_, _013760_);
  or g_086141_(out[293], _013760_, _013771_);
  and g_086142_(out[294], _013771_, _013782_);
  and g_086143_(out[295], _013782_, _013793_);
  or g_086144_(out[296], _013793_, _013804_);
  or g_086145_(out[297], _013804_, _013815_);
  or g_086146_(out[298], _013815_, _013826_);
  xor g_086147_(_004465_, _013826_, _013837_);
  xor g_086148_(out[299], _013826_, _013848_);
  and g_086149_(_013705_, _013837_, _013859_);
  or g_086150_(_013716_, _013848_, _013870_);
  and g_086151_(out[306], out[305], _013881_);
  not g_086152_(_013881_, _013892_);
  or g_086153_(out[307], _013881_, _013903_);
  or g_086154_(out[308], _013903_, _013914_);
  or g_086155_(out[309], _013914_, _013925_);
  and g_086156_(out[310], _013925_, _013936_);
  and g_086157_(out[311], _013936_, _013947_);
  or g_086158_(out[312], _013947_, _013958_);
  or g_086159_(out[313], _013958_, _013969_);
  or g_086160_(out[314], _013969_, _013980_);
  xor g_086161_(_004498_, _013980_, _013991_);
  xor g_086162_(out[315], _013980_, _014002_);
  and g_086163_(_013859_, _013991_, _014013_);
  or g_086164_(_013870_, _014002_, _014024_);
  and g_086165_(out[322], out[321], _014035_);
  or g_086166_(out[323], out[324], _014046_);
  or g_086167_(out[323], _014035_, _014057_);
  or g_086168_(_014035_, _014046_, _014068_);
  or g_086169_(out[325], _014068_, _014079_);
  and g_086170_(out[326], _014079_, _014090_);
  and g_086171_(out[327], _014090_, _014101_);
  or g_086172_(out[328], _014101_, _014112_);
  or g_086173_(out[329], _014112_, _014123_);
  or g_086174_(out[330], _014123_, _014134_);
  xor g_086175_(_004531_, _014134_, _014145_);
  xor g_086176_(out[331], _014134_, _014156_);
  and g_086177_(_014013_, _014145_, _014167_);
  or g_086178_(_014024_, _014156_, _014178_);
  and g_086179_(out[338], out[337], _014189_);
  or g_086180_(out[339], out[340], _014200_);
  or g_086181_(out[339], _014189_, _014211_);
  or g_086182_(_014189_, _014200_, _014222_);
  or g_086183_(out[341], _014222_, _014233_);
  and g_086184_(out[342], _014233_, _014244_);
  and g_086185_(out[343], _014244_, _014255_);
  or g_086186_(out[344], _014255_, _014266_);
  or g_086187_(out[345], _014266_, _014277_);
  or g_086188_(out[346], _014277_, _014288_);
  xor g_086189_(_004564_, _014288_, _014299_);
  xor g_086190_(out[347], _014288_, _014310_);
  and g_086191_(_014167_, _014299_, _014321_);
  or g_086192_(_014178_, _014310_, _014332_);
  and g_086193_(out[354], out[353], _014343_);
  or g_086194_(out[355], out[356], _014354_);
  or g_086195_(out[355], _014343_, _014365_);
  or g_086196_(_014343_, _014354_, _014376_);
  or g_086197_(out[357], _014376_, _014387_);
  and g_086198_(out[358], _014387_, _014398_);
  and g_086199_(out[359], _014398_, _014409_);
  or g_086200_(out[360], _014409_, _014420_);
  or g_086201_(out[361], _014420_, _014431_);
  or g_086202_(out[362], _014431_, _014442_);
  xor g_086203_(_004597_, _014442_, _014453_);
  xor g_086204_(out[363], _014442_, _014464_);
  and g_086205_(_014321_, _014453_, _014475_);
  or g_086206_(_014332_, _014464_, _014486_);
  and g_086207_(out[370], out[369], _014497_);
  or g_086208_(out[371], out[372], _014508_);
  or g_086209_(out[371], _014497_, _014519_);
  or g_086210_(_014497_, _014508_, _014530_);
  or g_086211_(out[373], _014530_, _014541_);
  and g_086212_(out[374], _014541_, _014552_);
  and g_086213_(out[375], _014552_, _014563_);
  or g_086214_(out[376], _014563_, _014574_);
  or g_086215_(out[377], _014574_, _014585_);
  or g_086216_(out[378], _014585_, _014596_);
  xor g_086217_(_004630_, _014596_, _014607_);
  xor g_086218_(out[379], _014596_, _014618_);
  and g_086219_(_014475_, _014607_, _014629_);
  or g_086220_(_014486_, _014618_, _014640_);
  and g_086221_(out[386], out[385], _014651_);
  or g_086222_(out[387], out[388], _014662_);
  or g_086223_(out[387], _014651_, _014673_);
  or g_086224_(_014651_, _014662_, _014684_);
  or g_086225_(out[389], _014684_, _014695_);
  and g_086226_(out[390], _014695_, _014706_);
  and g_086227_(out[391], _014706_, _014717_);
  or g_086228_(out[392], _014717_, _014728_);
  or g_086229_(out[393], _014728_, _014739_);
  or g_086230_(out[394], _014739_, _014750_);
  xor g_086231_(_004663_, _014750_, _014761_);
  xor g_086232_(out[395], _014750_, _014772_);
  and g_086233_(_014629_, _014761_, _014783_);
  or g_086234_(_014640_, _014772_, _014794_);
  and g_086235_(out[402], out[401], _014805_);
  or g_086236_(out[403], out[404], _014816_);
  or g_086237_(out[403], _014805_, _014827_);
  or g_086238_(_014805_, _014816_, _014838_);
  or g_086239_(out[405], _014838_, _014849_);
  and g_086240_(out[406], _014849_, _014860_);
  and g_086241_(out[407], _014860_, _014871_);
  or g_086242_(out[408], _014871_, _014882_);
  or g_086243_(out[409], _014882_, _014893_);
  or g_086244_(out[410], _014893_, _014904_);
  xor g_086245_(_004696_, _014904_, _014915_);
  xor g_086246_(out[411], _014904_, _014926_);
  and g_086247_(_014783_, _014915_, _014937_);
  or g_086248_(_014794_, _014926_, _014948_);
  and g_086249_(out[418], out[417], _014959_);
  or g_086250_(out[419], out[420], _014970_);
  or g_086251_(out[419], _014959_, _014981_);
  or g_086252_(_014959_, _014970_, _014992_);
  or g_086253_(out[421], _014992_, _015003_);
  and g_086254_(out[422], _015003_, _015014_);
  and g_086255_(out[423], _015014_, _015025_);
  or g_086256_(out[424], _015025_, _015036_);
  or g_086257_(out[425], _015036_, _015047_);
  or g_086258_(out[426], _015047_, _015058_);
  xor g_086259_(_004729_, _015058_, _015069_);
  xor g_086260_(out[427], _015058_, _015080_);
  and g_086261_(_014937_, _015069_, _015091_);
  or g_086262_(_014948_, _015080_, _015102_);
  and g_086263_(out[434], out[433], _015113_);
  or g_086264_(out[435], out[436], _015124_);
  or g_086265_(out[435], _015113_, _015135_);
  or g_086266_(_015113_, _015124_, _015146_);
  or g_086267_(out[437], _015146_, _015157_);
  and g_086268_(out[438], _015157_, _015168_);
  and g_086269_(out[439], _015168_, _015179_);
  or g_086270_(out[440], _015179_, _015190_);
  or g_086271_(out[441], _015190_, _015201_);
  or g_086272_(out[442], _015201_, _015212_);
  xor g_086273_(_004762_, _015212_, _015223_);
  xor g_086274_(out[443], _015212_, _015234_);
  or g_086275_(_015102_, _015234_, _015245_);
  not g_086276_(_015245_, _015256_);
  and g_086277_(out[450], out[449], _015267_);
  or g_086278_(out[451], out[452], _015278_);
  or g_086279_(out[451], _015267_, _015289_);
  or g_086280_(_015267_, _015278_, _015300_);
  or g_086281_(out[453], _015300_, _015311_);
  and g_086282_(out[454], _015311_, _015322_);
  and g_086283_(out[455], _015322_, _015333_);
  or g_086284_(out[456], _015333_, _015344_);
  or g_086285_(out[457], _015344_, _015355_);
  or g_086286_(out[458], _015355_, _015366_);
  xor g_086287_(out[459], _015366_, _015377_);
  not g_086288_(_015377_, _015388_);
  or g_086289_(_015245_, _015377_, _015399_);
  not g_086290_(_015399_, _015410_);
  and g_086291_(out[466], out[465], _015421_);
  or g_086292_(out[467], out[468], _015432_);
  or g_086293_(out[467], _015421_, _015443_);
  or g_086294_(_015421_, _015432_, _015454_);
  or g_086295_(out[469], _015454_, _015465_);
  and g_086296_(out[470], _015465_, _015476_);
  and g_086297_(out[471], _015476_, _015487_);
  or g_086298_(out[472], _015487_, _015498_);
  or g_086299_(out[473], _015498_, _015509_);
  or g_086300_(out[474], _015509_, _015520_);
  xor g_086301_(out[475], _015520_, _015531_);
  not g_086302_(_015531_, _015542_);
  or g_086303_(_015399_, _015531_, _015553_);
  and g_086304_(out[545], out[546], _015564_);
  or g_086305_(out[548], out[547], _015575_);
  or g_086306_(out[547], _015564_, _015586_);
  or g_086307_(_015564_, _015575_, _015597_);
  or g_086308_(out[549], _015597_, _015608_);
  and g_086309_(out[550], _015608_, _015619_);
  and g_086310_(out[551], _015619_, _015630_);
  or g_086311_(out[552], _015630_, _015641_);
  or g_086312_(out[553], _015641_, _015652_);
  or g_086313_(out[554], _015652_, _015663_);
  xor g_086314_(out[555], _015663_, _015674_);
  not g_086315_(_015674_, _015685_);
  and g_086316_(out[529], out[530], _015696_);
  or g_086317_(out[532], out[531], _015707_);
  or g_086318_(out[531], _015696_, _015718_);
  or g_086319_(_015696_, _015707_, _015729_);
  or g_086320_(out[533], _015729_, _015740_);
  and g_086321_(out[534], _015740_, _015751_);
  and g_086322_(out[535], _015751_, _015762_);
  or g_086323_(out[536], _015762_, _015773_);
  or g_086324_(out[537], _015773_, _015784_);
  or g_086325_(out[538], _015784_, _015795_);
  xor g_086326_(_054743_, _015795_, _015806_);
  xor g_086327_(out[539], _015795_, _015817_);
  and g_086328_(out[513], out[514], _015828_);
  or g_086329_(out[516], out[515], _015839_);
  or g_086330_(out[515], _015828_, _015850_);
  or g_086331_(_015828_, _015839_, _015861_);
  or g_086332_(out[517], _015861_, _015872_);
  and g_086333_(out[518], _015872_, _015883_);
  and g_086334_(out[519], _015883_, _015894_);
  or g_086335_(out[520], _015894_, _015905_);
  or g_086336_(out[521], _015905_, _015916_);
  or g_086337_(out[522], _015916_, _015927_);
  xor g_086338_(_054611_, _015927_, _015938_);
  xor g_086339_(out[523], _015927_, _015949_);
  and g_086340_(out[497], out[498], _015960_);
  or g_086341_(out[500], out[499], _015971_);
  or g_086342_(out[499], _015960_, _015982_);
  or g_086343_(_015960_, _015971_, _015993_);
  or g_086344_(out[501], _015993_, _016004_);
  and g_086345_(out[502], _016004_, _016015_);
  and g_086346_(out[503], _016015_, _016026_);
  or g_086347_(out[504], _016026_, _016037_);
  or g_086348_(out[505], _016037_, _016048_);
  or g_086349_(out[506], _016048_, _016059_);
  xor g_086350_(_054479_, _016059_, _016070_);
  xor g_086351_(out[507], _016059_, _016081_);
  and g_086352_(out[481], out[482], _016092_);
  or g_086353_(out[484], out[483], _016103_);
  or g_086354_(out[483], _016092_, _016114_);
  or g_086355_(_016092_, _016103_, _016125_);
  or g_086356_(out[485], _016125_, _016136_);
  and g_086357_(out[486], _016136_, _016147_);
  and g_086358_(out[487], _016147_, _016158_);
  or g_086359_(out[488], _016158_, _016169_);
  or g_086360_(out[489], _016169_, _016180_);
  or g_086361_(out[490], _016180_, _016191_);
  xor g_086362_(_054358_, _016191_, _016202_);
  xor g_086363_(out[491], _016191_, _016213_);
  xor g_086364_(out[486], _016136_, _016224_);
  not g_086365_(_016224_, _016235_);
  xor g_086366_(out[502], _016004_, _016246_);
  not g_086367_(_016246_, _016257_);
  and g_086368_(_016224_, _016257_, _016268_);
  or g_086369_(_016235_, _016246_, _016279_);
  xor g_086370_(out[483], _016092_, _016290_);
  xor g_086371_(_054435_, _016092_, _016301_);
  xor g_086372_(out[499], _015960_, _016312_);
  xor g_086373_(_054567_, _015960_, _016323_);
  and g_086374_(_016301_, _016312_, _016334_);
  or g_086375_(_016290_, _016323_, _016345_);
  or g_086376_(out[497], out[498], _016356_);
  xor g_086377_(out[497], out[498], _016367_);
  xor g_086378_(_054534_, out[498], _016378_);
  or g_086379_(out[481], out[482], _016389_);
  xor g_086380_(out[481], out[482], _016400_);
  xor g_086381_(_054413_, out[482], _016411_);
  and g_086382_(_016378_, _016400_, _016422_);
  or g_086383_(_016367_, _016411_, _016433_);
  and g_086384_(_016367_, _016411_, _016444_);
  or g_086385_(_016378_, _016400_, _016455_);
  and g_086386_(_016290_, _016323_, _016466_);
  or g_086387_(_016301_, _016312_, _016477_);
  and g_086388_(_016433_, _016477_, _016488_);
  or g_086389_(_016422_, _016466_, _016499_);
  and g_086390_(_016345_, _016455_, _016510_);
  or g_086391_(_016334_, _016444_, _016521_);
  and g_086392_(_016488_, _016510_, _016532_);
  or g_086393_(_016499_, _016521_, _016543_);
  and g_086394_(_054413_, out[497], _016554_);
  or g_086395_(out[481], _054534_, _016565_);
  and g_086396_(_054347_, out[496], _016576_);
  or g_086397_(out[480], _054545_, _016587_);
  and g_086398_(out[481], _054534_, _016598_);
  or g_086399_(_054413_, out[497], _016609_);
  and g_086400_(_016587_, _016609_, _016620_);
  or g_086401_(_016576_, _016598_, _016631_);
  and g_086402_(_016565_, _016620_, _016642_);
  or g_086403_(_016554_, _016631_, _016653_);
  and g_086404_(_016565_, _016653_, _016664_);
  or g_086405_(_016554_, _016642_, _016675_);
  and g_086406_(_016532_, _016675_, _016686_);
  or g_086407_(_016543_, _016664_, _016697_);
  and g_086408_(_016422_, _016477_, _016708_);
  or g_086409_(_016433_, _016466_, _016719_);
  or g_086410_(_016334_, _016708_, _016730_);
  and g_086411_(_016345_, _016719_, _016741_);
  and g_086412_(_016697_, _016741_, _016752_);
  or g_086413_(_016686_, _016730_, _016763_);
  xor g_086414_(out[484], _016114_, _016774_);
  xor g_086415_(_054402_, _016114_, _016785_);
  xor g_086416_(out[500], _015982_, _016796_);
  xor g_086417_(_054523_, _015982_, _016807_);
  and g_086418_(_016774_, _016807_, _016818_);
  or g_086419_(_016785_, _016796_, _016829_);
  and g_086420_(out[480], _054545_, _016840_);
  or g_086421_(_054347_, out[496], _016851_);
  and g_086422_(_016642_, _016851_, _016862_);
  or g_086423_(_016653_, _016840_, _016873_);
  and g_086424_(_016532_, _016862_, _016884_);
  or g_086425_(_016543_, _016873_, _016895_);
  and g_086426_(_016829_, _016895_, _016906_);
  or g_086427_(_016818_, _016884_, _016917_);
  and g_086428_(_016763_, _016906_, _016928_);
  or g_086429_(_016752_, _016917_, _016939_);
  xor g_086430_(out[485], _016125_, _016950_);
  xor g_086431_(_054391_, _016125_, _016961_);
  xor g_086432_(out[501], _015993_, _016972_);
  xor g_086433_(_054512_, _015993_, _016983_);
  and g_086434_(_016961_, _016972_, _016994_);
  or g_086435_(_016950_, _016983_, _017005_);
  and g_086436_(_016785_, _016796_, _017016_);
  or g_086437_(_016774_, _016807_, _017027_);
  and g_086438_(_017005_, _017027_, _017038_);
  or g_086439_(_016994_, _017016_, _017049_);
  and g_086440_(_016939_, _017038_, _017060_);
  or g_086441_(_016928_, _017049_, _017071_);
  and g_086442_(_016950_, _016983_, _017082_);
  or g_086443_(_016961_, _016972_, _017093_);
  xor g_086444_(out[487], _016147_, _017104_);
  not g_086445_(_017104_, _017115_);
  xor g_086446_(out[503], _016015_, _017126_);
  not g_086447_(_017126_, _017137_);
  and g_086448_(_017115_, _017126_, _017148_);
  or g_086449_(_017104_, _017137_, _017159_);
  and g_086450_(_016235_, _016246_, _017170_);
  or g_086451_(_016224_, _016257_, _017181_);
  and g_086452_(_017093_, _017181_, _017192_);
  or g_086453_(_017082_, _017170_, _017203_);
  and g_086454_(_017071_, _017192_, _017214_);
  or g_086455_(_017060_, _017203_, _017225_);
  and g_086456_(_016279_, _017225_, _017236_);
  or g_086457_(_016268_, _017214_, _017247_);
  and g_086458_(_017159_, _017247_, _017258_);
  or g_086459_(_017148_, _017236_, _017269_);
  and g_086460_(_017104_, _017137_, _017280_);
  or g_086461_(_017115_, _017126_, _017291_);
  xor g_086462_(out[488], _016158_, _017302_);
  xor g_086463_(_054446_, _016158_, _017313_);
  xor g_086464_(out[504], _016026_, _017324_);
  xor g_086465_(_054578_, _016026_, _017335_);
  and g_086466_(_017313_, _017324_, _017346_);
  or g_086467_(_017302_, _017335_, _017357_);
  and g_086468_(_017291_, _017357_, _017368_);
  or g_086469_(_017280_, _017346_, _017379_);
  and g_086470_(_017269_, _017368_, _017390_);
  or g_086471_(_017258_, _017379_, _017401_);
  and g_086472_(_017302_, _017335_, _017412_);
  or g_086473_(_017313_, _017324_, _017423_);
  xor g_086474_(out[505], _016037_, _017434_);
  xor g_086475_(_054589_, _016037_, _017445_);
  xor g_086476_(out[489], _016169_, _017456_);
  xor g_086477_(_054457_, _016169_, _017467_);
  and g_086478_(_017445_, _017456_, _017478_);
  or g_086479_(_017434_, _017467_, _017489_);
  and g_086480_(_017423_, _017489_, _017500_);
  or g_086481_(_017412_, _017478_, _017511_);
  and g_086482_(_017401_, _017500_, _017522_);
  or g_086483_(_017390_, _017511_, _017533_);
  xor g_086484_(out[490], _016180_, _017544_);
  xor g_086485_(_054468_, _016180_, _017555_);
  xor g_086486_(out[506], _016048_, _017566_);
  xor g_086487_(_054600_, _016048_, _017577_);
  and g_086488_(_017555_, _017566_, _017588_);
  or g_086489_(_017544_, _017577_, _017599_);
  and g_086490_(_017434_, _017467_, _017610_);
  or g_086491_(_017445_, _017456_, _017621_);
  and g_086492_(_017599_, _017621_, _017632_);
  or g_086493_(_017588_, _017610_, _017643_);
  and g_086494_(_017533_, _017632_, _017654_);
  or g_086495_(_017522_, _017643_, _017665_);
  and g_086496_(_016070_, _016213_, _017676_);
  or g_086497_(_016081_, _016202_, _017687_);
  and g_086498_(_017544_, _017577_, _017698_);
  or g_086499_(_017555_, _017566_, _017709_);
  and g_086500_(_017687_, _017709_, _017720_);
  or g_086501_(_017676_, _017698_, _017731_);
  and g_086502_(_017665_, _017720_, _017742_);
  or g_086503_(_017654_, _017731_, _017753_);
  and g_086504_(_016070_, _016202_, _017764_);
  or g_086505_(_016081_, _016213_, _017775_);
  and g_086506_(_015949_, _017764_, _017786_);
  or g_086507_(_015938_, _017775_, _017797_);
  and g_086508_(_016081_, _016202_, _017808_);
  or g_086509_(_016070_, _016213_, _017819_);
  and g_086510_(_017753_, _017819_, _017830_);
  or g_086511_(_017742_, _017808_, _017841_);
  and g_086512_(_017544_, _017830_, _017852_);
  and g_086513_(_017566_, _017841_, _017863_);
  or g_086514_(_017852_, _017863_, _017874_);
  xor g_086515_(out[522], _015916_, _017885_);
  not g_086516_(_017885_, _017896_);
  or g_086517_(_017874_, _017896_, _017907_);
  not g_086518_(_017907_, _017918_);
  and g_086519_(_017797_, _017907_, _017929_);
  or g_086520_(_017786_, _017918_, _017940_);
  and g_086521_(_017874_, _017896_, _017951_);
  and g_086522_(_015938_, _017775_, _017962_);
  or g_086523_(_015949_, _017764_, _017973_);
  xor g_086524_(out[521], _015905_, _017984_);
  xor g_086525_(_054721_, _015905_, _017995_);
  and g_086526_(_017456_, _017830_, _018006_);
  or g_086527_(_017467_, _017841_, _018017_);
  and g_086528_(_017434_, _017841_, _018028_);
  or g_086529_(_017445_, _017830_, _018039_);
  and g_086530_(_018017_, _018039_, _018050_);
  or g_086531_(_018006_, _018028_, _018061_);
  and g_086532_(_017995_, _018061_, _018072_);
  or g_086533_(_017984_, _018050_, _018083_);
  or g_086534_(_017962_, _018072_, _018094_);
  or g_086535_(_017951_, _018094_, _018105_);
  and g_086536_(_017797_, _017973_, _018116_);
  xor g_086537_(_017874_, _017896_, _018127_);
  and g_086538_(_018116_, _018127_, _018138_);
  and g_086539_(_018083_, _018138_, _018149_);
  or g_086540_(_017940_, _018105_, _018160_);
  and g_086541_(_017984_, _018050_, _018171_);
  or g_086542_(_017995_, _018061_, _018182_);
  xor g_086543_(out[520], _015894_, _018193_);
  xor g_086544_(_054710_, _015894_, _018204_);
  and g_086545_(_017324_, _017841_, _018215_);
  or g_086546_(_017335_, _017830_, _018226_);
  and g_086547_(_017302_, _017830_, _018237_);
  or g_086548_(_017313_, _017841_, _018248_);
  and g_086549_(_018226_, _018248_, _018259_);
  or g_086550_(_018215_, _018237_, _018270_);
  and g_086551_(_018193_, _018259_, _018281_);
  or g_086552_(_018204_, _018270_, _018292_);
  and g_086553_(_018182_, _018292_, _018303_);
  or g_086554_(_018171_, _018281_, _018314_);
  and g_086555_(_018204_, _018270_, _018325_);
  or g_086556_(_018193_, _018259_, _018336_);
  and g_086557_(_018303_, _018336_, _018347_);
  or g_086558_(_018314_, _018325_, _018358_);
  and g_086559_(_018149_, _018347_, _018369_);
  or g_086560_(_018160_, _018358_, _018380_);
  xor g_086561_(out[518], _015872_, _018391_);
  xor g_086562_(_054633_, _015872_, _018402_);
  or g_086563_(_016224_, _017841_, _018413_);
  or g_086564_(_016246_, _017830_, _018424_);
  and g_086565_(_018413_, _018424_, _018435_);
  and g_086566_(_018402_, _018435_, _018446_);
  xor g_086567_(out[519], _015883_, _018457_);
  xor g_086568_(_054622_, _015883_, _018468_);
  or g_086569_(_017104_, _017841_, _018479_);
  or g_086570_(_017126_, _017830_, _018490_);
  and g_086571_(_018479_, _018490_, _018501_);
  not g_086572_(_018501_, _018512_);
  or g_086573_(_018468_, _018501_, _018523_);
  and g_086574_(_018468_, _018501_, _018534_);
  xor g_086575_(_018402_, _018435_, _018545_);
  xor g_086576_(_018391_, _018435_, _018556_);
  xor g_086577_(_018468_, _018501_, _018567_);
  xor g_086578_(_018457_, _018501_, _018578_);
  and g_086579_(_018545_, _018567_, _018589_);
  or g_086580_(_018556_, _018578_, _018600_);
  xor g_086581_(out[517], _015861_, _018611_);
  xor g_086582_(_054644_, _015861_, _018622_);
  and g_086583_(_016950_, _017830_, _018633_);
  or g_086584_(_016961_, _017841_, _018644_);
  and g_086585_(_016972_, _017841_, _018655_);
  or g_086586_(_016983_, _017830_, _018666_);
  and g_086587_(_018644_, _018666_, _018677_);
  or g_086588_(_018633_, _018655_, _018688_);
  and g_086589_(_018611_, _018677_, _018699_);
  or g_086590_(_018622_, _018688_, _018710_);
  xor g_086591_(out[516], _015850_, _018721_);
  xor g_086592_(_054655_, _015850_, _018732_);
  and g_086593_(_016796_, _017841_, _018743_);
  or g_086594_(_016807_, _017830_, _018754_);
  and g_086595_(_016774_, _017830_, _018765_);
  or g_086596_(_016785_, _017841_, _018776_);
  and g_086597_(_018754_, _018776_, _018787_);
  or g_086598_(_018743_, _018765_, _018798_);
  and g_086599_(_018721_, _018787_, _018809_);
  or g_086600_(_018732_, _018798_, _018820_);
  and g_086601_(_018710_, _018820_, _018831_);
  or g_086602_(_018699_, _018809_, _018842_);
  and g_086603_(_018622_, _018688_, _018853_);
  or g_086604_(_018611_, _018677_, _018864_);
  and g_086605_(_018732_, _018798_, _018875_);
  or g_086606_(_018721_, _018787_, _018886_);
  and g_086607_(_018864_, _018886_, _018897_);
  or g_086608_(_018853_, _018875_, _018908_);
  and g_086609_(_018831_, _018897_, _018919_);
  or g_086610_(_018842_, _018908_, _018930_);
  and g_086611_(_018589_, _018919_, _018941_);
  or g_086612_(_018600_, _018930_, _018952_);
  and g_086613_(_018369_, _018941_, _018963_);
  or g_086614_(_018380_, _018952_, _018974_);
  xor g_086615_(out[515], _015828_, _018985_);
  xor g_086616_(_054699_, _015828_, _018996_);
  and g_086617_(_016312_, _017841_, _019007_);
  and g_086618_(_016290_, _017830_, _019018_);
  or g_086619_(_019007_, _019018_, _019029_);
  not g_086620_(_019029_, _019040_);
  and g_086621_(_018985_, _019040_, _019051_);
  or g_086622_(_018996_, _019029_, _019062_);
  or g_086623_(out[513], out[514], _019073_);
  xor g_086624_(out[513], out[514], _019084_);
  xor g_086625_(_054666_, out[514], _019095_);
  or g_086626_(_016367_, _017830_, _019106_);
  or g_086627_(_016400_, _017841_, _019117_);
  and g_086628_(_019106_, _019117_, _019128_);
  not g_086629_(_019128_, _019139_);
  and g_086630_(_019095_, _019128_, _019150_);
  or g_086631_(_019084_, _019139_, _019161_);
  and g_086632_(_019062_, _019161_, _019172_);
  or g_086633_(_019051_, _019150_, _019183_);
  and g_086634_(_018996_, _019029_, _019194_);
  or g_086635_(_018985_, _019040_, _019205_);
  and g_086636_(_019084_, _019139_, _019216_);
  or g_086637_(_019095_, _019128_, _019227_);
  and g_086638_(_019205_, _019227_, _019238_);
  or g_086639_(_019194_, _019216_, _019249_);
  and g_086640_(_019172_, _019238_, _019260_);
  or g_086641_(_019183_, _019249_, _019271_);
  or g_086642_(_054413_, _017841_, _019282_);
  or g_086643_(_054534_, _017830_, _019293_);
  and g_086644_(_019282_, _019293_, _019304_);
  and g_086645_(out[513], _019304_, _019315_);
  not g_086646_(_019315_, _019326_);
  and g_086647_(_054545_, _017841_, _019337_);
  or g_086648_(out[496], _017830_, _019348_);
  and g_086649_(_054347_, _017830_, _019359_);
  or g_086650_(out[480], _017841_, _019370_);
  and g_086651_(_019348_, _019370_, _019381_);
  or g_086652_(_019337_, _019359_, _019392_);
  and g_086653_(out[512], _019392_, _019403_);
  or g_086654_(_054677_, _019381_, _019414_);
  xor g_086655_(out[513], _019304_, _019425_);
  xor g_086656_(_054666_, _019304_, _019436_);
  and g_086657_(_019414_, _019425_, _019447_);
  or g_086658_(_019403_, _019436_, _019458_);
  and g_086659_(_019326_, _019458_, _019469_);
  or g_086660_(_019315_, _019447_, _019480_);
  and g_086661_(_019260_, _019480_, _019491_);
  or g_086662_(_019271_, _019469_, _019502_);
  and g_086663_(_019183_, _019205_, _019513_);
  or g_086664_(_019172_, _019194_, _019524_);
  and g_086665_(_019502_, _019524_, _019535_);
  or g_086666_(_019491_, _019513_, _019546_);
  and g_086667_(_018963_, _019546_, _019557_);
  or g_086668_(_018974_, _019535_, _019568_);
  and g_086669_(_018589_, _018842_, _019579_);
  or g_086670_(_018600_, _018831_, _019590_);
  and g_086671_(_018864_, _019579_, _019601_);
  or g_086672_(_018853_, _019590_, _019612_);
  and g_086673_(_018446_, _018523_, _019623_);
  or g_086674_(_018534_, _019623_, _019634_);
  not g_086675_(_019634_, _019645_);
  and g_086676_(_019612_, _019645_, _019656_);
  or g_086677_(_019601_, _019634_, _019667_);
  and g_086678_(_018369_, _019667_, _019678_);
  or g_086679_(_018380_, _019656_, _019689_);
  and g_086680_(_018149_, _018314_, _019700_);
  or g_086681_(_018160_, _018303_, _019711_);
  and g_086682_(_017940_, _017973_, _019722_);
  or g_086683_(_017929_, _017962_, _019733_);
  and g_086684_(_019568_, _019733_, _019744_);
  or g_086685_(_019557_, _019722_, _019755_);
  and g_086686_(_019689_, _019711_, _019766_);
  or g_086687_(_019678_, _019700_, _019777_);
  and g_086688_(_019744_, _019766_, _019788_);
  or g_086689_(_019755_, _019777_, _019799_);
  and g_086690_(_054677_, _019381_, _019810_);
  or g_086691_(out[512], _019392_, _019821_);
  and g_086692_(_019260_, _019821_, _019832_);
  or g_086693_(_019271_, _019810_, _019843_);
  and g_086694_(_019447_, _019832_, _019854_);
  or g_086695_(_019458_, _019843_, _019865_);
  and g_086696_(_018963_, _019854_, _019876_);
  or g_086697_(_018974_, _019865_, _019887_);
  and g_086698_(_019799_, _019887_, _019898_);
  or g_086699_(_019788_, _019876_, _019909_);
  and g_086700_(_015949_, _019898_, _019920_);
  or g_086701_(_015938_, _019909_, _019931_);
  and g_086702_(_017775_, _019909_, _019942_);
  or g_086703_(_017764_, _019898_, _019953_);
  and g_086704_(_019931_, _019953_, _019964_);
  or g_086705_(_019920_, _019942_, _019975_);
  and g_086706_(_015806_, _019975_, _019986_);
  or g_086707_(_015817_, _019964_, _019997_);
  xor g_086708_(out[538], _015784_, _020008_);
  xor g_086709_(_054864_, _015784_, _020019_);
  and g_086710_(_017874_, _019909_, _020030_);
  and g_086711_(_017885_, _019898_, _020041_);
  or g_086712_(_020030_, _020041_, _020052_);
  not g_086713_(_020052_, _020063_);
  and g_086714_(_020008_, _020063_, _020074_);
  or g_086715_(_020019_, _020052_, _020085_);
  and g_086716_(_015817_, _019964_, _020096_);
  or g_086717_(_015806_, _019975_, _020107_);
  xor g_086718_(out[537], _015773_, _020118_);
  xor g_086719_(_054853_, _015773_, _020129_);
  and g_086720_(_017984_, _019898_, _020140_);
  or g_086721_(_017995_, _019909_, _020151_);
  and g_086722_(_018061_, _019909_, _020162_);
  or g_086723_(_018050_, _019898_, _020173_);
  and g_086724_(_020151_, _020173_, _020184_);
  or g_086725_(_020140_, _020162_, _020195_);
  and g_086726_(_020129_, _020195_, _020206_);
  or g_086727_(_020118_, _020184_, _020217_);
  and g_086728_(_020118_, _020184_, _020228_);
  or g_086729_(_020129_, _020195_, _020239_);
  xor g_086730_(out[536], _015762_, _020250_);
  xor g_086731_(_054842_, _015762_, _020261_);
  and g_086732_(_018193_, _019898_, _020272_);
  or g_086733_(_018204_, _019909_, _020283_);
  and g_086734_(_018270_, _019909_, _020294_);
  or g_086735_(_018259_, _019898_, _020305_);
  and g_086736_(_020283_, _020305_, _020316_);
  or g_086737_(_020272_, _020294_, _020327_);
  and g_086738_(_020250_, _020316_, _020338_);
  or g_086739_(_020261_, _020327_, _020349_);
  and g_086740_(_020239_, _020349_, _020360_);
  or g_086741_(_020228_, _020338_, _020371_);
  xor g_086742_(out[534], _015740_, _020382_);
  xor g_086743_(_054765_, _015740_, _020393_);
  or g_086744_(_018391_, _019909_, _020404_);
  or g_086745_(_018435_, _019898_, _020415_);
  and g_086746_(_020404_, _020415_, _020426_);
  not g_086747_(_020426_, _020437_);
  and g_086748_(_020393_, _020426_, _020448_);
  or g_086749_(_020382_, _020437_, _020459_);
  xor g_086750_(out[535], _015751_, _020470_);
  xor g_086751_(_054754_, _015751_, _020481_);
  and g_086752_(_018457_, _019898_, _020492_);
  or g_086753_(_018468_, _019909_, _020503_);
  and g_086754_(_018501_, _019909_, _020514_);
  or g_086755_(_018512_, _019898_, _020525_);
  and g_086756_(_020503_, _020525_, _020536_);
  or g_086757_(_020492_, _020514_, _020547_);
  and g_086758_(_020481_, _020547_, _020558_);
  or g_086759_(_020470_, _020536_, _020569_);
  and g_086760_(_020459_, _020569_, _020580_);
  or g_086761_(_020448_, _020558_, _020591_);
  xor g_086762_(out[533], _015729_, _020602_);
  xor g_086763_(_054776_, _015729_, _020613_);
  and g_086764_(_018622_, _019898_, _020624_);
  or g_086765_(_018611_, _019909_, _020635_);
  and g_086766_(_018677_, _019909_, _020646_);
  or g_086767_(_018688_, _019898_, _020657_);
  and g_086768_(_020635_, _020657_, _020668_);
  or g_086769_(_020624_, _020646_, _020679_);
  and g_086770_(_020613_, _020668_, _020690_);
  or g_086771_(_020602_, _020679_, _020701_);
  and g_086772_(_020602_, _020679_, _020712_);
  or g_086773_(_020613_, _020668_, _020723_);
  xor g_086774_(out[532], _015718_, _020734_);
  xor g_086775_(_054787_, _015718_, _020745_);
  and g_086776_(_018721_, _019898_, _020756_);
  or g_086777_(_018732_, _019909_, _020767_);
  and g_086778_(_018798_, _019909_, _020778_);
  or g_086779_(_018787_, _019898_, _020789_);
  and g_086780_(_020767_, _020789_, _020800_);
  or g_086781_(_020756_, _020778_, _020811_);
  and g_086782_(_020734_, _020800_, _020822_);
  or g_086783_(_020745_, _020811_, _020833_);
  and g_086784_(_020723_, _020833_, _020844_);
  or g_086785_(_020712_, _020822_, _020855_);
  xor g_086786_(out[531], _015696_, _020866_);
  xor g_086787_(_054831_, _015696_, _020877_);
  or g_086788_(_019029_, _019898_, _020888_);
  not g_086789_(_020888_, _020899_);
  and g_086790_(_018996_, _019898_, _020910_);
  or g_086791_(_018985_, _019909_, _020921_);
  and g_086792_(_020888_, _020921_, _020932_);
  or g_086793_(_020899_, _020910_, _020943_);
  and g_086794_(_020866_, _020943_, _020954_);
  or g_086795_(_020877_, _020932_, _020965_);
  or g_086796_(out[529], out[530], _020976_);
  xor g_086797_(out[529], out[530], _020987_);
  xor g_086798_(_054798_, out[530], _020998_);
  or g_086799_(_019084_, _019909_, _021009_);
  or g_086800_(_019128_, _019898_, _021020_);
  and g_086801_(_021009_, _021020_, _021031_);
  not g_086802_(_021031_, _021042_);
  and g_086803_(_020998_, _021031_, _021053_);
  or g_086804_(_020987_, _021042_, _021064_);
  and g_086805_(_020965_, _021064_, _021075_);
  or g_086806_(_020954_, _021053_, _021086_);
  and g_086807_(_020877_, _020932_, _021097_);
  or g_086808_(_020866_, _020943_, _021108_);
  and g_086809_(_020987_, _021042_, _021119_);
  or g_086810_(_020998_, _021031_, _021130_);
  and g_086811_(_021108_, _021130_, _021141_);
  or g_086812_(_021097_, _021119_, _021152_);
  and g_086813_(_021075_, _021141_, _021163_);
  or g_086814_(_021086_, _021152_, _021174_);
  or g_086815_(_054666_, _019909_, _021185_);
  or g_086816_(_019304_, _019898_, _021196_);
  and g_086817_(_021185_, _021196_, _021207_);
  and g_086818_(out[529], _021207_, _021218_);
  not g_086819_(_021218_, _021229_);
  and g_086820_(_019392_, _019909_, _021240_);
  or g_086821_(_019381_, _019898_, _021251_);
  and g_086822_(_054677_, _019898_, _021262_);
  or g_086823_(out[512], _019909_, _021273_);
  and g_086824_(_021251_, _021273_, _021284_);
  or g_086825_(_021240_, _021262_, _021295_);
  and g_086826_(out[528], _021295_, _021306_);
  or g_086827_(_054809_, _021284_, _021317_);
  xor g_086828_(out[529], _021207_, _021328_);
  xor g_086829_(_054798_, _021207_, _021339_);
  and g_086830_(_021317_, _021328_, _021350_);
  or g_086831_(_021306_, _021339_, _021361_);
  and g_086832_(_021229_, _021361_, _021372_);
  or g_086833_(_021218_, _021350_, _021383_);
  and g_086834_(_021163_, _021383_, _021394_);
  or g_086835_(_021174_, _021372_, _021405_);
  and g_086836_(_021086_, _021108_, _021416_);
  or g_086837_(_021075_, _021097_, _021427_);
  and g_086838_(_021405_, _021427_, _021438_);
  or g_086839_(_021394_, _021416_, _021449_);
  and g_086840_(_020745_, _020811_, _021460_);
  or g_086841_(_020734_, _020800_, _021471_);
  and g_086842_(_020261_, _020327_, _021482_);
  or g_086843_(_020250_, _020316_, _021493_);
  and g_086844_(_020470_, _020536_, _021504_);
  or g_086845_(_020481_, _020547_, _021515_);
  xor g_086846_(_020019_, _020052_, _021526_);
  xor g_086847_(_020008_, _020052_, _021537_);
  and g_086848_(_019997_, _020107_, _021548_);
  or g_086849_(_019986_, _020096_, _021559_);
  and g_086850_(_021526_, _021548_, _021570_);
  or g_086851_(_021537_, _021559_, _021581_);
  and g_086852_(_020217_, _020371_, _021592_);
  or g_086853_(_020206_, _020360_, _021603_);
  and g_086854_(_021570_, _021592_, _021614_);
  or g_086855_(_021581_, _021603_, _021625_);
  and g_086856_(_020217_, _020360_, _021636_);
  or g_086857_(_020206_, _020371_, _021647_);
  and g_086858_(_021493_, _021570_, _021658_);
  or g_086859_(_021482_, _021581_, _021669_);
  and g_086860_(_021636_, _021658_, _021680_);
  or g_086861_(_021647_, _021669_, _021691_);
  xor g_086862_(_020393_, _020426_, _021702_);
  xor g_086863_(_020382_, _020426_, _021713_);
  and g_086864_(_020569_, _021515_, _021724_);
  or g_086865_(_020558_, _021504_, _021735_);
  and g_086866_(_021702_, _021724_, _021746_);
  or g_086867_(_021713_, _021735_, _021757_);
  and g_086868_(_020701_, _021471_, _021768_);
  or g_086869_(_020690_, _021460_, _021779_);
  and g_086870_(_020844_, _021768_, _021790_);
  or g_086871_(_020855_, _021779_, _021801_);
  and g_086872_(_021746_, _021790_, _021812_);
  or g_086873_(_021757_, _021801_, _021823_);
  and g_086874_(_021449_, _021812_, _021834_);
  or g_086875_(_021438_, _021823_, _021845_);
  and g_086876_(_020855_, _021746_, _021856_);
  or g_086877_(_020844_, _021757_, _021867_);
  and g_086878_(_020701_, _021856_, _021878_);
  or g_086879_(_020690_, _021867_, _021889_);
  and g_086880_(_020591_, _021515_, _021900_);
  or g_086881_(_020580_, _021504_, _021911_);
  and g_086882_(_021889_, _021911_, _021922_);
  or g_086883_(_021878_, _021900_, _021933_);
  and g_086884_(_021845_, _021922_, _021944_);
  or g_086885_(_021834_, _021933_, _021955_);
  and g_086886_(_021680_, _021955_, _021966_);
  or g_086887_(_021691_, _021944_, _021977_);
  and g_086888_(_019997_, _020074_, _021988_);
  or g_086889_(_019986_, _020085_, _021999_);
  and g_086890_(_020107_, _021625_, _022010_);
  or g_086891_(_020096_, _021614_, _022021_);
  and g_086892_(_021999_, _022010_, _022032_);
  or g_086893_(_021988_, _022021_, _022043_);
  and g_086894_(_021977_, _022032_, _022054_);
  or g_086895_(_021966_, _022043_, _022065_);
  and g_086896_(_054809_, _021284_, _022076_);
  or g_086897_(out[528], _021295_, _022087_);
  and g_086898_(_021350_, _022087_, _022098_);
  or g_086899_(_021361_, _022076_, _022109_);
  and g_086900_(_021163_, _022098_, _022120_);
  or g_086901_(_021174_, _022109_, _022131_);
  and g_086902_(_021812_, _022120_, _022142_);
  or g_086903_(_021823_, _022131_, _022153_);
  and g_086904_(_021680_, _022142_, _022164_);
  or g_086905_(_021691_, _022153_, _022175_);
  and g_086906_(_022065_, _022175_, _022186_);
  or g_086907_(_022054_, _022164_, _022197_);
  and g_086908_(_015817_, _022186_, _022208_);
  not g_086909_(_022208_, _022219_);
  or g_086910_(_019964_, _022186_, _022230_);
  not g_086911_(_022230_, _022241_);
  and g_086912_(_022219_, _022230_, _022252_);
  or g_086913_(_022208_, _022241_, _022263_);
  and g_086914_(_015685_, _022252_, _022274_);
  or g_086915_(_015674_, _022263_, _022285_);
  and g_086916_(out[561], out[562], _022296_);
  or g_086917_(out[564], out[563], _022307_);
  or g_086918_(out[563], _022296_, _022318_);
  or g_086919_(_022296_, _022307_, _022329_);
  or g_086920_(out[565], _022329_, _022340_);
  and g_086921_(out[566], _022340_, _022351_);
  and g_086922_(out[567], _022351_, _022362_);
  or g_086923_(out[568], _022362_, _022373_);
  or g_086924_(out[569], _022373_, _022384_);
  or g_086925_(out[570], _022384_, _022395_);
  xor g_086926_(_055007_, _022395_, _022406_);
  xor g_086927_(out[571], _022395_, _022417_);
  and g_086928_(_022274_, _022406_, _022428_);
  or g_086929_(_022285_, _022417_, _022439_);
  and g_086930_(out[577], out[578], _022450_);
  or g_086931_(out[580], out[579], _022461_);
  or g_086932_(out[579], _022450_, _022472_);
  or g_086933_(_022450_, _022461_, _022483_);
  or g_086934_(out[581], _022483_, _022494_);
  and g_086935_(out[582], _022494_, _022505_);
  and g_086936_(out[583], _022505_, _022516_);
  or g_086937_(out[584], _022516_, _022527_);
  or g_086938_(out[585], _022527_, _022538_);
  or g_086939_(out[586], _022538_, _022549_);
  xor g_086940_(_055139_, _022549_, _022560_);
  xor g_086941_(out[587], _022549_, _022571_);
  and g_086942_(_022428_, _022560_, _022582_);
  or g_086943_(_022439_, _022571_, _022593_);
  and g_086944_(out[593], out[594], _022604_);
  or g_086945_(out[596], out[595], _022615_);
  or g_086946_(out[595], _022604_, _022626_);
  or g_086947_(_022604_, _022615_, _022637_);
  or g_086948_(out[597], _022637_, _022648_);
  and g_086949_(out[598], _022648_, _022659_);
  and g_086950_(out[599], _022659_, _022670_);
  or g_086951_(out[600], _022670_, _022681_);
  or g_086952_(out[601], _022681_, _022692_);
  or g_086953_(out[602], _022692_, _022703_);
  xor g_086954_(_055271_, _022703_, _022714_);
  xor g_086955_(out[603], _022703_, _022725_);
  and g_086956_(_022582_, _022714_, _022736_);
  or g_086957_(_022593_, _022725_, _022747_);
  and g_086958_(out[609], out[610], _022758_);
  or g_086959_(out[612], out[611], _022769_);
  or g_086960_(out[611], _022758_, _022780_);
  or g_086961_(_022758_, _022769_, _022791_);
  or g_086962_(out[613], _022791_, _022802_);
  and g_086963_(out[614], _022802_, _022813_);
  and g_086964_(out[615], _022813_, _022824_);
  or g_086965_(out[616], _022824_, _022835_);
  or g_086966_(out[617], _022835_, _022846_);
  or g_086967_(out[618], _022846_, _022857_);
  xor g_086968_(_055403_, _022857_, _022868_);
  xor g_086969_(out[619], _022857_, _022879_);
  and g_086970_(_022736_, _022868_, _022890_);
  or g_086971_(_022747_, _022879_, _022901_);
  and g_086972_(out[625], out[626], _022912_);
  or g_086973_(out[628], out[627], _022923_);
  or g_086974_(out[627], _022912_, _022934_);
  or g_086975_(_022912_, _022923_, _022945_);
  or g_086976_(out[629], _022945_, _022956_);
  and g_086977_(out[630], _022956_, _022967_);
  and g_086978_(out[631], _022967_, _022978_);
  or g_086979_(out[632], _022978_, _022989_);
  or g_086980_(out[633], _022989_, _023000_);
  or g_086981_(out[634], _023000_, _023011_);
  xor g_086982_(_055535_, _023011_, _023022_);
  xor g_086983_(out[635], _023011_, _023033_);
  and g_086984_(_022890_, _023022_, _023044_);
  or g_086985_(_022901_, _023033_, _023055_);
  and g_086986_(out[641], out[642], _023066_);
  or g_086987_(out[644], out[643], _023077_);
  or g_086988_(out[643], _023066_, _023088_);
  or g_086989_(_023066_, _023077_, _023099_);
  or g_086990_(out[645], _023099_, _023110_);
  and g_086991_(out[646], _023110_, _023121_);
  and g_086992_(out[647], _023121_, _023132_);
  or g_086993_(out[648], _023132_, _023143_);
  or g_086994_(out[649], _023143_, _023154_);
  or g_086995_(out[650], _023154_, _023165_);
  xor g_086996_(_055667_, _023165_, _023176_);
  xor g_086997_(out[651], _023165_, _023187_);
  and g_086998_(_023044_, _023176_, _023198_);
  or g_086999_(_023055_, _023187_, _023209_);
  and g_087000_(out[657], out[658], _023220_);
  or g_087001_(out[660], out[659], _023231_);
  or g_087002_(out[659], _023220_, _023242_);
  or g_087003_(_023220_, _023231_, _023253_);
  or g_087004_(out[661], _023253_, _023264_);
  and g_087005_(out[662], _023264_, _023275_);
  and g_087006_(out[663], _023275_, _023286_);
  or g_087007_(out[664], _023286_, _023297_);
  or g_087008_(out[665], _023297_, _023308_);
  or g_087009_(out[666], _023308_, _023319_);
  xor g_087010_(out[667], _023319_, _023330_);
  or g_087011_(_023209_, _023330_, _023341_);
  not g_087012_(_023341_, _023352_);
  and g_087013_(out[673], out[674], _023363_);
  or g_087014_(out[676], out[675], _023374_);
  or g_087015_(out[675], _023363_, _023385_);
  or g_087016_(_023363_, _023374_, _023396_);
  or g_087017_(out[677], _023396_, _023407_);
  and g_087018_(out[678], _023407_, _023418_);
  and g_087019_(out[679], _023418_, _023429_);
  or g_087020_(out[680], _023429_, _023440_);
  or g_087021_(out[681], _023440_, _023451_);
  or g_087022_(out[682], _023451_, _023462_);
  xor g_087023_(_055931_, _023462_, _023473_);
  xor g_087024_(out[683], _023462_, _023484_);
  and g_087025_(_023352_, _023473_, _023495_);
  or g_087026_(_023341_, _023484_, _023506_);
  and g_087027_(out[689], out[690], _023517_);
  or g_087028_(out[692], out[691], _023528_);
  or g_087029_(out[691], _023517_, _023539_);
  or g_087030_(_023517_, _023528_, _023550_);
  or g_087031_(out[693], _023550_, _023561_);
  and g_087032_(out[694], _023561_, _023572_);
  and g_087033_(out[695], _023572_, _023583_);
  or g_087034_(out[696], _023583_, _023594_);
  or g_087035_(out[697], _023594_, _023605_);
  or g_087036_(out[698], _023605_, _023616_);
  xor g_087037_(_000098_, _023616_, _023627_);
  xor g_087038_(out[699], _023616_, _023638_);
  and g_087039_(_023495_, _023627_, _023649_);
  or g_087040_(_023506_, _023638_, _023660_);
  and g_087041_(out[705], out[706], _023671_);
  or g_087042_(out[708], out[707], _023682_);
  or g_087043_(out[707], _023671_, _023693_);
  or g_087044_(_023671_, _023682_, _023704_);
  or g_087045_(out[709], _023704_, _023715_);
  and g_087046_(out[710], _023715_, _023726_);
  and g_087047_(out[711], _023726_, _023737_);
  or g_087048_(out[712], _023737_, _023748_);
  or g_087049_(out[713], _023748_, _023759_);
  or g_087050_(out[714], _023759_, _023770_);
  xor g_087051_(_000230_, _023770_, _023781_);
  xor g_087052_(out[715], _023770_, _023792_);
  and g_087053_(_023649_, _023781_, _023803_);
  or g_087054_(_023660_, _023792_, _023814_);
  and g_087055_(out[721], out[722], _023825_);
  or g_087056_(out[724], out[723], _023836_);
  or g_087057_(out[723], _023825_, _023847_);
  or g_087058_(_023825_, _023836_, _023858_);
  or g_087059_(out[725], _023858_, _023869_);
  and g_087060_(out[726], _023869_, _023880_);
  and g_087061_(out[727], _023880_, _023891_);
  or g_087062_(out[728], _023891_, _023902_);
  or g_087063_(out[729], _023902_, _023913_);
  or g_087064_(out[730], _023913_, _023924_);
  xor g_087065_(_000362_, _023924_, _023935_);
  xor g_087066_(out[731], _023924_, _023946_);
  and g_087067_(_023803_, _023935_, _023957_);
  or g_087068_(_023814_, _023946_, _023968_);
  and g_087069_(out[737], out[738], _023979_);
  or g_087070_(out[740], out[739], _023990_);
  or g_087071_(out[739], _023979_, _024001_);
  or g_087072_(_023979_, _023990_, _024012_);
  or g_087073_(out[741], _024012_, _024023_);
  and g_087074_(out[742], _024023_, _024034_);
  and g_087075_(out[743], _024034_, _024045_);
  or g_087076_(out[744], _024045_, _024056_);
  or g_087077_(out[745], _024056_, _024067_);
  or g_087078_(out[746], _024067_, _024078_);
  xor g_087079_(_000494_, _024078_, _024089_);
  xor g_087080_(out[747], _024078_, _024100_);
  and g_087081_(_023957_, _024089_, _024111_);
  or g_087082_(_023968_, _024100_, _024122_);
  and g_087083_(out[753], out[754], _024133_);
  or g_087084_(out[756], out[755], _024144_);
  or g_087085_(out[755], _024133_, _024155_);
  or g_087086_(_024133_, _024144_, _024166_);
  or g_087087_(out[757], _024166_, _024177_);
  and g_087088_(out[758], _024177_, _024188_);
  and g_087089_(out[759], _024188_, _024199_);
  or g_087090_(out[760], _024199_, _024210_);
  or g_087091_(out[761], _024210_, _024221_);
  or g_087092_(out[762], _024221_, _024232_);
  xor g_087093_(_000626_, _024232_, _024243_);
  xor g_087094_(out[763], _024232_, _024254_);
  and g_087095_(_024111_, _024243_, _024265_);
  or g_087096_(_024122_, _024254_, _024276_);
  and g_087097_(out[769], out[770], _024287_);
  or g_087098_(out[772], out[771], _024298_);
  or g_087099_(out[771], _024287_, _024309_);
  or g_087100_(_024287_, _024298_, _024320_);
  or g_087101_(out[773], _024320_, _024331_);
  and g_087102_(out[774], _024331_, _024342_);
  and g_087103_(out[775], _024342_, _024353_);
  or g_087104_(out[776], _024353_, _024364_);
  or g_087105_(out[777], _024364_, _024375_);
  or g_087106_(out[778], _024375_, _024386_);
  xor g_087107_(_000758_, _024386_, _024397_);
  xor g_087108_(out[779], _024386_, _024408_);
  and g_087109_(_024265_, _024397_, _024419_);
  or g_087110_(_024276_, _024408_, _024430_);
  and g_087111_(out[785], out[786], _024441_);
  or g_087112_(out[788], out[787], _024452_);
  or g_087113_(out[787], _024441_, _024463_);
  or g_087114_(_024441_, _024452_, _024474_);
  or g_087115_(out[789], _024474_, _024485_);
  and g_087116_(out[790], _024485_, _024496_);
  and g_087117_(out[791], _024496_, _024507_);
  or g_087118_(out[792], _024507_, _024518_);
  or g_087119_(out[793], _024518_, _024529_);
  or g_087120_(out[794], _024529_, _024540_);
  xor g_087121_(_000890_, _024540_, _024551_);
  xor g_087122_(out[795], _024540_, _024562_);
  and g_087123_(_024419_, _024551_, _024573_);
  or g_087124_(_024430_, _024562_, _024584_);
  and g_087125_(out[801], out[802], _024595_);
  or g_087126_(out[804], out[803], _024606_);
  or g_087127_(out[803], _024595_, _024617_);
  or g_087128_(_024595_, _024606_, _024628_);
  or g_087129_(out[805], _024628_, _024639_);
  and g_087130_(out[806], _024639_, _024650_);
  and g_087131_(out[807], _024650_, _024661_);
  or g_087132_(out[808], _024661_, _024672_);
  or g_087133_(out[809], _024672_, _024683_);
  or g_087134_(out[810], _024683_, _024694_);
  xor g_087135_(_001022_, _024694_, _024705_);
  xor g_087136_(out[811], _024694_, _024716_);
  and g_087137_(_024573_, _024705_, _024727_);
  or g_087138_(_024584_, _024716_, _024738_);
  and g_087139_(out[817], out[818], _024749_);
  or g_087140_(out[820], out[819], _024760_);
  or g_087141_(out[819], _024749_, _024771_);
  or g_087142_(_024749_, _024760_, _024782_);
  or g_087143_(out[821], _024782_, _024793_);
  and g_087144_(out[822], _024793_, _024804_);
  and g_087145_(out[823], _024804_, _024815_);
  or g_087146_(out[824], _024815_, _024826_);
  or g_087147_(out[825], _024826_, _024837_);
  or g_087148_(out[826], _024837_, _024848_);
  xor g_087149_(_001154_, _024848_, _024859_);
  xor g_087150_(out[827], _024848_, _024870_);
  and g_087151_(_024727_, _024859_, _024881_);
  or g_087152_(_024738_, _024870_, _024892_);
  and g_087153_(out[833], out[834], _024903_);
  or g_087154_(out[836], out[835], _024914_);
  or g_087155_(out[835], _024903_, _024925_);
  or g_087156_(_024903_, _024914_, _024936_);
  or g_087157_(out[837], _024936_, _024947_);
  and g_087158_(out[838], _024947_, _024958_);
  and g_087159_(out[839], _024958_, _024969_);
  or g_087160_(out[840], _024969_, _024980_);
  or g_087161_(out[841], _024980_, _024991_);
  or g_087162_(out[842], _024991_, _025002_);
  xor g_087163_(_001286_, _025002_, _025013_);
  xor g_087164_(out[843], _025002_, _025024_);
  and g_087165_(_024881_, _025013_, _025035_);
  or g_087166_(_024892_, _025024_, _025046_);
  and g_087167_(out[849], out[850], _025057_);
  or g_087168_(out[852], out[851], _025068_);
  or g_087169_(out[851], _025057_, _025079_);
  or g_087170_(_025057_, _025068_, _025090_);
  or g_087171_(out[853], _025090_, _025101_);
  and g_087172_(out[854], _025101_, _025112_);
  and g_087173_(out[855], _025112_, _025123_);
  or g_087174_(out[856], _025123_, _025134_);
  or g_087175_(out[857], _025134_, _025145_);
  or g_087176_(out[858], _025145_, _025156_);
  xor g_087177_(_001418_, _025156_, _025167_);
  xor g_087178_(out[859], _025156_, _025178_);
  and g_087179_(_025035_, _025167_, _025189_);
  or g_087180_(_025046_, _025178_, _025200_);
  and g_087181_(out[865], out[866], _025211_);
  or g_087182_(out[868], out[867], _025222_);
  or g_087183_(out[867], _025211_, _025233_);
  or g_087184_(_025211_, _025222_, _025244_);
  or g_087185_(out[869], _025244_, _025255_);
  and g_087186_(out[870], _025255_, _025266_);
  and g_087187_(out[871], _025266_, _025277_);
  or g_087188_(out[872], _025277_, _025288_);
  or g_087189_(out[873], _025288_, _025299_);
  or g_087190_(out[874], _025299_, _025310_);
  xor g_087191_(out[875], _025310_, _025321_);
  not g_087192_(_025321_, _025332_);
  and g_087193_(_025189_, _025332_, _025343_);
  or g_087194_(_025200_, _025321_, _025354_);
  and g_087195_(out[881], out[882], _025365_);
  or g_087196_(out[884], out[883], _025376_);
  or g_087197_(out[883], _025365_, _025387_);
  or g_087198_(_025365_, _025376_, _025398_);
  or g_087199_(out[885], _025398_, _025409_);
  and g_087200_(out[886], _025409_, _025420_);
  and g_087201_(out[887], _025420_, _025431_);
  or g_087202_(out[888], _025431_, _025442_);
  or g_087203_(out[889], _025442_, _025453_);
  or g_087204_(out[890], _025453_, _025464_);
  xor g_087205_(_001682_, _025464_, _025475_);
  xor g_087206_(out[891], _025464_, _025486_);
  and g_087207_(_025343_, _025475_, _025497_);
  or g_087208_(_025354_, _025486_, _025508_);
  and g_087209_(out[897], out[898], _025519_);
  or g_087210_(out[900], out[899], _025530_);
  or g_087211_(out[899], _025519_, _025541_);
  or g_087212_(_025519_, _025530_, _025552_);
  or g_087213_(out[901], _025552_, _025563_);
  and g_087214_(out[902], _025563_, _025574_);
  and g_087215_(out[903], _025574_, _025585_);
  or g_087216_(out[904], _025585_, _025596_);
  or g_087217_(out[905], _025596_, _025607_);
  or g_087218_(out[906], _025607_, _025618_);
  xor g_087219_(_001814_, _025618_, _025629_);
  xor g_087220_(out[907], _025618_, _025640_);
  and g_087221_(_025497_, _025629_, _025651_);
  or g_087222_(_025508_, _025640_, _025662_);
  and g_087223_(out[913], out[914], _025673_);
  or g_087224_(out[916], out[915], _025684_);
  or g_087225_(out[915], _025673_, _025695_);
  or g_087226_(_025673_, _025684_, _025706_);
  or g_087227_(out[917], _025706_, _025717_);
  and g_087228_(out[918], _025717_, _025728_);
  and g_087229_(out[919], _025728_, _025739_);
  or g_087230_(out[920], _025739_, _025750_);
  or g_087231_(out[921], _025750_, _025761_);
  or g_087232_(out[922], _025761_, _025772_);
  xor g_087233_(_001946_, _025772_, _025783_);
  xor g_087234_(out[923], _025772_, _025794_);
  or g_087235_(_025662_, _025794_, _025805_);
  not g_087236_(_025805_, _025816_);
  and g_087237_(out[929], out[930], _025827_);
  or g_087238_(out[932], out[931], _025838_);
  or g_087239_(out[931], _025827_, _025849_);
  or g_087240_(_025827_, _025838_, _025860_);
  or g_087241_(out[933], _025860_, _025871_);
  and g_087242_(out[934], _025871_, _025882_);
  and g_087243_(out[935], _025882_, _025893_);
  or g_087244_(out[936], _025893_, _025904_);
  or g_087245_(out[937], _025904_, _025915_);
  or g_087246_(out[938], _025915_, _025926_);
  xor g_087247_(out[939], _025926_, _025937_);
  not g_087248_(_025937_, _025948_);
  or g_087249_(_025805_, _025937_, _025959_);
  not g_087250_(_025959_, _025970_);
  and g_087251_(out[945], out[946], _025981_);
  or g_087252_(out[947], _025981_, _025992_);
  or g_087253_(out[948], _025992_, _026003_);
  or g_087254_(out[949], _026003_, _026014_);
  and g_087255_(out[950], _026014_, _026025_);
  and g_087256_(out[951], _026025_, _026036_);
  or g_087257_(out[952], _026036_, _026047_);
  or g_087258_(out[953], _026047_, _026058_);
  or g_087259_(out[954], _026058_, _026069_);
  xor g_087260_(out[955], _026069_, _026080_);
  not g_087261_(_026080_, _026091_);
  or g_087262_(_025959_, _026080_, _026102_);
  xor g_087263_(_015553_, _026102_, _026113_);
  xor g_087264_(out[473], _015498_, _026124_);
  not g_087265_(_026124_, _026135_);
  xor g_087266_(out[474], _015509_, _026146_);
  not g_087267_(_026146_, _026157_);
  xor g_087268_(out[394], _014739_, _026168_);
  xor g_087269_(_004685_, _014739_, _026179_);
  xor g_087270_(out[388], _014673_, _026190_);
  xor g_087271_(_053797_, _014673_, _026201_);
  xor g_087272_(out[372], _014519_, _026212_);
  not g_087273_(_026212_, _026223_);
  xor g_087274_(out[375], _014552_, _026234_);
  xor g_087275_(_053643_, _014552_, _026245_);
  xor g_087276_(out[359], _014398_, _026256_);
  xor g_087277_(_053544_, _014398_, _026267_);
  and g_087278_(_014321_, _014464_, _026278_);
  or g_087279_(_014332_, _014453_, _026289_);
  xor g_087280_(out[330], _014123_, _026300_);
  xor g_087281_(_004553_, _014123_, _026311_);
  and g_087282_(_014024_, _014145_, _026322_);
  or g_087283_(_014013_, _014156_, _026333_);
  and g_087284_(_014013_, _014156_, _026344_);
  or g_087285_(_014024_, _014145_, _026355_);
  xor g_087286_(out[298], _013815_, _026366_);
  xor g_087287_(_004487_, _013815_, _026377_);
  and g_087288_(_013705_, _013848_, _026388_);
  or g_087289_(_013716_, _013837_, _026399_);
  xor g_087290_(out[202], _012891_, _026410_);
  xor g_087291_(out[202], _012902_, _026421_);
  and g_087292_(_012781_, _012935_, _026432_);
  or g_087293_(_012792_, _012924_, _026443_);
  xor g_087294_(out[154], _012429_, _026454_);
  xor g_087295_(_003607_, _012429_, _026465_);
  and g_087296_(_012319_, _012462_, _026476_);
  or g_087297_(_012330_, _012451_, _026487_);
  xor g_087298_(out[138], _012275_, _026498_);
  not g_087299_(_026498_, _026509_);
  xor g_087300_(out[106], _011967_, _026520_);
  xor g_087301_(out[100], _011901_, _026531_);
  xor g_087302_(_003134_, _011901_, _026542_);
  xor g_087303_(out[84], _011747_, _026553_);
  xor g_087304_(_003002_, _011747_, _026564_);
  or g_087305_(out[81], out[82], _026575_);
  xor g_087306_(out[81], out[82], _026586_);
  xor g_087307_(_003013_, out[82], _026597_);
  or g_087308_(out[65], out[66], _026608_);
  xor g_087309_(out[65], out[66], _026619_);
  xor g_087310_(_002881_, out[66], _026630_);
  xor g_087311_(out[68], _004872_, _026641_);
  xor g_087312_(_002870_, _004872_, _026652_);
  and g_087313_(_010493_, _011615_, _026663_);
  or g_087314_(_010504_, _011626_, _026674_);
  and g_087315_(_010570_, _011626_, _026685_);
  or g_087316_(_010559_, _011615_, _026696_);
  and g_087317_(_026674_, _026696_, _026707_);
  or g_087318_(_026663_, _026685_, _026718_);
  and g_087319_(_026652_, _026718_, _026729_);
  or g_087320_(_026641_, _026707_, _026740_);
  or g_087321_(_010801_, _011615_, _026751_);
  not g_087322_(_026751_, _026762_);
  and g_087323_(_010768_, _011615_, _026773_);
  not g_087324_(_026773_, _026784_);
  and g_087325_(_026751_, _026784_, _026795_);
  or g_087326_(_026762_, _026773_, _026806_);
  xor g_087327_(out[67], _004850_, _026817_);
  xor g_087328_(_002914_, _004850_, _026828_);
  and g_087329_(_026795_, _026828_, _026839_);
  or g_087330_(_026806_, _026817_, _026850_);
  xor g_087331_(out[69], _004883_, _026861_);
  xor g_087332_(_002859_, _004883_, _026872_);
  and g_087333_(_010394_, _011615_, _026883_);
  or g_087334_(_010383_, _011626_, _026894_);
  and g_087335_(_010460_, _011626_, _026905_);
  or g_087336_(_010449_, _011615_, _026916_);
  and g_087337_(_026894_, _026916_, _026927_);
  or g_087338_(_026883_, _026905_, _026938_);
  and g_087339_(_026861_, _026938_, _026949_);
  or g_087340_(_026872_, _026927_, _026960_);
  and g_087341_(_026641_, _026707_, _026971_);
  or g_087342_(_026652_, _026718_, _026982_);
  and g_087343_(_026960_, _026982_, _026993_);
  or g_087344_(_026949_, _026971_, _027004_);
  xor g_087345_(out[74], _004938_, _027015_);
  not g_087346_(_027015_, _027026_);
  or g_087347_(_009459_, _011615_, _027037_);
  or g_087348_(_005125_, _011626_, _027048_);
  and g_087349_(_027037_, _027048_, _027059_);
  not g_087350_(_027059_, _027070_);
  and g_087351_(_009822_, _011615_, _027081_);
  or g_087352_(_009811_, _011626_, _027092_);
  and g_087353_(_009877_, _011626_, _027103_);
  or g_087354_(_009888_, _011615_, _027114_);
  and g_087355_(_027092_, _027114_, _027125_);
  or g_087356_(_027081_, _027103_, _027136_);
  xor g_087357_(out[73], _004927_, _027147_);
  xor g_087358_(_002936_, _004927_, _027158_);
  and g_087359_(_027125_, _027158_, _027169_);
  or g_087360_(_027136_, _027147_, _027180_);
  or g_087361_(_010878_, _011615_, _027191_);
  not g_087362_(_027191_, _027202_);
  and g_087363_(_010845_, _011615_, _027213_);
  not g_087364_(_027213_, _027224_);
  and g_087365_(_027191_, _027224_, _027235_);
  or g_087366_(_027202_, _027213_, _027246_);
  and g_087367_(_026630_, _027235_, _027257_);
  or g_087368_(_026619_, _027246_, _027268_);
  and g_087369_(_026806_, _026817_, _027279_);
  or g_087370_(_026795_, _026828_, _027290_);
  and g_087371_(_027268_, _027290_, _027301_);
  or g_087372_(_027257_, _027279_, _027312_);
  xor g_087373_(out[72], _004916_, _027323_);
  xor g_087374_(_002925_, _004916_, _027334_);
  and g_087375_(_009701_, _011615_, _027345_);
  or g_087376_(_009712_, _011626_, _027356_);
  and g_087377_(_009778_, _011626_, _027367_);
  or g_087378_(_009767_, _011615_, _027378_);
  and g_087379_(_027356_, _027378_, _027389_);
  or g_087380_(_027345_, _027367_, _027400_);
  and g_087381_(_027334_, _027400_, _027411_);
  or g_087382_(_027323_, _027389_, _027422_);
  and g_087383_(_027136_, _027147_, _027433_);
  or g_087384_(_027125_, _027158_, _027444_);
  and g_087385_(_027323_, _027389_, _027455_);
  or g_087386_(_027334_, _027400_, _027466_);
  and g_087387_(_027444_, _027466_, _027477_);
  or g_087388_(_027433_, _027455_, _027488_);
  and g_087389_(_027015_, _027059_, _027499_);
  and g_087390_(_004971_, _011681_, _027510_);
  and g_087391_(_026872_, _026927_, _027521_);
  or g_087392_(_026861_, _026938_, _027532_);
  xor g_087393_(out[70], _004894_, _027543_);
  not g_087394_(_027543_, _027554_);
  and g_087395_(_010196_, _011615_, _027565_);
  or g_087396_(_010185_, _011626_, _027576_);
  and g_087397_(_010262_, _011626_, _027587_);
  or g_087398_(_010251_, _011615_, _027598_);
  and g_087399_(_027576_, _027598_, _027609_);
  or g_087400_(_027565_, _027587_, _027620_);
  or g_087401_(_027543_, _027620_, _027631_);
  xor g_087402_(_027554_, _027609_, _027642_);
  xor g_087403_(_027543_, _027609_, _027653_);
  xor g_087404_(out[71], _004905_, _027664_);
  not g_087405_(_027664_, _027675_);
  or g_087406_(_009998_, _011626_, _027686_);
  or g_087407_(_010053_, _011615_, _027697_);
  and g_087408_(_027686_, _027697_, _027708_);
  not g_087409_(_027708_, _027719_);
  or g_087410_(_027664_, _027708_, _027730_);
  and g_087411_(_027664_, _027708_, _027741_);
  or g_087412_(_004971_, _011681_, _027752_);
  xor g_087413_(_026630_, _027235_, _027763_);
  xor g_087414_(_026619_, _027235_, _027774_);
  xor g_087415_(_027015_, _027059_, _027785_);
  xor g_087416_(_027026_, _027059_, _027796_);
  xor g_087417_(_004971_, _011681_, _027807_);
  xor g_087418_(_004960_, _011681_, _027818_);
  and g_087419_(_027785_, _027807_, _027829_);
  or g_087420_(_027796_, _027818_, _027840_);
  and g_087421_(_027422_, _027477_, _027851_);
  or g_087422_(_027411_, _027488_, _027862_);
  and g_087423_(_027180_, _027851_, _027873_);
  or g_087424_(_027169_, _027862_, _027884_);
  and g_087425_(_027829_, _027873_, _027895_);
  or g_087426_(_027840_, _027884_, _027906_);
  xor g_087427_(_027664_, _027708_, _027917_);
  xor g_087428_(_027675_, _027708_, _027928_);
  and g_087429_(_027642_, _027917_, _027939_);
  or g_087430_(_027653_, _027928_, _027950_);
  and g_087431_(_027532_, _027939_, _027961_);
  or g_087432_(_027521_, _027950_, _027972_);
  and g_087433_(_026740_, _026993_, _027983_);
  or g_087434_(_026729_, _027004_, _027994_);
  and g_087435_(_027961_, _027983_, _028005_);
  or g_087436_(_027972_, _027994_, _028016_);
  and g_087437_(_027895_, _028005_, _028027_);
  or g_087438_(_027906_, _028016_, _028038_);
  and g_087439_(_026850_, _027290_, _028049_);
  or g_087440_(_026839_, _027279_, _028060_);
  and g_087441_(_028027_, _028049_, _028071_);
  or g_087442_(_028038_, _028060_, _028082_);
  and g_087443_(_027763_, _028071_, _028093_);
  or g_087444_(_027774_, _028082_, _028104_);
  or g_087445_(_002749_, _011626_, _028115_);
  or g_087446_(_011010_, _011615_, _028126_);
  and g_087447_(_028115_, _028126_, _028137_);
  and g_087448_(out[65], _028137_, _028148_);
  not g_087449_(_028148_, _028159_);
  and g_087450_(_028093_, _028148_, _028170_);
  or g_087451_(_028104_, _028159_, _028181_);
  and g_087452_(_027631_, _027730_, _028192_);
  and g_087453_(_027004_, _027961_, _028203_);
  or g_087454_(_026993_, _027972_, _028214_);
  or g_087455_(_027741_, _028192_, _028225_);
  not g_087456_(_028225_, _028236_);
  and g_087457_(_028214_, _028225_, _028247_);
  or g_087458_(_028203_, _028236_, _028258_);
  and g_087459_(_027895_, _028258_, _028269_);
  or g_087460_(_027906_, _028247_, _028280_);
  and g_087461_(_027499_, _027752_, _028291_);
  or g_087462_(_027510_, _028291_, _028302_);
  not g_087463_(_028302_, _028313_);
  and g_087464_(_028280_, _028313_, _028324_);
  or g_087465_(_028269_, _028302_, _028335_);
  or g_087466_(_026839_, _027301_, _028346_);
  and g_087467_(_026850_, _027312_, _028357_);
  and g_087468_(_028027_, _028357_, _028368_);
  or g_087469_(_028038_, _028346_, _028379_);
  and g_087470_(_027488_, _027829_, _028390_);
  or g_087471_(_027477_, _027840_, _028401_);
  and g_087472_(_027180_, _028390_, _028412_);
  or g_087473_(_027169_, _028401_, _028423_);
  and g_087474_(_028379_, _028423_, _028434_);
  or g_087475_(_028368_, _028412_, _028445_);
  or g_087476_(_028335_, _028445_, _028456_);
  and g_087477_(_028324_, _028434_, _028467_);
  and g_087478_(_028181_, _028467_, _028478_);
  or g_087479_(_028170_, _028456_, _028489_);
  or g_087480_(_011087_, _011615_, _028500_);
  not g_087481_(_028500_, _028511_);
  and g_087482_(_002760_, _011615_, _028522_);
  not g_087483_(_028522_, _028533_);
  and g_087484_(_028500_, _028533_, _028544_);
  or g_087485_(_028511_, _028522_, _028555_);
  and g_087486_(out[64], _028555_, _028566_);
  or g_087487_(_002892_, _028544_, _028577_);
  xor g_087488_(out[65], _028137_, _028588_);
  xor g_087489_(_002881_, _028137_, _028599_);
  and g_087490_(_028577_, _028588_, _028610_);
  or g_087491_(_028566_, _028599_, _028621_);
  and g_087492_(_028093_, _028610_, _028632_);
  or g_087493_(_028104_, _028621_, _028643_);
  and g_087494_(_002892_, _028544_, _028654_);
  or g_087495_(out[64], _028555_, _028665_);
  and g_087496_(_028632_, _028654_, _028676_);
  or g_087497_(_028643_, _028665_, _028687_);
  and g_087498_(_028478_, _028687_, _028698_);
  or g_087499_(_028489_, _028676_, _028709_);
  and g_087500_(_026630_, _028709_, _028720_);
  not g_087501_(_028720_, _028731_);
  or g_087502_(_027235_, _028709_, _028742_);
  not g_087503_(_028742_, _028753_);
  and g_087504_(_028731_, _028742_, _028764_);
  or g_087505_(_028720_, _028753_, _028775_);
  and g_087506_(_026597_, _028764_, _028786_);
  or g_087507_(_026586_, _028775_, _028797_);
  or g_087508_(_026795_, _028709_, _028808_);
  not g_087509_(_028808_, _028819_);
  and g_087510_(_026828_, _028709_, _028830_);
  not g_087511_(_028830_, _028841_);
  and g_087512_(_028808_, _028841_, _028852_);
  or g_087513_(_028819_, _028830_, _028863_);
  xor g_087514_(out[83], _011725_, _028874_);
  xor g_087515_(_003046_, _011725_, _028885_);
  and g_087516_(_028863_, _028874_, _028896_);
  or g_087517_(_028852_, _028885_, _028907_);
  and g_087518_(_028797_, _028907_, _028918_);
  or g_087519_(_028786_, _028896_, _028929_);
  or g_087520_(_028137_, _028709_, _028940_);
  or g_087521_(_002881_, _028698_, _028951_);
  and g_087522_(_028940_, _028951_, _028962_);
  and g_087523_(out[81], _028962_, _028973_);
  not g_087524_(_028973_, _028984_);
  and g_087525_(out[64], _028489_, _028995_);
  not g_087526_(_028995_, _029006_);
  or g_087527_(_028555_, _028709_, _029017_);
  not g_087528_(_029017_, _029028_);
  and g_087529_(_029006_, _029017_, _029039_);
  or g_087530_(_028995_, _029028_, _029050_);
  and g_087531_(out[80], _029039_, _029061_);
  or g_087532_(_003024_, _029050_, _029072_);
  xor g_087533_(out[81], _028962_, _029083_);
  xor g_087534_(_003013_, _028962_, _029094_);
  and g_087535_(_029072_, _029083_, _029105_);
  or g_087536_(_029061_, _029094_, _029116_);
  and g_087537_(_028984_, _029116_, _029127_);
  or g_087538_(_028973_, _029105_, _029138_);
  xor g_087539_(_026597_, _028764_, _029149_);
  xor g_087540_(_026586_, _028764_, _029160_);
  or g_087541_(_029127_, _029160_, _029171_);
  and g_087542_(_028918_, _029171_, _029182_);
  and g_087543_(_028852_, _028885_, _029193_);
  or g_087544_(_028863_, _028874_, _029204_);
  and g_087545_(_011703_, _011846_, _029215_);
  or g_087546_(_011714_, _011835_, _029226_);
  xor g_087547_(out[90], _011813_, _029237_);
  xor g_087548_(_003079_, _011813_, _029248_);
  and g_087549_(_027070_, _028698_, _029259_);
  or g_087550_(_027059_, _028709_, _029270_);
  and g_087551_(_027015_, _028709_, _029281_);
  or g_087552_(_027026_, _028698_, _029292_);
  and g_087553_(_029270_, _029292_, _029303_);
  or g_087554_(_029259_, _029281_, _029314_);
  and g_087555_(_029237_, _029303_, _029325_);
  or g_087556_(_029248_, _029314_, _029336_);
  and g_087557_(_029226_, _029336_, _029347_);
  or g_087558_(_029215_, _029325_, _029358_);
  and g_087559_(_029248_, _029314_, _029369_);
  or g_087560_(_029237_, _029303_, _029380_);
  and g_087561_(_011714_, _011835_, _029391_);
  or g_087562_(_011703_, _011846_, _029402_);
  and g_087563_(_029380_, _029402_, _029413_);
  or g_087564_(_029369_, _029391_, _029424_);
  and g_087565_(_029347_, _029413_, _029435_);
  or g_087566_(_029358_, _029424_, _029446_);
  xor g_087567_(out[88], _011791_, _029457_);
  xor g_087568_(_003057_, _011791_, _029468_);
  and g_087569_(_027323_, _028709_, _029479_);
  not g_087570_(_029479_, _029490_);
  or g_087571_(_027389_, _028709_, _029501_);
  not g_087572_(_029501_, _029512_);
  and g_087573_(_029490_, _029501_, _029523_);
  or g_087574_(_029479_, _029512_, _029534_);
  and g_087575_(_029457_, _029523_, _029545_);
  or g_087576_(_029468_, _029534_, _029556_);
  xor g_087577_(out[89], _011802_, _029567_);
  xor g_087578_(_003068_, _011802_, _029578_);
  and g_087579_(_027158_, _028709_, _029589_);
  not g_087580_(_029589_, _029600_);
  or g_087581_(_027125_, _028709_, _029611_);
  not g_087582_(_029611_, _029622_);
  and g_087583_(_029600_, _029611_, _029633_);
  or g_087584_(_029589_, _029622_, _029644_);
  and g_087585_(_029567_, _029644_, _029655_);
  or g_087586_(_029578_, _029633_, _029666_);
  and g_087587_(_029556_, _029666_, _029677_);
  or g_087588_(_029545_, _029655_, _029688_);
  and g_087589_(_029578_, _029633_, _029699_);
  or g_087590_(_029567_, _029644_, _029710_);
  and g_087591_(_029468_, _029534_, _029721_);
  or g_087592_(_029457_, _029523_, _029732_);
  and g_087593_(_029710_, _029732_, _029743_);
  or g_087594_(_029699_, _029721_, _029754_);
  and g_087595_(_029677_, _029743_, _029765_);
  or g_087596_(_029688_, _029754_, _029776_);
  and g_087597_(_029435_, _029765_, _029787_);
  or g_087598_(_029446_, _029776_, _029798_);
  xor g_087599_(out[85], _011758_, _029809_);
  xor g_087600_(_002991_, _011758_, _029820_);
  and g_087601_(_026872_, _028709_, _029831_);
  or g_087602_(_026861_, _028698_, _029842_);
  and g_087603_(_026938_, _028698_, _029853_);
  or g_087604_(_026927_, _028709_, _029864_);
  and g_087605_(_029842_, _029864_, _029875_);
  or g_087606_(_029831_, _029853_, _029886_);
  and g_087607_(_029820_, _029875_, _029897_);
  or g_087608_(_029809_, _029886_, _029908_);
  xor g_087609_(out[86], _011769_, _029919_);
  xor g_087610_(_002980_, _011769_, _029930_);
  and g_087611_(_027554_, _028709_, _029941_);
  or g_087612_(_027543_, _028698_, _029952_);
  and g_087613_(_027620_, _028698_, _029963_);
  or g_087614_(_027609_, _028709_, _029974_);
  and g_087615_(_029952_, _029974_, _029985_);
  or g_087616_(_029941_, _029963_, _029996_);
  and g_087617_(_029919_, _029996_, _030007_);
  or g_087618_(_029930_, _029985_, _030018_);
  and g_087619_(_029908_, _030018_, _030029_);
  or g_087620_(_029897_, _030007_, _030040_);
  xor g_087621_(out[87], _011780_, _030051_);
  xor g_087622_(_002969_, _011780_, _030062_);
  and g_087623_(_027664_, _028709_, _030073_);
  or g_087624_(_027675_, _028698_, _030084_);
  and g_087625_(_027719_, _028698_, _030095_);
  or g_087626_(_027708_, _028709_, _030106_);
  and g_087627_(_030084_, _030106_, _030117_);
  or g_087628_(_030073_, _030095_, _030128_);
  and g_087629_(_030051_, _030117_, _030139_);
  or g_087630_(_030062_, _030128_, _030150_);
  and g_087631_(_026718_, _028698_, _030161_);
  or g_087632_(_026707_, _028709_, _030172_);
  and g_087633_(_026641_, _028709_, _030183_);
  or g_087634_(_026652_, _028698_, _030194_);
  and g_087635_(_030172_, _030194_, _030205_);
  or g_087636_(_030161_, _030183_, _030216_);
  and g_087637_(_026564_, _030216_, _030227_);
  or g_087638_(_026553_, _030205_, _030238_);
  and g_087639_(_030150_, _030238_, _030249_);
  or g_087640_(_030139_, _030227_, _030260_);
  and g_087641_(_030029_, _030249_, _030271_);
  or g_087642_(_030040_, _030260_, _030282_);
  and g_087643_(_029930_, _029985_, _030293_);
  or g_087644_(_029919_, _029996_, _030304_);
  and g_087645_(_030062_, _030128_, _030315_);
  or g_087646_(_030051_, _030117_, _030326_);
  and g_087647_(_030304_, _030326_, _030337_);
  or g_087648_(_030293_, _030315_, _030348_);
  and g_087649_(_026553_, _030205_, _030359_);
  or g_087650_(_026564_, _030216_, _030370_);
  and g_087651_(_029809_, _029886_, _030381_);
  or g_087652_(_029820_, _029875_, _030392_);
  and g_087653_(_030370_, _030392_, _030403_);
  or g_087654_(_030359_, _030381_, _030414_);
  and g_087655_(_030337_, _030403_, _030425_);
  or g_087656_(_030348_, _030414_, _030436_);
  and g_087657_(_030271_, _030425_, _030447_);
  or g_087658_(_030282_, _030436_, _030458_);
  and g_087659_(_029787_, _030447_, _030469_);
  or g_087660_(_029798_, _030458_, _030480_);
  or g_087661_(_029193_, _030480_, _030491_);
  and g_087662_(_028907_, _029204_, _030502_);
  and g_087663_(_029149_, _030502_, _030513_);
  and g_087664_(_029138_, _030513_, _030524_);
  and g_087665_(_028929_, _029204_, _030535_);
  or g_087666_(_030524_, _030535_, _030546_);
  and g_087667_(_030469_, _030546_, _030557_);
  or g_087668_(_029182_, _030491_, _030568_);
  and g_087669_(_030029_, _030414_, _030579_);
  or g_087670_(_030040_, _030403_, _030590_);
  and g_087671_(_030337_, _030590_, _030601_);
  or g_087672_(_030348_, _030579_, _030612_);
  and g_087673_(_030150_, _030612_, _030623_);
  or g_087674_(_030139_, _030601_, _030634_);
  and g_087675_(_029787_, _030623_, _030645_);
  or g_087676_(_029798_, _030634_, _030656_);
  and g_087677_(_029435_, _029688_, _030667_);
  or g_087678_(_029446_, _029677_, _030678_);
  and g_087679_(_029710_, _030667_, _030689_);
  or g_087680_(_029699_, _030678_, _030700_);
  and g_087681_(_029358_, _029402_, _030711_);
  or g_087682_(_029347_, _029391_, _030722_);
  and g_087683_(_030700_, _030722_, _030733_);
  or g_087684_(_030689_, _030711_, _030744_);
  and g_087685_(_030656_, _030733_, _030755_);
  or g_087686_(_030645_, _030744_, _030766_);
  and g_087687_(_030568_, _030755_, _030777_);
  or g_087688_(_030557_, _030766_, _030788_);
  or g_087689_(out[80], _029039_, _030799_);
  and g_087690_(_029105_, _030799_, _030810_);
  and g_087691_(_029787_, _030513_, _030821_);
  and g_087692_(_030447_, _030821_, _030832_);
  and g_087693_(_030810_, _030832_, _030843_);
  not g_087694_(_030843_, _030854_);
  and g_087695_(_030788_, _030854_, _030865_);
  or g_087696_(_030777_, _030843_, _030876_);
  and g_087697_(_026553_, _030865_, _030887_);
  or g_087698_(_026564_, _030876_, _030898_);
  and g_087699_(_030216_, _030876_, _030909_);
  or g_087700_(_030205_, _030865_, _030920_);
  and g_087701_(_030898_, _030920_, _030931_);
  or g_087702_(_030887_, _030909_, _030942_);
  and g_087703_(_026531_, _030931_, _030953_);
  or g_087704_(_026542_, _030942_, _030964_);
  xor g_087705_(out[101], _011912_, _030975_);
  xor g_087706_(_003123_, _011912_, _030986_);
  and g_087707_(_029820_, _030865_, _030997_);
  or g_087708_(_029809_, _030876_, _031008_);
  and g_087709_(_029886_, _030876_, _031019_);
  or g_087710_(_029875_, _030865_, _031030_);
  and g_087711_(_031008_, _031030_, _031041_);
  or g_087712_(_030997_, _031019_, _031052_);
  and g_087713_(_030975_, _031052_, _031063_);
  or g_087714_(_030986_, _031041_, _031074_);
  and g_087715_(_030964_, _031074_, _031085_);
  or g_087716_(_030953_, _031063_, _031096_);
  and g_087717_(_028863_, _030876_, _031107_);
  or g_087718_(_028852_, _030865_, _031118_);
  and g_087719_(_028885_, _030865_, _031129_);
  or g_087720_(_028874_, _030876_, _031140_);
  and g_087721_(_031118_, _031140_, _031151_);
  or g_087722_(_031107_, _031129_, _031162_);
  xor g_087723_(out[99], _011879_, _031173_);
  and g_087724_(_031162_, _031173_, _031184_);
  or g_087725_(out[97], out[98], _031195_);
  xor g_087726_(out[97], out[98], _031206_);
  xor g_087727_(_003145_, out[98], _031217_);
  or g_087728_(_028764_, _030865_, _031228_);
  or g_087729_(_026586_, _030876_, _031239_);
  and g_087730_(_031228_, _031239_, _031250_);
  and g_087731_(_031217_, _031250_, _031261_);
  or g_087732_(_031184_, _031261_, _031272_);
  or g_087733_(_031162_, _031173_, _031283_);
  xor g_087734_(_031162_, _031173_, _031294_);
  xor g_087735_(_031151_, _031173_, _031305_);
  xor g_087736_(_031217_, _031250_, _031316_);
  xor g_087737_(_031206_, _031250_, _031327_);
  and g_087738_(_031294_, _031316_, _031338_);
  or g_087739_(_031305_, _031327_, _031349_);
  or g_087740_(_003013_, _030876_, _031360_);
  or g_087741_(_028962_, _030865_, _031371_);
  and g_087742_(_031360_, _031371_, _031382_);
  and g_087743_(out[97], _031382_, _031393_);
  not g_087744_(_031393_, _031404_);
  and g_087745_(_029039_, _030876_, _031415_);
  or g_087746_(_029050_, _030865_, _031426_);
  and g_087747_(_003024_, _030865_, _031437_);
  or g_087748_(out[80], _030876_, _031448_);
  and g_087749_(_031426_, _031448_, _031459_);
  or g_087750_(_031415_, _031437_, _031470_);
  and g_087751_(out[96], _031470_, _031481_);
  or g_087752_(_003156_, _031459_, _031492_);
  xor g_087753_(out[97], _031382_, _031503_);
  xor g_087754_(_003145_, _031382_, _031514_);
  and g_087755_(_031492_, _031503_, _031525_);
  or g_087756_(_031481_, _031514_, _031536_);
  and g_087757_(_031404_, _031536_, _031547_);
  or g_087758_(_031393_, _031525_, _031558_);
  and g_087759_(_031338_, _031558_, _031569_);
  or g_087760_(_031349_, _031547_, _031580_);
  and g_087761_(_031272_, _031283_, _031591_);
  not g_087762_(_031591_, _031602_);
  and g_087763_(_031580_, _031602_, _031613_);
  or g_087764_(_031569_, _031591_, _031624_);
  and g_087765_(_026542_, _030942_, _031635_);
  or g_087766_(_026531_, _030931_, _031646_);
  and g_087767_(_031624_, _031646_, _031657_);
  or g_087768_(_031613_, _031635_, _031668_);
  and g_087769_(_031085_, _031668_, _031679_);
  or g_087770_(_031096_, _031657_, _031690_);
  and g_087771_(_029314_, _030876_, _031701_);
  or g_087772_(_029303_, _030865_, _031712_);
  and g_087773_(_029237_, _030865_, _031723_);
  or g_087774_(_029248_, _030876_, _031734_);
  and g_087775_(_031712_, _031734_, _031745_);
  or g_087776_(_031701_, _031723_, _031756_);
  and g_087777_(_026520_, _031745_, _031767_);
  and g_087778_(_011857_, _011989_, _031778_);
  or g_087779_(_031767_, _031778_, _031789_);
  xor g_087780_(out[105], _011956_, _031800_);
  xor g_087781_(_003200_, _011956_, _031811_);
  and g_087782_(_029578_, _030865_, _031822_);
  or g_087783_(_029567_, _030876_, _031833_);
  and g_087784_(_029644_, _030876_, _031844_);
  or g_087785_(_029633_, _030865_, _031855_);
  and g_087786_(_031833_, _031855_, _031866_);
  or g_087787_(_031822_, _031844_, _031877_);
  and g_087788_(_031811_, _031866_, _031888_);
  or g_087789_(_031800_, _031877_, _031899_);
  or g_087790_(_011857_, _011989_, _031910_);
  xor g_087791_(_026520_, _031745_, _031921_);
  xor g_087792_(_026520_, _031756_, _031932_);
  xor g_087793_(_011868_, _012000_, _031943_);
  xor g_087794_(_011857_, _012000_, _031954_);
  and g_087795_(_031921_, _031943_, _031965_);
  or g_087796_(_031932_, _031954_, _031976_);
  and g_087797_(_031899_, _031965_, _031987_);
  or g_087798_(_031888_, _031976_, _031998_);
  and g_087799_(_031800_, _031877_, _032009_);
  or g_087800_(_031811_, _031866_, _032020_);
  xor g_087801_(out[104], _011945_, _032031_);
  xor g_087802_(_003189_, _011945_, _032042_);
  and g_087803_(_029457_, _030865_, _032053_);
  or g_087804_(_029468_, _030876_, _032064_);
  and g_087805_(_029534_, _030876_, _032075_);
  or g_087806_(_029523_, _030865_, _032086_);
  and g_087807_(_032064_, _032086_, _032097_);
  or g_087808_(_032053_, _032075_, _032108_);
  and g_087809_(_032031_, _032097_, _032119_);
  or g_087810_(_032042_, _032108_, _032130_);
  and g_087811_(_032020_, _032130_, _032141_);
  or g_087812_(_032009_, _032119_, _032152_);
  and g_087813_(_032042_, _032108_, _032163_);
  or g_087814_(_032031_, _032097_, _032174_);
  and g_087815_(_032141_, _032174_, _032185_);
  or g_087816_(_032152_, _032163_, _032196_);
  and g_087817_(_031987_, _032185_, _032207_);
  or g_087818_(_031998_, _032196_, _032218_);
  xor g_087819_(out[102], _011923_, _032229_);
  xor g_087820_(_003112_, _011923_, _032240_);
  and g_087821_(_029930_, _030865_, _032251_);
  or g_087822_(_029919_, _030876_, _032262_);
  and g_087823_(_029996_, _030876_, _032273_);
  not g_087824_(_032273_, _032284_);
  and g_087825_(_032262_, _032284_, _032295_);
  or g_087826_(_032251_, _032273_, _032306_);
  and g_087827_(_032240_, _032295_, _032317_);
  or g_087828_(_032229_, _032306_, _032328_);
  xor g_087829_(out[103], _011934_, _032339_);
  xor g_087830_(_003101_, _011934_, _032350_);
  or g_087831_(_030062_, _030876_, _032361_);
  or g_087832_(_030117_, _030865_, _032372_);
  and g_087833_(_032361_, _032372_, _032383_);
  not g_087834_(_032383_, _032394_);
  and g_087835_(_032350_, _032394_, _032405_);
  or g_087836_(_032339_, _032383_, _032416_);
  and g_087837_(_032328_, _032416_, _032427_);
  or g_087838_(_032317_, _032405_, _032438_);
  and g_087839_(_030986_, _031041_, _032449_);
  or g_087840_(_030975_, _031052_, _032460_);
  and g_087841_(_032339_, _032383_, _032471_);
  or g_087842_(_032350_, _032394_, _032482_);
  and g_087843_(_032229_, _032306_, _032493_);
  or g_087844_(_032240_, _032295_, _032504_);
  and g_087845_(_032460_, _032482_, _032515_);
  or g_087846_(_032449_, _032471_, _032526_);
  or g_087847_(_032493_, _032526_, _032537_);
  and g_087848_(_032427_, _032504_, _032548_);
  and g_087849_(_032515_, _032548_, _032559_);
  or g_087850_(_032438_, _032537_, _032570_);
  and g_087851_(_032207_, _032559_, _032581_);
  or g_087852_(_032218_, _032570_, _032592_);
  and g_087853_(_031690_, _032581_, _032603_);
  or g_087854_(_031679_, _032592_, _032614_);
  and g_087855_(_031987_, _032152_, _032625_);
  and g_087856_(_031789_, _031910_, _032636_);
  or g_087857_(_032625_, _032636_, _032647_);
  not g_087858_(_032647_, _032658_);
  and g_087859_(_032438_, _032482_, _032669_);
  or g_087860_(_032427_, _032471_, _032680_);
  and g_087861_(_032207_, _032669_, _032691_);
  or g_087862_(_032218_, _032680_, _032702_);
  and g_087863_(_032658_, _032702_, _032713_);
  or g_087864_(_032647_, _032691_, _032724_);
  and g_087865_(_032614_, _032713_, _032735_);
  or g_087866_(_032603_, _032724_, _032746_);
  and g_087867_(_003156_, _031459_, _032757_);
  or g_087868_(out[96], _031470_, _032768_);
  and g_087869_(_031646_, _032768_, _032779_);
  or g_087870_(_031635_, _032757_, _032790_);
  and g_087871_(_031085_, _032779_, _032801_);
  or g_087872_(_031096_, _032790_, _032812_);
  and g_087873_(_031338_, _032801_, _032823_);
  or g_087874_(_031349_, _032812_, _032834_);
  and g_087875_(_031525_, _032823_, _032845_);
  or g_087876_(_031536_, _032834_, _032856_);
  and g_087877_(_032581_, _032845_, _032867_);
  or g_087878_(_032592_, _032856_, _032878_);
  and g_087879_(_032746_, _032878_, _032889_);
  or g_087880_(_032735_, _032867_, _032900_);
  and g_087881_(_026520_, _032889_, _032911_);
  not g_087882_(_032911_, _032922_);
  and g_087883_(_031756_, _032900_, _032933_);
  or g_087884_(_031745_, _032889_, _032944_);
  and g_087885_(_032922_, _032944_, _032955_);
  or g_087886_(_032911_, _032933_, _032966_);
  and g_087887_(_012011_, _012154_, _032977_);
  or g_087888_(_012022_, _012143_, _032988_);
  xor g_087889_(out[122], _012121_, _032999_);
  xor g_087890_(_003343_, _012121_, _033010_);
  and g_087891_(_032955_, _032999_, _033021_);
  or g_087892_(_032966_, _033010_, _033032_);
  and g_087893_(_032988_, _033032_, _033043_);
  or g_087894_(_032977_, _033021_, _033054_);
  and g_087895_(_012022_, _012143_, _033065_);
  or g_087896_(_012011_, _012154_, _033076_);
  and g_087897_(_032966_, _033010_, _033087_);
  or g_087898_(_032955_, _032999_, _033098_);
  and g_087899_(_033076_, _033098_, _033109_);
  or g_087900_(_033065_, _033087_, _033120_);
  xor g_087901_(out[121], _012110_, _033131_);
  xor g_087902_(_003332_, _012110_, _033142_);
  and g_087903_(_031877_, _032900_, _033153_);
  or g_087904_(_031866_, _032889_, _033164_);
  and g_087905_(_031811_, _032889_, _033175_);
  or g_087906_(_031800_, _032900_, _033186_);
  and g_087907_(_033164_, _033186_, _033197_);
  or g_087908_(_033153_, _033175_, _033208_);
  and g_087909_(_033142_, _033197_, _033219_);
  or g_087910_(_033131_, _033208_, _033230_);
  xor g_087911_(out[120], _012099_, _033241_);
  xor g_087912_(_003321_, _012099_, _033252_);
  and g_087913_(_032108_, _032900_, _033263_);
  or g_087914_(_032097_, _032889_, _033274_);
  and g_087915_(_032031_, _032889_, _033285_);
  or g_087916_(_032042_, _032900_, _033296_);
  and g_087917_(_033274_, _033296_, _033307_);
  or g_087918_(_033263_, _033285_, _033318_);
  and g_087919_(_033252_, _033318_, _033329_);
  or g_087920_(_033241_, _033307_, _033340_);
  and g_087921_(_033131_, _033208_, _033351_);
  or g_087922_(_033142_, _033197_, _033362_);
  and g_087923_(_033241_, _033307_, _033373_);
  or g_087924_(_033252_, _033318_, _033384_);
  and g_087925_(_033362_, _033384_, _033395_);
  or g_087926_(_033351_, _033373_, _033406_);
  and g_087927_(_033230_, _033395_, _033417_);
  or g_087928_(_033219_, _033406_, _033428_);
  and g_087929_(_033043_, _033109_, _033439_);
  or g_087930_(_033054_, _033120_, _033450_);
  and g_087931_(_033340_, _033439_, _033461_);
  or g_087932_(_033329_, _033450_, _033472_);
  and g_087933_(_033417_, _033461_, _033483_);
  or g_087934_(_033428_, _033472_, _033494_);
  xor g_087935_(out[118], _012077_, _033505_);
  not g_087936_(_033505_, _033516_);
  and g_087937_(_032306_, _032900_, _033527_);
  or g_087938_(_032295_, _032889_, _033538_);
  and g_087939_(_032240_, _032889_, _033549_);
  or g_087940_(_032229_, _032900_, _033560_);
  and g_087941_(_033538_, _033560_, _033571_);
  or g_087942_(_033527_, _033549_, _033582_);
  or g_087943_(_033505_, _033582_, _033593_);
  xor g_087944_(out[119], _012088_, _033604_);
  not g_087945_(_033604_, _033615_);
  or g_087946_(_032383_, _032889_, _033626_);
  or g_087947_(_032350_, _032900_, _033637_);
  and g_087948_(_033626_, _033637_, _033648_);
  or g_087949_(_033604_, _033648_, _033659_);
  and g_087950_(_033593_, _033659_, _033670_);
  and g_087951_(_033604_, _033648_, _033681_);
  xor g_087952_(out[117], _012066_, _033692_);
  xor g_087953_(_003255_, _012066_, _033703_);
  and g_087954_(_031052_, _032900_, _033714_);
  or g_087955_(_031041_, _032889_, _033725_);
  and g_087956_(_030986_, _032889_, _033736_);
  or g_087957_(_030975_, _032900_, _033747_);
  and g_087958_(_033725_, _033747_, _033758_);
  or g_087959_(_033714_, _033736_, _033769_);
  and g_087960_(_033703_, _033758_, _033780_);
  xor g_087961_(_033505_, _033571_, _033791_);
  xor g_087962_(_033615_, _033648_, _033802_);
  or g_087963_(_033791_, _033802_, _033813_);
  or g_087964_(_033780_, _033813_, _033824_);
  not g_087965_(_033824_, _033835_);
  xor g_087966_(out[116], _012055_, _033846_);
  xor g_087967_(_003266_, _012055_, _033857_);
  and g_087968_(_026531_, _032889_, _033868_);
  or g_087969_(_026542_, _032900_, _033879_);
  and g_087970_(_030942_, _032900_, _033890_);
  or g_087971_(_030931_, _032889_, _033901_);
  and g_087972_(_033879_, _033901_, _033912_);
  or g_087973_(_033868_, _033890_, _033923_);
  or g_087974_(_033846_, _033912_, _033934_);
  or g_087975_(_033703_, _033758_, _033945_);
  or g_087976_(_033857_, _033923_, _033956_);
  and g_087977_(_033945_, _033956_, _033967_);
  and g_087978_(_033934_, _033967_, _033978_);
  not g_087979_(_033978_, _033989_);
  and g_087980_(_033835_, _033978_, _034000_);
  or g_087981_(_033824_, _033989_, _034011_);
  or g_087982_(_031151_, _032889_, _034022_);
  or g_087983_(_031173_, _032900_, _034033_);
  and g_087984_(_034022_, _034033_, _034044_);
  not g_087985_(_034044_, _034055_);
  xor g_087986_(out[115], _012033_, _034066_);
  xor g_087987_(_003310_, _012033_, _034077_);
  and g_087988_(_034055_, _034066_, _034088_);
  or g_087989_(_034044_, _034077_, _034099_);
  or g_087990_(out[113], out[114], _034110_);
  xor g_087991_(out[113], out[114], _034121_);
  xor g_087992_(_003277_, out[114], _034132_);
  or g_087993_(_031250_, _032889_, _034143_);
  or g_087994_(_031206_, _032900_, _034154_);
  and g_087995_(_034143_, _034154_, _034165_);
  not g_087996_(_034165_, _034176_);
  and g_087997_(_034132_, _034165_, _034187_);
  or g_087998_(_034121_, _034176_, _034198_);
  and g_087999_(_034099_, _034198_, _034209_);
  or g_088000_(_034088_, _034187_, _034220_);
  and g_088001_(_034044_, _034077_, _034231_);
  or g_088002_(_034055_, _034066_, _034242_);
  and g_088003_(_034121_, _034176_, _034253_);
  or g_088004_(_034132_, _034165_, _034264_);
  and g_088005_(_034242_, _034264_, _034275_);
  or g_088006_(_034231_, _034253_, _034286_);
  and g_088007_(_034209_, _034275_, _034297_);
  or g_088008_(_034220_, _034286_, _034308_);
  or g_088009_(_003145_, _032900_, _034319_);
  or g_088010_(_031382_, _032889_, _034330_);
  and g_088011_(_034319_, _034330_, _034341_);
  and g_088012_(out[113], _034341_, _034352_);
  not g_088013_(_034352_, _034363_);
  and g_088014_(_031470_, _032900_, _034374_);
  or g_088015_(_031459_, _032889_, _034385_);
  and g_088016_(_003156_, _032889_, _034396_);
  or g_088017_(out[96], _032900_, _034407_);
  and g_088018_(_034385_, _034407_, _034418_);
  or g_088019_(_034374_, _034396_, _034429_);
  and g_088020_(out[112], _034429_, _034440_);
  or g_088021_(_003288_, _034418_, _034451_);
  xor g_088022_(out[113], _034341_, _034462_);
  xor g_088023_(_003277_, _034341_, _034473_);
  and g_088024_(_034451_, _034462_, _034484_);
  or g_088025_(_034440_, _034473_, _034495_);
  and g_088026_(_034363_, _034495_, _034506_);
  or g_088027_(_034352_, _034484_, _034517_);
  and g_088028_(_034297_, _034517_, _034528_);
  or g_088029_(_034308_, _034506_, _034539_);
  and g_088030_(_034220_, _034242_, _034550_);
  or g_088031_(_034209_, _034231_, _034561_);
  and g_088032_(_034539_, _034561_, _034572_);
  or g_088033_(_034528_, _034550_, _034583_);
  and g_088034_(_034000_, _034583_, _034594_);
  or g_088035_(_034011_, _034572_, _034605_);
  or g_088036_(_033824_, _033967_, _034616_);
  or g_088037_(_033670_, _033681_, _034627_);
  and g_088038_(_034616_, _034627_, _034638_);
  not g_088039_(_034638_, _034649_);
  and g_088040_(_034605_, _034638_, _034660_);
  or g_088041_(_034594_, _034649_, _034671_);
  and g_088042_(_033483_, _034671_, _034682_);
  or g_088043_(_033494_, _034660_, _034693_);
  and g_088044_(_033054_, _033076_, _034704_);
  or g_088045_(_033043_, _033065_, _034715_);
  and g_088046_(_033230_, _033406_, _034726_);
  or g_088047_(_033219_, _033395_, _034737_);
  and g_088048_(_033439_, _034726_, _034748_);
  or g_088049_(_033450_, _034737_, _034759_);
  and g_088050_(_034715_, _034759_, _034770_);
  or g_088051_(_034704_, _034748_, _034781_);
  and g_088052_(_034693_, _034770_, _034792_);
  or g_088053_(_034682_, _034781_, _034803_);
  and g_088054_(_003288_, _034418_, _034814_);
  not g_088055_(_034814_, _034825_);
  and g_088056_(_034484_, _034825_, _034836_);
  not g_088057_(_034836_, _034847_);
  and g_088058_(_034297_, _034836_, _034858_);
  or g_088059_(_034308_, _034847_, _034869_);
  and g_088060_(_034000_, _034858_, _034880_);
  or g_088061_(_034011_, _034869_, _034891_);
  and g_088062_(_033483_, _034880_, _034902_);
  or g_088063_(_033494_, _034891_, _034913_);
  and g_088064_(_034803_, _034913_, _034924_);
  or g_088065_(_034792_, _034902_, _034935_);
  or g_088066_(_032955_, _034924_, _034946_);
  not g_088067_(_034946_, _034957_);
  and g_088068_(_032999_, _034924_, _034968_);
  not g_088069_(_034968_, _034979_);
  and g_088070_(_034946_, _034979_, _034990_);
  or g_088071_(_034957_, _034968_, _035001_);
  and g_088072_(_026509_, _035001_, _035012_);
  and g_088073_(_012165_, _012308_, _035023_);
  or g_088074_(_012176_, _012297_, _035034_);
  and g_088075_(_012176_, _012297_, _035045_);
  or g_088076_(_012165_, _012308_, _035056_);
  and g_088077_(_035034_, _035056_, _035067_);
  and g_088078_(_026498_, _034990_, _035078_);
  or g_088079_(_026509_, _035001_, _035089_);
  or g_088080_(_035012_, _035023_, _035100_);
  or g_088081_(_035045_, _035078_, _035111_);
  xor g_088082_(_026498_, _034990_, _035122_);
  and g_088083_(_035067_, _035122_, _035133_);
  or g_088084_(_035100_, _035111_, _035144_);
  xor g_088085_(out[137], _012264_, _035155_);
  xor g_088086_(_003464_, _012264_, _035166_);
  and g_088087_(_033142_, _034924_, _035177_);
  or g_088088_(_033131_, _034935_, _035188_);
  and g_088089_(_033208_, _034935_, _035199_);
  or g_088090_(_033197_, _034924_, _035210_);
  and g_088091_(_035188_, _035210_, _035221_);
  or g_088092_(_035177_, _035199_, _035232_);
  and g_088093_(_035155_, _035232_, _035243_);
  or g_088094_(_035166_, _035221_, _035254_);
  xor g_088095_(out[136], _012253_, _035265_);
  xor g_088096_(_003453_, _012253_, _035276_);
  and g_088097_(_033241_, _034924_, _035287_);
  or g_088098_(_033252_, _034935_, _035298_);
  and g_088099_(_033318_, _034935_, _035309_);
  or g_088100_(_033307_, _034924_, _035320_);
  and g_088101_(_035298_, _035320_, _035331_);
  or g_088102_(_035287_, _035309_, _035342_);
  and g_088103_(_035265_, _035331_, _035353_);
  or g_088104_(_035276_, _035342_, _035364_);
  and g_088105_(_035254_, _035364_, _035375_);
  or g_088106_(_035243_, _035353_, _035386_);
  and g_088107_(_035166_, _035221_, _035397_);
  or g_088108_(_035155_, _035232_, _035408_);
  and g_088109_(_035386_, _035408_, _035419_);
  or g_088110_(_035375_, _035397_, _035430_);
  and g_088111_(_035133_, _035419_, _035441_);
  or g_088112_(_035144_, _035430_, _035452_);
  and g_088113_(_035056_, _035078_, _035463_);
  or g_088114_(_035045_, _035089_, _035474_);
  and g_088115_(_035034_, _035474_, _035485_);
  or g_088116_(_035023_, _035463_, _035496_);
  and g_088117_(_035452_, _035485_, _035507_);
  and g_088118_(_035276_, _035342_, _035518_);
  or g_088119_(_035265_, _035331_, _035529_);
  and g_088120_(_035408_, _035529_, _035540_);
  or g_088121_(_035397_, _035518_, _035551_);
  and g_088122_(_035375_, _035540_, _035562_);
  or g_088123_(_035386_, _035551_, _035573_);
  and g_088124_(_035133_, _035562_, _035584_);
  or g_088125_(_035144_, _035573_, _035595_);
  xor g_088126_(out[135], _012242_, _035606_);
  not g_088127_(_035606_, _035617_);
  or g_088128_(_033615_, _034935_, _035628_);
  or g_088129_(_033648_, _034924_, _035639_);
  and g_088130_(_035628_, _035639_, _035650_);
  not g_088131_(_035650_, _035661_);
  and g_088132_(_035606_, _035650_, _035672_);
  or g_088133_(_035606_, _035650_, _035683_);
  xor g_088134_(out[134], _012231_, _035694_);
  not g_088135_(_035694_, _035705_);
  and g_088136_(_033516_, _034924_, _035716_);
  or g_088137_(_033505_, _034935_, _035727_);
  and g_088138_(_033582_, _034935_, _035738_);
  or g_088139_(_033571_, _034924_, _035749_);
  and g_088140_(_035727_, _035749_, _035760_);
  or g_088141_(_035716_, _035738_, _035771_);
  or g_088142_(_035694_, _035771_, _035782_);
  and g_088143_(_035683_, _035782_, _035793_);
  or g_088144_(_035672_, _035793_, _035804_);
  not g_088145_(_035804_, _035815_);
  xor g_088146_(_035606_, _035650_, _035826_);
  xor g_088147_(_035617_, _035650_, _035837_);
  xor g_088148_(out[133], _012220_, _035848_);
  xor g_088149_(_003387_, _012220_, _035859_);
  and g_088150_(_033703_, _034924_, _035870_);
  or g_088151_(_033692_, _034935_, _035881_);
  and g_088152_(_033769_, _034935_, _035892_);
  or g_088153_(_033758_, _034924_, _035903_);
  and g_088154_(_035881_, _035903_, _035914_);
  or g_088155_(_035870_, _035892_, _035925_);
  and g_088156_(_035859_, _035914_, _035936_);
  or g_088157_(_035848_, _035925_, _035947_);
  xor g_088158_(_035705_, _035760_, _035958_);
  xor g_088159_(_035694_, _035760_, _035969_);
  and g_088160_(_035826_, _035958_, _035980_);
  or g_088161_(_035837_, _035969_, _035991_);
  and g_088162_(_035947_, _035980_, _036002_);
  or g_088163_(_035936_, _035991_, _036013_);
  and g_088164_(_035848_, _035925_, _036024_);
  or g_088165_(_035859_, _035914_, _036035_);
  xor g_088166_(out[132], _012209_, _036046_);
  xor g_088167_(_003398_, _012209_, _036057_);
  and g_088168_(_033846_, _034924_, _036068_);
  or g_088169_(_033857_, _034935_, _036079_);
  and g_088170_(_033923_, _034935_, _036090_);
  or g_088171_(_033912_, _034924_, _036101_);
  and g_088172_(_036079_, _036101_, _036112_);
  or g_088173_(_036068_, _036090_, _036123_);
  and g_088174_(_036046_, _036112_, _036134_);
  or g_088175_(_036057_, _036123_, _036145_);
  and g_088176_(_036035_, _036145_, _036156_);
  or g_088177_(_036024_, _036134_, _036167_);
  or g_088178_(out[129], out[130], _036178_);
  xor g_088179_(out[129], out[130], _036189_);
  xor g_088180_(_003409_, out[130], _036200_);
  or g_088181_(_034165_, _034924_, _036211_);
  not g_088182_(_036211_, _036222_);
  and g_088183_(_034132_, _034924_, _036233_);
  not g_088184_(_036233_, _036244_);
  and g_088185_(_036211_, _036244_, _036255_);
  or g_088186_(_036222_, _036233_, _036266_);
  and g_088187_(_036200_, _036255_, _036277_);
  or g_088188_(_036189_, _036266_, _036288_);
  or g_088189_(_034044_, _034924_, _036299_);
  not g_088190_(_036299_, _036310_);
  and g_088191_(_034077_, _034924_, _036321_);
  not g_088192_(_036321_, _036332_);
  and g_088193_(_036299_, _036332_, _036343_);
  or g_088194_(_036310_, _036321_, _036354_);
  xor g_088195_(out[131], _012187_, _036365_);
  xor g_088196_(_003442_, _012187_, _036376_);
  and g_088197_(_036354_, _036365_, _036387_);
  or g_088198_(_036343_, _036376_, _036398_);
  and g_088199_(_036288_, _036398_, _036409_);
  or g_088200_(_036277_, _036387_, _036420_);
  or g_088201_(_003277_, _034935_, _036431_);
  or g_088202_(_034341_, _034924_, _036442_);
  and g_088203_(_036431_, _036442_, _036453_);
  not g_088204_(_036453_, _036464_);
  or g_088205_(_003409_, _036464_, _036475_);
  not g_088206_(_036475_, _036486_);
  and g_088207_(_036189_, _036266_, _036497_);
  or g_088208_(_036200_, _036255_, _036508_);
  or g_088209_(_036475_, _036497_, _036519_);
  and g_088210_(_036409_, _036519_, _036530_);
  and g_088211_(_036343_, _036376_, _036541_);
  or g_088212_(_036354_, _036365_, _036552_);
  and g_088213_(_036057_, _036123_, _036563_);
  or g_088214_(_036046_, _036112_, _036574_);
  or g_088215_(_036541_, _036563_, _036585_);
  or g_088216_(_036530_, _036585_, _036596_);
  and g_088217_(_036156_, _036596_, _036607_);
  or g_088218_(_036013_, _036607_, _036618_);
  and g_088219_(_035804_, _036618_, _036629_);
  or g_088220_(_035595_, _036629_, _036640_);
  and g_088221_(_036002_, _036167_, _036651_);
  or g_088222_(_035815_, _036651_, _036662_);
  and g_088223_(_035584_, _036662_, _036673_);
  or g_088224_(_035496_, _036673_, _036684_);
  and g_088225_(_036156_, _036574_, _036695_);
  or g_088226_(_036167_, _036563_, _036706_);
  and g_088227_(_036002_, _036695_, _036717_);
  or g_088228_(_036013_, _036706_, _036728_);
  and g_088229_(_035584_, _036717_, _036739_);
  or g_088230_(_035595_, _036728_, _036750_);
  and g_088231_(_036420_, _036552_, _036761_);
  and g_088232_(_036739_, _036761_, _036772_);
  or g_088233_(_035441_, _036772_, _036783_);
  or g_088234_(_036684_, _036783_, _036794_);
  and g_088235_(_036398_, _036552_, _036805_);
  or g_088236_(_036387_, _036541_, _036816_);
  and g_088237_(_036288_, _036805_, _036827_);
  or g_088238_(_036277_, _036816_, _036838_);
  and g_088239_(_036508_, _036739_, _036849_);
  or g_088240_(_036497_, _036750_, _036860_);
  and g_088241_(_036827_, _036849_, _036871_);
  or g_088242_(_036838_, _036860_, _036882_);
  and g_088243_(_036486_, _036871_, _036893_);
  and g_088244_(_035507_, _036640_, _036904_);
  or g_088245_(_036794_, _036893_, _036915_);
  or g_088246_(_034418_, _034924_, _036926_);
  not g_088247_(_036926_, _036937_);
  and g_088248_(_003288_, _034924_, _036948_);
  not g_088249_(_036948_, _036959_);
  and g_088250_(_036926_, _036959_, _036970_);
  or g_088251_(_036937_, _036948_, _036981_);
  and g_088252_(out[128], _036981_, _036992_);
  or g_088253_(_003420_, _036970_, _037003_);
  xor g_088254_(out[129], _036453_, _037014_);
  xor g_088255_(_003409_, _036453_, _037025_);
  and g_088256_(_037003_, _037014_, _037036_);
  or g_088257_(_036992_, _037025_, _037047_);
  and g_088258_(_036871_, _037036_, _037058_);
  or g_088259_(_036882_, _037047_, _037069_);
  and g_088260_(_003420_, _036970_, _037080_);
  or g_088261_(out[128], _036981_, _037091_);
  and g_088262_(_037058_, _037080_, _037102_);
  or g_088263_(_037069_, _037091_, _037113_);
  and g_088264_(_036904_, _037113_, _037124_);
  or g_088265_(_036915_, _037102_, _037135_);
  and g_088266_(_026498_, _037135_, _037146_);
  not g_088267_(_037146_, _037157_);
  and g_088268_(_035001_, _037124_, _037168_);
  or g_088269_(_034990_, _037135_, _037179_);
  and g_088270_(_037157_, _037179_, _037190_);
  or g_088271_(_037146_, _037168_, _037201_);
  and g_088272_(_026454_, _037190_, _037212_);
  or g_088273_(_026465_, _037201_, _037223_);
  and g_088274_(_026487_, _037223_, _037234_);
  or g_088275_(_026476_, _037212_, _037245_);
  and g_088276_(_012330_, _012451_, _037256_);
  or g_088277_(_012319_, _012462_, _037267_);
  and g_088278_(_026465_, _037201_, _037278_);
  or g_088279_(_026454_, _037190_, _037289_);
  and g_088280_(_037267_, _037289_, _037300_);
  or g_088281_(_037256_, _037278_, _037311_);
  and g_088282_(_037234_, _037300_, _037322_);
  or g_088283_(_037245_, _037311_, _037333_);
  xor g_088284_(out[153], _012418_, _037344_);
  xor g_088285_(_003596_, _012418_, _037355_);
  and g_088286_(_035232_, _037124_, _037366_);
  or g_088287_(_035221_, _037135_, _037377_);
  and g_088288_(_035166_, _037135_, _037388_);
  or g_088289_(_035155_, _037124_, _037399_);
  and g_088290_(_037377_, _037399_, _037410_);
  or g_088291_(_037366_, _037388_, _037421_);
  and g_088292_(_037344_, _037421_, _037432_);
  or g_088293_(_037355_, _037410_, _037443_);
  xor g_088294_(out[152], _012407_, _037454_);
  xor g_088295_(_003585_, _012407_, _037465_);
  and g_088296_(_035342_, _037124_, _037476_);
  or g_088297_(_035331_, _037135_, _037487_);
  and g_088298_(_035265_, _037135_, _037498_);
  or g_088299_(_035276_, _037124_, _037509_);
  and g_088300_(_037487_, _037509_, _037520_);
  or g_088301_(_037476_, _037498_, _037531_);
  and g_088302_(_037454_, _037520_, _037542_);
  or g_088303_(_037465_, _037531_, _037553_);
  and g_088304_(_037443_, _037553_, _037564_);
  or g_088305_(_037432_, _037542_, _037575_);
  or g_088306_(_037454_, _037520_, _037586_);
  and g_088307_(_037355_, _037410_, _037597_);
  or g_088308_(_037344_, _037421_, _037608_);
  and g_088309_(_037586_, _037608_, _037619_);
  and g_088310_(_037564_, _037619_, _037630_);
  and g_088311_(_037322_, _037630_, _037641_);
  not g_088312_(_037641_, _037652_);
  xor g_088313_(out[150], _012385_, _037663_);
  not g_088314_(_037663_, _037674_);
  and g_088315_(_035771_, _037124_, _037685_);
  or g_088316_(_035760_, _037135_, _037696_);
  and g_088317_(_035705_, _037135_, _037707_);
  or g_088318_(_035694_, _037124_, _037718_);
  and g_088319_(_037696_, _037718_, _037729_);
  or g_088320_(_037685_, _037707_, _037740_);
  and g_088321_(_037674_, _037729_, _037751_);
  or g_088322_(_037663_, _037740_, _037762_);
  xor g_088323_(out[151], _012396_, _037773_);
  xor g_088324_(_003497_, _012396_, _037784_);
  and g_088325_(_035661_, _037124_, _037795_);
  or g_088326_(_035650_, _037135_, _037806_);
  and g_088327_(_035606_, _037135_, _037817_);
  or g_088328_(_035617_, _037124_, _037828_);
  and g_088329_(_037806_, _037828_, _037839_);
  or g_088330_(_037795_, _037817_, _037850_);
  and g_088331_(_037784_, _037850_, _037861_);
  or g_088332_(_037773_, _037839_, _037872_);
  and g_088333_(_037762_, _037872_, _037883_);
  or g_088334_(_037751_, _037861_, _037894_);
  and g_088335_(_037663_, _037740_, _037905_);
  or g_088336_(_037674_, _037729_, _037916_);
  and g_088337_(_037773_, _037839_, _037927_);
  or g_088338_(_037784_, _037850_, _037938_);
  and g_088339_(_037916_, _037938_, _037949_);
  or g_088340_(_037905_, _037927_, _037960_);
  and g_088341_(_037883_, _037949_, _037971_);
  or g_088342_(_037894_, _037960_, _037982_);
  xor g_088343_(out[148], _012363_, _037993_);
  xor g_088344_(_003530_, _012363_, _038004_);
  and g_088345_(_036123_, _037124_, _038015_);
  or g_088346_(_036112_, _037135_, _038026_);
  and g_088347_(_036046_, _037135_, _038037_);
  or g_088348_(_036057_, _037124_, _038048_);
  and g_088349_(_038026_, _038048_, _038059_);
  or g_088350_(_038015_, _038037_, _038070_);
  and g_088351_(_037993_, _038059_, _038081_);
  or g_088352_(_038004_, _038070_, _038092_);
  xor g_088353_(out[149], _012374_, _038103_);
  xor g_088354_(_003519_, _012374_, _038114_);
  and g_088355_(_035925_, _037124_, _038125_);
  or g_088356_(_035914_, _037135_, _038136_);
  and g_088357_(_035859_, _037135_, _038147_);
  or g_088358_(_035848_, _037124_, _038158_);
  and g_088359_(_038136_, _038158_, _038169_);
  or g_088360_(_038125_, _038147_, _038180_);
  and g_088361_(_038103_, _038180_, _038191_);
  or g_088362_(_038114_, _038169_, _038202_);
  and g_088363_(_038092_, _038202_, _038213_);
  or g_088364_(_038081_, _038191_, _038224_);
  and g_088365_(_038004_, _038070_, _038235_);
  or g_088366_(_037993_, _038059_, _038246_);
  and g_088367_(_038114_, _038169_, _038257_);
  or g_088368_(_038103_, _038180_, _038268_);
  and g_088369_(_038246_, _038268_, _038279_);
  or g_088370_(_038235_, _038257_, _038290_);
  and g_088371_(_038213_, _038279_, _038301_);
  or g_088372_(_038224_, _038290_, _038312_);
  and g_088373_(_037971_, _038301_, _038323_);
  or g_088374_(_037982_, _038312_, _038334_);
  and g_088375_(_036354_, _037124_, _038345_);
  or g_088376_(_036343_, _037135_, _038356_);
  and g_088377_(_036376_, _037135_, _038367_);
  or g_088378_(_036365_, _037124_, _038378_);
  and g_088379_(_038356_, _038378_, _038389_);
  or g_088380_(_038345_, _038367_, _038400_);
  xor g_088381_(out[147], _012341_, _038411_);
  xor g_088382_(_003574_, _012341_, _038422_);
  and g_088383_(_038400_, _038411_, _038433_);
  or g_088384_(_038389_, _038422_, _038444_);
  or g_088385_(out[145], out[146], _038455_);
  xor g_088386_(out[145], out[146], _038466_);
  xor g_088387_(_003541_, out[146], _038477_);
  and g_088388_(_036266_, _037124_, _038488_);
  or g_088389_(_036255_, _037135_, _038499_);
  and g_088390_(_036200_, _037135_, _038510_);
  or g_088391_(_036189_, _037124_, _038521_);
  and g_088392_(_038499_, _038521_, _038532_);
  or g_088393_(_038488_, _038510_, _038543_);
  and g_088394_(_038477_, _038532_, _038554_);
  or g_088395_(_038466_, _038543_, _038565_);
  and g_088396_(_038389_, _038422_, _038576_);
  or g_088397_(_038400_, _038411_, _038587_);
  xor g_088398_(_038477_, _038532_, _038598_);
  xor g_088399_(_038466_, _038532_, _038609_);
  and g_088400_(_038444_, _038587_, _038620_);
  or g_088401_(_038433_, _038576_, _038631_);
  and g_088402_(_038598_, _038620_, _038642_);
  or g_088403_(_038609_, _038631_, _038653_);
  or g_088404_(_036453_, _037135_, _038664_);
  or g_088405_(_003409_, _037124_, _038675_);
  and g_088406_(_038664_, _038675_, _038686_);
  and g_088407_(out[145], _038686_, _038697_);
  not g_088408_(_038697_, _038708_);
  and g_088409_(out[128], _036915_, _038719_);
  or g_088410_(_003420_, _036904_, _038730_);
  and g_088411_(_036970_, _037124_, _038741_);
  or g_088412_(_036981_, _037135_, _038752_);
  and g_088413_(_038730_, _038752_, _038763_);
  or g_088414_(_038719_, _038741_, _038774_);
  and g_088415_(out[144], _038763_, _038785_);
  or g_088416_(_003552_, _038774_, _038796_);
  xor g_088417_(out[145], _038686_, _038807_);
  xor g_088418_(_003541_, _038686_, _038818_);
  and g_088419_(_038796_, _038807_, _038829_);
  or g_088420_(_038785_, _038818_, _038840_);
  and g_088421_(_038708_, _038840_, _038851_);
  or g_088422_(_038697_, _038829_, _038862_);
  and g_088423_(_038642_, _038862_, _038873_);
  or g_088424_(_038653_, _038851_, _038884_);
  and g_088425_(_038554_, _038587_, _038895_);
  or g_088426_(_038565_, _038576_, _038906_);
  and g_088427_(_038444_, _038906_, _038917_);
  or g_088428_(_038433_, _038895_, _038928_);
  and g_088429_(_038884_, _038917_, _038939_);
  or g_088430_(_038873_, _038928_, _038950_);
  and g_088431_(_038323_, _038950_, _038961_);
  or g_088432_(_038334_, _038939_, _038972_);
  or g_088433_(_037883_, _037927_, _038983_);
  not g_088434_(_038983_, _038994_);
  and g_088435_(_038224_, _038268_, _039005_);
  or g_088436_(_038213_, _038257_, _039016_);
  and g_088437_(_037971_, _039005_, _039027_);
  or g_088438_(_037982_, _039016_, _039038_);
  and g_088439_(_038983_, _039038_, _039049_);
  or g_088440_(_038994_, _039027_, _039060_);
  and g_088441_(_038972_, _039049_, _039071_);
  or g_088442_(_038961_, _039060_, _039082_);
  and g_088443_(_037641_, _039082_, _039093_);
  or g_088444_(_037652_, _039071_, _039104_);
  and g_088445_(_037245_, _037267_, _039115_);
  or g_088446_(_037234_, _037256_, _039126_);
  and g_088447_(_037575_, _037608_, _039137_);
  or g_088448_(_037564_, _037597_, _039148_);
  and g_088449_(_037322_, _039137_, _039159_);
  or g_088450_(_037333_, _039148_, _039170_);
  and g_088451_(_039126_, _039170_, _039181_);
  or g_088452_(_039115_, _039159_, _039192_);
  and g_088453_(_039104_, _039181_, _039203_);
  or g_088454_(_039093_, _039192_, _039214_);
  and g_088455_(_037641_, _038323_, _039225_);
  or g_088456_(out[144], _038763_, _039236_);
  and g_088457_(_038642_, _038829_, _039247_);
  and g_088458_(_039236_, _039247_, _039258_);
  and g_088459_(_039225_, _039258_, _039269_);
  not g_088460_(_039269_, _039280_);
  and g_088461_(_039214_, _039280_, _039291_);
  or g_088462_(_039203_, _039269_, _039302_);
  and g_088463_(_026454_, _039291_, _039313_);
  and g_088464_(_037201_, _039302_, _039324_);
  or g_088465_(_039313_, _039324_, _039335_);
  not g_088466_(_039335_, _039346_);
  xor g_088467_(out[166], _012539_, _039357_);
  or g_088468_(_037729_, _039291_, _039368_);
  or g_088469_(_037663_, _039302_, _039379_);
  and g_088470_(_039368_, _039379_, _039390_);
  not g_088471_(_039390_, _039401_);
  or g_088472_(_039357_, _039401_, _039412_);
  xor g_088473_(out[167], _012550_, _039423_);
  not g_088474_(_039423_, _039434_);
  or g_088475_(_037839_, _039291_, _039445_);
  or g_088476_(_037784_, _039302_, _039456_);
  and g_088477_(_039445_, _039456_, _039467_);
  or g_088478_(_039423_, _039467_, _039478_);
  and g_088479_(_039412_, _039478_, _039489_);
  xor g_088480_(out[165], _012528_, _039500_);
  xor g_088481_(_003651_, _012528_, _039511_);
  or g_088482_(_038169_, _039291_, _039522_);
  not g_088483_(_039522_, _039533_);
  and g_088484_(_038114_, _039291_, _039544_);
  not g_088485_(_039544_, _039555_);
  and g_088486_(_039522_, _039555_, _039566_);
  or g_088487_(_039533_, _039544_, _039577_);
  and g_088488_(_039511_, _039566_, _039588_);
  or g_088489_(_039500_, _039577_, _039599_);
  and g_088490_(_039423_, _039467_, _039610_);
  xor g_088491_(_039423_, _039467_, _039621_);
  xor g_088492_(_039434_, _039467_, _039632_);
  xor g_088493_(_039357_, _039401_, _039643_);
  xor g_088494_(_039357_, _039390_, _039654_);
  and g_088495_(_039621_, _039643_, _039665_);
  or g_088496_(_039632_, _039654_, _039676_);
  or g_088497_(_039588_, _039676_, _039687_);
  xor g_088498_(out[170], _012583_, _039698_);
  not g_088499_(_039698_, _039709_);
  and g_088500_(_039346_, _039698_, _039720_);
  and g_088501_(_012473_, _012605_, _039731_);
  or g_088502_(_039720_, _039731_, _039742_);
  and g_088503_(_039335_, _039709_, _039753_);
  and g_088504_(_012484_, _012616_, _039764_);
  or g_088505_(_012473_, _012605_, _039775_);
  or g_088506_(_039753_, _039764_, _039786_);
  xor g_088507_(_039335_, _039709_, _039797_);
  xor g_088508_(_012484_, _012616_, _039808_);
  and g_088509_(_039797_, _039808_, _039819_);
  or g_088510_(_039742_, _039786_, _039830_);
  xor g_088511_(out[168], _012561_, _039841_);
  xor g_088512_(_003717_, _012561_, _039852_);
  or g_088513_(_037520_, _039291_, _039863_);
  not g_088514_(_039863_, _039874_);
  and g_088515_(_037454_, _039291_, _039885_);
  not g_088516_(_039885_, _039896_);
  and g_088517_(_039863_, _039896_, _039907_);
  or g_088518_(_039874_, _039885_, _039918_);
  and g_088519_(_039852_, _039918_, _039929_);
  or g_088520_(_039841_, _039907_, _039940_);
  xor g_088521_(out[169], _012572_, _039951_);
  not g_088522_(_039951_, _039962_);
  or g_088523_(_037410_, _039291_, _039973_);
  not g_088524_(_039973_, _039984_);
  and g_088525_(_037355_, _039291_, _039995_);
  not g_088526_(_039995_, _040006_);
  and g_088527_(_039973_, _040006_, _040017_);
  or g_088528_(_039984_, _039995_, _040028_);
  and g_088529_(_039962_, _040017_, _040039_);
  or g_088530_(_039951_, _040028_, _040050_);
  and g_088531_(_039940_, _040050_, _040061_);
  or g_088532_(_039929_, _040039_, _040072_);
  and g_088533_(_039951_, _040028_, _040083_);
  or g_088534_(_039962_, _040017_, _040094_);
  and g_088535_(_039841_, _039907_, _040105_);
  or g_088536_(_039852_, _039918_, _040116_);
  and g_088537_(_040094_, _040116_, _040127_);
  or g_088538_(_040083_, _040105_, _040138_);
  and g_088539_(_040061_, _040127_, _040149_);
  or g_088540_(_040072_, _040138_, _040160_);
  and g_088541_(_039819_, _040149_, _040171_);
  or g_088542_(_039830_, _040160_, _040182_);
  and g_088543_(_039500_, _039577_, _040193_);
  or g_088544_(_039511_, _039566_, _040204_);
  xor g_088545_(out[164], _012517_, _040215_);
  xor g_088546_(_003662_, _012517_, _040226_);
  or g_088547_(_038059_, _039291_, _040237_);
  not g_088548_(_040237_, _040248_);
  and g_088549_(_037993_, _039291_, _040259_);
  not g_088550_(_040259_, _040270_);
  and g_088551_(_040237_, _040270_, _040281_);
  or g_088552_(_040248_, _040259_, _040292_);
  and g_088553_(_040215_, _040281_, _040303_);
  or g_088554_(_040226_, _040292_, _040314_);
  and g_088555_(_040204_, _040314_, _040325_);
  or g_088556_(_040193_, _040303_, _040336_);
  and g_088557_(_040226_, _040292_, _040347_);
  or g_088558_(_040215_, _040281_, _040358_);
  or g_088559_(_040336_, _040347_, _040369_);
  or g_088560_(_040182_, _040369_, _040380_);
  and g_088561_(_039599_, _040358_, _040391_);
  and g_088562_(_039665_, _040391_, _040402_);
  and g_088563_(_040325_, _040402_, _040413_);
  and g_088564_(_040171_, _040413_, _040424_);
  or g_088565_(_039687_, _040380_, _040435_);
  xor g_088566_(out[163], _012495_, _040446_);
  xor g_088567_(_003706_, _012495_, _040457_);
  or g_088568_(_038389_, _039291_, _040468_);
  not g_088569_(_040468_, _040479_);
  and g_088570_(_038422_, _039291_, _040490_);
  not g_088571_(_040490_, _040501_);
  and g_088572_(_040468_, _040501_, _040512_);
  or g_088573_(_040479_, _040490_, _040523_);
  and g_088574_(_040457_, _040512_, _040534_);
  or g_088575_(_040446_, _040523_, _040545_);
  or g_088576_(out[161], out[162], _040556_);
  xor g_088577_(out[161], out[162], _040567_);
  xor g_088578_(_003673_, out[162], _040578_);
  or g_088579_(_038532_, _039291_, _040589_);
  not g_088580_(_040589_, _040600_);
  and g_088581_(_038477_, _039291_, _040611_);
  not g_088582_(_040611_, _040622_);
  and g_088583_(_040589_, _040622_, _040633_);
  or g_088584_(_040600_, _040611_, _040644_);
  and g_088585_(_040578_, _040633_, _040655_);
  or g_088586_(_040567_, _040644_, _040666_);
  and g_088587_(_040446_, _040523_, _040677_);
  or g_088588_(_040457_, _040512_, _040688_);
  and g_088589_(_040666_, _040688_, _040699_);
  or g_088590_(_040655_, _040677_, _040710_);
  or g_088591_(_003541_, _039302_, _040721_);
  or g_088592_(_038686_, _039291_, _040732_);
  and g_088593_(_040721_, _040732_, _040743_);
  and g_088594_(out[161], _040743_, _040754_);
  not g_088595_(_040754_, _040765_);
  and g_088596_(_003552_, _039291_, _040776_);
  and g_088597_(_038763_, _039302_, _040787_);
  or g_088598_(_040776_, _040787_, _040798_);
  and g_088599_(out[160], _040798_, _040809_);
  not g_088600_(_040809_, _040820_);
  xor g_088601_(out[161], _040743_, _040831_);
  xor g_088602_(_003673_, _040743_, _040842_);
  and g_088603_(_040820_, _040831_, _040853_);
  or g_088604_(_040809_, _040842_, _040864_);
  and g_088605_(_040765_, _040864_, _040875_);
  or g_088606_(_040754_, _040853_, _040886_);
  xor g_088607_(_040578_, _040633_, _040897_);
  xor g_088608_(_040567_, _040633_, _040908_);
  and g_088609_(_040886_, _040897_, _040919_);
  or g_088610_(_040875_, _040908_, _040930_);
  and g_088611_(_040699_, _040930_, _040941_);
  or g_088612_(_040710_, _040919_, _040952_);
  or g_088613_(_040534_, _040908_, _040963_);
  and g_088614_(_040545_, _040952_, _040974_);
  or g_088615_(_040534_, _040941_, _040985_);
  and g_088616_(_040424_, _040974_, _040996_);
  or g_088617_(_040435_, _040985_, _041007_);
  or g_088618_(_039687_, _040325_, _041018_);
  or g_088619_(_039489_, _039610_, _041029_);
  and g_088620_(_041018_, _041029_, _041040_);
  or g_088621_(_040182_, _041040_, _041051_);
  or g_088622_(_040039_, _040127_, _041062_);
  or g_088623_(_039830_, _041062_, _041073_);
  and g_088624_(_039742_, _039775_, _041084_);
  not g_088625_(_041084_, _041095_);
  and g_088626_(_041073_, _041095_, _041106_);
  and g_088627_(_041051_, _041106_, _041117_);
  not g_088628_(_041117_, _041128_);
  and g_088629_(_041007_, _041117_, _041139_);
  or g_088630_(_040996_, _041128_, _041150_);
  or g_088631_(out[160], _040798_, _041161_);
  not g_088632_(_041161_, _041172_);
  or g_088633_(_040677_, _041172_, _041183_);
  or g_088634_(_040963_, _041183_, _041194_);
  or g_088635_(_040435_, _041194_, _041205_);
  not g_088636_(_041205_, _041216_);
  and g_088637_(_040853_, _041216_, _041227_);
  or g_088638_(_040864_, _041205_, _041238_);
  and g_088639_(_041150_, _041238_, _041249_);
  or g_088640_(_041139_, _041227_, _041260_);
  and g_088641_(_039335_, _041260_, _041271_);
  not g_088642_(_041271_, _041282_);
  or g_088643_(_039709_, _041260_, _041293_);
  not g_088644_(_041293_, _041304_);
  and g_088645_(_041282_, _041293_, _041315_);
  or g_088646_(_041271_, _041304_, _041326_);
  and g_088647_(_012638_, _012759_, _041337_);
  or g_088648_(_012627_, _012770_, _041348_);
  and g_088649_(_012627_, _012770_, _041359_);
  or g_088650_(_012638_, _012759_, _041370_);
  xor g_088651_(out[186], _012737_, _041381_);
  xor g_088652_(_003871_, _012737_, _041392_);
  and g_088653_(_041315_, _041381_, _041403_);
  or g_088654_(_041326_, _041392_, _041414_);
  and g_088655_(_041370_, _041414_, _041425_);
  or g_088656_(_041359_, _041403_, _041436_);
  and g_088657_(_041348_, _041436_, _041447_);
  or g_088658_(_041337_, _041425_, _041458_);
  and g_088659_(_041326_, _041392_, _041469_);
  or g_088660_(_041315_, _041381_, _041480_);
  and g_088661_(_041348_, _041480_, _041491_);
  or g_088662_(_041337_, _041469_, _041502_);
  xor g_088663_(out[185], _012726_, _041513_);
  xor g_088664_(_003860_, _012726_, _041524_);
  or g_088665_(_040017_, _041249_, _041535_);
  or g_088666_(_039951_, _041260_, _041546_);
  and g_088667_(_041535_, _041546_, _041557_);
  not g_088668_(_041557_, _041568_);
  and g_088669_(_041524_, _041557_, _041579_);
  or g_088670_(_041513_, _041568_, _041590_);
  and g_088671_(_041491_, _041590_, _041601_);
  or g_088672_(_041502_, _041579_, _041612_);
  and g_088673_(_041425_, _041601_, _041623_);
  or g_088674_(_041436_, _041612_, _041634_);
  xor g_088675_(out[184], _012715_, _041645_);
  not g_088676_(_041645_, _041656_);
  and g_088677_(_039918_, _041260_, _041667_);
  not g_088678_(_041667_, _041678_);
  or g_088679_(_039852_, _041260_, _041689_);
  not g_088680_(_041689_, _041700_);
  and g_088681_(_041678_, _041689_, _041711_);
  or g_088682_(_041667_, _041700_, _041722_);
  and g_088683_(_041645_, _041711_, _041733_);
  or g_088684_(_041656_, _041722_, _041744_);
  and g_088685_(_041513_, _041568_, _041755_);
  or g_088686_(_041524_, _041557_, _041766_);
  and g_088687_(_041744_, _041766_, _041777_);
  or g_088688_(_041733_, _041755_, _041788_);
  and g_088689_(_040743_, _041260_, _041799_);
  not g_088690_(_041799_, _041810_);
  and g_088691_(_003673_, _041249_, _041821_);
  or g_088692_(out[161], _041260_, _041832_);
  or g_088693_(_041799_, _041821_, _041843_);
  and g_088694_(_041810_, _041832_, _041854_);
  and g_088695_(out[177], _041843_, _041865_);
  or g_088696_(_003805_, _041854_, _041876_);
  and g_088697_(_040798_, _041260_, _041887_);
  not g_088698_(_041887_, _041898_);
  or g_088699_(out[160], _041260_, _041909_);
  and g_088700_(_041898_, _041909_, _041920_);
  not g_088701_(_041920_, _041931_);
  and g_088702_(out[176], _041931_, _041942_);
  or g_088703_(_003816_, _041920_, _041953_);
  xor g_088704_(out[177], _041843_, _041964_);
  xor g_088705_(_003805_, _041843_, _041975_);
  and g_088706_(_041953_, _041964_, _041986_);
  or g_088707_(_041942_, _041975_, _041997_);
  and g_088708_(_041876_, _041997_, _042008_);
  or g_088709_(_041865_, _041986_, _042019_);
  xor g_088710_(out[182], _012693_, _042030_);
  xor g_088711_(_003772_, _012693_, _042041_);
  or g_088712_(_039390_, _041249_, _042052_);
  or g_088713_(_039357_, _041260_, _042063_);
  and g_088714_(_042052_, _042063_, _042074_);
  not g_088715_(_042074_, _042085_);
  or g_088716_(_042030_, _042085_, _042096_);
  xor g_088717_(out[183], _012704_, _042107_);
  or g_088718_(_039467_, _041249_, _042118_);
  or g_088719_(_039434_, _041260_, _042129_);
  and g_088720_(_042118_, _042129_, _042140_);
  and g_088721_(_042107_, _042140_, _042151_);
  xor g_088722_(_042041_, _042074_, _042162_);
  xor g_088723_(_042030_, _042074_, _042173_);
  or g_088724_(_042151_, _042173_, _042184_);
  xor g_088725_(out[181], _012682_, _042195_);
  xor g_088726_(_003783_, _012682_, _042206_);
  and g_088727_(_039577_, _041260_, _042217_);
  or g_088728_(_039566_, _041249_, _042228_);
  and g_088729_(_039511_, _041249_, _042239_);
  or g_088730_(_039500_, _041260_, _042250_);
  and g_088731_(_042228_, _042250_, _042261_);
  or g_088732_(_042217_, _042239_, _042272_);
  and g_088733_(_042206_, _042261_, _042283_);
  not g_088734_(_042283_, _042294_);
  xor g_088735_(out[180], _012671_, _042305_);
  not g_088736_(_042305_, _042316_);
  and g_088737_(_040292_, _041260_, _042327_);
  or g_088738_(_040281_, _041249_, _042338_);
  and g_088739_(_040215_, _041249_, _042349_);
  or g_088740_(_040226_, _041260_, _042360_);
  and g_088741_(_042338_, _042360_, _042371_);
  or g_088742_(_042327_, _042349_, _042382_);
  and g_088743_(_042305_, _042371_, _042393_);
  or g_088744_(_042316_, _042382_, _042404_);
  or g_088745_(_042283_, _042393_, _042415_);
  and g_088746_(_042316_, _042382_, _042426_);
  or g_088747_(_042305_, _042371_, _042437_);
  and g_088748_(_042195_, _042272_, _042448_);
  or g_088749_(_042206_, _042261_, _042459_);
  or g_088750_(_042107_, _042140_, _042470_);
  not g_088751_(_042470_, _042481_);
  xor g_088752_(_042107_, _042140_, _042492_);
  and g_088753_(_042162_, _042492_, _042503_);
  or g_088754_(_042184_, _042481_, _042514_);
  and g_088755_(_042404_, _042459_, _042525_);
  and g_088756_(_042437_, _042525_, _042536_);
  or g_088757_(_042426_, _042448_, _042547_);
  and g_088758_(_042294_, _042536_, _042558_);
  or g_088759_(_042415_, _042547_, _042569_);
  and g_088760_(_042503_, _042558_, _042580_);
  or g_088761_(_042514_, _042569_, _042591_);
  xor g_088762_(out[179], _012649_, _042602_);
  xor g_088763_(_003838_, _012649_, _042613_);
  or g_088764_(_040512_, _041249_, _042624_);
  or g_088765_(_040446_, _041260_, _042635_);
  and g_088766_(_042624_, _042635_, _042646_);
  not g_088767_(_042646_, _042657_);
  and g_088768_(_042602_, _042657_, _042668_);
  or g_088769_(out[177], out[178], _042679_);
  xor g_088770_(out[177], out[178], _042690_);
  xor g_088771_(_003805_, out[178], _042701_);
  or g_088772_(_040633_, _041249_, _042712_);
  or g_088773_(_040567_, _041260_, _042723_);
  and g_088774_(_042712_, _042723_, _042734_);
  and g_088775_(_042701_, _042734_, _042745_);
  or g_088776_(_042668_, _042745_, _042756_);
  or g_088777_(_042602_, _042657_, _042767_);
  xor g_088778_(_042613_, _042646_, _042778_);
  xor g_088779_(_042602_, _042646_, _042789_);
  xor g_088780_(_042701_, _042734_, _042800_);
  xor g_088781_(_042690_, _042734_, _042811_);
  and g_088782_(_042778_, _042800_, _042822_);
  or g_088783_(_042789_, _042811_, _042833_);
  and g_088784_(_042580_, _042822_, _042844_);
  or g_088785_(_042591_, _042833_, _042855_);
  and g_088786_(_042019_, _042844_, _042866_);
  or g_088787_(_042008_, _042855_, _042877_);
  and g_088788_(_042756_, _042767_, _042888_);
  and g_088789_(_042580_, _042888_, _042899_);
  not g_088790_(_042899_, _042910_);
  and g_088791_(_042096_, _042470_, _042921_);
  or g_088792_(_042151_, _042921_, _042932_);
  or g_088793_(_042283_, _042525_, _042943_);
  or g_088794_(_042184_, _042943_, _042954_);
  and g_088795_(_042932_, _042954_, _042965_);
  not g_088796_(_042965_, _042976_);
  and g_088797_(_042910_, _042965_, _042987_);
  or g_088798_(_042899_, _042976_, _042998_);
  and g_088799_(_042877_, _042987_, _043009_);
  or g_088800_(_042866_, _042998_, _043020_);
  and g_088801_(_041656_, _041722_, _043031_);
  or g_088802_(_041645_, _041711_, _043042_);
  and g_088803_(_043020_, _043042_, _043053_);
  or g_088804_(_043009_, _043031_, _043064_);
  and g_088805_(_041777_, _043064_, _043075_);
  or g_088806_(_041788_, _043053_, _043086_);
  and g_088807_(_041623_, _043086_, _043097_);
  or g_088808_(_041634_, _043075_, _043108_);
  and g_088809_(_041458_, _043108_, _043119_);
  or g_088810_(_041447_, _043097_, _043130_);
  or g_088811_(out[176], _041931_, _043141_);
  and g_088812_(_043042_, _043141_, _043152_);
  and g_088813_(_041777_, _043152_, _043163_);
  and g_088814_(_041623_, _041986_, _043174_);
  or g_088815_(_041634_, _041997_, _043185_);
  and g_088816_(_042844_, _043163_, _043196_);
  not g_088817_(_043196_, _043207_);
  and g_088818_(_043174_, _043196_, _043218_);
  or g_088819_(_043185_, _043207_, _043229_);
  and g_088820_(_043130_, _043229_, _043240_);
  or g_088821_(_043119_, _043218_, _043251_);
  and g_088822_(_041326_, _043251_, _043262_);
  or g_088823_(_041315_, _043240_, _043273_);
  and g_088824_(_041381_, _043240_, _043284_);
  or g_088825_(_041392_, _043251_, _043295_);
  and g_088826_(_043273_, _043295_, _043306_);
  or g_088827_(_043262_, _043284_, _043317_);
  and g_088828_(_026410_, _043306_, _043328_);
  or g_088829_(_026421_, _043317_, _043339_);
  and g_088830_(_026443_, _043339_, _043350_);
  or g_088831_(_026432_, _043328_, _043361_);
  and g_088832_(_026421_, _043317_, _043372_);
  or g_088833_(_026410_, _043306_, _043383_);
  and g_088834_(_012792_, _012924_, _043394_);
  or g_088835_(_012781_, _012935_, _043405_);
  and g_088836_(_043383_, _043405_, _043416_);
  or g_088837_(_043372_, _043394_, _043427_);
  and g_088838_(_043350_, _043416_, _043438_);
  or g_088839_(_043361_, _043427_, _043449_);
  and g_088840_(out[201], _012880_, _043460_);
  xor g_088841_(out[201], _012880_, _043471_);
  or g_088842_(_012902_, _043460_, _043482_);
  and g_088843_(_041524_, _043240_, _043493_);
  not g_088844_(_043493_, _043504_);
  or g_088845_(_041557_, _043240_, _043515_);
  not g_088846_(_043515_, _043526_);
  and g_088847_(_043504_, _043515_, _043537_);
  or g_088848_(_043493_, _043526_, _043548_);
  and g_088849_(_043471_, _043548_, _043559_);
  or g_088850_(_043482_, _043537_, _043570_);
  xor g_088851_(out[200], _012869_, _043581_);
  xor g_088852_(_003981_, _012869_, _043592_);
  and g_088853_(_041645_, _043240_, _043603_);
  not g_088854_(_043603_, _043614_);
  or g_088855_(_041711_, _043240_, _043625_);
  not g_088856_(_043625_, _043636_);
  and g_088857_(_043614_, _043625_, _043647_);
  or g_088858_(_043603_, _043636_, _043658_);
  and g_088859_(_043581_, _043647_, _043669_);
  or g_088860_(_043592_, _043658_, _043680_);
  and g_088861_(_043570_, _043680_, _043691_);
  or g_088862_(_043559_, _043669_, _043702_);
  and g_088863_(_043482_, _043537_, _043713_);
  or g_088864_(_043471_, _043548_, _043724_);
  and g_088865_(_043592_, _043658_, _043735_);
  or g_088866_(_043581_, _043647_, _043746_);
  and g_088867_(_043724_, _043746_, _043757_);
  or g_088868_(_043713_, _043735_, _043768_);
  and g_088869_(_043691_, _043757_, _043779_);
  or g_088870_(_043702_, _043768_, _043790_);
  and g_088871_(_043438_, _043779_, _043801_);
  or g_088872_(_043449_, _043790_, _043812_);
  and g_088873_(_042041_, _043240_, _043823_);
  not g_088874_(_043823_, _043834_);
  or g_088875_(_042074_, _043240_, _043845_);
  not g_088876_(_043845_, _043856_);
  and g_088877_(_043834_, _043845_, _043867_);
  or g_088878_(_043823_, _043856_, _043878_);
  xor g_088879_(out[198], _012847_, _043889_);
  or g_088880_(_043878_, _043889_, _043900_);
  xor g_088881_(out[199], _012858_, _043911_);
  xor g_088882_(_003893_, _012858_, _043922_);
  and g_088883_(_042107_, _043240_, _043933_);
  not g_088884_(_043933_, _043944_);
  or g_088885_(_042140_, _043240_, _043955_);
  not g_088886_(_043955_, _043966_);
  and g_088887_(_043944_, _043955_, _043977_);
  or g_088888_(_043933_, _043966_, _043988_);
  or g_088889_(_043911_, _043977_, _043999_);
  and g_088890_(_043900_, _043999_, _044010_);
  xor g_088891_(out[197], _012836_, _044021_);
  xor g_088892_(_003915_, _012836_, _044032_);
  and g_088893_(_042206_, _043240_, _044043_);
  not g_088894_(_044043_, _044054_);
  or g_088895_(_042261_, _043240_, _044065_);
  not g_088896_(_044065_, _044076_);
  and g_088897_(_044054_, _044065_, _044087_);
  or g_088898_(_044043_, _044076_, _044098_);
  and g_088899_(_044032_, _044087_, _044109_);
  or g_088900_(_044021_, _044098_, _044120_);
  and g_088901_(_043911_, _043977_, _044131_);
  xor g_088902_(_043878_, _043889_, _044142_);
  xor g_088903_(_043867_, _043889_, _044153_);
  xor g_088904_(_043911_, _043977_, _044164_);
  xor g_088905_(_043922_, _043977_, _044175_);
  and g_088906_(_044142_, _044164_, _044186_);
  or g_088907_(_044153_, _044175_, _044197_);
  and g_088908_(_044120_, _044186_, _044208_);
  or g_088909_(_044109_, _044197_, _044219_);
  and g_088910_(_044021_, _044098_, _044230_);
  or g_088911_(_044032_, _044087_, _044241_);
  xor g_088912_(out[196], _012825_, _044252_);
  xor g_088913_(_003926_, _012825_, _044263_);
  and g_088914_(_042305_, _043240_, _044274_);
  not g_088915_(_044274_, _044285_);
  or g_088916_(_042371_, _043240_, _044296_);
  not g_088917_(_044296_, _044307_);
  and g_088918_(_044285_, _044296_, _044318_);
  or g_088919_(_044274_, _044307_, _044329_);
  and g_088920_(_044252_, _044318_, _044340_);
  or g_088921_(_044263_, _044329_, _044351_);
  and g_088922_(_044241_, _044351_, _044362_);
  or g_088923_(_044230_, _044340_, _044373_);
  xor g_088924_(out[195], _012803_, _044384_);
  xor g_088925_(_003970_, _012803_, _044395_);
  and g_088926_(_042613_, _043240_, _044406_);
  not g_088927_(_044406_, _044417_);
  or g_088928_(_042646_, _043240_, _044428_);
  not g_088929_(_044428_, _044439_);
  and g_088930_(_044417_, _044428_, _044450_);
  or g_088931_(_044406_, _044439_, _044461_);
  and g_088932_(_044395_, _044450_, _044472_);
  or g_088933_(_044384_, _044461_, _044483_);
  and g_088934_(_044263_, _044329_, _044494_);
  or g_088935_(_044252_, _044318_, _044505_);
  or g_088936_(out[193], out[194], _044516_);
  xor g_088937_(out[193], out[194], _044527_);
  xor g_088938_(_003937_, out[194], _044538_);
  or g_088939_(_042734_, _043240_, _044549_);
  not g_088940_(_044549_, _044560_);
  and g_088941_(_042701_, _043240_, _044571_);
  not g_088942_(_044571_, _044582_);
  and g_088943_(_044549_, _044582_, _044593_);
  or g_088944_(_044560_, _044571_, _044604_);
  and g_088945_(_044538_, _044593_, _044615_);
  or g_088946_(_044527_, _044604_, _044626_);
  xor g_088947_(_044538_, _044593_, _044637_);
  xor g_088948_(_044527_, _044593_, _044648_);
  and g_088949_(_044384_, _044461_, _044659_);
  or g_088950_(_044395_, _044450_, _044670_);
  and g_088951_(_044483_, _044670_, _044681_);
  or g_088952_(_044472_, _044659_, _044692_);
  and g_088953_(_044362_, _044505_, _044703_);
  or g_088954_(_044373_, _044494_, _044714_);
  and g_088955_(_044208_, _044703_, _044725_);
  or g_088956_(_044219_, _044714_, _044736_);
  and g_088957_(_043801_, _044725_, _044747_);
  or g_088958_(_043812_, _044736_, _044758_);
  and g_088959_(_044681_, _044747_, _044769_);
  or g_088960_(_044692_, _044758_, _044780_);
  and g_088961_(_044637_, _044769_, _044791_);
  or g_088962_(_044648_, _044780_, _044802_);
  or g_088963_(_041843_, _043240_, _044813_);
  not g_088964_(_044813_, _044824_);
  and g_088965_(out[177], _043240_, _044835_);
  not g_088966_(_044835_, _044846_);
  and g_088967_(_044813_, _044846_, _044857_);
  or g_088968_(_044824_, _044835_, _044868_);
  and g_088969_(out[193], _044857_, _044879_);
  or g_088970_(_003937_, _044868_, _044890_);
  and g_088971_(_044791_, _044879_, _044901_);
  or g_088972_(_044802_, _044890_, _044912_);
  and g_088973_(_044208_, _044373_, _044923_);
  or g_088974_(_044219_, _044362_, _044934_);
  or g_088975_(_044010_, _044131_, _044945_);
  not g_088976_(_044945_, _044956_);
  and g_088977_(_044934_, _044945_, _044967_);
  or g_088978_(_044923_, _044956_, _044978_);
  and g_088979_(_043801_, _044978_, _044989_);
  or g_088980_(_043812_, _044967_, _045000_);
  and g_088981_(_043361_, _043405_, _045011_);
  or g_088982_(_043350_, _043394_, _045022_);
  and g_088983_(_043702_, _043724_, _045033_);
  or g_088984_(_043691_, _043713_, _045044_);
  and g_088985_(_043438_, _045033_, _045055_);
  or g_088986_(_043449_, _045044_, _045066_);
  and g_088987_(_045022_, _045066_, _045077_);
  or g_088988_(_045011_, _045055_, _045088_);
  and g_088989_(_044626_, _044670_, _045099_);
  or g_088990_(_044615_, _044659_, _045110_);
  or g_088991_(_044472_, _045099_, _045121_);
  and g_088992_(_044483_, _045110_, _045132_);
  and g_088993_(_044747_, _045132_, _045143_);
  or g_088994_(_044758_, _045121_, _045154_);
  and g_088995_(_045077_, _045154_, _045165_);
  or g_088996_(_045088_, _045143_, _045176_);
  and g_088997_(_045000_, _045165_, _045187_);
  or g_088998_(_044989_, _045176_, _045198_);
  and g_088999_(_044912_, _045187_, _045209_);
  or g_089000_(_044901_, _045198_, _045220_);
  or g_089001_(_041920_, _043240_, _045231_);
  not g_089002_(_045231_, _045242_);
  and g_089003_(_003816_, _043240_, _045253_);
  not g_089004_(_045253_, _045264_);
  and g_089005_(_045231_, _045264_, _045275_);
  or g_089006_(_045242_, _045253_, _045286_);
  and g_089007_(out[192], _045286_, _045297_);
  or g_089008_(_003948_, _045275_, _045308_);
  xor g_089009_(out[193], _044857_, _045319_);
  xor g_089010_(_003937_, _044857_, _045330_);
  and g_089011_(_045308_, _045319_, _045341_);
  or g_089012_(_045297_, _045330_, _045352_);
  and g_089013_(_044791_, _045341_, _045363_);
  or g_089014_(_044802_, _045352_, _045374_);
  and g_089015_(_003948_, _045275_, _045385_);
  or g_089016_(out[192], _045286_, _045396_);
  and g_089017_(_045363_, _045385_, _045407_);
  or g_089018_(_045374_, _045396_, _045418_);
  and g_089019_(_045209_, _045418_, _045429_);
  or g_089020_(_045220_, _045407_, _045440_);
  and g_089021_(_026410_, _045440_, _045451_);
  or g_089022_(_026421_, _045429_, _045462_);
  and g_089023_(_043317_, _045429_, _045473_);
  or g_089024_(_043306_, _045440_, _045484_);
  and g_089025_(_045462_, _045484_, _045495_);
  or g_089026_(_045451_, _045473_, _045506_);
  and g_089027_(_012946_, _013089_, _045517_);
  or g_089028_(_012957_, _013078_, _045528_);
  xor g_089029_(out[218], _013056_, _045539_);
  xor g_089030_(_004113_, _013056_, _045550_);
  and g_089031_(_045495_, _045539_, _045561_);
  or g_089032_(_045506_, _045550_, _045572_);
  and g_089033_(_045528_, _045572_, _045583_);
  or g_089034_(_045517_, _045561_, _045594_);
  and g_089035_(_045506_, _045550_, _045605_);
  or g_089036_(_045495_, _045539_, _045616_);
  and g_089037_(_012957_, _013078_, _045627_);
  or g_089038_(_012946_, _013089_, _045638_);
  and g_089039_(_045616_, _045638_, _045649_);
  or g_089040_(_045605_, _045627_, _045660_);
  and g_089041_(_045583_, _045649_, _045671_);
  or g_089042_(_045594_, _045660_, _045682_);
  xor g_089043_(out[216], _013034_, _045693_);
  not g_089044_(_045693_, _045704_);
  and g_089045_(_043658_, _045429_, _045715_);
  or g_089046_(_043647_, _045440_, _045726_);
  and g_089047_(_043581_, _045440_, _045737_);
  or g_089048_(_043592_, _045429_, _045748_);
  and g_089049_(_045726_, _045748_, _045759_);
  or g_089050_(_045715_, _045737_, _045770_);
  and g_089051_(_045693_, _045759_, _045781_);
  or g_089052_(_045704_, _045770_, _045792_);
  xor g_089053_(out[217], _013045_, _045803_);
  xor g_089054_(_004102_, _013045_, _045814_);
  or g_089055_(_043537_, _045440_, _045825_);
  or g_089056_(_043471_, _045429_, _045836_);
  and g_089057_(_045825_, _045836_, _045847_);
  not g_089058_(_045847_, _045858_);
  and g_089059_(_045803_, _045858_, _045869_);
  or g_089060_(_045814_, _045847_, _045880_);
  and g_089061_(_045792_, _045880_, _045891_);
  or g_089062_(_045781_, _045869_, _045902_);
  and g_089063_(_045704_, _045770_, _045913_);
  or g_089064_(_045693_, _045759_, _045924_);
  and g_089065_(_045814_, _045847_, _045935_);
  or g_089066_(_045803_, _045858_, _045946_);
  and g_089067_(_045924_, _045946_, _045957_);
  or g_089068_(_045913_, _045935_, _045968_);
  and g_089069_(_045891_, _045957_, _045979_);
  or g_089070_(_045902_, _045968_, _045990_);
  and g_089071_(_045671_, _045979_, _046001_);
  or g_089072_(_045682_, _045990_, _046012_);
  and g_089073_(_043878_, _045429_, _046023_);
  or g_089074_(_043867_, _045440_, _046034_);
  or g_089075_(_043889_, _045429_, _046045_);
  not g_089076_(_046045_, _046056_);
  and g_089077_(_046034_, _046045_, _046067_);
  or g_089078_(_046023_, _046056_, _046078_);
  xor g_089079_(out[214], _013012_, _046089_);
  not g_089080_(_046089_, _046100_);
  or g_089081_(_046078_, _046089_, _046111_);
  xor g_089082_(out[215], _013023_, _046122_);
  and g_089083_(_043988_, _045429_, _046133_);
  or g_089084_(_043977_, _045440_, _046144_);
  and g_089085_(_043911_, _045440_, _046155_);
  or g_089086_(_043922_, _045429_, _046166_);
  and g_089087_(_046144_, _046166_, _046177_);
  or g_089088_(_046133_, _046155_, _046188_);
  or g_089089_(_046122_, _046177_, _046199_);
  and g_089090_(_046111_, _046199_, _046210_);
  and g_089091_(_046122_, _046177_, _046221_);
  xor g_089092_(_046067_, _046100_, _046232_);
  xor g_089093_(_046067_, _046089_, _046243_);
  xor g_089094_(_046122_, _046177_, _046254_);
  xor g_089095_(_046122_, _046188_, _046265_);
  and g_089096_(_046232_, _046254_, _046276_);
  or g_089097_(_046243_, _046265_, _046287_);
  xor g_089098_(out[213], _013001_, _046298_);
  xor g_089099_(_004025_, _013001_, _046309_);
  and g_089100_(_044098_, _045429_, _046320_);
  or g_089101_(_044087_, _045440_, _046331_);
  and g_089102_(_044032_, _045440_, _046342_);
  or g_089103_(_044021_, _045429_, _046353_);
  and g_089104_(_046331_, _046353_, _046364_);
  or g_089105_(_046320_, _046342_, _046375_);
  and g_089106_(_046298_, _046375_, _046386_);
  or g_089107_(_046309_, _046364_, _046397_);
  xor g_089108_(out[212], _012990_, _046408_);
  xor g_089109_(_004036_, _012990_, _046419_);
  and g_089110_(_044329_, _045429_, _046430_);
  or g_089111_(_044318_, _045440_, _046441_);
  and g_089112_(_044252_, _045440_, _046452_);
  or g_089113_(_044263_, _045429_, _046463_);
  and g_089114_(_046441_, _046463_, _046474_);
  or g_089115_(_046430_, _046452_, _046485_);
  and g_089116_(_046408_, _046474_, _046496_);
  or g_089117_(_046419_, _046485_, _046507_);
  and g_089118_(_046397_, _046507_, _046518_);
  or g_089119_(_046386_, _046496_, _046529_);
  and g_089120_(_046419_, _046485_, _046540_);
  or g_089121_(_046408_, _046474_, _046551_);
  and g_089122_(_046309_, _046364_, _046562_);
  or g_089123_(_046298_, _046375_, _046573_);
  and g_089124_(_046551_, _046573_, _046584_);
  or g_089125_(_046540_, _046562_, _046595_);
  and g_089126_(_046518_, _046584_, _046606_);
  or g_089127_(_046529_, _046595_, _046617_);
  and g_089128_(_046276_, _046606_, _046628_);
  or g_089129_(_046287_, _046617_, _046639_);
  and g_089130_(_046001_, _046628_, _046650_);
  or g_089131_(_046012_, _046639_, _046661_);
  and g_089132_(_044868_, _045429_, _046672_);
  or g_089133_(_044857_, _045440_, _046683_);
  and g_089134_(out[193], _045440_, _046694_);
  or g_089135_(_003937_, _045429_, _046705_);
  and g_089136_(_046683_, _046705_, _046716_);
  or g_089137_(_046672_, _046694_, _046727_);
  and g_089138_(out[192], _045220_, _046738_);
  and g_089139_(_045275_, _045429_, _046749_);
  or g_089140_(_046738_, _046749_, _046760_);
  not g_089141_(_046760_, _046771_);
  and g_089142_(out[208], _046771_, _046782_);
  or g_089143_(_004058_, _046760_, _046793_);
  and g_089144_(out[209], _046716_, _046804_);
  or g_089145_(_004047_, _046727_, _046815_);
  xor g_089146_(out[209], _046716_, _046826_);
  xor g_089147_(_004047_, _046716_, _046837_);
  and g_089148_(_046793_, _046826_, _046848_);
  or g_089149_(_046782_, _046837_, _046859_);
  or g_089150_(out[209], out[210], _046870_);
  xor g_089151_(out[209], out[210], _046881_);
  xor g_089152_(_004047_, out[210], _046892_);
  and g_089153_(_044604_, _045429_, _046903_);
  or g_089154_(_044593_, _045440_, _046914_);
  and g_089155_(_044538_, _045440_, _046925_);
  or g_089156_(_044527_, _045429_, _046936_);
  and g_089157_(_046914_, _046936_, _046947_);
  or g_089158_(_046903_, _046925_, _046958_);
  and g_089159_(_046892_, _046947_, _046969_);
  or g_089160_(_046881_, _046958_, _046980_);
  xor g_089161_(_046892_, _046947_, _046991_);
  xor g_089162_(_046881_, _046947_, _047002_);
  xor g_089163_(out[211], _012968_, _047013_);
  xor g_089164_(_004080_, _012968_, _047024_);
  or g_089165_(_044450_, _045440_, _047035_);
  or g_089166_(_044384_, _045429_, _047046_);
  and g_089167_(_047035_, _047046_, _047057_);
  not g_089168_(_047057_, _047068_);
  and g_089169_(_047013_, _047068_, _047079_);
  or g_089170_(_047024_, _047057_, _047090_);
  and g_089171_(_047024_, _047057_, _047101_);
  or g_089172_(_047013_, _047068_, _047112_);
  and g_089173_(_004058_, _046760_, _047123_);
  or g_089174_(out[208], _046771_, _047134_);
  and g_089175_(_046991_, _047112_, _047145_);
  or g_089176_(_047002_, _047101_, _047156_);
  and g_089177_(_047090_, _047134_, _047167_);
  or g_089178_(_047079_, _047123_, _047178_);
  and g_089179_(_047145_, _047167_, _047189_);
  or g_089180_(_047156_, _047178_, _047200_);
  and g_089181_(_046848_, _047189_, _047211_);
  or g_089182_(_046859_, _047200_, _047222_);
  and g_089183_(_046650_, _047211_, _047233_);
  or g_089184_(_046661_, _047222_, _047244_);
  and g_089185_(_046815_, _046859_, _047255_);
  or g_089186_(_046804_, _046848_, _047266_);
  and g_089187_(_046969_, _047112_, _047277_);
  or g_089188_(_046980_, _047101_, _047288_);
  and g_089189_(_047145_, _047266_, _047299_);
  or g_089190_(_047156_, _047255_, _047310_);
  and g_089191_(_047288_, _047310_, _047321_);
  or g_089192_(_047277_, _047299_, _047332_);
  and g_089193_(_047090_, _047321_, _047343_);
  or g_089194_(_047079_, _047332_, _047354_);
  and g_089195_(_046650_, _047354_, _047365_);
  or g_089196_(_046661_, _047343_, _047376_);
  or g_089197_(_046210_, _046221_, _047387_);
  not g_089198_(_047387_, _047398_);
  and g_089199_(_046276_, _046529_, _047409_);
  or g_089200_(_046287_, _046518_, _047420_);
  and g_089201_(_046573_, _047409_, _047431_);
  or g_089202_(_046562_, _047420_, _047442_);
  and g_089203_(_047387_, _047442_, _047453_);
  or g_089204_(_047398_, _047431_, _047464_);
  and g_089205_(_046001_, _047464_, _047475_);
  or g_089206_(_046012_, _047453_, _047486_);
  or g_089207_(_045891_, _045935_, _047497_);
  and g_089208_(_045671_, _045902_, _047508_);
  and g_089209_(_045946_, _047508_, _047519_);
  or g_089210_(_045682_, _047497_, _047530_);
  and g_089211_(_045594_, _045638_, _047541_);
  or g_089212_(_045583_, _045627_, _047552_);
  and g_089213_(_047530_, _047552_, _047563_);
  or g_089214_(_047519_, _047541_, _047574_);
  and g_089215_(_047486_, _047563_, _047585_);
  or g_089216_(_047475_, _047574_, _047596_);
  and g_089217_(_047376_, _047585_, _047607_);
  or g_089218_(_047365_, _047596_, _047618_);
  and g_089219_(_047244_, _047618_, _047629_);
  or g_089220_(_047233_, _047607_, _047640_);
  and g_089221_(_045506_, _047640_, _047651_);
  or g_089222_(_045495_, _047629_, _047662_);
  and g_089223_(_045539_, _047629_, _047673_);
  or g_089224_(_045550_, _047640_, _047684_);
  and g_089225_(_047662_, _047684_, _047695_);
  or g_089226_(_047651_, _047673_, _047706_);
  xor g_089227_(out[227], _013122_, _047717_);
  or g_089228_(_047057_, _047629_, _047728_);
  not g_089229_(_047728_, _047739_);
  and g_089230_(_047024_, _047629_, _047750_);
  not g_089231_(_047750_, _047761_);
  and g_089232_(_047728_, _047761_, _047772_);
  or g_089233_(_047739_, _047750_, _047783_);
  and g_089234_(_047717_, _047783_, _047794_);
  or g_089235_(out[225], out[226], _047805_);
  xor g_089236_(out[225], out[226], _047816_);
  xor g_089237_(_004179_, out[226], _047827_);
  or g_089238_(_046947_, _047629_, _047838_);
  or g_089239_(_046881_, _047640_, _047849_);
  and g_089240_(_047838_, _047849_, _047860_);
  and g_089241_(_047827_, _047860_, _047871_);
  or g_089242_(_047794_, _047871_, _047882_);
  or g_089243_(_047717_, _047783_, _047893_);
  xor g_089244_(_047717_, _047783_, _047904_);
  xor g_089245_(_047717_, _047772_, _047915_);
  xor g_089246_(_047827_, _047860_, _047926_);
  xor g_089247_(_047816_, _047860_, _047937_);
  and g_089248_(_047904_, _047926_, _047948_);
  or g_089249_(_047915_, _047937_, _047959_);
  and g_089250_(out[209], _047629_, _047970_);
  and g_089251_(_046727_, _047640_, _047981_);
  or g_089252_(_047970_, _047981_, _047992_);
  or g_089253_(_004179_, _047992_, _048003_);
  and g_089254_(_004058_, _047629_, _048014_);
  not g_089255_(_048014_, _048025_);
  or g_089256_(_046760_, _047629_, _048036_);
  not g_089257_(_048036_, _048047_);
  and g_089258_(_048025_, _048036_, _048058_);
  or g_089259_(_048014_, _048047_, _048069_);
  and g_089260_(out[224], _048069_, _048080_);
  or g_089261_(_004190_, _048058_, _048091_);
  xor g_089262_(_004179_, _047992_, _048102_);
  xor g_089263_(out[225], _047992_, _048113_);
  and g_089264_(_048091_, _048102_, _048124_);
  or g_089265_(_048080_, _048113_, _048135_);
  and g_089266_(_048003_, _048135_, _048146_);
  or g_089267_(_047959_, _048146_, _048157_);
  and g_089268_(_047882_, _047893_, _048168_);
  not g_089269_(_048168_, _048179_);
  and g_089270_(_048157_, _048179_, _048190_);
  and g_089271_(_013100_, _013243_, _048201_);
  or g_089272_(_013111_, _013232_, _048212_);
  xor g_089273_(out[234], _013210_, _048223_);
  xor g_089274_(_004234_, _013210_, _048234_);
  and g_089275_(_047695_, _048223_, _048245_);
  or g_089276_(_047706_, _048234_, _048256_);
  and g_089277_(_048212_, _048256_, _048267_);
  or g_089278_(_048201_, _048245_, _048278_);
  and g_089279_(_013111_, _013232_, _048289_);
  or g_089280_(_013100_, _013243_, _048300_);
  and g_089281_(_047706_, _048234_, _048311_);
  not g_089282_(_048311_, _048322_);
  or g_089283_(_048289_, _048311_, _048333_);
  and g_089284_(_048267_, _048322_, _048344_);
  and g_089285_(_048300_, _048344_, _048355_);
  or g_089286_(_048278_, _048333_, _048366_);
  xor g_089287_(out[233], _013199_, _048377_);
  not g_089288_(_048377_, _048388_);
  and g_089289_(_045814_, _047629_, _048399_);
  not g_089290_(_048399_, _048410_);
  or g_089291_(_045847_, _047629_, _048421_);
  not g_089292_(_048421_, _048432_);
  and g_089293_(_048410_, _048421_, _048443_);
  or g_089294_(_048399_, _048432_, _048454_);
  or g_089295_(_048388_, _048443_, _048465_);
  xor g_089296_(out[232], _013188_, _048476_);
  not g_089297_(_048476_, _048487_);
  and g_089298_(_045693_, _047629_, _048498_);
  not g_089299_(_048498_, _048509_);
  or g_089300_(_045759_, _047629_, _048520_);
  not g_089301_(_048520_, _048531_);
  and g_089302_(_048509_, _048520_, _048542_);
  or g_089303_(_048498_, _048531_, _048553_);
  or g_089304_(_048487_, _048553_, _048564_);
  and g_089305_(_048465_, _048564_, _048575_);
  or g_089306_(_048476_, _048542_, _048586_);
  not g_089307_(_048586_, _048597_);
  or g_089308_(_048377_, _048454_, _048608_);
  not g_089309_(_048608_, _048619_);
  xor g_089310_(out[231], _013177_, _048630_);
  xor g_089311_(_004135_, _013177_, _048641_);
  and g_089312_(_046122_, _047629_, _048652_);
  and g_089313_(_046188_, _047640_, _048663_);
  or g_089314_(_048652_, _048663_, _048674_);
  not g_089315_(_048674_, _048685_);
  and g_089316_(_048630_, _048685_, _048696_);
  or g_089317_(_048641_, _048674_, _048707_);
  and g_089318_(_046100_, _047629_, _048718_);
  or g_089319_(_046089_, _047640_, _048729_);
  or g_089320_(_046067_, _047629_, _048740_);
  not g_089321_(_048740_, _048751_);
  and g_089322_(_048729_, _048740_, _048762_);
  or g_089323_(_048718_, _048751_, _048773_);
  xor g_089324_(out[230], _013166_, _048784_);
  not g_089325_(_048784_, _048795_);
  and g_089326_(_048762_, _048795_, _048806_);
  or g_089327_(_048773_, _048784_, _048817_);
  and g_089328_(_048641_, _048674_, _048828_);
  or g_089329_(_048630_, _048685_, _048839_);
  and g_089330_(_048817_, _048839_, _048850_);
  or g_089331_(_048806_, _048828_, _048861_);
  and g_089332_(_048773_, _048784_, _048872_);
  not g_089333_(_048872_, _048883_);
  and g_089334_(_048850_, _048883_, _048894_);
  or g_089335_(_048861_, _048872_, _048905_);
  xor g_089336_(out[228], _013144_, _048916_);
  xor g_089337_(_004168_, _013144_, _048927_);
  and g_089338_(_046408_, _047629_, _048938_);
  not g_089339_(_048938_, _048949_);
  and g_089340_(_046485_, _047640_, _048960_);
  or g_089341_(_046474_, _047629_, _048971_);
  and g_089342_(_048949_, _048971_, _048982_);
  or g_089343_(_048938_, _048960_, _048993_);
  and g_089344_(_048916_, _048982_, _049004_);
  or g_089345_(_048927_, _048993_, _049015_);
  xor g_089346_(out[229], _013155_, _049026_);
  not g_089347_(_049026_, _049037_);
  and g_089348_(_046309_, _047629_, _049048_);
  or g_089349_(_046298_, _047640_, _049059_);
  or g_089350_(_046364_, _047629_, _049070_);
  not g_089351_(_049070_, _049081_);
  and g_089352_(_049059_, _049070_, _049092_);
  or g_089353_(_049048_, _049081_, _049103_);
  and g_089354_(_049026_, _049103_, _049114_);
  or g_089355_(_049037_, _049092_, _049125_);
  and g_089356_(_049015_, _049125_, _049136_);
  or g_089357_(_049004_, _049114_, _049147_);
  and g_089358_(_049037_, _049092_, _049158_);
  or g_089359_(_049026_, _049103_, _049169_);
  or g_089360_(_048916_, _048982_, _049180_);
  and g_089361_(_049169_, _049180_, _049191_);
  not g_089362_(_049191_, _049202_);
  and g_089363_(_049136_, _049191_, _049213_);
  or g_089364_(_049147_, _049202_, _049224_);
  and g_089365_(_048575_, _048608_, _049235_);
  not g_089366_(_049235_, _049246_);
  and g_089367_(_048355_, _048586_, _049257_);
  or g_089368_(_048366_, _048597_, _049268_);
  and g_089369_(_049235_, _049257_, _049279_);
  or g_089370_(_049246_, _049268_, _049290_);
  and g_089371_(_048707_, _048894_, _049301_);
  or g_089372_(_048696_, _048905_, _049312_);
  and g_089373_(_049213_, _049301_, _049323_);
  or g_089374_(_049224_, _049312_, _049334_);
  and g_089375_(_049279_, _049323_, _049345_);
  or g_089376_(_049290_, _049334_, _049356_);
  or g_089377_(_048190_, _049356_, _049367_);
  or g_089378_(_049136_, _049158_, _049378_);
  or g_089379_(_048905_, _049378_, _049389_);
  and g_089380_(_048850_, _049389_, _049400_);
  or g_089381_(_048696_, _049400_, _049411_);
  or g_089382_(_049290_, _049411_, _049422_);
  or g_089383_(_048267_, _048289_, _049433_);
  or g_089384_(_048366_, _048575_, _049444_);
  or g_089385_(_048619_, _049444_, _049455_);
  and g_089386_(_049433_, _049455_, _049466_);
  and g_089387_(_049422_, _049466_, _049477_);
  and g_089388_(_049367_, _049477_, _049488_);
  or g_089389_(out[224], _048069_, _049499_);
  and g_089390_(_047948_, _049499_, _049510_);
  and g_089391_(_048124_, _049510_, _049521_);
  and g_089392_(_049345_, _049521_, _049532_);
  or g_089393_(_049488_, _049532_, _049543_);
  not g_089394_(_049543_, _049554_);
  and g_089395_(_047706_, _049543_, _049565_);
  not g_089396_(_049565_, _049576_);
  and g_089397_(_048223_, _049554_, _049587_);
  or g_089398_(_048234_, _049543_, _049598_);
  and g_089399_(_049576_, _049598_, _049609_);
  or g_089400_(_049565_, _049587_, _049620_);
  or g_089401_(_013265_, _013375_, _049631_);
  xor g_089402_(out[250], _013353_, _049642_);
  not g_089403_(_049642_, _049653_);
  or g_089404_(_049620_, _049653_, _049664_);
  and g_089405_(_049631_, _049664_, _049675_);
  xor g_089406_(out[249], _013342_, _049686_);
  or g_089407_(_048377_, _049543_, _049697_);
  not g_089408_(_049697_, _049708_);
  and g_089409_(_048454_, _049543_, _049719_);
  or g_089410_(_048443_, _049554_, _049730_);
  and g_089411_(_049697_, _049730_, _049741_);
  or g_089412_(_049708_, _049719_, _049752_);
  or g_089413_(_049686_, _049752_, _049763_);
  and g_089414_(_049686_, _049752_, _049774_);
  xor g_089415_(_049686_, _049752_, _049785_);
  xor g_089416_(_049686_, _049741_, _049796_);
  xor g_089417_(out[248], _013331_, _049807_);
  not g_089418_(_049807_, _049818_);
  or g_089419_(_048487_, _049543_, _049829_);
  or g_089420_(_048542_, _049554_, _049840_);
  and g_089421_(_049829_, _049840_, _049851_);
  and g_089422_(_049807_, _049851_, _049862_);
  xor g_089423_(_049807_, _049851_, _049873_);
  xor g_089424_(_049818_, _049851_, _049884_);
  and g_089425_(_049785_, _049873_, _049895_);
  or g_089426_(_049796_, _049884_, _049906_);
  xor g_089427_(out[247], _013320_, _049917_);
  and g_089428_(_048630_, _049554_, _049928_);
  or g_089429_(_048641_, _049543_, _049939_);
  and g_089430_(_048674_, _049543_, _049950_);
  not g_089431_(_049950_, _049961_);
  and g_089432_(_049939_, _049961_, _049972_);
  or g_089433_(_049928_, _049950_, _049983_);
  or g_089434_(_049917_, _049972_, _049994_);
  and g_089435_(_049917_, _049972_, _050005_);
  xor g_089436_(_049917_, _049972_, _050016_);
  xor g_089437_(_049917_, _049983_, _050027_);
  and g_089438_(_048795_, _049554_, _050038_);
  and g_089439_(_048773_, _049543_, _050049_);
  or g_089440_(_050038_, _050049_, _050060_);
  not g_089441_(_050060_, _050071_);
  xor g_089442_(out[246], _013309_, _050082_);
  or g_089443_(_050060_, _050082_, _050093_);
  xor g_089444_(_050060_, _050082_, _050104_);
  xor g_089445_(_050071_, _050082_, _050115_);
  xor g_089446_(out[245], _013298_, _050126_);
  xor g_089447_(_004278_, _013298_, _050137_);
  or g_089448_(_049026_, _049543_, _050148_);
  or g_089449_(_049092_, _049554_, _050159_);
  and g_089450_(_050148_, _050159_, _050170_);
  not g_089451_(_050170_, _050181_);
  and g_089452_(_050137_, _050170_, _050192_);
  or g_089453_(_050126_, _050181_, _050203_);
  and g_089454_(_050104_, _050203_, _050214_);
  or g_089455_(_050027_, _050192_, _050225_);
  and g_089456_(_050016_, _050214_, _050236_);
  or g_089457_(_050115_, _050225_, _050247_);
  xor g_089458_(out[244], _013287_, _050258_);
  not g_089459_(_050258_, _050269_);
  and g_089460_(_048916_, _049554_, _050280_);
  and g_089461_(_048993_, _049543_, _050291_);
  or g_089462_(_050280_, _050291_, _050302_);
  not g_089463_(_050302_, _050313_);
  or g_089464_(_050269_, _050302_, _050324_);
  or g_089465_(_050137_, _050170_, _050335_);
  and g_089466_(_050324_, _050335_, _050346_);
  xor g_089467_(out[243], _013276_, _050357_);
  not g_089468_(_050357_, _050368_);
  and g_089469_(_047783_, _049543_, _050379_);
  or g_089470_(_047772_, _049554_, _050390_);
  or g_089471_(_047717_, _049543_, _050401_);
  not g_089472_(_050401_, _050412_);
  and g_089473_(_050390_, _050401_, _050423_);
  or g_089474_(_050379_, _050412_, _050434_);
  and g_089475_(_050368_, _050423_, _050445_);
  or g_089476_(_050368_, _050423_, _050456_);
  or g_089477_(out[241], out[242], _050467_);
  xor g_089478_(out[241], out[242], _050478_);
  xor g_089479_(_053038_, out[242], _050489_);
  and g_089480_(_047860_, _049543_, _050500_);
  not g_089481_(_050500_, _050511_);
  or g_089482_(_047827_, _049543_, _050522_);
  not g_089483_(_050522_, _050533_);
  or g_089484_(_050500_, _050533_, _050544_);
  and g_089485_(_050511_, _050522_, _050555_);
  or g_089486_(_050478_, _050555_, _050566_);
  and g_089487_(_050456_, _050566_, _050577_);
  or g_089488_(_050445_, _050577_, _050588_);
  xor g_089489_(_050368_, _050423_, _050599_);
  xor g_089490_(_050357_, _050423_, _050610_);
  xor g_089491_(_050489_, _050544_, _050621_);
  xor g_089492_(_050478_, _050544_, _050632_);
  and g_089493_(_050599_, _050621_, _050643_);
  or g_089494_(_050610_, _050632_, _050654_);
  and g_089495_(out[225], _049554_, _050665_);
  and g_089496_(_047992_, _049543_, _050676_);
  or g_089497_(_050665_, _050676_, _050687_);
  not g_089498_(_050687_, _050698_);
  or g_089499_(_053038_, _050687_, _050709_);
  and g_089500_(_048069_, _049543_, _050720_);
  and g_089501_(_004190_, _049554_, _050731_);
  or g_089502_(_050720_, _050731_, _050742_);
  and g_089503_(out[240], _050742_, _050753_);
  not g_089504_(_050753_, _050764_);
  and g_089505_(_053038_, _050687_, _050775_);
  or g_089506_(out[241], _050698_, _050786_);
  and g_089507_(_050764_, _050786_, _050797_);
  or g_089508_(_050753_, _050775_, _050808_);
  and g_089509_(_050709_, _050808_, _050819_);
  or g_089510_(_050654_, _050819_, _050830_);
  and g_089511_(_050588_, _050830_, _050841_);
  and g_089512_(_050269_, _050302_, _050852_);
  or g_089513_(_050258_, _050313_, _050863_);
  or g_089514_(_050841_, _050852_, _050874_);
  and g_089515_(_050346_, _050874_, _050885_);
  or g_089516_(_050247_, _050885_, _050896_);
  and g_089517_(_049994_, _050093_, _050907_);
  or g_089518_(_050005_, _050907_, _050918_);
  and g_089519_(_050896_, _050918_, _050929_);
  or g_089520_(_049906_, _050929_, _050940_);
  and g_089521_(_049763_, _049862_, _050951_);
  or g_089522_(_049774_, _050951_, _050962_);
  not g_089523_(_050962_, _050973_);
  and g_089524_(_050940_, _050973_, _050984_);
  and g_089525_(_049620_, _049653_, _050995_);
  or g_089526_(_049609_, _049642_, _051006_);
  or g_089527_(_050984_, _050995_, _051017_);
  and g_089528_(_049675_, _051017_, _051028_);
  and g_089529_(_013265_, _013375_, _051039_);
  and g_089530_(_050709_, _050863_, _051050_);
  or g_089531_(out[240], _050742_, _051061_);
  and g_089532_(_051006_, _051061_, _051072_);
  and g_089533_(_051050_, _051072_, _051083_);
  and g_089534_(_049895_, _051083_, _051094_);
  and g_089535_(_050643_, _051094_, _051105_);
  and g_089536_(_049675_, _050346_, _051116_);
  and g_089537_(_050797_, _051116_, _051127_);
  and g_089538_(_050236_, _051127_, _051138_);
  and g_089539_(_051105_, _051138_, _051149_);
  or g_089540_(_051039_, _051149_, _051160_);
  or g_089541_(_051028_, _051160_, _051171_);
  not g_089542_(_051171_, _051182_);
  and g_089543_(_049620_, _051171_, _051193_);
  or g_089544_(_049609_, _051182_, _051204_);
  and g_089545_(_049642_, _051182_, _051215_);
  or g_089546_(_049653_, _051171_, _051226_);
  and g_089547_(_051204_, _051226_, _051237_);
  or g_089548_(_051193_, _051215_, _051248_);
  xor g_089549_(out[265], _013496_, _051259_);
  xor g_089550_(_004410_, _013496_, _051270_);
  or g_089551_(_049686_, _051171_, _051281_);
  not g_089552_(_051281_, _051292_);
  and g_089553_(_049752_, _051171_, _051303_);
  or g_089554_(_049741_, _051182_, _051314_);
  and g_089555_(_051281_, _051314_, _051325_);
  or g_089556_(_051292_, _051303_, _051336_);
  and g_089557_(_051259_, _051336_, _051347_);
  xor g_089558_(out[264], _013485_, _051357_);
  and g_089559_(_049851_, _051171_, _051361_);
  not g_089560_(_051361_, _051362_);
  or g_089561_(_049807_, _051171_, _051363_);
  not g_089562_(_051363_, _051364_);
  or g_089563_(_051361_, _051364_, _051365_);
  and g_089564_(_051362_, _051363_, _051366_);
  and g_089565_(_051357_, _051365_, _051367_);
  or g_089566_(_051347_, _051367_, _051368_);
  xor g_089567_(out[263], _013474_, _051369_);
  xor g_089568_(_004377_, _013474_, _051370_);
  and g_089569_(_049972_, _051171_, _051371_);
  or g_089570_(_049983_, _051182_, _051372_);
  or g_089571_(_049917_, _051171_, _051373_);
  not g_089572_(_051373_, _051374_);
  or g_089573_(_051371_, _051374_, _051375_);
  and g_089574_(_051372_, _051373_, _051376_);
  and g_089575_(_051369_, _051375_, _051377_);
  or g_089576_(_051370_, _051376_, _051378_);
  and g_089577_(_051370_, _051376_, _051379_);
  or g_089578_(_051369_, _051375_, _051380_);
  or g_089579_(_050082_, _051171_, _051381_);
  or g_089580_(_050071_, _051182_, _051382_);
  and g_089581_(_051381_, _051382_, _051383_);
  not g_089582_(_051383_, _051384_);
  xor g_089583_(out[262], _013463_, _051385_);
  not g_089584_(_051385_, _051386_);
  and g_089585_(_051383_, _051386_, _051387_);
  or g_089586_(_051384_, _051385_, _051388_);
  and g_089587_(_051380_, _051388_, _051389_);
  or g_089588_(_051379_, _051387_, _051390_);
  and g_089589_(_051378_, _051390_, _051391_);
  or g_089590_(_051377_, _051389_, _051392_);
  and g_089591_(_051378_, _051380_, _051393_);
  or g_089592_(_051377_, _051379_, _051394_);
  xor g_089593_(out[261], _013452_, _051395_);
  xor g_089594_(_052972_, _013452_, _051396_);
  or g_089595_(_050126_, _051171_, _051397_);
  not g_089596_(_051397_, _051398_);
  and g_089597_(_050181_, _051171_, _051399_);
  or g_089598_(_050170_, _051182_, _051400_);
  and g_089599_(_051397_, _051400_, _051401_);
  or g_089600_(_051398_, _051399_, _051402_);
  and g_089601_(_051396_, _051401_, _051403_);
  or g_089602_(_051395_, _051402_, _051404_);
  xor g_089603_(_051383_, _051386_, _051405_);
  xor g_089604_(_051383_, _051385_, _051406_);
  and g_089605_(_051404_, _051405_, _051407_);
  or g_089606_(_051403_, _051406_, _051408_);
  and g_089607_(_051393_, _051407_, _051409_);
  or g_089608_(_051394_, _051408_, _051410_);
  and g_089609_(_051395_, _051402_, _051411_);
  or g_089610_(_051396_, _051401_, _051412_);
  xor g_089611_(out[260], _013441_, _051413_);
  xor g_089612_(_052994_, _013441_, _051414_);
  and g_089613_(_050258_, _051182_, _051415_);
  or g_089614_(_050269_, _051171_, _051416_);
  and g_089615_(_050302_, _051171_, _051417_);
  not g_089616_(_051417_, _051418_);
  and g_089617_(_051416_, _051418_, _051419_);
  or g_089618_(_051415_, _051417_, _051420_);
  and g_089619_(_051413_, _051419_, _051421_);
  or g_089620_(_051414_, _051420_, _051422_);
  and g_089621_(_051412_, _051422_, _051423_);
  or g_089622_(_051411_, _051421_, _051424_);
  or g_089623_(out[258], out[257], _051425_);
  and g_089624_(_013430_, _051425_, _051426_);
  xor g_089625_(_053016_, out[257], _051427_);
  or g_089626_(_050489_, _051171_, _051428_);
  not g_089627_(_051428_, _051429_);
  and g_089628_(_050544_, _051171_, _051430_);
  not g_089629_(_051430_, _051431_);
  or g_089630_(_051429_, _051430_, _051432_);
  and g_089631_(_051428_, _051431_, _051433_);
  and g_089632_(_051427_, _051432_, _051434_);
  or g_089633_(_051426_, _051433_, _051435_);
  xor g_089634_(out[259], _013419_, _051436_);
  xor g_089635_(_053005_, _013419_, _051437_);
  and g_089636_(_050434_, _051171_, _051438_);
  or g_089637_(_050423_, _051182_, _051439_);
  or g_089638_(_050357_, _051171_, _051440_);
  not g_089639_(_051440_, _051441_);
  and g_089640_(_051439_, _051440_, _051442_);
  or g_089641_(_051438_, _051441_, _051443_);
  and g_089642_(_051436_, _051443_, _051444_);
  or g_089643_(_051437_, _051442_, _051445_);
  and g_089644_(_051435_, _051445_, _051446_);
  or g_089645_(_051434_, _051444_, _051447_);
  and g_089646_(_051437_, _051442_, _051448_);
  or g_089647_(_051436_, _051443_, _051449_);
  and g_089648_(_051414_, _051420_, _051450_);
  or g_089649_(_051413_, _051419_, _051451_);
  xor g_089650_(out[266], _013507_, _051452_);
  and g_089651_(_051237_, _051452_, _051453_);
  and g_089652_(_013397_, _013529_, _051454_);
  or g_089653_(_051453_, _051454_, _051455_);
  or g_089654_(_013397_, _013529_, _051456_);
  xor g_089655_(_051237_, _051452_, _051457_);
  xor g_089656_(_051248_, _051452_, _051458_);
  xor g_089657_(_013408_, _013540_, _051459_);
  xor g_089658_(_013397_, _013540_, _051460_);
  and g_089659_(_051457_, _051459_, _051461_);
  or g_089660_(_051458_, _051460_, _051462_);
  or g_089661_(_051259_, _051336_, _051463_);
  and g_089662_(_051455_, _051456_, _051464_);
  not g_089663_(_051464_, _051465_);
  and g_089664_(_051445_, _051449_, _051466_);
  or g_089665_(_051444_, _051448_, _051467_);
  xor g_089666_(_051357_, _051365_, _051468_);
  xor g_089667_(_051357_, _051366_, _051469_);
  xor g_089668_(_051270_, _051325_, _051470_);
  xor g_089669_(_051259_, _051325_, _051471_);
  and g_089670_(_051461_, _051470_, _051472_);
  or g_089671_(_051462_, _051471_, _051473_);
  and g_089672_(_051468_, _051472_, _051474_);
  or g_089673_(_051469_, _051473_, _051475_);
  and g_089674_(_051423_, _051451_, _051476_);
  or g_089675_(_051424_, _051450_, _051477_);
  or g_089676_(_051410_, _051477_, _051478_);
  and g_089677_(_051474_, _051476_, _051479_);
  and g_089678_(_051409_, _051479_, _051480_);
  or g_089679_(_051475_, _051478_, _051481_);
  xor g_089680_(_051427_, _051432_, _051482_);
  xor g_089681_(_051426_, _051432_, _051483_);
  and g_089682_(_051466_, _051480_, _051484_);
  or g_089683_(_051467_, _051481_, _051485_);
  and g_089684_(_051482_, _051484_, _051486_);
  or g_089685_(_051483_, _051485_, _051487_);
  and g_089686_(out[241], _051182_, _051488_);
  or g_089687_(_053038_, _051171_, _051489_);
  and g_089688_(_050687_, _051171_, _051490_);
  not g_089689_(_051490_, _051491_);
  and g_089690_(_051489_, _051491_, _051492_);
  or g_089691_(_051488_, _051490_, _051493_);
  and g_089692_(out[257], _051492_, _051494_);
  or g_089693_(_053027_, _051493_, _051495_);
  and g_089694_(_051486_, _051494_, _051496_);
  or g_089695_(_051487_, _051495_, _051497_);
  and g_089696_(_051409_, _051424_, _051498_);
  or g_089697_(_051410_, _051423_, _051499_);
  and g_089698_(_051392_, _051499_, _051500_);
  or g_089699_(_051391_, _051498_, _051501_);
  and g_089700_(_051474_, _051501_, _051502_);
  or g_089701_(_051475_, _051500_, _051503_);
  and g_089702_(_051368_, _051461_, _051504_);
  and g_089703_(_051463_, _051504_, _051505_);
  not g_089704_(_051505_, _051506_);
  and g_089705_(_051503_, _051506_, _051507_);
  or g_089706_(_051502_, _051505_, _051508_);
  or g_089707_(_051446_, _051448_, _051509_);
  and g_089708_(_051447_, _051449_, _051510_);
  and g_089709_(_051480_, _051510_, _051511_);
  or g_089710_(_051481_, _051509_, _051512_);
  and g_089711_(_051465_, _051512_, _051513_);
  or g_089712_(_051464_, _051511_, _051514_);
  and g_089713_(_051507_, _051513_, _051515_);
  or g_089714_(_051508_, _051514_, _051516_);
  and g_089715_(_051497_, _051515_, _051517_);
  or g_089716_(_051496_, _051516_, _051518_);
  and g_089717_(_050742_, _051171_, _051519_);
  not g_089718_(_051519_, _051520_);
  or g_089719_(out[240], _051171_, _051521_);
  not g_089720_(_051521_, _051522_);
  and g_089721_(_051520_, _051521_, _051523_);
  or g_089722_(_051519_, _051522_, _051524_);
  and g_089723_(out[256], _051524_, _051525_);
  xor g_089724_(_053027_, _051492_, _051526_);
  or g_089725_(_051525_, _051526_, _051527_);
  not g_089726_(_051527_, _051528_);
  and g_089727_(_051486_, _051528_, _051529_);
  or g_089728_(_051487_, _051527_, _051530_);
  and g_089729_(_004388_, _051523_, _051531_);
  or g_089730_(out[256], _051524_, _051532_);
  and g_089731_(_051529_, _051531_, _051533_);
  or g_089732_(_051530_, _051532_, _051534_);
  and g_089733_(_051517_, _051534_, _051535_);
  or g_089734_(_051518_, _051533_, _051536_);
  and g_089735_(_051248_, _051535_, _051537_);
  or g_089736_(_051237_, _051536_, _051538_);
  and g_089737_(_051452_, _051536_, _051539_);
  not g_089738_(_051539_, _051540_);
  and g_089739_(_051538_, _051540_, _051541_);
  or g_089740_(_051537_, _051539_, _051542_);
  and g_089741_(_013551_, _013694_, _051543_);
  or g_089742_(_013562_, _013683_, _051544_);
  xor g_089743_(out[282], _013661_, _051545_);
  xor g_089744_(_004454_, _013661_, _051546_);
  and g_089745_(_051541_, _051545_, _051547_);
  or g_089746_(_051542_, _051546_, _051548_);
  and g_089747_(_051544_, _051548_, _051549_);
  or g_089748_(_051543_, _051547_, _051550_);
  and g_089749_(_013562_, _013683_, _051551_);
  or g_089750_(_013551_, _013694_, _051552_);
  and g_089751_(_051542_, _051546_, _051553_);
  or g_089752_(_051541_, _051545_, _051554_);
  and g_089753_(_051552_, _051554_, _051555_);
  or g_089754_(_051551_, _051553_, _051556_);
  xor g_089755_(out[281], _013650_, _051557_);
  xor g_089756_(_053137_, _013650_, _051558_);
  and g_089757_(_051270_, _051536_, _051559_);
  or g_089758_(_051259_, _051535_, _051560_);
  and g_089759_(_051336_, _051535_, _051561_);
  or g_089760_(_051325_, _051536_, _051562_);
  and g_089761_(_051560_, _051562_, _051563_);
  or g_089762_(_051559_, _051561_, _051564_);
  and g_089763_(_051558_, _051563_, _051565_);
  or g_089764_(_051557_, _051564_, _051566_);
  or g_089765_(_051556_, _051565_, _051567_);
  and g_089766_(_051549_, _051555_, _051568_);
  and g_089767_(_051566_, _051568_, _051569_);
  or g_089768_(_051550_, _051567_, _051570_);
  xor g_089769_(out[280], _013639_, _051571_);
  xor g_089770_(_053060_, _013639_, _051572_);
  and g_089771_(_051357_, _051536_, _051573_);
  not g_089772_(_051573_, _051574_);
  and g_089773_(_051366_, _051535_, _051575_);
  or g_089774_(_051365_, _051536_, _051576_);
  and g_089775_(_051574_, _051576_, _051577_);
  or g_089776_(_051573_, _051575_, _051578_);
  and g_089777_(_051572_, _051578_, _051579_);
  or g_089778_(_051571_, _051577_, _051580_);
  and g_089779_(_051557_, _051564_, _051581_);
  or g_089780_(_051558_, _051563_, _051582_);
  and g_089781_(_051571_, _051577_, _051583_);
  or g_089782_(_051572_, _051578_, _051584_);
  and g_089783_(_051582_, _051584_, _051585_);
  or g_089784_(_051581_, _051583_, _051586_);
  and g_089785_(_051580_, _051585_, _051587_);
  or g_089786_(_051579_, _051586_, _051588_);
  and g_089787_(_051569_, _051587_, _051589_);
  or g_089788_(_051570_, _051588_, _051590_);
  xor g_089789_(out[279], _013628_, _051591_);
  xor g_089790_(_053049_, _013628_, _051592_);
  and g_089791_(_051369_, _051536_, _051593_);
  or g_089792_(_051370_, _051535_, _051594_);
  and g_089793_(_051376_, _051535_, _051595_);
  or g_089794_(_051375_, _051536_, _051596_);
  and g_089795_(_051594_, _051596_, _051597_);
  or g_089796_(_051593_, _051595_, _051598_);
  or g_089797_(_051592_, _051598_, _051599_);
  or g_089798_(_051385_, _051535_, _051600_);
  or g_089799_(_051383_, _051536_, _051601_);
  and g_089800_(_051600_, _051601_, _051602_);
  xor g_089801_(out[278], _013617_, _051603_);
  xor g_089802_(_053082_, _013617_, _051604_);
  and g_089803_(_051602_, _051604_, _051605_);
  and g_089804_(_051592_, _051598_, _051606_);
  xor g_089805_(_051591_, _051597_, _051607_);
  xor g_089806_(_051592_, _051597_, _051608_);
  xor g_089807_(_051602_, _051604_, _051609_);
  xor g_089808_(_051602_, _051603_, _051610_);
  and g_089809_(_051607_, _051609_, _051611_);
  or g_089810_(_051608_, _051610_, _051612_);
  xor g_089811_(out[276], _013595_, _051613_);
  and g_089812_(_051420_, _051535_, _051614_);
  or g_089813_(_051419_, _051536_, _051615_);
  and g_089814_(_051413_, _051536_, _051616_);
  or g_089815_(_051414_, _051535_, _051617_);
  and g_089816_(_051615_, _051617_, _051618_);
  or g_089817_(_051614_, _051616_, _051619_);
  and g_089818_(_051613_, _051618_, _051620_);
  xor g_089819_(_051613_, _051618_, _051621_);
  xor g_089820_(_051613_, _051619_, _051622_);
  xor g_089821_(out[277], _013606_, _051623_);
  and g_089822_(_051396_, _051536_, _051624_);
  or g_089823_(_051395_, _051535_, _051625_);
  and g_089824_(_051402_, _051535_, _051626_);
  or g_089825_(_051401_, _051536_, _051627_);
  and g_089826_(_051625_, _051627_, _051628_);
  or g_089827_(_051624_, _051626_, _051629_);
  and g_089828_(_051623_, _051629_, _051630_);
  or g_089829_(_051623_, _051629_, _051631_);
  xor g_089830_(_051623_, _051629_, _051632_);
  xor g_089831_(_051623_, _051628_, _051633_);
  and g_089832_(_051621_, _051632_, _051634_);
  or g_089833_(_051622_, _051633_, _051635_);
  and g_089834_(_051611_, _051634_, _051636_);
  or g_089835_(_051612_, _051635_, _051637_);
  and g_089836_(_051589_, _051636_, _051638_);
  or g_089837_(_051590_, _051637_, _051639_);
  or g_089838_(out[274], out[273], _051640_);
  xor g_089839_(out[274], out[273], _051641_);
  xor g_089840_(_053115_, out[273], _051642_);
  and g_089841_(_051427_, _051536_, _051643_);
  or g_089842_(_051426_, _051535_, _051644_);
  and g_089843_(_051433_, _051535_, _051645_);
  or g_089844_(_051432_, _051536_, _051646_);
  and g_089845_(_051644_, _051646_, _051647_);
  or g_089846_(_051643_, _051645_, _051648_);
  and g_089847_(_051642_, _051647_, _051649_);
  xor g_089848_(out[275], _013573_, _051650_);
  xor g_089849_(_053093_, _013573_, _051651_);
  and g_089850_(_051443_, _051535_, _051652_);
  or g_089851_(_051442_, _051536_, _051653_);
  and g_089852_(_051437_, _051536_, _051654_);
  or g_089853_(_051436_, _051535_, _051655_);
  and g_089854_(_051653_, _051655_, _051656_);
  or g_089855_(_051652_, _051654_, _051657_);
  and g_089856_(_051651_, _051656_, _051658_);
  or g_089857_(_051650_, _051657_, _051659_);
  or g_089858_(_051649_, _051658_, _051660_);
  and g_089859_(_051641_, _051648_, _051661_);
  and g_089860_(_051650_, _051657_, _051662_);
  or g_089861_(_051661_, _051662_, _051663_);
  or g_089862_(_051660_, _051663_, _051664_);
  xor g_089863_(_051642_, _051647_, _051665_);
  xor g_089864_(_051651_, _051656_, _051666_);
  and g_089865_(_051638_, _051666_, _051667_);
  and g_089866_(_051665_, _051667_, _051668_);
  or g_089867_(_051639_, _051664_, _051669_);
  and g_089868_(out[257], _051536_, _051670_);
  not g_089869_(_051670_, _051671_);
  and g_089870_(_051493_, _051535_, _051672_);
  or g_089871_(_051492_, _051536_, _051673_);
  and g_089872_(_051671_, _051673_, _051674_);
  or g_089873_(_051670_, _051672_, _051675_);
  and g_089874_(out[256], _051518_, _051676_);
  not g_089875_(_051676_, _051677_);
  and g_089876_(_051523_, _051535_, _051678_);
  or g_089877_(_051524_, _051536_, _051679_);
  and g_089878_(_051677_, _051679_, _051680_);
  or g_089879_(_051676_, _051678_, _051681_);
  and g_089880_(out[272], _051680_, _051682_);
  or g_089881_(_004443_, _051681_, _051683_);
  and g_089882_(out[273], _051674_, _051684_);
  xor g_089883_(_053126_, _051675_, _051685_);
  xor g_089884_(out[273], _051675_, _051686_);
  and g_089885_(_051683_, _051685_, _051687_);
  or g_089886_(_051682_, _051686_, _051688_);
  and g_089887_(_004443_, _051681_, _051689_);
  or g_089888_(_051688_, _051689_, _051690_);
  or g_089889_(_051669_, _051690_, _051691_);
  or g_089890_(_051684_, _051687_, _051692_);
  and g_089891_(_051668_, _051692_, _051693_);
  or g_089892_(_051649_, _051662_, _051694_);
  and g_089893_(_051659_, _051694_, _051695_);
  and g_089894_(_051638_, _051695_, _051696_);
  or g_089895_(_051620_, _051630_, _051697_);
  and g_089896_(_051611_, _051697_, _051698_);
  and g_089897_(_051631_, _051698_, _051699_);
  or g_089898_(_051605_, _051606_, _051700_);
  and g_089899_(_051599_, _051700_, _051701_);
  or g_089900_(_051699_, _051701_, _051702_);
  and g_089901_(_051589_, _051702_, _051703_);
  and g_089902_(_051569_, _051586_, _051704_);
  and g_089903_(_051550_, _051552_, _051705_);
  or g_089904_(_051704_, _051705_, _051706_);
  or g_089905_(_051703_, _051706_, _051707_);
  or g_089906_(_051696_, _051707_, _051708_);
  or g_089907_(_051693_, _051708_, _051709_);
  and g_089908_(_051691_, _051709_, _051710_);
  not g_089909_(_051710_, _051711_);
  and g_089910_(_051542_, _051711_, _051712_);
  or g_089911_(_051541_, _051710_, _051713_);
  and g_089912_(_051545_, _051710_, _051714_);
  or g_089913_(_051546_, _051711_, _051715_);
  and g_089914_(_051713_, _051715_, _051716_);
  or g_089915_(_051712_, _051714_, _051717_);
  and g_089916_(_026366_, _051716_, _051718_);
  or g_089917_(_026377_, _051717_, _051719_);
  and g_089918_(_026399_, _051719_, _051720_);
  or g_089919_(_026388_, _051718_, _051721_);
  and g_089920_(_013716_, _013837_, _051722_);
  or g_089921_(_013705_, _013848_, _051723_);
  and g_089922_(_026377_, _051717_, _051724_);
  or g_089923_(_026366_, _051716_, _051725_);
  and g_089924_(_051723_, _051725_, _051726_);
  or g_089925_(_051722_, _051724_, _051727_);
  xor g_089926_(out[297], _013804_, _051728_);
  xor g_089927_(_053236_, _013804_, _051729_);
  or g_089928_(_051557_, _051711_, _051730_);
  or g_089929_(_051563_, _051710_, _051731_);
  and g_089930_(_051730_, _051731_, _051732_);
  not g_089931_(_051732_, _051733_);
  and g_089932_(_051729_, _051732_, _051734_);
  or g_089933_(_051728_, _051733_, _051735_);
  and g_089934_(_051726_, _051735_, _051736_);
  and g_089935_(_051720_, _051736_, _051737_);
  xor g_089936_(out[296], _013793_, _051738_);
  not g_089937_(_051738_, _051739_);
  and g_089938_(_051571_, _051710_, _051740_);
  not g_089939_(_051740_, _051741_);
  and g_089940_(_051578_, _051711_, _051742_);
  or g_089941_(_051577_, _051710_, _051743_);
  and g_089942_(_051741_, _051743_, _051744_);
  or g_089943_(_051740_, _051742_, _051745_);
  and g_089944_(_051739_, _051745_, _051746_);
  or g_089945_(_051738_, _051744_, _051747_);
  and g_089946_(_051728_, _051733_, _051748_);
  or g_089947_(_051729_, _051732_, _051749_);
  and g_089948_(_051738_, _051744_, _051750_);
  or g_089949_(_051739_, _051745_, _051751_);
  and g_089950_(_051749_, _051751_, _051752_);
  or g_089951_(_051748_, _051750_, _051753_);
  and g_089952_(_051747_, _051752_, _051754_);
  or g_089953_(_051734_, _051753_, _051755_);
  or g_089954_(_051721_, _051727_, _051756_);
  or g_089955_(_051746_, _051756_, _051757_);
  and g_089956_(_051737_, _051754_, _051758_);
  or g_089957_(_051755_, _051757_, _051759_);
  xor g_089958_(out[294], _013771_, _051760_);
  or g_089959_(_051603_, _051711_, _051761_);
  or g_089960_(_051602_, _051710_, _051762_);
  and g_089961_(_051761_, _051762_, _051763_);
  not g_089962_(_051763_, _051764_);
  or g_089963_(_051760_, _051764_, _051765_);
  xor g_089964_(out[295], _013782_, _051766_);
  and g_089965_(_051591_, _051710_, _051767_);
  not g_089966_(_051767_, _051768_);
  and g_089967_(_051598_, _051711_, _051769_);
  or g_089968_(_051597_, _051710_, _051770_);
  and g_089969_(_051768_, _051770_, _051771_);
  or g_089970_(_051767_, _051769_, _051772_);
  or g_089971_(_051766_, _051771_, _051773_);
  and g_089972_(_051765_, _051773_, _051774_);
  and g_089973_(_051766_, _051771_, _051775_);
  xor g_089974_(_051760_, _051764_, _051776_);
  xor g_089975_(_051760_, _051763_, _051777_);
  xor g_089976_(_051766_, _051771_, _051778_);
  xor g_089977_(_051766_, _051772_, _051779_);
  and g_089978_(_051776_, _051778_, _051780_);
  or g_089979_(_051777_, _051779_, _051781_);
  xor g_089980_(out[292], _013749_, _051782_);
  not g_089981_(_051782_, _051783_);
  and g_089982_(_051613_, _051710_, _051784_);
  not g_089983_(_051784_, _051785_);
  and g_089984_(_051619_, _051711_, _051786_);
  or g_089985_(_051618_, _051710_, _051787_);
  and g_089986_(_051785_, _051787_, _051788_);
  or g_089987_(_051784_, _051786_, _051789_);
  or g_089988_(_051783_, _051789_, _051790_);
  xor g_089989_(out[293], _013760_, _051791_);
  xor g_089990_(_053170_, _013760_, _051792_);
  or g_089991_(_051623_, _051711_, _051793_);
  or g_089992_(_051628_, _051710_, _051794_);
  and g_089993_(_051793_, _051794_, _051795_);
  or g_089994_(_051792_, _051795_, _051796_);
  and g_089995_(_051790_, _051796_, _051797_);
  and g_089996_(_051792_, _051795_, _051798_);
  not g_089997_(_051798_, _051799_);
  or g_089998_(_051782_, _051788_, _051800_);
  and g_089999_(_051799_, _051800_, _051801_);
  and g_090000_(_051797_, _051801_, _051802_);
  and g_090001_(_051780_, _051802_, _051803_);
  xor g_090002_(_051791_, _051795_, _051804_);
  xor g_090003_(_051783_, _051788_, _051805_);
  or g_090004_(_051781_, _051805_, _051806_);
  or g_090005_(_051759_, _051806_, _051807_);
  and g_090006_(_051758_, _051803_, _051808_);
  or g_090007_(_051804_, _051807_, _051809_);
  xor g_090008_(_053192_, _013727_, _051810_);
  or g_090009_(_051656_, _051710_, _051811_);
  or g_090010_(_051650_, _051711_, _051812_);
  and g_090011_(_051811_, _051812_, _051813_);
  or g_090012_(_051810_, _051813_, _051814_);
  or g_090013_(out[290], out[289], _051815_);
  xor g_090014_(out[290], out[289], _051816_);
  xor g_090015_(_053214_, out[289], _051817_);
  and g_090016_(_051648_, _051711_, _051818_);
  or g_090017_(_051647_, _051710_, _051819_);
  and g_090018_(_051642_, _051710_, _051820_);
  not g_090019_(_051820_, _051821_);
  and g_090020_(_051819_, _051821_, _051822_);
  or g_090021_(_051818_, _051820_, _051823_);
  and g_090022_(_051810_, _051813_, _051824_);
  or g_090023_(_051816_, _051823_, _051825_);
  xor g_090024_(_051810_, _051813_, _051826_);
  xor g_090025_(_051817_, _051822_, _051827_);
  and g_090026_(_051826_, _051827_, _051828_);
  or g_090027_(_053126_, _051711_, _051829_);
  or g_090028_(_051674_, _051710_, _051830_);
  and g_090029_(_051829_, _051830_, _051831_);
  and g_090030_(out[289], _051831_, _051832_);
  and g_090031_(_004443_, _051710_, _051833_);
  or g_090032_(out[272], _051711_, _051834_);
  and g_090033_(_051680_, _051711_, _051835_);
  or g_090034_(_051681_, _051710_, _051836_);
  and g_090035_(_051834_, _051836_, _051837_);
  or g_090036_(_051833_, _051835_, _051838_);
  or g_090037_(_004476_, _051837_, _051839_);
  xor g_090038_(out[289], _051831_, _051840_);
  and g_090039_(_051839_, _051840_, _051841_);
  or g_090040_(_051832_, _051841_, _051842_);
  and g_090041_(_051828_, _051842_, _051843_);
  or g_090042_(_051824_, _051825_, _051844_);
  and g_090043_(_051814_, _051844_, _051845_);
  not g_090044_(_051845_, _051846_);
  or g_090045_(_051843_, _051846_, _051847_);
  not g_090046_(_051847_, _051848_);
  and g_090047_(_051808_, _051847_, _051849_);
  or g_090048_(_051809_, _051848_, _051850_);
  or g_090049_(_051781_, _051797_, _051851_);
  or g_090050_(_051798_, _051851_, _051852_);
  or g_090051_(_051774_, _051775_, _051853_);
  and g_090052_(_051852_, _051853_, _051854_);
  or g_090053_(_051759_, _051854_, _051855_);
  and g_090054_(_051721_, _051723_, _051856_);
  or g_090055_(_051720_, _051722_, _051857_);
  or g_090056_(_051734_, _051752_, _051858_);
  or g_090057_(_051756_, _051858_, _051859_);
  and g_090058_(_051850_, _051857_, _051860_);
  or g_090059_(_051849_, _051856_, _051861_);
  and g_090060_(_051855_, _051859_, _051862_);
  not g_090061_(_051862_, _051863_);
  and g_090062_(_051860_, _051862_, _051864_);
  or g_090063_(_051861_, _051863_, _051865_);
  or g_090064_(out[288], _051838_, _051866_);
  and g_090065_(_051828_, _051866_, _051867_);
  and g_090066_(_051841_, _051867_, _051868_);
  and g_090067_(_051808_, _051868_, _051869_);
  not g_090068_(_051869_, _051870_);
  and g_090069_(_051865_, _051870_, _051871_);
  or g_090070_(_051864_, _051869_, _051872_);
  and g_090071_(_026366_, _051871_, _051873_);
  or g_090072_(_026377_, _051872_, _051874_);
  and g_090073_(_051717_, _051872_, _051875_);
  or g_090074_(_051716_, _051871_, _051876_);
  and g_090075_(_051874_, _051876_, _051877_);
  or g_090076_(_051873_, _051875_, _051878_);
  xor g_090077_(_053247_, _013936_, _051879_);
  and g_090078_(_051772_, _051872_, _051880_);
  and g_090079_(_051766_, _051871_, _051881_);
  or g_090080_(_051880_, _051881_, _051882_);
  not g_090081_(_051882_, _051883_);
  or g_090082_(_051879_, _051882_, _051884_);
  and g_090083_(_051879_, _051882_, _051885_);
  xor g_090084_(_051879_, _051882_, _051886_);
  xor g_090085_(_051879_, _051883_, _051887_);
  xor g_090086_(out[309], _013914_, _051888_);
  xor g_090087_(_053269_, _013914_, _051889_);
  or g_090088_(_051795_, _051871_, _051890_);
  not g_090089_(_051890_, _051891_);
  and g_090090_(_051792_, _051871_, _051892_);
  not g_090091_(_051892_, _051893_);
  and g_090092_(_051890_, _051893_, _051894_);
  or g_090093_(_051891_, _051892_, _051895_);
  and g_090094_(_051889_, _051894_, _051896_);
  or g_090095_(_051888_, _051895_, _051897_);
  xor g_090096_(out[310], _013925_, _051898_);
  not g_090097_(_051898_, _051899_);
  or g_090098_(_051763_, _051871_, _051900_);
  or g_090099_(_051760_, _051872_, _051901_);
  and g_090100_(_051900_, _051901_, _051902_);
  and g_090101_(_051899_, _051902_, _051903_);
  xor g_090102_(_051899_, _051902_, _051904_);
  xor g_090103_(_051898_, _051902_, _051905_);
  or g_090104_(_051896_, _051905_, _051906_);
  and g_090105_(_051886_, _051904_, _051907_);
  and g_090106_(_051897_, _051907_, _051908_);
  or g_090107_(_051887_, _051906_, _051909_);
  and g_090108_(_013859_, _014002_, _051910_);
  or g_090109_(_013870_, _013991_, _051911_);
  xor g_090110_(out[314], _013969_, _051912_);
  xor g_090111_(_004520_, _013969_, _051913_);
  and g_090112_(_051877_, _051912_, _051914_);
  or g_090113_(_051878_, _051913_, _051915_);
  and g_090114_(_051911_, _051915_, _051916_);
  or g_090115_(_051910_, _051914_, _051917_);
  and g_090116_(_013870_, _013991_, _051918_);
  or g_090117_(_013859_, _014002_, _051919_);
  and g_090118_(_051878_, _051913_, _051920_);
  not g_090119_(_051920_, _051921_);
  or g_090120_(_051918_, _051920_, _051922_);
  and g_090121_(_051916_, _051921_, _051923_);
  and g_090122_(_051919_, _051923_, _051924_);
  or g_090123_(_051917_, _051922_, _051925_);
  xor g_090124_(out[312], _013947_, _051926_);
  xor g_090125_(_053258_, _013947_, _051927_);
  or g_090126_(_051744_, _051871_, _051928_);
  not g_090127_(_051928_, _051929_);
  and g_090128_(_051738_, _051871_, _051930_);
  not g_090129_(_051930_, _051931_);
  and g_090130_(_051928_, _051931_, _051932_);
  or g_090131_(_051929_, _051930_, _051933_);
  and g_090132_(_051926_, _051932_, _051934_);
  xor g_090133_(out[313], _013958_, _051935_);
  not g_090134_(_051935_, _051936_);
  or g_090135_(_051732_, _051871_, _051937_);
  not g_090136_(_051937_, _051938_);
  and g_090137_(_051729_, _051871_, _051939_);
  not g_090138_(_051939_, _051940_);
  and g_090139_(_051937_, _051940_, _051941_);
  or g_090140_(_051938_, _051939_, _051942_);
  and g_090141_(_051935_, _051942_, _051943_);
  or g_090142_(_051934_, _051943_, _051944_);
  and g_090143_(_051927_, _051933_, _051945_);
  and g_090144_(_051936_, _051941_, _051946_);
  or g_090145_(_051935_, _051942_, _051947_);
  or g_090146_(_051945_, _051946_, _051948_);
  or g_090147_(_051944_, _051948_, _051949_);
  xor g_090148_(_051926_, _051932_, _051950_);
  xor g_090149_(_051936_, _051941_, _051951_);
  and g_090150_(_051924_, _051951_, _051952_);
  and g_090151_(_051950_, _051952_, _051953_);
  or g_090152_(_051925_, _051949_, _051954_);
  and g_090153_(_051908_, _051953_, _051955_);
  or g_090154_(out[306], out[305], _051956_);
  and g_090155_(_013892_, _051956_, _051957_);
  xor g_090156_(_053313_, out[305], _051958_);
  or g_090157_(_051822_, _051871_, _051959_);
  or g_090158_(_051816_, _051872_, _051960_);
  and g_090159_(_051959_, _051960_, _051961_);
  not g_090160_(_051961_, _051962_);
  or g_090161_(_051958_, _051961_, _051963_);
  xor g_090162_(out[307], _013881_, _051964_);
  not g_090163_(_051964_, _051965_);
  and g_090164_(_051810_, _051871_, _051966_);
  not g_090165_(_051966_, _051967_);
  or g_090166_(_051813_, _051871_, _051968_);
  not g_090167_(_051968_, _051969_);
  and g_090168_(_051967_, _051968_, _051970_);
  or g_090169_(_051966_, _051969_, _051971_);
  and g_090170_(_051964_, _051971_, _051972_);
  or g_090171_(_051965_, _051970_, _051973_);
  and g_090172_(_051963_, _051973_, _051974_);
  or g_090173_(_051837_, _051871_, _051975_);
  or g_090174_(out[288], _051872_, _051976_);
  and g_090175_(_051975_, _051976_, _051977_);
  not g_090176_(_051977_, _051978_);
  and g_090177_(out[304], _051978_, _051979_);
  or g_090178_(_004509_, _051977_, _051980_);
  and g_090179_(out[289], _051871_, _051981_);
  or g_090180_(_051831_, _051871_, _051982_);
  not g_090181_(_051982_, _051983_);
  or g_090182_(_051981_, _051983_, _051984_);
  not g_090183_(_051984_, _051985_);
  or g_090184_(out[305], _051985_, _051986_);
  and g_090185_(_051980_, _051986_, _051987_);
  and g_090186_(_051974_, _051987_, _051988_);
  and g_090187_(_051888_, _051895_, _051989_);
  or g_090188_(_051889_, _051894_, _051990_);
  xor g_090189_(out[308], _013903_, _051991_);
  xor g_090190_(_053291_, _013903_, _051992_);
  or g_090191_(_051788_, _051871_, _051993_);
  not g_090192_(_051993_, _051994_);
  and g_090193_(_051782_, _051871_, _051995_);
  not g_090194_(_051995_, _051996_);
  and g_090195_(_051993_, _051996_, _051997_);
  or g_090196_(_051994_, _051995_, _051998_);
  and g_090197_(_051991_, _051997_, _051999_);
  or g_090198_(_051992_, _051998_, _052000_);
  and g_090199_(_051990_, _052000_, _052001_);
  or g_090200_(_051989_, _051999_, _052002_);
  or g_090201_(_053324_, _051984_, _052003_);
  not g_090202_(_052003_, _052004_);
  and g_090203_(_051958_, _051961_, _052005_);
  or g_090204_(_051957_, _051962_, _052006_);
  and g_090205_(_052003_, _052006_, _052007_);
  and g_090206_(_051992_, _051998_, _052008_);
  or g_090207_(_051991_, _051997_, _052009_);
  or g_090208_(_051964_, _051971_, _052010_);
  and g_090209_(_052009_, _052010_, _052011_);
  and g_090210_(_052007_, _052011_, _052012_);
  and g_090211_(_052001_, _052012_, _052013_);
  and g_090212_(_051988_, _052013_, _052014_);
  xor g_090213_(out[305], _051984_, _052015_);
  or g_090214_(_051979_, _052015_, _052016_);
  and g_090215_(_051963_, _052006_, _052017_);
  and g_090216_(_052010_, _052017_, _052018_);
  not g_090217_(_052018_, _052019_);
  or g_090218_(_052002_, _052008_, _052020_);
  or g_090219_(_051909_, _052020_, _052021_);
  or g_090220_(_051954_, _052021_, _052022_);
  or g_090221_(_051972_, _052022_, _052023_);
  or g_090222_(_052019_, _052023_, _052024_);
  and g_090223_(_051955_, _052014_, _052025_);
  or g_090224_(_052016_, _052024_, _052026_);
  and g_090225_(_004509_, _051977_, _052027_);
  or g_090226_(out[304], _051978_, _052028_);
  and g_090227_(_052025_, _052027_, _052029_);
  or g_090228_(_052026_, _052028_, _052030_);
  or g_090229_(_051972_, _052005_, _052031_);
  and g_090230_(_051963_, _052004_, _052032_);
  or g_090231_(_052031_, _052032_, _052033_);
  and g_090232_(_052011_, _052033_, _052034_);
  or g_090233_(_052002_, _052034_, _052035_);
  and g_090234_(_051955_, _052035_, _052036_);
  and g_090235_(_051944_, _051947_, _052037_);
  and g_090236_(_051924_, _052037_, _052038_);
  or g_090237_(_051916_, _051918_, _052039_);
  not g_090238_(_052039_, _052040_);
  or g_090239_(_052038_, _052040_, _052041_);
  or g_090240_(_051885_, _051903_, _052042_);
  and g_090241_(_051884_, _052042_, _052043_);
  and g_090242_(_051953_, _052043_, _052044_);
  or g_090243_(_052041_, _052044_, _052045_);
  or g_090244_(_052036_, _052045_, _052046_);
  not g_090245_(_052046_, _052047_);
  and g_090246_(_052030_, _052047_, _052048_);
  or g_090247_(_052029_, _052046_, _052049_);
  and g_090248_(_051878_, _052048_, _052050_);
  not g_090249_(_052050_, _052051_);
  or g_090250_(_051913_, _052048_, _052052_);
  not g_090251_(_052052_, _052053_);
  and g_090252_(_052051_, _052052_, _052054_);
  or g_090253_(_052050_, _052053_, _052055_);
  and g_090254_(_026300_, _052054_, _052056_);
  or g_090255_(_026311_, _052055_, _052057_);
  and g_090256_(_026355_, _052057_, _052058_);
  or g_090257_(_026344_, _052056_, _052059_);
  and g_090258_(_026333_, _052059_, _052060_);
  or g_090259_(_026322_, _052058_, _052061_);
  and g_090260_(_026311_, _052055_, _052062_);
  or g_090261_(_026300_, _052054_, _052063_);
  and g_090262_(_026333_, _052063_, _052064_);
  or g_090263_(_026322_, _052062_, _052065_);
  xor g_090264_(out[329], _014112_, _052066_);
  xor g_090265_(_053434_, _014112_, _052067_);
  or g_090266_(_051935_, _052048_, _052068_);
  or g_090267_(_051941_, _052049_, _052069_);
  and g_090268_(_052068_, _052069_, _052070_);
  not g_090269_(_052070_, _052071_);
  and g_090270_(_052067_, _052070_, _052072_);
  or g_090271_(_052066_, _052071_, _052073_);
  and g_090272_(_052064_, _052073_, _052074_);
  or g_090273_(_052065_, _052072_, _052075_);
  and g_090274_(_052058_, _052074_, _052076_);
  or g_090275_(_052059_, _052075_, _052077_);
  xor g_090276_(out[328], _014101_, _052078_);
  not g_090277_(_052078_, _052079_);
  or g_090278_(_051927_, _052048_, _052080_);
  not g_090279_(_052080_, _052081_);
  and g_090280_(_051933_, _052048_, _052082_);
  not g_090281_(_052082_, _052083_);
  and g_090282_(_052080_, _052083_, _052084_);
  or g_090283_(_052081_, _052082_, _052085_);
  and g_090284_(_052078_, _052084_, _052086_);
  or g_090285_(_052079_, _052085_, _052087_);
  and g_090286_(_052066_, _052071_, _052088_);
  or g_090287_(_052067_, _052070_, _052089_);
  and g_090288_(_052087_, _052089_, _052090_);
  or g_090289_(_052086_, _052088_, _052091_);
  or g_090290_(_053324_, _052048_, _052092_);
  not g_090291_(_052092_, _052093_);
  and g_090292_(_051984_, _052048_, _052094_);
  not g_090293_(_052094_, _052095_);
  and g_090294_(_052092_, _052095_, _052096_);
  or g_090295_(_052093_, _052094_, _052097_);
  and g_090296_(out[321], _052096_, _052098_);
  or g_090297_(_053423_, _052097_, _052099_);
  or g_090298_(_004509_, _052047_, _052100_);
  not g_090299_(_052100_, _052101_);
  and g_090300_(_051977_, _052048_, _052102_);
  or g_090301_(_052101_, _052102_, _052103_);
  not g_090302_(_052103_, _052104_);
  and g_090303_(out[320], _052104_, _052105_);
  or g_090304_(_004542_, _052103_, _052106_);
  xor g_090305_(out[321], _052096_, _052107_);
  xor g_090306_(_053423_, _052096_, _052108_);
  and g_090307_(_052106_, _052107_, _052109_);
  or g_090308_(_052105_, _052108_, _052110_);
  and g_090309_(_052099_, _052110_, _052111_);
  or g_090310_(_052098_, _052109_, _052112_);
  xor g_090311_(out[326], _014079_, _052113_);
  xor g_090312_(_053379_, _014079_, _052114_);
  or g_090313_(_051898_, _052048_, _052115_);
  or g_090314_(_051902_, _052049_, _052116_);
  and g_090315_(_052115_, _052116_, _052117_);
  and g_090316_(_052114_, _052117_, _052118_);
  xor g_090317_(out[327], _014090_, _052119_);
  not g_090318_(_052119_, _052120_);
  or g_090319_(_051879_, _052048_, _052121_);
  not g_090320_(_052121_, _052122_);
  and g_090321_(_051882_, _052048_, _052123_);
  not g_090322_(_052123_, _052124_);
  and g_090323_(_052121_, _052124_, _052125_);
  or g_090324_(_052122_, _052123_, _052126_);
  and g_090325_(_052120_, _052126_, _052127_);
  or g_090326_(_052118_, _052127_, _052128_);
  or g_090327_(_052120_, _052126_, _052129_);
  xor g_090328_(_052114_, _052117_, _052130_);
  xor g_090329_(_052113_, _052117_, _052131_);
  xor g_090330_(_052119_, _052125_, _052132_);
  xor g_090331_(_052120_, _052125_, _052133_);
  and g_090332_(_052130_, _052132_, _052134_);
  or g_090333_(_052131_, _052133_, _052135_);
  xor g_090334_(out[325], _014068_, _052136_);
  xor g_090335_(_053368_, _014068_, _052137_);
  or g_090336_(_051888_, _052048_, _052138_);
  or g_090337_(_051894_, _052049_, _052139_);
  and g_090338_(_052138_, _052139_, _052140_);
  and g_090339_(_052137_, _052140_, _052141_);
  or g_090340_(_052137_, _052140_, _052142_);
  xor g_090341_(_052137_, _052140_, _052143_);
  xor g_090342_(_052136_, _052140_, _052144_);
  xor g_090343_(out[324], _014057_, _052145_);
  not g_090344_(_052145_, _052146_);
  and g_090345_(_051998_, _052048_, _052147_);
  or g_090346_(_051997_, _052049_, _052148_);
  and g_090347_(_051991_, _052049_, _052149_);
  or g_090348_(_051992_, _052048_, _052150_);
  and g_090349_(_052148_, _052150_, _052151_);
  or g_090350_(_052147_, _052149_, _052152_);
  or g_090351_(_052146_, _052152_, _052153_);
  xor g_090352_(_052145_, _052151_, _052154_);
  xor g_090353_(_052146_, _052151_, _052155_);
  and g_090354_(_052143_, _052154_, _052156_);
  or g_090355_(_052144_, _052155_, _052157_);
  and g_090356_(_052134_, _052156_, _052158_);
  or g_090357_(_052135_, _052157_, _052159_);
  xor g_090358_(_053390_, _014035_, _052160_);
  or g_090359_(_051964_, _052048_, _052161_);
  or g_090360_(_051970_, _052049_, _052162_);
  and g_090361_(_052161_, _052162_, _052163_);
  not g_090362_(_052163_, _052164_);
  and g_090363_(_052160_, _052163_, _052165_);
  or g_090364_(out[322], out[321], _052166_);
  xor g_090365_(out[322], out[321], _052167_);
  xor g_090366_(_053412_, out[321], _052168_);
  and g_090367_(_051962_, _052048_, _052169_);
  and g_090368_(_051958_, _052049_, _052170_);
  or g_090369_(_052169_, _052170_, _052171_);
  or g_090370_(_052167_, _052171_, _052172_);
  or g_090371_(_052160_, _052163_, _052173_);
  xor g_090372_(_052167_, _052171_, _052174_);
  xor g_090373_(_052168_, _052171_, _052175_);
  xor g_090374_(_052160_, _052163_, _052176_);
  xor g_090375_(_052160_, _052164_, _052177_);
  and g_090376_(_052174_, _052176_, _052178_);
  or g_090377_(_052175_, _052177_, _052179_);
  and g_090378_(_052158_, _052178_, _052180_);
  or g_090379_(_052159_, _052179_, _052181_);
  and g_090380_(_052112_, _052180_, _052182_);
  or g_090381_(_052111_, _052181_, _052183_);
  and g_090382_(_052172_, _052173_, _052184_);
  or g_090383_(_052165_, _052184_, _052185_);
  or g_090384_(_052159_, _052185_, _052186_);
  and g_090385_(_052128_, _052129_, _052187_);
  not g_090386_(_052187_, _052188_);
  or g_090387_(_052141_, _052153_, _052189_);
  and g_090388_(_052142_, _052189_, _052190_);
  or g_090389_(_052135_, _052190_, _052191_);
  and g_090390_(_052186_, _052191_, _052192_);
  not g_090391_(_052192_, _052193_);
  and g_090392_(_052188_, _052192_, _052194_);
  or g_090393_(_052187_, _052193_, _052195_);
  and g_090394_(_052183_, _052194_, _052196_);
  or g_090395_(_052182_, _052195_, _052197_);
  and g_090396_(_052079_, _052085_, _052198_);
  or g_090397_(_052078_, _052084_, _052199_);
  and g_090398_(_052197_, _052199_, _052200_);
  or g_090399_(_052196_, _052198_, _052201_);
  and g_090400_(_052090_, _052201_, _052202_);
  or g_090401_(_052091_, _052200_, _052203_);
  and g_090402_(_052076_, _052203_, _052204_);
  or g_090403_(_052077_, _052202_, _052205_);
  and g_090404_(_052061_, _052205_, _052206_);
  or g_090405_(_052060_, _052204_, _052207_);
  and g_090406_(_004542_, _052103_, _052208_);
  or g_090407_(out[320], _052104_, _052209_);
  and g_090408_(_052199_, _052209_, _052210_);
  or g_090409_(_052198_, _052208_, _052211_);
  and g_090410_(_052090_, _052210_, _052212_);
  or g_090411_(_052091_, _052211_, _052213_);
  and g_090412_(_052109_, _052212_, _052214_);
  or g_090413_(_052110_, _052213_, _052215_);
  and g_090414_(_052076_, _052214_, _052216_);
  or g_090415_(_052077_, _052215_, _052217_);
  and g_090416_(_052180_, _052216_, _052218_);
  or g_090417_(_052181_, _052217_, _052219_);
  and g_090418_(_052207_, _052219_, _052220_);
  or g_090419_(_052206_, _052218_, _052221_);
  and g_090420_(_026300_, _052220_, _052222_);
  or g_090421_(_026311_, _052221_, _052223_);
  and g_090422_(_052055_, _052221_, _052224_);
  or g_090423_(_052054_, _052220_, _052225_);
  and g_090424_(_052223_, _052225_, _052226_);
  or g_090425_(_052222_, _052224_, _052227_);
  xor g_090426_(out[346], _014277_, _052228_);
  xor g_090427_(_004586_, _014277_, _052229_);
  and g_090428_(_052227_, _052229_, _052230_);
  or g_090429_(_052226_, _052228_, _052231_);
  xor g_090430_(out[345], _014266_, _052232_);
  xor g_090431_(_053533_, _014266_, _052233_);
  or g_090432_(_052070_, _052220_, _052234_);
  not g_090433_(_052234_, _052235_);
  and g_090434_(_052067_, _052220_, _052236_);
  not g_090435_(_052236_, _052237_);
  and g_090436_(_052234_, _052237_, _052238_);
  or g_090437_(_052235_, _052236_, _052239_);
  and g_090438_(_052233_, _052238_, _052240_);
  or g_090439_(_052232_, _052239_, _052241_);
  xor g_090440_(out[343], _014244_, _052242_);
  xor g_090441_(_053445_, _014244_, _052243_);
  or g_090442_(_052125_, _052220_, _052244_);
  not g_090443_(_052244_, _052245_);
  and g_090444_(_052119_, _052220_, _052246_);
  not g_090445_(_052246_, _052247_);
  and g_090446_(_052244_, _052247_, _052248_);
  or g_090447_(_052245_, _052246_, _052249_);
  and g_090448_(_052242_, _052248_, _052250_);
  or g_090449_(_052243_, _052249_, _052251_);
  and g_090450_(_014167_, _014310_, _052252_);
  or g_090451_(_014178_, _014299_, _052253_);
  and g_090452_(_052226_, _052228_, _052254_);
  or g_090453_(_052227_, _052229_, _052255_);
  and g_090454_(_052253_, _052255_, _052256_);
  or g_090455_(_052252_, _052254_, _052257_);
  and g_090456_(_052232_, _052239_, _052258_);
  or g_090457_(_052233_, _052238_, _052259_);
  or g_090458_(_052084_, _052220_, _052260_);
  not g_090459_(_052260_, _052261_);
  and g_090460_(_052078_, _052220_, _052262_);
  not g_090461_(_052262_, _052263_);
  and g_090462_(_052260_, _052263_, _052264_);
  or g_090463_(_052261_, _052262_, _052265_);
  xor g_090464_(out[344], _014255_, _052266_);
  xor g_090465_(_053456_, _014255_, _052267_);
  and g_090466_(_052264_, _052266_, _052268_);
  or g_090467_(_052265_, _052267_, _052269_);
  and g_090468_(_052259_, _052269_, _052270_);
  or g_090469_(_052258_, _052268_, _052271_);
  and g_090470_(_014178_, _014299_, _052272_);
  or g_090471_(_014167_, _014310_, _052273_);
  and g_090472_(_052265_, _052267_, _052274_);
  or g_090473_(_052264_, _052266_, _052275_);
  and g_090474_(_052231_, _052273_, _052276_);
  or g_090475_(_052230_, _052272_, _052277_);
  and g_090476_(_052256_, _052276_, _052278_);
  or g_090477_(_052257_, _052277_, _052279_);
  xor g_090478_(out[340], _014211_, _052280_);
  xor g_090479_(_053500_, _014211_, _052281_);
  and g_090480_(_052145_, _052220_, _052282_);
  not g_090481_(_052282_, _052283_);
  or g_090482_(_052151_, _052220_, _052284_);
  not g_090483_(_052284_, _052285_);
  and g_090484_(_052283_, _052284_, _052286_);
  or g_090485_(_052282_, _052285_, _052287_);
  and g_090486_(_052280_, _052286_, _052288_);
  or g_090487_(_052281_, _052287_, _052289_);
  xor g_090488_(out[341], _014222_, _052290_);
  xor g_090489_(_053467_, _014222_, _052291_);
  or g_090490_(_052140_, _052220_, _052292_);
  not g_090491_(_052292_, _052293_);
  and g_090492_(_052137_, _052220_, _052294_);
  not g_090493_(_052294_, _052295_);
  and g_090494_(_052292_, _052295_, _052296_);
  or g_090495_(_052293_, _052294_, _052297_);
  and g_090496_(_052290_, _052297_, _052298_);
  or g_090497_(_052291_, _052296_, _052299_);
  and g_090498_(_052281_, _052287_, _052300_);
  or g_090499_(_052280_, _052286_, _052301_);
  and g_090500_(_052299_, _052301_, _052302_);
  or g_090501_(_052298_, _052300_, _052303_);
  xor g_090502_(out[342], _014233_, _052304_);
  xor g_090503_(_053478_, _014233_, _052305_);
  or g_090504_(_052117_, _052220_, _052306_);
  not g_090505_(_052306_, _052307_);
  and g_090506_(_052114_, _052220_, _052308_);
  not g_090507_(_052308_, _052309_);
  and g_090508_(_052306_, _052309_, _052310_);
  or g_090509_(_052307_, _052308_, _052311_);
  and g_090510_(_052305_, _052310_, _052312_);
  or g_090511_(_052304_, _052311_, _052313_);
  and g_090512_(_052243_, _052249_, _052314_);
  or g_090513_(_052242_, _052248_, _052315_);
  and g_090514_(_052313_, _052315_, _052316_);
  or g_090515_(_052312_, _052314_, _052317_);
  and g_090516_(_052291_, _052296_, _052318_);
  or g_090517_(_052290_, _052297_, _052319_);
  and g_090518_(_052304_, _052311_, _052320_);
  or g_090519_(_052305_, _052310_, _052321_);
  and g_090520_(_052319_, _052321_, _052322_);
  or g_090521_(_052318_, _052320_, _052323_);
  and g_090522_(_052316_, _052321_, _052324_);
  or g_090523_(_052317_, _052320_, _052325_);
  and g_090524_(_052302_, _052319_, _052326_);
  or g_090525_(_052303_, _052318_, _052327_);
  and g_090526_(_052289_, _052326_, _052328_);
  or g_090527_(_052288_, _052327_, _052329_);
  and g_090528_(_052259_, _052275_, _052330_);
  or g_090529_(_052258_, _052274_, _052331_);
  and g_090530_(_052241_, _052269_, _052332_);
  or g_090531_(_052240_, _052268_, _052333_);
  and g_090532_(_052330_, _052332_, _052334_);
  or g_090533_(_052331_, _052333_, _052335_);
  and g_090534_(_052278_, _052334_, _052336_);
  or g_090535_(_052279_, _052335_, _052337_);
  and g_090536_(_052251_, _052324_, _052338_);
  or g_090537_(_052250_, _052325_, _052339_);
  and g_090538_(_052336_, _052338_, _052340_);
  or g_090539_(_052337_, _052339_, _052341_);
  and g_090540_(_052328_, _052340_, _052342_);
  or g_090541_(_052329_, _052341_, _052343_);
  xor g_090542_(out[339], _014189_, _052344_);
  xor g_090543_(_053489_, _014189_, _052345_);
  or g_090544_(_052163_, _052220_, _052346_);
  not g_090545_(_052346_, _052347_);
  and g_090546_(_052160_, _052220_, _052348_);
  not g_090547_(_052348_, _052349_);
  and g_090548_(_052346_, _052349_, _052350_);
  or g_090549_(_052347_, _052348_, _052351_);
  and g_090550_(_052344_, _052351_, _052352_);
  or g_090551_(out[338], out[337], _052353_);
  xor g_090552_(out[338], out[337], _052354_);
  xor g_090553_(_053511_, out[337], _052355_);
  and g_090554_(_052171_, _052221_, _052356_);
  and g_090555_(_052168_, _052220_, _052357_);
  or g_090556_(_052356_, _052357_, _052358_);
  not g_090557_(_052358_, _052359_);
  and g_090558_(_052355_, _052359_, _052360_);
  or g_090559_(_052352_, _052360_, _052361_);
  and g_090560_(_052345_, _052350_, _052362_);
  or g_090561_(_052344_, _052351_, _052363_);
  and g_090562_(_052354_, _052358_, _052364_);
  or g_090563_(_052362_, _052364_, _052365_);
  xor g_090564_(_052345_, _052350_, _052366_);
  xor g_090565_(_052354_, _052358_, _052367_);
  and g_090566_(_052366_, _052367_, _052368_);
  or g_090567_(_052361_, _052365_, _052369_);
  or g_090568_(_053423_, _052221_, _052370_);
  or g_090569_(_052096_, _052220_, _052371_);
  and g_090570_(_052370_, _052371_, _052372_);
  and g_090571_(out[337], _052372_, _052373_);
  or g_090572_(_052103_, _052220_, _052374_);
  not g_090573_(_052374_, _052375_);
  and g_090574_(_004542_, _052220_, _052376_);
  not g_090575_(_052376_, _052377_);
  and g_090576_(_052374_, _052377_, _052378_);
  or g_090577_(_052375_, _052376_, _052379_);
  and g_090578_(out[336], _052379_, _052380_);
  or g_090579_(_004575_, _052378_, _052381_);
  xor g_090580_(out[337], _052372_, _052382_);
  xor g_090581_(_053522_, _052372_, _052383_);
  and g_090582_(_052381_, _052382_, _052384_);
  or g_090583_(_052380_, _052383_, _052385_);
  or g_090584_(_052373_, _052384_, _052386_);
  and g_090585_(_052368_, _052386_, _052387_);
  and g_090586_(_052361_, _052363_, _052388_);
  or g_090587_(_052387_, _052388_, _052389_);
  not g_090588_(_052389_, _052390_);
  and g_090589_(_052342_, _052389_, _052391_);
  or g_090590_(_052343_, _052390_, _052392_);
  and g_090591_(_052289_, _052299_, _052393_);
  or g_090592_(_052288_, _052298_, _052394_);
  and g_090593_(_052322_, _052394_, _052395_);
  or g_090594_(_052323_, _052393_, _052396_);
  and g_090595_(_052316_, _052396_, _052397_);
  or g_090596_(_052317_, _052395_, _052398_);
  and g_090597_(_052251_, _052398_, _052399_);
  or g_090598_(_052250_, _052397_, _052400_);
  and g_090599_(_052336_, _052399_, _052401_);
  or g_090600_(_052337_, _052400_, _052402_);
  and g_090601_(_052231_, _052241_, _052403_);
  or g_090602_(_052230_, _052240_, _052404_);
  and g_090603_(_052271_, _052403_, _052405_);
  or g_090604_(_052270_, _052404_, _052406_);
  and g_090605_(_052256_, _052406_, _052407_);
  or g_090606_(_052257_, _052405_, _052408_);
  and g_090607_(_052273_, _052408_, _052409_);
  or g_090608_(_052272_, _052407_, _052410_);
  and g_090609_(_052402_, _052410_, _052411_);
  or g_090610_(_052401_, _052409_, _052412_);
  and g_090611_(_052392_, _052411_, _052413_);
  or g_090612_(_052391_, _052412_, _052414_);
  and g_090613_(_004575_, _052378_, _052415_);
  or g_090614_(out[336], _052379_, _052416_);
  and g_090615_(_052368_, _052416_, _052417_);
  or g_090616_(_052369_, _052415_, _052418_);
  and g_090617_(_052384_, _052417_, _052419_);
  or g_090618_(_052385_, _052418_, _052420_);
  and g_090619_(_052342_, _052419_, _052421_);
  or g_090620_(_052343_, _052420_, _052422_);
  and g_090621_(_052414_, _052422_, _052423_);
  or g_090622_(_052413_, _052421_, _052424_);
  or g_090623_(_052226_, _052423_, _052425_);
  not g_090624_(_052425_, _052426_);
  and g_090625_(_052228_, _052423_, _052427_);
  not g_090626_(_052427_, _052428_);
  and g_090627_(_052425_, _052428_, _052429_);
  or g_090628_(_052426_, _052427_, _052430_);
  xor g_090629_(out[362], _014431_, _052431_);
  xor g_090630_(_004619_, _014431_, _052432_);
  and g_090631_(_052429_, _052431_, _052433_);
  or g_090632_(_052430_, _052432_, _052434_);
  and g_090633_(_026289_, _052434_, _052435_);
  or g_090634_(_026278_, _052433_, _052436_);
  and g_090635_(_052430_, _052432_, _052437_);
  or g_090636_(_052429_, _052431_, _052438_);
  and g_090637_(_014332_, _014453_, _052439_);
  or g_090638_(_014321_, _014464_, _052440_);
  xor g_090639_(out[361], _014420_, _052441_);
  xor g_090640_(_053632_, _014420_, _052442_);
  and g_090641_(_052233_, _052423_, _052443_);
  or g_090642_(_052232_, _052424_, _052444_);
  and g_090643_(_052239_, _052424_, _052445_);
  or g_090644_(_052238_, _052423_, _052446_);
  and g_090645_(_052444_, _052446_, _052447_);
  or g_090646_(_052443_, _052445_, _052448_);
  and g_090647_(_052442_, _052447_, _052449_);
  or g_090648_(_052441_, _052448_, _052450_);
  and g_090649_(_052440_, _052450_, _052451_);
  or g_090650_(_052439_, _052449_, _052452_);
  and g_090651_(_052438_, _052451_, _052453_);
  or g_090652_(_052437_, _052452_, _052454_);
  and g_090653_(_052435_, _052453_, _052455_);
  or g_090654_(_052436_, _052454_, _052456_);
  and g_090655_(_052266_, _052423_, _052457_);
  not g_090656_(_052457_, _052458_);
  or g_090657_(_052264_, _052423_, _052459_);
  not g_090658_(_052459_, _052460_);
  and g_090659_(_052458_, _052459_, _052461_);
  or g_090660_(_052457_, _052460_, _052462_);
  xor g_090661_(out[360], _014409_, _052463_);
  xor g_090662_(_053555_, _014409_, _052464_);
  and g_090663_(_052461_, _052463_, _052465_);
  or g_090664_(_052462_, _052464_, _052466_);
  and g_090665_(_052441_, _052448_, _052467_);
  or g_090666_(_052442_, _052447_, _052468_);
  and g_090667_(_052466_, _052468_, _052469_);
  or g_090668_(_052465_, _052467_, _052470_);
  and g_090669_(_052462_, _052464_, _052471_);
  or g_090670_(_052461_, _052463_, _052472_);
  and g_090671_(_052469_, _052472_, _052473_);
  or g_090672_(_052470_, _052471_, _052474_);
  and g_090673_(_052455_, _052473_, _052475_);
  or g_090674_(_052456_, _052474_, _052476_);
  xor g_090675_(out[358], _014387_, _052477_);
  xor g_090676_(_053577_, _014387_, _052478_);
  and g_090677_(_052305_, _052423_, _052479_);
  not g_090678_(_052479_, _052480_);
  or g_090679_(_052310_, _052423_, _052481_);
  not g_090680_(_052481_, _052482_);
  and g_090681_(_052480_, _052481_, _052483_);
  or g_090682_(_052479_, _052482_, _052484_);
  and g_090683_(_052478_, _052483_, _052485_);
  or g_090684_(_052477_, _052484_, _052486_);
  and g_090685_(_052242_, _052423_, _052487_);
  not g_090686_(_052487_, _052488_);
  or g_090687_(_052248_, _052423_, _052489_);
  not g_090688_(_052489_, _052490_);
  and g_090689_(_052488_, _052489_, _052491_);
  or g_090690_(_052487_, _052490_, _052492_);
  and g_090691_(_026267_, _052492_, _052493_);
  or g_090692_(_026256_, _052491_, _052494_);
  and g_090693_(_052486_, _052494_, _052495_);
  or g_090694_(_052485_, _052493_, _052496_);
  and g_090695_(_026256_, _052491_, _052497_);
  or g_090696_(_026267_, _052492_, _052498_);
  and g_090697_(_052477_, _052484_, _052499_);
  or g_090698_(_052478_, _052483_, _052500_);
  and g_090699_(_052498_, _052500_, _052501_);
  or g_090700_(_052497_, _052499_, _052502_);
  and g_090701_(_052495_, _052501_, _052503_);
  or g_090702_(_052496_, _052502_, _052504_);
  xor g_090703_(out[357], _014376_, _052505_);
  xor g_090704_(_053566_, _014376_, _052506_);
  and g_090705_(_052291_, _052423_, _052507_);
  not g_090706_(_052507_, _052508_);
  or g_090707_(_052296_, _052423_, _052509_);
  not g_090708_(_052509_, _052510_);
  and g_090709_(_052508_, _052509_, _052511_);
  or g_090710_(_052507_, _052510_, _052512_);
  and g_090711_(_052505_, _052512_, _052513_);
  or g_090712_(_052506_, _052511_, _052514_);
  xor g_090713_(out[356], _014365_, _052515_);
  xor g_090714_(_053599_, _014365_, _052516_);
  and g_090715_(_052280_, _052423_, _052517_);
  not g_090716_(_052517_, _052518_);
  or g_090717_(_052286_, _052423_, _052519_);
  not g_090718_(_052519_, _052520_);
  and g_090719_(_052518_, _052519_, _052521_);
  or g_090720_(_052517_, _052520_, _052522_);
  and g_090721_(_052515_, _052521_, _052523_);
  or g_090722_(_052516_, _052522_, _052524_);
  and g_090723_(_052514_, _052524_, _052525_);
  or g_090724_(_052513_, _052523_, _052526_);
  and g_090725_(_052506_, _052511_, _052527_);
  or g_090726_(_052505_, _052512_, _052528_);
  and g_090727_(_052516_, _052522_, _052529_);
  or g_090728_(_052515_, _052521_, _052530_);
  and g_090729_(_052528_, _052530_, _052531_);
  or g_090730_(_052527_, _052529_, _052532_);
  and g_090731_(_052525_, _052531_, _052533_);
  or g_090732_(_052526_, _052532_, _052534_);
  and g_090733_(_052503_, _052533_, _052535_);
  or g_090734_(_052504_, _052534_, _052536_);
  and g_090735_(_052475_, _052535_, _052537_);
  or g_090736_(_052476_, _052536_, _052538_);
  xor g_090737_(out[355], _014343_, _052539_);
  or g_090738_(_052350_, _052423_, _052540_);
  not g_090739_(_052540_, _052541_);
  and g_090740_(_052345_, _052423_, _052542_);
  not g_090741_(_052542_, _052543_);
  and g_090742_(_052540_, _052543_, _052544_);
  or g_090743_(_052541_, _052542_, _052545_);
  and g_090744_(_052539_, _052545_, _052546_);
  or g_090745_(out[354], out[353], _052547_);
  xor g_090746_(out[354], out[353], _052548_);
  xor g_090747_(_053610_, out[353], _052549_);
  and g_090748_(_052358_, _052424_, _052550_);
  and g_090749_(_052355_, _052423_, _052551_);
  or g_090750_(_052550_, _052551_, _052552_);
  not g_090751_(_052552_, _052553_);
  and g_090752_(_052549_, _052553_, _052554_);
  or g_090753_(_052539_, _052545_, _052555_);
  not g_090754_(_052555_, _052556_);
  xor g_090755_(_052548_, _052552_, _052557_);
  xor g_090756_(_052549_, _052552_, _052558_);
  xor g_090757_(_052539_, _052545_, _052559_);
  or g_090758_(_052546_, _052556_, _052560_);
  and g_090759_(_052557_, _052559_, _052561_);
  or g_090760_(_052558_, _052560_, _052562_);
  and g_090761_(out[337], _052423_, _052563_);
  not g_090762_(_052563_, _052564_);
  or g_090763_(_052372_, _052423_, _052565_);
  not g_090764_(_052565_, _052566_);
  and g_090765_(_052564_, _052565_, _052567_);
  or g_090766_(_052563_, _052566_, _052568_);
  and g_090767_(out[353], _052567_, _052569_);
  or g_090768_(_053621_, _052568_, _052570_);
  or g_090769_(_052378_, _052423_, _052571_);
  not g_090770_(_052571_, _052572_);
  and g_090771_(_004575_, _052423_, _052573_);
  not g_090772_(_052573_, _052574_);
  and g_090773_(_052571_, _052574_, _052575_);
  or g_090774_(_052572_, _052573_, _052576_);
  and g_090775_(out[352], _052576_, _052577_);
  or g_090776_(_004608_, _052575_, _052578_);
  xor g_090777_(out[353], _052567_, _052579_);
  xor g_090778_(_053621_, _052567_, _052580_);
  and g_090779_(_052578_, _052579_, _052581_);
  or g_090780_(_052577_, _052580_, _052582_);
  and g_090781_(_052570_, _052582_, _052583_);
  or g_090782_(_052569_, _052581_, _052584_);
  and g_090783_(_052561_, _052584_, _052585_);
  or g_090784_(_052562_, _052583_, _052586_);
  and g_090785_(_052554_, _052555_, _052587_);
  or g_090786_(_052546_, _052587_, _052588_);
  not g_090787_(_052588_, _052589_);
  and g_090788_(_052586_, _052589_, _052590_);
  or g_090789_(_052585_, _052588_, _052591_);
  and g_090790_(_052537_, _052591_, _052592_);
  or g_090791_(_052538_, _052590_, _052593_);
  and g_090792_(_052496_, _052498_, _052594_);
  or g_090793_(_052495_, _052497_, _052595_);
  and g_090794_(_052526_, _052528_, _052596_);
  or g_090795_(_052525_, _052527_, _052597_);
  and g_090796_(_052503_, _052596_, _052598_);
  or g_090797_(_052504_, _052597_, _052599_);
  and g_090798_(_052595_, _052599_, _052600_);
  or g_090799_(_052594_, _052598_, _052601_);
  and g_090800_(_052475_, _052601_, _052602_);
  or g_090801_(_052476_, _052600_, _052603_);
  and g_090802_(_052436_, _052440_, _052604_);
  or g_090803_(_052435_, _052439_, _052605_);
  and g_090804_(_052455_, _052470_, _052606_);
  or g_090805_(_052456_, _052469_, _052607_);
  and g_090806_(_052605_, _052607_, _052608_);
  or g_090807_(_052604_, _052606_, _052609_);
  and g_090808_(_052603_, _052608_, _052610_);
  or g_090809_(_052602_, _052609_, _052611_);
  and g_090810_(_052593_, _052610_, _052612_);
  or g_090811_(_052592_, _052611_, _052613_);
  and g_090812_(_004608_, _052575_, _052614_);
  or g_090813_(out[352], _052576_, _052615_);
  or g_090814_(_052562_, _052582_, _052616_);
  not g_090815_(_052616_, _052617_);
  and g_090816_(_052615_, _052617_, _052618_);
  or g_090817_(_052614_, _052616_, _052619_);
  and g_090818_(_052537_, _052618_, _052620_);
  or g_090819_(_052538_, _052619_, _052621_);
  and g_090820_(_052613_, _052621_, _052622_);
  or g_090821_(_052612_, _052620_, _052623_);
  and g_090822_(_026256_, _052622_, _052624_);
  not g_090823_(_052624_, _052625_);
  or g_090824_(_052491_, _052622_, _052626_);
  not g_090825_(_052626_, _052627_);
  and g_090826_(_052625_, _052626_, _052628_);
  or g_090827_(_052624_, _052627_, _052629_);
  and g_090828_(_026245_, _052629_, _052630_);
  or g_090829_(_026234_, _052628_, _052631_);
  xor g_090830_(out[374], _014541_, _052632_);
  xor g_090831_(_053676_, _014541_, _052633_);
  and g_090832_(_052478_, _052622_, _052634_);
  not g_090833_(_052634_, _052635_);
  or g_090834_(_052483_, _052622_, _052636_);
  not g_090835_(_052636_, _052637_);
  and g_090836_(_052635_, _052636_, _052638_);
  or g_090837_(_052634_, _052637_, _052639_);
  and g_090838_(_052633_, _052638_, _052640_);
  or g_090839_(_052632_, _052639_, _052641_);
  and g_090840_(_052631_, _052641_, _052642_);
  xor g_090841_(out[373], _014530_, _052643_);
  xor g_090842_(_053665_, _014530_, _052644_);
  or g_090843_(_052505_, _052623_, _052645_);
  or g_090844_(_052511_, _052622_, _052646_);
  and g_090845_(_052645_, _052646_, _052647_);
  not g_090846_(_052647_, _052648_);
  and g_090847_(_052643_, _052648_, _052649_);
  or g_090848_(_052644_, _052647_, _052650_);
  and g_090849_(_052515_, _052622_, _052651_);
  not g_090850_(_052651_, _052652_);
  or g_090851_(_052521_, _052622_, _052653_);
  not g_090852_(_052653_, _052654_);
  and g_090853_(_052652_, _052653_, _052655_);
  or g_090854_(_052651_, _052654_, _052656_);
  or g_090855_(_026223_, _052656_, _052657_);
  and g_090856_(_052650_, _052657_, _052658_);
  and g_090857_(_052644_, _052647_, _052659_);
  or g_090858_(_052643_, _052648_, _052660_);
  and g_090859_(_052632_, _052639_, _052661_);
  or g_090860_(_052633_, _052638_, _052662_);
  and g_090861_(_052631_, _052662_, _052663_);
  or g_090862_(_052630_, _052661_, _052664_);
  or g_090863_(_052658_, _052664_, _052665_);
  or g_090864_(_052659_, _052665_, _052666_);
  and g_090865_(_052642_, _052666_, _052667_);
  and g_090866_(_014475_, _014618_, _052668_);
  or g_090867_(_014486_, _014607_, _052669_);
  and g_090868_(_052430_, _052623_, _052670_);
  or g_090869_(_052429_, _052622_, _052671_);
  and g_090870_(_052431_, _052622_, _052672_);
  or g_090871_(_052432_, _052623_, _052673_);
  and g_090872_(_052671_, _052673_, _052674_);
  or g_090873_(_052670_, _052672_, _052675_);
  xor g_090874_(out[378], _014585_, _052676_);
  xor g_090875_(_004652_, _014585_, _052677_);
  and g_090876_(_052674_, _052676_, _052678_);
  or g_090877_(_052675_, _052677_, _052679_);
  and g_090878_(_052669_, _052679_, _052680_);
  or g_090879_(_052668_, _052678_, _052681_);
  and g_090880_(_014486_, _014607_, _052682_);
  or g_090881_(_014475_, _014618_, _052683_);
  and g_090882_(_052675_, _052677_, _052684_);
  or g_090883_(_052674_, _052676_, _052685_);
  and g_090884_(_052683_, _052685_, _052686_);
  or g_090885_(_052682_, _052684_, _052687_);
  xor g_090886_(out[377], _014574_, _052688_);
  xor g_090887_(_053731_, _014574_, _052689_);
  and g_090888_(_052442_, _052622_, _052690_);
  not g_090889_(_052690_, _052691_);
  or g_090890_(_052447_, _052622_, _052692_);
  not g_090891_(_052692_, _052693_);
  and g_090892_(_052691_, _052692_, _052694_);
  or g_090893_(_052690_, _052693_, _052695_);
  and g_090894_(_052689_, _052694_, _052696_);
  or g_090895_(_052688_, _052695_, _052697_);
  and g_090896_(_052686_, _052697_, _052698_);
  or g_090897_(_052687_, _052696_, _052699_);
  and g_090898_(_052680_, _052698_, _052700_);
  or g_090899_(_052681_, _052699_, _052701_);
  and g_090900_(_052463_, _052622_, _052702_);
  not g_090901_(_052702_, _052703_);
  or g_090902_(_052461_, _052622_, _052704_);
  not g_090903_(_052704_, _052705_);
  and g_090904_(_052703_, _052704_, _052706_);
  or g_090905_(_052702_, _052705_, _052707_);
  xor g_090906_(out[376], _014563_, _052708_);
  not g_090907_(_052708_, _052709_);
  and g_090908_(_052706_, _052708_, _052710_);
  or g_090909_(_052707_, _052709_, _052711_);
  or g_090910_(_052689_, _052694_, _052712_);
  not g_090911_(_052712_, _052713_);
  and g_090912_(_052711_, _052712_, _052714_);
  or g_090913_(_052710_, _052713_, _052715_);
  and g_090914_(_052707_, _052709_, _052716_);
  or g_090915_(_052706_, _052708_, _052717_);
  and g_090916_(_052714_, _052717_, _052718_);
  or g_090917_(_052701_, _052716_, _052719_);
  and g_090918_(_052700_, _052718_, _052720_);
  or g_090919_(_052715_, _052719_, _052721_);
  and g_090920_(_026234_, _052628_, _052722_);
  or g_090921_(_026245_, _052629_, _052723_);
  or g_090922_(_052667_, _052721_, _052724_);
  or g_090923_(_052722_, _052724_, _052725_);
  not g_090924_(_052725_, _052726_);
  and g_090925_(_052641_, _052660_, _052727_);
  or g_090926_(_026212_, _052655_, _052728_);
  and g_090927_(_052723_, _052728_, _052729_);
  and g_090928_(_052727_, _052729_, _052730_);
  and g_090929_(_052658_, _052663_, _052731_);
  xor g_090930_(_026223_, _052655_, _052732_);
  or g_090931_(_052659_, _052732_, _052733_);
  or g_090932_(_052649_, _052733_, _052734_);
  or g_090933_(_052640_, _052664_, _052735_);
  or g_090934_(_052722_, _052735_, _052736_);
  and g_090935_(_052730_, _052731_, _052737_);
  or g_090936_(_052734_, _052736_, _052738_);
  and g_090937_(_052720_, _052737_, _052739_);
  or g_090938_(_052721_, _052738_, _052740_);
  or g_090939_(out[370], out[369], _052741_);
  xor g_090940_(out[370], out[369], _052742_);
  xor g_090941_(_053709_, out[369], _052743_);
  and g_090942_(_052552_, _052623_, _052744_);
  and g_090943_(_052549_, _052622_, _052745_);
  or g_090944_(_052744_, _052745_, _052746_);
  or g_090945_(_052742_, _052746_, _052747_);
  xor g_090946_(out[371], _014497_, _052748_);
  xor g_090947_(_053687_, _014497_, _052749_);
  or g_090948_(_052544_, _052622_, _052750_);
  or g_090949_(_052539_, _052623_, _052751_);
  and g_090950_(_052750_, _052751_, _052752_);
  or g_090951_(_052749_, _052752_, _052753_);
  and g_090952_(_052749_, _052752_, _052754_);
  xor g_090953_(_052742_, _052746_, _052755_);
  xor g_090954_(_052743_, _052746_, _052756_);
  xor g_090955_(_052749_, _052752_, _052757_);
  xor g_090956_(_052748_, _052752_, _052758_);
  and g_090957_(_052755_, _052757_, _052759_);
  or g_090958_(_052756_, _052758_, _052760_);
  or g_090959_(_053621_, _052623_, _052761_);
  or g_090960_(_052567_, _052622_, _052762_);
  and g_090961_(_052761_, _052762_, _052763_);
  and g_090962_(out[369], _052763_, _052764_);
  or g_090963_(_052575_, _052622_, _052765_);
  or g_090964_(out[352], _052623_, _052766_);
  and g_090965_(_052765_, _052766_, _052767_);
  or g_090966_(_004641_, _052767_, _052768_);
  xor g_090967_(out[369], _052763_, _052769_);
  and g_090968_(_052768_, _052769_, _052770_);
  or g_090969_(_052764_, _052770_, _052771_);
  and g_090970_(_052759_, _052771_, _052772_);
  or g_090971_(_052747_, _052754_, _052773_);
  and g_090972_(_052753_, _052773_, _052774_);
  not g_090973_(_052774_, _052775_);
  or g_090974_(_052772_, _052775_, _052776_);
  not g_090975_(_052776_, _052777_);
  and g_090976_(_052739_, _052776_, _052778_);
  or g_090977_(_052740_, _052777_, _052779_);
  and g_090978_(_052681_, _052683_, _052780_);
  or g_090979_(_052680_, _052682_, _052781_);
  or g_090980_(_052701_, _052714_, _052782_);
  not g_090981_(_052782_, _052783_);
  and g_090982_(_052781_, _052782_, _052784_);
  or g_090983_(_052780_, _052783_, _052785_);
  and g_090984_(_052779_, _052784_, _052786_);
  or g_090985_(_052778_, _052785_, _052787_);
  and g_090986_(_052725_, _052786_, _052788_);
  or g_090987_(_052726_, _052787_, _052789_);
  and g_090988_(_004641_, _052767_, _052790_);
  or g_090989_(_052760_, _052790_, _052791_);
  not g_090990_(_052791_, _052792_);
  and g_090991_(_052770_, _052792_, _052793_);
  not g_090992_(_052793_, _052794_);
  or g_090993_(_052740_, _052794_, _052795_);
  not g_090994_(_052795_, _052796_);
  and g_090995_(_052789_, _052795_, _052797_);
  or g_090996_(_052788_, _052796_, _052798_);
  and g_090997_(_026212_, _052797_, _052799_);
  not g_090998_(_052799_, _052800_);
  or g_090999_(_052655_, _052797_, _052801_);
  not g_091000_(_052801_, _052802_);
  and g_091001_(_052800_, _052801_, _052803_);
  or g_091002_(_052799_, _052802_, _052804_);
  and g_091003_(_026190_, _052803_, _052805_);
  or g_091004_(_026201_, _052804_, _052806_);
  xor g_091005_(out[389], _014684_, _052807_);
  xor g_091006_(_053764_, _014684_, _052808_);
  and g_091007_(_052644_, _052797_, _052809_);
  not g_091008_(_052809_, _052810_);
  or g_091009_(_052647_, _052797_, _052811_);
  not g_091010_(_052811_, _052812_);
  and g_091011_(_052810_, _052811_, _052813_);
  or g_091012_(_052809_, _052812_, _052814_);
  and g_091013_(_052807_, _052814_, _052815_);
  or g_091014_(_052808_, _052813_, _052816_);
  and g_091015_(_052806_, _052816_, _052817_);
  or g_091016_(_052805_, _052815_, _052818_);
  and g_091017_(_026201_, _052804_, _052819_);
  or g_091018_(_026190_, _052803_, _052820_);
  and g_091019_(_052817_, _052820_, _052821_);
  or g_091020_(_052818_, _052819_, _052822_);
  and g_091021_(_014629_, _014772_, _052823_);
  or g_091022_(_014640_, _014761_, _052824_);
  and g_091023_(_052675_, _052798_, _052825_);
  or g_091024_(_052674_, _052797_, _052826_);
  and g_091025_(_052676_, _052797_, _052827_);
  or g_091026_(_052677_, _052798_, _052828_);
  and g_091027_(_052826_, _052828_, _052829_);
  or g_091028_(_052825_, _052827_, _052830_);
  and g_091029_(_026168_, _052829_, _052831_);
  or g_091030_(_026179_, _052830_, _052832_);
  and g_091031_(_052824_, _052832_, _052833_);
  or g_091032_(_052823_, _052831_, _052834_);
  and g_091033_(_014640_, _014761_, _052835_);
  or g_091034_(_014629_, _014772_, _052836_);
  and g_091035_(_026179_, _052830_, _052837_);
  or g_091036_(_026168_, _052829_, _052838_);
  and g_091037_(_052836_, _052838_, _052839_);
  or g_091038_(_052835_, _052837_, _052840_);
  and g_091039_(_052833_, _052839_, _052841_);
  or g_091040_(_052834_, _052840_, _052842_);
  xor g_091041_(out[393], _014728_, _052843_);
  xor g_091042_(_053830_, _014728_, _052844_);
  and g_091043_(_052689_, _052797_, _052845_);
  not g_091044_(_052845_, _052846_);
  or g_091045_(_052694_, _052797_, _052847_);
  not g_091046_(_052847_, _052848_);
  and g_091047_(_052846_, _052847_, _052849_);
  or g_091048_(_052845_, _052848_, _052850_);
  and g_091049_(_052843_, _052850_, _052851_);
  or g_091050_(_052844_, _052849_, _052852_);
  and g_091051_(_052708_, _052797_, _052853_);
  not g_091052_(_052853_, _052854_);
  or g_091053_(_052706_, _052797_, _052855_);
  not g_091054_(_052855_, _052856_);
  and g_091055_(_052854_, _052855_, _052857_);
  or g_091056_(_052853_, _052856_, _052858_);
  xor g_091057_(out[392], _014717_, _052859_);
  xor g_091058_(_053753_, _014717_, _052860_);
  and g_091059_(_052857_, _052859_, _052861_);
  or g_091060_(_052858_, _052860_, _052862_);
  and g_091061_(_052852_, _052862_, _052863_);
  or g_091062_(_052851_, _052861_, _052864_);
  and g_091063_(_052844_, _052849_, _052865_);
  or g_091064_(_052843_, _052850_, _052866_);
  and g_091065_(_052858_, _052860_, _052867_);
  or g_091066_(_052857_, _052859_, _052868_);
  and g_091067_(_052866_, _052868_, _052869_);
  or g_091068_(_052865_, _052867_, _052870_);
  and g_091069_(_052863_, _052869_, _052871_);
  or g_091070_(_052864_, _052870_, _052872_);
  and g_091071_(_052841_, _052871_, _052873_);
  or g_091072_(_052842_, _052872_, _052874_);
  xor g_091073_(out[390], _014695_, _052875_);
  not g_091074_(_052875_, _052876_);
  and g_091075_(_052633_, _052797_, _052877_);
  not g_091076_(_052877_, _052878_);
  or g_091077_(_052638_, _052797_, _052879_);
  not g_091078_(_052879_, _052880_);
  and g_091079_(_052878_, _052879_, _052881_);
  or g_091080_(_052877_, _052880_, _052882_);
  or g_091081_(_052875_, _052882_, _052883_);
  and g_091082_(_052808_, _052813_, _052884_);
  or g_091083_(_052807_, _052814_, _052885_);
  xor g_091084_(out[391], _014706_, _052886_);
  xor g_091085_(_053742_, _014706_, _052887_);
  and g_091086_(_026234_, _052797_, _052888_);
  or g_091087_(_026245_, _052798_, _052889_);
  and g_091088_(_052629_, _052798_, _052890_);
  or g_091089_(_052628_, _052797_, _052891_);
  and g_091090_(_052889_, _052891_, _052892_);
  or g_091091_(_052888_, _052890_, _052893_);
  and g_091092_(_052886_, _052892_, _052894_);
  or g_091093_(_052886_, _052892_, _052895_);
  xor g_091094_(_052876_, _052881_, _052896_);
  xor g_091095_(_052875_, _052881_, _052897_);
  xor g_091096_(_052886_, _052892_, _052898_);
  xor g_091097_(_052887_, _052892_, _052899_);
  and g_091098_(_052896_, _052898_, _052900_);
  or g_091099_(_052897_, _052899_, _052901_);
  and g_091100_(_052885_, _052900_, _052902_);
  or g_091101_(_052884_, _052901_, _052903_);
  and g_091102_(_052821_, _052902_, _052904_);
  or g_091103_(_052822_, _052903_, _052905_);
  and g_091104_(_052873_, _052904_, _052906_);
  or g_091105_(_052874_, _052905_, _052907_);
  xor g_091106_(out[387], _014651_, _052908_);
  xor g_091107_(_053786_, _014651_, _052909_);
  or g_091108_(_052752_, _052797_, _052910_);
  not g_091109_(_052910_, _052911_);
  and g_091110_(_052749_, _052797_, _052912_);
  not g_091111_(_052912_, _052913_);
  and g_091112_(_052910_, _052913_, _052914_);
  or g_091113_(_052911_, _052912_, _052915_);
  and g_091114_(_052908_, _052915_, _052916_);
  and g_091115_(_052743_, _052797_, _052917_);
  and g_091116_(_052746_, _052798_, _052918_);
  or g_091117_(_052917_, _052918_, _052919_);
  not g_091118_(_052919_, _052920_);
  or g_091119_(out[386], out[385], _052921_);
  xor g_091120_(out[386], out[385], _052922_);
  xor g_091121_(_053808_, out[385], _052923_);
  and g_091122_(_052920_, _052923_, _052924_);
  or g_091123_(_052916_, _052924_, _052925_);
  and g_091124_(_052909_, _052914_, _052926_);
  or g_091125_(_052908_, _052915_, _052927_);
  and g_091126_(_052919_, _052922_, _052928_);
  or g_091127_(_052926_, _052928_, _052929_);
  xor g_091128_(_052909_, _052914_, _052930_);
  xor g_091129_(_052919_, _052922_, _052931_);
  and g_091130_(_052930_, _052931_, _052932_);
  or g_091131_(_052925_, _052929_, _052933_);
  or g_091132_(_053720_, _052798_, _052934_);
  or g_091133_(_052763_, _052797_, _052935_);
  and g_091134_(_052934_, _052935_, _052936_);
  and g_091135_(out[385], _052936_, _052937_);
  or g_091136_(_052767_, _052797_, _052938_);
  not g_091137_(_052938_, _052939_);
  and g_091138_(_004641_, _052797_, _052940_);
  not g_091139_(_052940_, _052941_);
  and g_091140_(_052938_, _052941_, _052942_);
  or g_091141_(_052939_, _052940_, _052943_);
  and g_091142_(out[384], _052943_, _052944_);
  or g_091143_(_004674_, _052942_, _052945_);
  xor g_091144_(out[385], _052936_, _052946_);
  xor g_091145_(_053819_, _052936_, _052947_);
  and g_091146_(_052945_, _052946_, _052948_);
  or g_091147_(_052944_, _052947_, _052949_);
  or g_091148_(_052937_, _052948_, _052950_);
  and g_091149_(_052932_, _052950_, _052951_);
  and g_091150_(_052925_, _052927_, _052952_);
  or g_091151_(_052951_, _052952_, _052953_);
  not g_091152_(_052953_, _052954_);
  and g_091153_(_052906_, _052953_, _052955_);
  or g_091154_(_052907_, _052954_, _052956_);
  and g_091155_(_052883_, _052895_, _052957_);
  or g_091156_(_052894_, _052957_, _052958_);
  not g_091157_(_052958_, _052959_);
  and g_091158_(_052834_, _052836_, _052960_);
  or g_091159_(_052833_, _052835_, _052961_);
  and g_091160_(_052841_, _052864_, _052962_);
  or g_091161_(_052842_, _052863_, _052963_);
  and g_091162_(_052866_, _052962_, _052964_);
  or g_091163_(_052865_, _052963_, _052965_);
  and g_091164_(_052818_, _052902_, _052966_);
  or g_091165_(_052817_, _052903_, _052967_);
  and g_091166_(_052958_, _052967_, _052968_);
  or g_091167_(_052959_, _052966_, _052969_);
  and g_091168_(_052873_, _052969_, _052970_);
  or g_091169_(_052874_, _052968_, _052971_);
  and g_091170_(_052961_, _052971_, _052973_);
  or g_091171_(_052960_, _052970_, _052974_);
  and g_091172_(_052956_, _052973_, _052975_);
  or g_091173_(_052955_, _052964_, _052976_);
  and g_091174_(_052965_, _052975_, _052977_);
  or g_091175_(_052974_, _052976_, _052978_);
  and g_091176_(_004674_, _052942_, _052979_);
  or g_091177_(out[384], _052943_, _052980_);
  and g_091178_(_052932_, _052980_, _052981_);
  or g_091179_(_052949_, _052979_, _052982_);
  and g_091180_(_052948_, _052981_, _052984_);
  or g_091181_(_052933_, _052982_, _052985_);
  and g_091182_(_052906_, _052984_, _052986_);
  or g_091183_(_052907_, _052985_, _052987_);
  and g_091184_(_052978_, _052987_, _052988_);
  or g_091185_(_052977_, _052986_, _052989_);
  and g_091186_(_026168_, _052988_, _052990_);
  not g_091187_(_052990_, _052991_);
  or g_091188_(_052829_, _052988_, _052992_);
  not g_091189_(_052992_, _052993_);
  and g_091190_(_052991_, _052992_, _052995_);
  or g_091191_(_052990_, _052993_, _052996_);
  xor g_091192_(out[403], _014805_, _052997_);
  or g_091193_(_052914_, _052988_, _052998_);
  not g_091194_(_052998_, _052999_);
  and g_091195_(_052909_, _052988_, _053000_);
  not g_091196_(_053000_, _053001_);
  and g_091197_(_052998_, _053001_, _053002_);
  or g_091198_(_052999_, _053000_, _053003_);
  and g_091199_(_052997_, _053003_, _053004_);
  or g_091200_(_052920_, _052988_, _053006_);
  or g_091201_(_052922_, _052989_, _053007_);
  and g_091202_(_053006_, _053007_, _053008_);
  or g_091203_(out[402], out[401], _053009_);
  xor g_091204_(out[402], out[401], _053010_);
  xor g_091205_(_053907_, out[401], _053011_);
  and g_091206_(_053008_, _053011_, _053012_);
  or g_091207_(_053004_, _053012_, _053013_);
  or g_091208_(_052997_, _053003_, _053014_);
  xor g_091209_(_052997_, _053003_, _053015_);
  xor g_091210_(_052997_, _053002_, _053017_);
  xor g_091211_(_053008_, _053011_, _053018_);
  xor g_091212_(_053008_, _053010_, _053019_);
  and g_091213_(_053015_, _053018_, _053020_);
  or g_091214_(_053017_, _053019_, _053021_);
  and g_091215_(out[385], _052988_, _053022_);
  not g_091216_(_053022_, _053023_);
  or g_091217_(_052936_, _052988_, _053024_);
  not g_091218_(_053024_, _053025_);
  and g_091219_(_053023_, _053024_, _053026_);
  or g_091220_(_053022_, _053025_, _053028_);
  and g_091221_(out[401], _053026_, _053029_);
  or g_091222_(_052942_, _052988_, _053030_);
  not g_091223_(_053030_, _053031_);
  and g_091224_(_004674_, _052988_, _053032_);
  not g_091225_(_053032_, _053033_);
  and g_091226_(_053030_, _053033_, _053034_);
  or g_091227_(_053031_, _053032_, _053035_);
  and g_091228_(out[400], _053035_, _053036_);
  or g_091229_(_004707_, _053034_, _053037_);
  xor g_091230_(out[401], _053026_, _053039_);
  xor g_091231_(_053918_, _053026_, _053040_);
  and g_091232_(_053037_, _053039_, _053041_);
  or g_091233_(_053036_, _053040_, _053042_);
  or g_091234_(_053029_, _053041_, _053043_);
  and g_091235_(_053020_, _053043_, _053044_);
  and g_091236_(_053013_, _053014_, _053045_);
  or g_091237_(_053044_, _053045_, _053046_);
  xor g_091238_(out[410], _014893_, _053047_);
  xor g_091239_(_004718_, _014893_, _053048_);
  and g_091240_(_052995_, _053047_, _053050_);
  or g_091241_(_052996_, _053048_, _053051_);
  and g_091242_(_014783_, _014926_, _053052_);
  or g_091243_(_014794_, _014915_, _053053_);
  and g_091244_(_053051_, _053053_, _053054_);
  or g_091245_(_053050_, _053052_, _053055_);
  and g_091246_(_052996_, _053048_, _053056_);
  or g_091247_(_052995_, _053047_, _053057_);
  and g_091248_(_053054_, _053057_, _053058_);
  or g_091249_(_053055_, _053056_, _053059_);
  xor g_091250_(out[409], _014882_, _053061_);
  xor g_091251_(_053929_, _014882_, _053062_);
  or g_091252_(_052849_, _052988_, _053063_);
  not g_091253_(_053063_, _053064_);
  and g_091254_(_052844_, _052988_, _053065_);
  not g_091255_(_053065_, _053066_);
  and g_091256_(_053063_, _053066_, _053067_);
  or g_091257_(_053064_, _053065_, _053068_);
  and g_091258_(_053061_, _053068_, _053069_);
  or g_091259_(_053062_, _053067_, _053070_);
  and g_091260_(_052858_, _052989_, _053072_);
  or g_091261_(_052857_, _052988_, _053073_);
  and g_091262_(_052859_, _052988_, _053074_);
  or g_091263_(_052860_, _052989_, _053075_);
  and g_091264_(_053073_, _053075_, _053076_);
  or g_091265_(_053072_, _053074_, _053077_);
  xor g_091266_(out[408], _014871_, _053078_);
  xor g_091267_(_053852_, _014871_, _053079_);
  and g_091268_(_053076_, _053078_, _053080_);
  or g_091269_(_053077_, _053079_, _053081_);
  and g_091270_(_053070_, _053081_, _053083_);
  or g_091271_(_053069_, _053080_, _053084_);
  and g_091272_(_053062_, _053067_, _053085_);
  or g_091273_(_053061_, _053068_, _053086_);
  and g_091274_(_014794_, _014915_, _053087_);
  or g_091275_(_014783_, _014926_, _053088_);
  and g_091276_(_053077_, _053079_, _053089_);
  or g_091277_(_053076_, _053078_, _053090_);
  and g_091278_(_053088_, _053090_, _053091_);
  or g_091279_(_053087_, _053089_, _053092_);
  and g_091280_(_053086_, _053091_, _053094_);
  or g_091281_(_053085_, _053092_, _053095_);
  and g_091282_(_053083_, _053094_, _053096_);
  or g_091283_(_053084_, _053095_, _053097_);
  and g_091284_(_053058_, _053096_, _053098_);
  or g_091285_(_053059_, _053097_, _053099_);
  xor g_091286_(out[407], _014860_, _053100_);
  xor g_091287_(_053841_, _014860_, _053101_);
  and g_091288_(_052893_, _052989_, _053102_);
  or g_091289_(_052892_, _052988_, _053103_);
  and g_091290_(_052886_, _052988_, _053105_);
  or g_091291_(_052887_, _052989_, _053106_);
  and g_091292_(_053103_, _053106_, _053107_);
  or g_091293_(_053102_, _053105_, _053108_);
  and g_091294_(_053100_, _053107_, _053109_);
  xor g_091295_(out[406], _014849_, _053110_);
  or g_091296_(_052881_, _052988_, _053111_);
  not g_091297_(_053111_, _053112_);
  and g_091298_(_052876_, _052988_, _053113_);
  not g_091299_(_053113_, _053114_);
  and g_091300_(_053111_, _053114_, _053116_);
  or g_091301_(_053112_, _053113_, _053117_);
  xor g_091302_(out[405], _014838_, _053118_);
  xor g_091303_(_053863_, _014838_, _053119_);
  or g_091304_(_052813_, _052988_, _053120_);
  not g_091305_(_053120_, _053121_);
  and g_091306_(_052808_, _052988_, _053122_);
  not g_091307_(_053122_, _053123_);
  and g_091308_(_053120_, _053123_, _053124_);
  or g_091309_(_053121_, _053122_, _053125_);
  and g_091310_(_053119_, _053124_, _053127_);
  or g_091311_(_053118_, _053125_, _053128_);
  xor g_091312_(out[404], _014827_, _053129_);
  xor g_091313_(_053896_, _014827_, _053130_);
  or g_091314_(_052803_, _052988_, _053131_);
  not g_091315_(_053131_, _053132_);
  and g_091316_(_026190_, _052988_, _053133_);
  not g_091317_(_053133_, _053134_);
  and g_091318_(_053131_, _053134_, _053135_);
  or g_091319_(_053132_, _053133_, _053136_);
  and g_091320_(_053130_, _053136_, _053138_);
  or g_091321_(_053129_, _053135_, _053139_);
  and g_091322_(_053128_, _053139_, _053140_);
  or g_091323_(_053127_, _053138_, _053141_);
  and g_091324_(_053118_, _053125_, _053142_);
  or g_091325_(_053119_, _053124_, _053143_);
  and g_091326_(_053129_, _053135_, _053144_);
  or g_091327_(_053130_, _053136_, _053145_);
  and g_091328_(_053143_, _053145_, _053146_);
  or g_091329_(_053142_, _053144_, _053147_);
  or g_091330_(_053110_, _053117_, _053149_);
  or g_091331_(_053100_, _053107_, _053150_);
  and g_091332_(_053149_, _053150_, _053151_);
  xor g_091333_(_053100_, _053107_, _053152_);
  xor g_091334_(_053101_, _053107_, _053153_);
  xor g_091335_(_053110_, _053117_, _053154_);
  xor g_091336_(_053110_, _053116_, _053155_);
  and g_091337_(_053152_, _053154_, _053156_);
  or g_091338_(_053153_, _053155_, _053157_);
  and g_091339_(_053140_, _053156_, _053158_);
  or g_091340_(_053141_, _053157_, _053160_);
  and g_091341_(_053146_, _053158_, _053161_);
  or g_091342_(_053147_, _053160_, _053162_);
  and g_091343_(_053098_, _053161_, _053163_);
  or g_091344_(_053099_, _053162_, _053164_);
  and g_091345_(_053046_, _053163_, _053165_);
  or g_091346_(_053109_, _053151_, _053166_);
  not g_091347_(_053166_, _053167_);
  and g_091348_(_053128_, _053156_, _053168_);
  and g_091349_(_053147_, _053168_, _053169_);
  or g_091350_(_053167_, _053169_, _053171_);
  and g_091351_(_053098_, _053171_, _053172_);
  and g_091352_(_053084_, _053086_, _053173_);
  and g_091353_(_053058_, _053173_, _053174_);
  or g_091354_(_053055_, _053174_, _053175_);
  and g_091355_(_053088_, _053175_, _053176_);
  or g_091356_(_053172_, _053176_, _053177_);
  or g_091357_(_053165_, _053177_, _053178_);
  not g_091358_(_053178_, _053179_);
  and g_091359_(_004707_, _053034_, _053180_);
  or g_091360_(out[400], _053035_, _053182_);
  and g_091361_(_053020_, _053182_, _053183_);
  or g_091362_(_053021_, _053180_, _053184_);
  and g_091363_(_053041_, _053183_, _053185_);
  or g_091364_(_053042_, _053184_, _053186_);
  and g_091365_(_053163_, _053185_, _053187_);
  or g_091366_(_053164_, _053186_, _053188_);
  and g_091367_(_053178_, _053188_, _053189_);
  or g_091368_(_053179_, _053187_, _053190_);
  and g_091369_(_052996_, _053190_, _053191_);
  not g_091370_(_053191_, _053193_);
  or g_091371_(_053048_, _053190_, _053194_);
  not g_091372_(_053194_, _053195_);
  and g_091373_(_053193_, _053194_, _053196_);
  or g_091374_(_053191_, _053195_, _053197_);
  or g_091375_(_014937_, _015080_, _053198_);
  xor g_091376_(out[426], _015047_, _053199_);
  xor g_091377_(_004751_, _015047_, _053200_);
  and g_091378_(_053196_, _053199_, _053201_);
  or g_091379_(_053197_, _053200_, _053202_);
  and g_091380_(_014937_, _015080_, _053204_);
  or g_091381_(_014948_, _015069_, _053205_);
  and g_091382_(_053202_, _053205_, _053206_);
  or g_091383_(_053201_, _053204_, _053207_);
  and g_091384_(_053198_, _053207_, _053208_);
  or g_091385_(_053196_, _053199_, _053209_);
  and g_091386_(_053198_, _053209_, _053210_);
  and g_091387_(_053206_, _053210_, _053211_);
  xor g_091388_(out[422], _015003_, _053212_);
  xor g_091389_(_053973_, _015003_, _053213_);
  or g_091390_(_053110_, _053190_, _053215_);
  not g_091391_(_053215_, _053216_);
  and g_091392_(_053117_, _053190_, _053217_);
  not g_091393_(_053217_, _053218_);
  and g_091394_(_053215_, _053218_, _053219_);
  or g_091395_(_053216_, _053217_, _053220_);
  and g_091396_(_053213_, _053219_, _053221_);
  xor g_091397_(out[423], _015014_, _053222_);
  xor g_091398_(_053940_, _015014_, _053223_);
  or g_091399_(_053101_, _053190_, _053224_);
  not g_091400_(_053224_, _053226_);
  and g_091401_(_053108_, _053190_, _053227_);
  not g_091402_(_053227_, _053228_);
  and g_091403_(_053224_, _053228_, _053229_);
  or g_091404_(_053226_, _053227_, _053230_);
  and g_091405_(_053223_, _053230_, _053231_);
  or g_091406_(_053221_, _053231_, _053232_);
  xor g_091407_(out[420], _014981_, _053233_);
  xor g_091408_(_053995_, _014981_, _053234_);
  or g_091409_(_053130_, _053190_, _053235_);
  not g_091410_(_053235_, _053237_);
  and g_091411_(_053136_, _053190_, _053238_);
  not g_091412_(_053238_, _053239_);
  and g_091413_(_053235_, _053239_, _053240_);
  or g_091414_(_053237_, _053238_, _053241_);
  and g_091415_(_053233_, _053240_, _053242_);
  xor g_091416_(out[421], _014992_, _053243_);
  xor g_091417_(_053962_, _014992_, _053244_);
  or g_091418_(_053118_, _053190_, _053245_);
  not g_091419_(_053245_, _053246_);
  and g_091420_(_053125_, _053190_, _053248_);
  not g_091421_(_053248_, _053249_);
  and g_091422_(_053245_, _053249_, _053250_);
  or g_091423_(_053246_, _053248_, _053251_);
  and g_091424_(_053243_, _053251_, _053252_);
  or g_091425_(_053242_, _053252_, _053253_);
  xor g_091426_(out[419], _014959_, _053254_);
  xor g_091427_(_053984_, _014959_, _053255_);
  and g_091428_(_053003_, _053190_, _053256_);
  not g_091429_(_053256_, _053257_);
  or g_091430_(_052997_, _053190_, _053259_);
  not g_091431_(_053259_, _053260_);
  and g_091432_(_053257_, _053259_, _053261_);
  or g_091433_(_053256_, _053260_, _053262_);
  and g_091434_(_053255_, _053261_, _053263_);
  or g_091435_(_053254_, _053262_, _053264_);
  and g_091436_(_053254_, _053262_, _053265_);
  or g_091437_(_053008_, _053189_, _053266_);
  or g_091438_(_053010_, _053190_, _053267_);
  and g_091439_(_053266_, _053267_, _053268_);
  or g_091440_(out[418], out[417], _053270_);
  xor g_091441_(out[418], out[417], _053271_);
  xor g_091442_(_054006_, out[417], _053272_);
  and g_091443_(_053268_, _053272_, _053273_);
  or g_091444_(_053265_, _053273_, _053274_);
  and g_091445_(_053264_, _053274_, _053275_);
  or g_091446_(_053918_, _053190_, _053276_);
  not g_091447_(_053276_, _053277_);
  and g_091448_(_053028_, _053190_, _053278_);
  or g_091449_(_053026_, _053189_, _053279_);
  and g_091450_(_053276_, _053279_, _053281_);
  or g_091451_(_053277_, _053278_, _053282_);
  and g_091452_(out[417], _053281_, _053283_);
  and g_091453_(_053035_, _053190_, _053284_);
  or g_091454_(_053034_, _053189_, _053285_);
  or g_091455_(out[400], _053190_, _053286_);
  not g_091456_(_053286_, _053287_);
  and g_091457_(_053285_, _053286_, _053288_);
  or g_091458_(_053284_, _053287_, _053289_);
  and g_091459_(out[416], _053289_, _053290_);
  or g_091460_(_004740_, _053288_, _053292_);
  or g_091461_(out[417], _053281_, _053293_);
  and g_091462_(_053292_, _053293_, _053294_);
  xor g_091463_(_054017_, _053281_, _053295_);
  or g_091464_(_053290_, _053295_, _053296_);
  or g_091465_(_053283_, _053294_, _053297_);
  xor g_091466_(_053268_, _053272_, _053298_);
  xor g_091467_(_053268_, _053271_, _053299_);
  and g_091468_(_053264_, _053298_, _053300_);
  or g_091469_(_053263_, _053299_, _053301_);
  and g_091470_(_053297_, _053300_, _053303_);
  or g_091471_(_053275_, _053303_, _053304_);
  and g_091472_(_053234_, _053241_, _053305_);
  or g_091473_(_053233_, _053240_, _053306_);
  and g_091474_(_053304_, _053306_, _053307_);
  or g_091475_(_053253_, _053307_, _053308_);
  and g_091476_(_053244_, _053250_, _053309_);
  or g_091477_(_053243_, _053251_, _053310_);
  and g_091478_(_053212_, _053220_, _053311_);
  or g_091479_(_053213_, _053219_, _053312_);
  and g_091480_(_053310_, _053312_, _053314_);
  and g_091481_(_053308_, _053314_, _053315_);
  or g_091482_(_053232_, _053315_, _053316_);
  xor g_091483_(out[425], _015036_, _053317_);
  or g_091484_(_053061_, _053190_, _053318_);
  not g_091485_(_053318_, _053319_);
  and g_091486_(_053068_, _053190_, _053320_);
  not g_091487_(_053320_, _053321_);
  and g_091488_(_053318_, _053321_, _053322_);
  or g_091489_(_053319_, _053320_, _053323_);
  or g_091490_(_053317_, _053323_, _053325_);
  and g_091491_(_053317_, _053323_, _053326_);
  xor g_091492_(_053317_, _053323_, _053327_);
  xor g_091493_(_053317_, _053322_, _053328_);
  or g_091494_(_053079_, _053190_, _053329_);
  not g_091495_(_053329_, _053330_);
  and g_091496_(_053077_, _053190_, _053331_);
  not g_091497_(_053331_, _053332_);
  and g_091498_(_053329_, _053332_, _053333_);
  or g_091499_(_053330_, _053331_, _053334_);
  xor g_091500_(out[424], _015025_, _053336_);
  and g_091501_(_053333_, _053336_, _053337_);
  xor g_091502_(_053333_, _053336_, _053338_);
  xor g_091503_(_053334_, _053336_, _053339_);
  and g_091504_(_053327_, _053338_, _053340_);
  or g_091505_(_053328_, _053339_, _053341_);
  and g_091506_(_053222_, _053229_, _053342_);
  or g_091507_(_053223_, _053230_, _053343_);
  and g_091508_(_053340_, _053343_, _053344_);
  or g_091509_(_053309_, _053342_, _053345_);
  or g_091510_(_053232_, _053311_, _053347_);
  or g_091511_(_053345_, _053347_, _053348_);
  and g_091512_(_053316_, _053344_, _053349_);
  and g_091513_(_053325_, _053337_, _053350_);
  or g_091514_(_053326_, _053350_, _053351_);
  or g_091515_(_053349_, _053351_, _053352_);
  and g_091516_(_053211_, _053352_, _053353_);
  or g_091517_(_053208_, _053353_, _053354_);
  or g_091518_(out[416], _053289_, _053355_);
  or g_091519_(_053265_, _053296_, _053356_);
  or g_091520_(_053305_, _053356_, _053358_);
  or g_091521_(_053253_, _053341_, _053359_);
  or g_091522_(_053301_, _053359_, _053360_);
  or g_091523_(_053358_, _053360_, _053361_);
  and g_091524_(_053211_, _053355_, _053362_);
  not g_091525_(_053362_, _053363_);
  or g_091526_(_053361_, _053363_, _053364_);
  or g_091527_(_053348_, _053364_, _053365_);
  and g_091528_(_053354_, _053365_, _053366_);
  not g_091529_(_053366_, _053367_);
  or g_091530_(_053196_, _053366_, _053369_);
  or g_091531_(_053200_, _053367_, _053370_);
  and g_091532_(_053369_, _053370_, _053371_);
  xor g_091533_(out[435], _015113_, _053372_);
  xor g_091534_(_054083_, _015113_, _053373_);
  and g_091535_(_053254_, _053366_, _053374_);
  not g_091536_(_053374_, _053375_);
  and g_091537_(_053261_, _053367_, _053376_);
  or g_091538_(_053262_, _053366_, _053377_);
  or g_091539_(_053374_, _053376_, _053378_);
  and g_091540_(_053375_, _053377_, _053380_);
  or g_091541_(_053373_, _053378_, _053381_);
  not g_091542_(_053381_, _053382_);
  or g_091543_(_053268_, _053366_, _053383_);
  or g_091544_(_053271_, _053367_, _053384_);
  and g_091545_(_053383_, _053384_, _053385_);
  or g_091546_(out[434], out[433], _053386_);
  xor g_091547_(out[434], out[433], _053387_);
  xor g_091548_(_054105_, out[433], _053388_);
  or g_091549_(_053372_, _053380_, _053389_);
  and g_091550_(_053385_, _053388_, _053391_);
  and g_091551_(_053381_, _053389_, _053392_);
  xor g_091552_(_053372_, _053378_, _053393_);
  xor g_091553_(_053385_, _053388_, _053394_);
  xor g_091554_(_053385_, _053387_, _053395_);
  and g_091555_(_053392_, _053394_, _053396_);
  or g_091556_(_053393_, _053395_, _053397_);
  and g_091557_(out[417], _053366_, _053398_);
  and g_091558_(_053282_, _053367_, _053399_);
  or g_091559_(_053398_, _053399_, _053400_);
  or g_091560_(_053288_, _053366_, _053402_);
  or g_091561_(out[416], _053367_, _053403_);
  and g_091562_(_053402_, _053403_, _053404_);
  not g_091563_(_053404_, _053405_);
  and g_091564_(out[432], _053405_, _053406_);
  or g_091565_(_004773_, _053404_, _053407_);
  or g_091566_(_054116_, _053400_, _053408_);
  not g_091567_(_053408_, _053409_);
  xor g_091568_(_054116_, _053400_, _053410_);
  xor g_091569_(out[433], _053400_, _053411_);
  and g_091570_(_053407_, _053410_, _053413_);
  or g_091571_(_053406_, _053411_, _053414_);
  and g_091572_(_004773_, _053404_, _053415_);
  or g_091573_(_053414_, _053415_, _053416_);
  or g_091574_(_053397_, _053416_, _053417_);
  and g_091575_(_015091_, _015234_, _053418_);
  or g_091576_(_015102_, _015223_, _053419_);
  xor g_091577_(out[442], _015201_, _053420_);
  and g_091578_(_053371_, _053420_, _053421_);
  not g_091579_(_053421_, _053422_);
  and g_091580_(_053419_, _053422_, _053424_);
  or g_091581_(_053418_, _053421_, _053425_);
  or g_091582_(_053371_, _053420_, _053426_);
  or g_091583_(_015091_, _015234_, _053427_);
  and g_091584_(_053426_, _053427_, _053428_);
  not g_091585_(_053428_, _053429_);
  and g_091586_(_053424_, _053428_, _053430_);
  or g_091587_(_053425_, _053429_, _053431_);
  xor g_091588_(out[441], _015190_, _053432_);
  xor g_091589_(_054127_, _015190_, _053433_);
  or g_091590_(_053317_, _053367_, _053435_);
  or g_091591_(_053322_, _053366_, _053436_);
  and g_091592_(_053435_, _053436_, _053437_);
  not g_091593_(_053437_, _053438_);
  and g_091594_(_053432_, _053438_, _053439_);
  or g_091595_(_053433_, _053437_, _053440_);
  and g_091596_(_053336_, _053366_, _053441_);
  not g_091597_(_053441_, _053442_);
  and g_091598_(_053334_, _053367_, _053443_);
  or g_091599_(_053333_, _053366_, _053444_);
  and g_091600_(_053442_, _053444_, _053446_);
  or g_091601_(_053441_, _053443_, _053447_);
  xor g_091602_(out[440], _015179_, _053448_);
  not g_091603_(_053448_, _053449_);
  and g_091604_(_053446_, _053448_, _053450_);
  or g_091605_(_053447_, _053449_, _053451_);
  and g_091606_(_053440_, _053451_, _053452_);
  or g_091607_(_053439_, _053450_, _053453_);
  and g_091608_(_053447_, _053449_, _053454_);
  or g_091609_(_053446_, _053448_, _053455_);
  and g_091610_(_053433_, _053437_, _053457_);
  or g_091611_(_053432_, _053438_, _053458_);
  and g_091612_(_053455_, _053458_, _053459_);
  or g_091613_(_053454_, _053457_, _053460_);
  and g_091614_(_053452_, _053459_, _053461_);
  or g_091615_(_053453_, _053460_, _053462_);
  and g_091616_(_053430_, _053461_, _053463_);
  or g_091617_(_053431_, _053462_, _053464_);
  xor g_091618_(out[438], _015157_, _053465_);
  and g_091619_(_053219_, _053367_, _053466_);
  or g_091620_(_053220_, _053366_, _053468_);
  and g_091621_(_053212_, _053366_, _053469_);
  not g_091622_(_053469_, _053470_);
  or g_091623_(_053466_, _053469_, _053471_);
  and g_091624_(_053468_, _053470_, _053472_);
  or g_091625_(_053465_, _053472_, _053473_);
  xor g_091626_(out[439], _015168_, _053474_);
  and g_091627_(_053222_, _053366_, _053475_);
  not g_091628_(_053475_, _053476_);
  and g_091629_(_053230_, _053367_, _053477_);
  or g_091630_(_053229_, _053366_, _053479_);
  and g_091631_(_053476_, _053479_, _053480_);
  or g_091632_(_053475_, _053477_, _053481_);
  or g_091633_(_053474_, _053480_, _053482_);
  and g_091634_(_053473_, _053482_, _053483_);
  and g_091635_(_053474_, _053480_, _053484_);
  xor g_091636_(_053465_, _053472_, _053485_);
  xor g_091637_(_053465_, _053471_, _053486_);
  xor g_091638_(_053474_, _053480_, _053487_);
  xor g_091639_(_053474_, _053481_, _053488_);
  and g_091640_(_053485_, _053487_, _053490_);
  or g_091641_(_053486_, _053488_, _053491_);
  xor g_091642_(out[437], _015146_, _053492_);
  xor g_091643_(_054061_, _015146_, _053493_);
  or g_091644_(_053243_, _053367_, _053494_);
  or g_091645_(_053250_, _053366_, _053495_);
  and g_091646_(_053494_, _053495_, _053496_);
  not g_091647_(_053496_, _053497_);
  and g_091648_(_053492_, _053497_, _053498_);
  or g_091649_(_053493_, _053496_, _053499_);
  xor g_091650_(out[436], _015135_, _053501_);
  or g_091651_(_053234_, _053367_, _053502_);
  or g_091652_(_053240_, _053366_, _053503_);
  and g_091653_(_053502_, _053503_, _053504_);
  and g_091654_(_053501_, _053504_, _053505_);
  not g_091655_(_053505_, _053506_);
  and g_091656_(_053499_, _053506_, _053507_);
  or g_091657_(_053498_, _053505_, _053508_);
  and g_091658_(_053493_, _053496_, _053509_);
  or g_091659_(_053492_, _053497_, _053510_);
  or g_091660_(_053501_, _053504_, _053512_);
  not g_091661_(_053512_, _053513_);
  and g_091662_(_053510_, _053512_, _053514_);
  or g_091663_(_053509_, _053513_, _053515_);
  and g_091664_(_053507_, _053514_, _053516_);
  or g_091665_(_053508_, _053515_, _053517_);
  and g_091666_(_053490_, _053516_, _053518_);
  or g_091667_(_053491_, _053517_, _053519_);
  or g_091668_(_053417_, _053464_, _053520_);
  or g_091669_(_053519_, _053520_, _053521_);
  or g_091670_(_053409_, _053413_, _053523_);
  and g_091671_(_053396_, _053523_, _053524_);
  and g_091672_(_053389_, _053391_, _053525_);
  or g_091673_(_053382_, _053525_, _053526_);
  or g_091674_(_053524_, _053526_, _053527_);
  and g_091675_(_053518_, _053527_, _053528_);
  or g_091676_(_053483_, _053484_, _053529_);
  not g_091677_(_053529_, _053530_);
  and g_091678_(_053490_, _053510_, _053531_);
  and g_091679_(_053508_, _053531_, _053532_);
  or g_091680_(_053530_, _053532_, _053534_);
  or g_091681_(_053528_, _053534_, _053535_);
  and g_091682_(_053463_, _053535_, _053536_);
  and g_091683_(_053425_, _053427_, _053537_);
  and g_091684_(_053453_, _053458_, _053538_);
  and g_091685_(_053430_, _053538_, _053539_);
  or g_091686_(_053537_, _053539_, _053540_);
  or g_091687_(_053536_, _053540_, _053541_);
  and g_091688_(_053521_, _053541_, _053542_);
  not g_091689_(_053542_, _053543_);
  or g_091690_(_053371_, _053542_, _053545_);
  not g_091691_(_053545_, _053546_);
  and g_091692_(_053420_, _053542_, _053547_);
  not g_091693_(_053547_, _053548_);
  and g_091694_(_053545_, _053548_, _053549_);
  or g_091695_(_053546_, _053547_, _053550_);
  xor g_091696_(out[451], _015267_, _053551_);
  or g_091697_(_053378_, _053542_, _053552_);
  not g_091698_(_053552_, _053553_);
  and g_091699_(_053373_, _053542_, _053554_);
  not g_091700_(_053554_, _053556_);
  and g_091701_(_053552_, _053556_, _053557_);
  or g_091702_(_053553_, _053554_, _053558_);
  and g_091703_(_053551_, _053558_, _053559_);
  or g_091704_(out[450], out[449], _053560_);
  xor g_091705_(out[450], out[449], _053561_);
  xor g_091706_(_054204_, out[449], _053562_);
  or g_091707_(_053385_, _053542_, _053563_);
  or g_091708_(_053387_, _053543_, _053564_);
  and g_091709_(_053563_, _053564_, _053565_);
  and g_091710_(_053562_, _053565_, _053567_);
  or g_091711_(_053559_, _053567_, _053568_);
  or g_091712_(_053551_, _053558_, _053569_);
  xor g_091713_(_053551_, _053558_, _053570_);
  xor g_091714_(_053551_, _053557_, _053571_);
  xor g_091715_(_053562_, _053565_, _053572_);
  xor g_091716_(_053561_, _053565_, _053573_);
  and g_091717_(_053570_, _053572_, _053574_);
  or g_091718_(_053571_, _053573_, _053575_);
  and g_091719_(out[433], _053542_, _053576_);
  and g_091720_(_053400_, _053543_, _053578_);
  or g_091721_(_053576_, _053578_, _053579_);
  not g_091722_(_053579_, _053580_);
  and g_091723_(out[449], _053580_, _053581_);
  or g_091724_(_054215_, _053579_, _053582_);
  or g_091725_(_053404_, _053542_, _053583_);
  or g_091726_(out[432], _053543_, _053584_);
  and g_091727_(_053583_, _053584_, _053585_);
  not g_091728_(_053585_, _053586_);
  and g_091729_(out[448], _053586_, _053587_);
  or g_091730_(_004806_, _053585_, _053589_);
  xor g_091731_(_054215_, _053579_, _053590_);
  xor g_091732_(out[449], _053579_, _053591_);
  and g_091733_(_053589_, _053590_, _053592_);
  or g_091734_(_053587_, _053591_, _053593_);
  and g_091735_(_053582_, _053593_, _053594_);
  or g_091736_(_053581_, _053592_, _053595_);
  and g_091737_(_053574_, _053595_, _053596_);
  or g_091738_(_053575_, _053594_, _053597_);
  and g_091739_(_053568_, _053569_, _053598_);
  not g_091740_(_053598_, _053600_);
  and g_091741_(_053597_, _053600_, _053601_);
  or g_091742_(_053596_, _053598_, _053602_);
  and g_091743_(_015245_, _015388_, _053603_);
  or g_091744_(_015256_, _015377_, _053604_);
  xor g_091745_(out[457], _015344_, _053605_);
  xor g_091746_(_054226_, _015344_, _053606_);
  and g_091747_(_053433_, _053542_, _053607_);
  or g_091748_(_053432_, _053543_, _053608_);
  or g_091749_(_053437_, _053542_, _053609_);
  not g_091750_(_053609_, _053611_);
  and g_091751_(_053608_, _053609_, _053612_);
  or g_091752_(_053607_, _053611_, _053613_);
  and g_091753_(_053606_, _053612_, _053614_);
  or g_091754_(_053605_, _053613_, _053615_);
  and g_091755_(_053604_, _053615_, _053616_);
  or g_091756_(_053603_, _053614_, _053617_);
  xor g_091757_(out[458], _015355_, _053618_);
  xor g_091758_(_004817_, _015355_, _053619_);
  and g_091759_(_053550_, _053619_, _053620_);
  or g_091760_(_053549_, _053618_, _053622_);
  and g_091761_(_053448_, _053542_, _053623_);
  not g_091762_(_053623_, _053624_);
  and g_091763_(_053447_, _053543_, _053625_);
  or g_091764_(_053446_, _053542_, _053626_);
  and g_091765_(_053624_, _053626_, _053627_);
  or g_091766_(_053623_, _053625_, _053628_);
  xor g_091767_(out[456], _015333_, _053629_);
  xor g_091768_(_054149_, _015333_, _053630_);
  and g_091769_(_053628_, _053630_, _053631_);
  or g_091770_(_053627_, _053629_, _053633_);
  and g_091771_(_053622_, _053633_, _053634_);
  or g_091772_(_053620_, _053631_, _053635_);
  and g_091773_(_053616_, _053634_, _053636_);
  or g_091774_(_053617_, _053635_, _053637_);
  and g_091775_(_015256_, _015377_, _053638_);
  or g_091776_(_015245_, _015388_, _053639_);
  and g_091777_(_053549_, _053618_, _053640_);
  or g_091778_(_053550_, _053619_, _053641_);
  and g_091779_(_053639_, _053641_, _053642_);
  or g_091780_(_053638_, _053640_, _053644_);
  and g_091781_(_053605_, _053613_, _053645_);
  or g_091782_(_053606_, _053612_, _053646_);
  and g_091783_(_053627_, _053629_, _053647_);
  or g_091784_(_053628_, _053630_, _053648_);
  and g_091785_(_053646_, _053648_, _053649_);
  or g_091786_(_053645_, _053647_, _053650_);
  and g_091787_(_053642_, _053649_, _053651_);
  or g_091788_(_053644_, _053650_, _053652_);
  and g_091789_(_053636_, _053651_, _053653_);
  or g_091790_(_053637_, _053652_, _053655_);
  xor g_091791_(out[454], _015311_, _053656_);
  or g_091792_(_053465_, _053543_, _053657_);
  or g_091793_(_053471_, _053542_, _053658_);
  and g_091794_(_053657_, _053658_, _053659_);
  not g_091795_(_053659_, _053660_);
  xor g_091796_(out[455], _015322_, _053661_);
  not g_091797_(_053661_, _053662_);
  and g_091798_(_053474_, _053542_, _053663_);
  not g_091799_(_053663_, _053664_);
  and g_091800_(_053481_, _053543_, _053666_);
  or g_091801_(_053480_, _053542_, _053667_);
  and g_091802_(_053664_, _053667_, _053668_);
  or g_091803_(_053663_, _053666_, _053669_);
  and g_091804_(_053661_, _053668_, _053670_);
  xor g_091805_(out[453], _015300_, _053671_);
  xor g_091806_(_054160_, _015300_, _053672_);
  and g_091807_(_053493_, _053542_, _053673_);
  or g_091808_(_053492_, _053543_, _053674_);
  or g_091809_(_053496_, _053542_, _053675_);
  not g_091810_(_053675_, _053677_);
  and g_091811_(_053674_, _053675_, _053678_);
  or g_091812_(_053673_, _053677_, _053679_);
  and g_091813_(_053672_, _053678_, _053680_);
  or g_091814_(_053671_, _053679_, _053681_);
  xor g_091815_(out[452], _015289_, _053682_);
  xor g_091816_(_054193_, _015289_, _053683_);
  and g_091817_(_053501_, _053542_, _053684_);
  not g_091818_(_053684_, _053685_);
  or g_091819_(_053504_, _053542_, _053686_);
  not g_091820_(_053686_, _053688_);
  and g_091821_(_053685_, _053686_, _053689_);
  or g_091822_(_053684_, _053688_, _053690_);
  and g_091823_(_053683_, _053690_, _053691_);
  or g_091824_(_053682_, _053689_, _053692_);
  or g_091825_(_053656_, _053660_, _053693_);
  or g_091826_(_053661_, _053668_, _053694_);
  and g_091827_(_053693_, _053694_, _053695_);
  and g_091828_(_053671_, _053679_, _053696_);
  or g_091829_(_053672_, _053678_, _053697_);
  and g_091830_(_053682_, _053689_, _053699_);
  or g_091831_(_053683_, _053690_, _053700_);
  and g_091832_(_053697_, _053700_, _053701_);
  or g_091833_(_053696_, _053699_, _053702_);
  xor g_091834_(_053656_, _053660_, _053703_);
  xor g_091835_(_053656_, _053659_, _053704_);
  xor g_091836_(_053661_, _053668_, _053705_);
  xor g_091837_(_053662_, _053668_, _053706_);
  and g_091838_(_053703_, _053705_, _053707_);
  or g_091839_(_053704_, _053706_, _053708_);
  and g_091840_(_053692_, _053701_, _053710_);
  or g_091841_(_053691_, _053702_, _053711_);
  and g_091842_(_053681_, _053710_, _053712_);
  or g_091843_(_053680_, _053711_, _053713_);
  and g_091844_(_053707_, _053712_, _053714_);
  or g_091845_(_053708_, _053713_, _053715_);
  and g_091846_(_053653_, _053714_, _053716_);
  or g_091847_(_053655_, _053715_, _053717_);
  and g_091848_(_053602_, _053716_, _053718_);
  or g_091849_(_053601_, _053717_, _053719_);
  or g_091850_(_053670_, _053695_, _053721_);
  not g_091851_(_053721_, _053722_);
  and g_091852_(_053702_, _053707_, _053723_);
  or g_091853_(_053701_, _053708_, _053724_);
  and g_091854_(_053681_, _053723_, _053725_);
  or g_091855_(_053680_, _053724_, _053726_);
  and g_091856_(_053721_, _053726_, _053727_);
  or g_091857_(_053722_, _053725_, _053728_);
  and g_091858_(_053653_, _053728_, _053729_);
  or g_091859_(_053655_, _053727_, _053730_);
  and g_091860_(_053615_, _053622_, _053732_);
  or g_091861_(_053614_, _053620_, _053733_);
  and g_091862_(_053650_, _053732_, _053734_);
  or g_091863_(_053649_, _053733_, _053735_);
  and g_091864_(_053642_, _053735_, _053736_);
  or g_091865_(_053644_, _053734_, _053737_);
  and g_091866_(_053604_, _053737_, _053738_);
  or g_091867_(_053603_, _053736_, _053739_);
  and g_091868_(_053730_, _053739_, _053740_);
  or g_091869_(_053729_, _053738_, _053741_);
  and g_091870_(_053719_, _053740_, _053743_);
  or g_091871_(_053718_, _053741_, _053744_);
  and g_091872_(_004806_, _053585_, _053745_);
  or g_091873_(out[448], _053586_, _053746_);
  and g_091874_(_053574_, _053746_, _053747_);
  or g_091875_(_053575_, _053745_, _053748_);
  and g_091876_(_053592_, _053747_, _053749_);
  or g_091877_(_053593_, _053748_, _053750_);
  and g_091878_(_053716_, _053749_, _053751_);
  or g_091879_(_053717_, _053750_, _053752_);
  and g_091880_(_053744_, _053752_, _053754_);
  or g_091881_(_053743_, _053751_, _053755_);
  and g_091882_(_053550_, _053755_, _053756_);
  or g_091883_(_053549_, _053754_, _053757_);
  and g_091884_(_053618_, _053754_, _053758_);
  or g_091885_(_053619_, _053755_, _053759_);
  and g_091886_(_053757_, _053759_, _053760_);
  or g_091887_(_053756_, _053758_, _053761_);
  and g_091888_(_026157_, _053761_, _053762_);
  not g_091889_(_053762_, _053763_);
  and g_091890_(_015399_, _015542_, _053765_);
  or g_091891_(_015410_, _015531_, _053766_);
  or g_091892_(_053762_, _053765_, _053767_);
  and g_091893_(_053629_, _053754_, _053768_);
  or g_091894_(_053630_, _053755_, _053769_);
  and g_091895_(_053628_, _053755_, _053770_);
  or g_091896_(_053627_, _053754_, _053771_);
  and g_091897_(_053769_, _053771_, _053772_);
  or g_091898_(_053768_, _053770_, _053773_);
  xor g_091899_(out[472], _015487_, _053774_);
  xor g_091900_(_054248_, _015487_, _053776_);
  and g_091901_(_053773_, _053776_, _053777_);
  or g_091902_(_053772_, _053774_, _053778_);
  and g_091903_(_053606_, _053754_, _053779_);
  or g_091904_(_053605_, _053755_, _053780_);
  and g_091905_(_053613_, _053755_, _053781_);
  or g_091906_(_053612_, _053754_, _053782_);
  and g_091907_(_053780_, _053782_, _053783_);
  or g_091908_(_053779_, _053781_, _053784_);
  and g_091909_(_026135_, _053783_, _053785_);
  not g_091910_(_053785_, _053787_);
  or g_091911_(_053777_, _053785_, _053788_);
  or g_091912_(_053767_, _053788_, _053789_);
  and g_091913_(_015410_, _015531_, _053790_);
  or g_091914_(_015399_, _015542_, _053791_);
  and g_091915_(_026146_, _053760_, _053792_);
  or g_091916_(_026157_, _053761_, _053793_);
  and g_091917_(_053791_, _053793_, _053794_);
  or g_091918_(_053790_, _053792_, _053795_);
  and g_091919_(_026124_, _053784_, _053796_);
  or g_091920_(_026135_, _053783_, _053798_);
  and g_091921_(_053772_, _053774_, _053799_);
  or g_091922_(_053773_, _053776_, _053800_);
  and g_091923_(_053798_, _053800_, _053801_);
  or g_091924_(_053796_, _053799_, _053802_);
  or g_091925_(_053795_, _053802_, _053803_);
  and g_091926_(_053763_, _053794_, _053804_);
  and g_091927_(_053766_, _053804_, _053805_);
  and g_091928_(_053787_, _053801_, _053806_);
  and g_091929_(_053778_, _053806_, _053807_);
  and g_091930_(_053805_, _053807_, _053809_);
  or g_091931_(_053789_, _053803_, _053810_);
  xor g_091932_(out[470], _015465_, _053811_);
  not g_091933_(_053811_, _053812_);
  or g_091934_(_053656_, _053755_, _053813_);
  or g_091935_(_053659_, _053754_, _053814_);
  and g_091936_(_053813_, _053814_, _053815_);
  xor g_091937_(out[471], _015476_, _053816_);
  xor g_091938_(_054237_, _015476_, _053817_);
  and g_091939_(_053661_, _053754_, _053818_);
  or g_091940_(_053662_, _053755_, _053820_);
  and g_091941_(_053669_, _053755_, _053821_);
  or g_091942_(_053668_, _053754_, _053822_);
  and g_091943_(_053820_, _053822_, _053823_);
  or g_091944_(_053818_, _053821_, _053824_);
  or g_091945_(_053817_, _053824_, _053825_);
  xor g_091946_(out[468], _015443_, _053826_);
  not g_091947_(_053826_, _053827_);
  and g_091948_(_053682_, _053754_, _053828_);
  or g_091949_(_053683_, _053755_, _053829_);
  and g_091950_(_053690_, _053755_, _053831_);
  or g_091951_(_053689_, _053754_, _053832_);
  and g_091952_(_053829_, _053832_, _053833_);
  or g_091953_(_053828_, _053831_, _053834_);
  and g_091954_(_053827_, _053834_, _053835_);
  or g_091955_(_053826_, _053833_, _053836_);
  xor g_091956_(out[469], _015454_, _053837_);
  xor g_091957_(_054259_, _015454_, _053838_);
  and g_091958_(_053672_, _053754_, _053839_);
  or g_091959_(_053671_, _053755_, _053840_);
  and g_091960_(_053679_, _053755_, _053842_);
  or g_091961_(_053678_, _053754_, _053843_);
  and g_091962_(_053840_, _053843_, _053844_);
  or g_091963_(_053839_, _053842_, _053845_);
  and g_091964_(_053838_, _053844_, _053846_);
  or g_091965_(_053837_, _053845_, _053847_);
  and g_091966_(_053836_, _053847_, _053848_);
  or g_091967_(_053835_, _053846_, _053849_);
  and g_091968_(_053812_, _053815_, _053850_);
  and g_091969_(_053817_, _053824_, _053851_);
  or g_091970_(_053850_, _053851_, _053853_);
  and g_091971_(_053837_, _053845_, _053854_);
  or g_091972_(_053838_, _053844_, _053855_);
  and g_091973_(_053826_, _053833_, _053856_);
  or g_091974_(_053827_, _053834_, _053857_);
  and g_091975_(_053855_, _053857_, _053858_);
  or g_091976_(_053854_, _053856_, _053859_);
  xor g_091977_(_053811_, _053815_, _053860_);
  xor g_091978_(_053817_, _053823_, _053861_);
  or g_091979_(_053860_, _053861_, _053862_);
  not g_091980_(_053862_, _053864_);
  and g_091981_(_053848_, _053855_, _053865_);
  or g_091982_(_053849_, _053854_, _053866_);
  and g_091983_(_053864_, _053865_, _053867_);
  or g_091984_(_053862_, _053866_, _053868_);
  and g_091985_(_053857_, _053867_, _053869_);
  or g_091986_(_053856_, _053868_, _053870_);
  and g_091987_(_053809_, _053869_, _053871_);
  or g_091988_(_053810_, _053870_, _053872_);
  and g_091989_(out[449], _053754_, _053873_);
  and g_091990_(_053579_, _053755_, _053875_);
  or g_091991_(_053873_, _053875_, _053876_);
  not g_091992_(_053876_, _053877_);
  and g_091993_(out[465], _053877_, _053878_);
  or g_091994_(_054314_, _053876_, _053879_);
  or g_091995_(out[466], out[465], _053880_);
  xor g_091996_(out[466], out[465], _053881_);
  xor g_091997_(_054303_, out[465], _053882_);
  or g_091998_(_053565_, _053754_, _053883_);
  or g_091999_(_053561_, _053755_, _053884_);
  and g_092000_(_053883_, _053884_, _053886_);
  not g_092001_(_053886_, _053887_);
  and g_092002_(_053882_, _053886_, _053888_);
  or g_092003_(_053881_, _053887_, _053889_);
  xor g_092004_(_053882_, _053886_, _053890_);
  xor g_092005_(_053881_, _053886_, _053891_);
  xor g_092006_(out[467], _015421_, _053892_);
  xor g_092007_(_054281_, _015421_, _053893_);
  or g_092008_(_053557_, _053754_, _053894_);
  or g_092009_(_053551_, _053755_, _053895_);
  and g_092010_(_053894_, _053895_, _053897_);
  not g_092011_(_053897_, _053898_);
  and g_092012_(_053892_, _053898_, _053899_);
  or g_092013_(_053893_, _053897_, _053900_);
  and g_092014_(_053893_, _053897_, _053901_);
  or g_092015_(_053892_, _053898_, _053902_);
  xor g_092016_(_053893_, _053897_, _053903_);
  xor g_092017_(_053892_, _053897_, _053904_);
  and g_092018_(_053890_, _053903_, _053905_);
  or g_092019_(_053891_, _053904_, _053906_);
  and g_092020_(_053878_, _053905_, _053908_);
  or g_092021_(_053879_, _053906_, _053909_);
  and g_092022_(_054314_, _053876_, _053910_);
  or g_092023_(out[465], _053877_, _053911_);
  or g_092024_(_053585_, _053754_, _053912_);
  or g_092025_(out[448], _053755_, _053913_);
  and g_092026_(_053912_, _053913_, _053914_);
  not g_092027_(_053914_, _053915_);
  and g_092028_(out[464], _053915_, _053916_);
  or g_092029_(_004839_, _053914_, _053917_);
  and g_092030_(_053911_, _053917_, _053919_);
  or g_092031_(_053910_, _053916_, _053920_);
  and g_092032_(_053879_, _053905_, _053921_);
  or g_092033_(_053878_, _053906_, _053922_);
  and g_092034_(_053919_, _053921_, _053923_);
  or g_092035_(_053920_, _053922_, _053924_);
  and g_092036_(_053889_, _053900_, _053925_);
  or g_092037_(_053888_, _053899_, _053926_);
  and g_092038_(_053902_, _053926_, _053927_);
  or g_092039_(_053901_, _053925_, _053928_);
  and g_092040_(_053909_, _053928_, _053930_);
  or g_092041_(_053908_, _053927_, _053931_);
  and g_092042_(_053924_, _053930_, _053932_);
  or g_092043_(_053923_, _053931_, _053933_);
  and g_092044_(_053871_, _053933_, _053934_);
  or g_092045_(_053872_, _053932_, _053935_);
  and g_092046_(_053825_, _053853_, _053936_);
  not g_092047_(_053936_, _053937_);
  and g_092048_(_053847_, _053859_, _053938_);
  or g_092049_(_053846_, _053858_, _053939_);
  and g_092050_(_053864_, _053938_, _053941_);
  or g_092051_(_053862_, _053939_, _053942_);
  and g_092052_(_053937_, _053942_, _053943_);
  or g_092053_(_053936_, _053941_, _053944_);
  and g_092054_(_053809_, _053944_, _053945_);
  or g_092055_(_053810_, _053943_, _053946_);
  or g_092056_(_053762_, _053785_, _053947_);
  or g_092057_(_053801_, _053947_, _053948_);
  and g_092058_(_053794_, _053948_, _053949_);
  not g_092059_(_053949_, _053950_);
  and g_092060_(_053766_, _053950_, _053952_);
  or g_092061_(_053765_, _053949_, _053953_);
  and g_092062_(_053946_, _053953_, _053954_);
  or g_092063_(_053945_, _053952_, _053955_);
  and g_092064_(_053935_, _053954_, _053956_);
  or g_092065_(_053934_, _053955_, _053957_);
  and g_092066_(_004839_, _053914_, _053958_);
  or g_092067_(out[464], _053915_, _053959_);
  and g_092068_(_053923_, _053959_, _053960_);
  or g_092069_(_053924_, _053958_, _053961_);
  and g_092070_(_053871_, _053960_, _053963_);
  or g_092071_(_053872_, _053961_, _053964_);
  and g_092072_(_053957_, _053964_, _053965_);
  or g_092073_(_053956_, _053963_, _053966_);
  or g_092074_(_026124_, _053966_, _053967_);
  or g_092075_(_053783_, _053965_, _053968_);
  and g_092076_(_053967_, _053968_, _053969_);
  xor g_092077_(out[937], _025904_, _053970_);
  not g_092078_(_053970_, _053971_);
  and g_092079_(_025816_, _025937_, _053972_);
  or g_092080_(_025805_, _025948_, _053974_);
  xor g_092081_(out[938], _025915_, _053975_);
  not g_092082_(_053975_, _053976_);
  xor g_092083_(out[922], _025761_, _053977_);
  xor g_092084_(_002067_, _025761_, _053978_);
  xor g_092085_(out[874], _025299_, _053979_);
  and g_092086_(_025189_, _025321_, _053980_);
  xor g_092087_(out[794], _024529_, _053981_);
  xor g_092088_(_001011_, _024529_, _053982_);
  xor g_092089_(out[730], _023913_, _053983_);
  xor g_092090_(_000483_, _023913_, _053985_);
  and g_092091_(_023803_, _023946_, _053986_);
  or g_092092_(_023814_, _023935_, _053987_);
  xor g_092093_(out[714], _023759_, _053988_);
  and g_092094_(_023649_, _023792_, _053989_);
  xor g_092095_(out[666], _023308_, _053990_);
  xor g_092096_(_055920_, _023308_, _053991_);
  xor g_092097_(out[659], _023220_, _053992_);
  xor g_092098_(_055887_, _023220_, _053993_);
  xor g_092099_(out[611], _022758_, _053994_);
  xor g_092100_(_055491_, _022758_, _053996_);
  xor g_092101_(out[618], _022846_, _053997_);
  not g_092102_(_053997_, _053998_);
  and g_092103_(_020008_, _022186_, _053999_);
  and g_092104_(_020052_, _022197_, _054000_);
  or g_092105_(_053999_, _054000_, _054001_);
  not g_092106_(_054001_, _054002_);
  or g_092107_(out[545], out[546], _054003_);
  xor g_092108_(out[545], out[546], _054004_);
  xor g_092109_(_054930_, out[546], _054005_);
  or g_092110_(_021031_, _022186_, _054007_);
  not g_092111_(_054007_, _054008_);
  and g_092112_(_020998_, _022186_, _054009_);
  not g_092113_(_054009_, _054010_);
  and g_092114_(_054007_, _054010_, _054011_);
  or g_092115_(_054008_, _054009_, _054012_);
  and g_092116_(_054005_, _054011_, _054013_);
  or g_092117_(_054004_, _054012_, _054014_);
  xor g_092118_(out[547], _015564_, _054015_);
  xor g_092119_(_054963_, _015564_, _054016_);
  or g_092120_(_020932_, _022186_, _054018_);
  not g_092121_(_054018_, _054019_);
  and g_092122_(_020877_, _022186_, _054020_);
  or g_092123_(_020866_, _022197_, _054021_);
  and g_092124_(_054018_, _054021_, _054022_);
  or g_092125_(_054019_, _054020_, _054023_);
  and g_092126_(_054015_, _054023_, _054024_);
  or g_092127_(_054016_, _054022_, _054025_);
  and g_092128_(_054014_, _054025_, _054026_);
  or g_092129_(_054798_, _022197_, _054027_);
  or g_092130_(_021207_, _022186_, _054029_);
  and g_092131_(_054027_, _054029_, _054030_);
  and g_092132_(out[545], _054030_, _054031_);
  not g_092133_(_054031_, _054032_);
  or g_092134_(_021284_, _022186_, _054033_);
  not g_092135_(_054033_, _054034_);
  and g_092136_(_054809_, _022186_, _054035_);
  or g_092137_(out[528], _022197_, _054036_);
  and g_092138_(_054033_, _054036_, _054037_);
  or g_092139_(_054034_, _054035_, _054038_);
  and g_092140_(out[544], _054038_, _054040_);
  or g_092141_(_054941_, _054037_, _054041_);
  xor g_092142_(out[545], _054030_, _054042_);
  xor g_092143_(_054930_, _054030_, _054043_);
  and g_092144_(_054041_, _054042_, _054044_);
  or g_092145_(_054040_, _054043_, _054045_);
  and g_092146_(_054032_, _054045_, _054046_);
  or g_092147_(_054031_, _054044_, _054047_);
  xor g_092148_(_054005_, _054011_, _054048_);
  xor g_092149_(_054004_, _054011_, _054049_);
  or g_092150_(_054046_, _054049_, _054051_);
  and g_092151_(_054026_, _054051_, _054052_);
  xor g_092152_(out[554], _015652_, _054053_);
  xor g_092153_(_054996_, _015652_, _054054_);
  and g_092154_(_054002_, _054053_, _054055_);
  and g_092155_(_015674_, _022252_, _054056_);
  or g_092156_(_054055_, _054056_, _054057_);
  and g_092157_(_054001_, _054054_, _054058_);
  and g_092158_(_015685_, _022263_, _054059_);
  or g_092159_(_015674_, _022252_, _054060_);
  or g_092160_(_054058_, _054059_, _054062_);
  xor g_092161_(_054001_, _054054_, _054063_);
  xor g_092162_(_015674_, _022252_, _054064_);
  and g_092163_(_054063_, _054064_, _054065_);
  or g_092164_(_054057_, _054062_, _054066_);
  and g_092165_(_020184_, _022197_, _054067_);
  or g_092166_(_020195_, _022186_, _054068_);
  and g_092167_(_020129_, _022186_, _054069_);
  or g_092168_(_020118_, _022197_, _054070_);
  and g_092169_(_054068_, _054070_, _054071_);
  or g_092170_(_054067_, _054069_, _054073_);
  xor g_092171_(out[553], _015641_, _054074_);
  xor g_092172_(_054985_, _015641_, _054075_);
  and g_092173_(_054073_, _054074_, _054076_);
  or g_092174_(_054071_, _054075_, _054077_);
  xor g_092175_(out[552], _015630_, _054078_);
  xor g_092176_(_054974_, _015630_, _054079_);
  and g_092177_(_020327_, _022197_, _054080_);
  or g_092178_(_020316_, _022186_, _054081_);
  and g_092179_(_020250_, _022186_, _054082_);
  or g_092180_(_020261_, _022197_, _054084_);
  and g_092181_(_054081_, _054084_, _054085_);
  or g_092182_(_054080_, _054082_, _054086_);
  and g_092183_(_054078_, _054085_, _054087_);
  or g_092184_(_054079_, _054086_, _054088_);
  and g_092185_(_054077_, _054088_, _054089_);
  or g_092186_(_054076_, _054087_, _054090_);
  and g_092187_(_054071_, _054075_, _054091_);
  or g_092188_(_054073_, _054074_, _054092_);
  and g_092189_(_054079_, _054086_, _054093_);
  or g_092190_(_054078_, _054085_, _054095_);
  and g_092191_(_054092_, _054095_, _054096_);
  or g_092192_(_054091_, _054093_, _054097_);
  and g_092193_(_054089_, _054096_, _054098_);
  or g_092194_(_054090_, _054097_, _054099_);
  and g_092195_(_054065_, _054098_, _054100_);
  or g_092196_(_054066_, _054099_, _054101_);
  xor g_092197_(out[550], _015608_, _054102_);
  not g_092198_(_054102_, _054103_);
  and g_092199_(_020437_, _022197_, _054104_);
  or g_092200_(_020426_, _022186_, _054106_);
  and g_092201_(_020393_, _022186_, _054107_);
  or g_092202_(_020382_, _022197_, _054108_);
  and g_092203_(_054106_, _054108_, _054109_);
  or g_092204_(_054104_, _054107_, _054110_);
  and g_092205_(_054103_, _054109_, _054111_);
  or g_092206_(_054102_, _054110_, _054112_);
  xor g_092207_(out[551], _015619_, _054113_);
  xor g_092208_(_054886_, _015619_, _054114_);
  and g_092209_(_020547_, _022197_, _054115_);
  or g_092210_(_020536_, _022186_, _054117_);
  and g_092211_(_020470_, _022186_, _054118_);
  or g_092212_(_020481_, _022197_, _054119_);
  and g_092213_(_054117_, _054119_, _054120_);
  or g_092214_(_054115_, _054118_, _054121_);
  and g_092215_(_054114_, _054121_, _054122_);
  or g_092216_(_054113_, _054120_, _054123_);
  and g_092217_(_054112_, _054123_, _054124_);
  or g_092218_(_054111_, _054122_, _054125_);
  and g_092219_(_054113_, _054120_, _054126_);
  or g_092220_(_054114_, _054121_, _054128_);
  xor g_092221_(out[548], _015586_, _054129_);
  xor g_092222_(_054919_, _015586_, _054130_);
  and g_092223_(_020734_, _022186_, _054131_);
  or g_092224_(_020745_, _022197_, _054132_);
  and g_092225_(_020811_, _022197_, _054133_);
  or g_092226_(_020800_, _022186_, _054134_);
  and g_092227_(_054132_, _054134_, _054135_);
  or g_092228_(_054131_, _054133_, _054136_);
  and g_092229_(_054130_, _054136_, _054137_);
  or g_092230_(_054129_, _054135_, _054139_);
  and g_092231_(_054128_, _054139_, _054140_);
  or g_092232_(_054126_, _054137_, _054141_);
  and g_092233_(_054124_, _054140_, _054142_);
  or g_092234_(_054125_, _054141_, _054143_);
  xor g_092235_(out[549], _015597_, _054144_);
  xor g_092236_(_054908_, _015597_, _054145_);
  and g_092237_(_020679_, _022197_, _054146_);
  or g_092238_(_020668_, _022186_, _054147_);
  and g_092239_(_020613_, _022186_, _054148_);
  or g_092240_(_020602_, _022197_, _054150_);
  and g_092241_(_054147_, _054150_, _054151_);
  or g_092242_(_054146_, _054148_, _054152_);
  and g_092243_(_054144_, _054152_, _054153_);
  or g_092244_(_054145_, _054151_, _054154_);
  and g_092245_(_054129_, _054135_, _054155_);
  or g_092246_(_054130_, _054136_, _054156_);
  and g_092247_(_054154_, _054156_, _054157_);
  or g_092248_(_054153_, _054155_, _054158_);
  and g_092249_(_054102_, _054110_, _054159_);
  or g_092250_(_054103_, _054109_, _054161_);
  and g_092251_(_054145_, _054151_, _054162_);
  or g_092252_(_054144_, _054152_, _054163_);
  and g_092253_(_054161_, _054163_, _054164_);
  or g_092254_(_054159_, _054162_, _054165_);
  and g_092255_(_054157_, _054164_, _054166_);
  or g_092256_(_054158_, _054165_, _054167_);
  and g_092257_(_054142_, _054166_, _054168_);
  or g_092258_(_054143_, _054167_, _054169_);
  and g_092259_(_054100_, _054168_, _054170_);
  or g_092260_(_054101_, _054169_, _054172_);
  and g_092261_(_054016_, _054022_, _054173_);
  or g_092262_(_054015_, _054023_, _054174_);
  or g_092263_(_054172_, _054173_, _054175_);
  and g_092264_(_054013_, _054174_, _054176_);
  and g_092265_(_054048_, _054174_, _054177_);
  or g_092266_(_054049_, _054173_, _054178_);
  and g_092267_(_054047_, _054177_, _054179_);
  or g_092268_(_054176_, _054179_, _054180_);
  or g_092269_(_054024_, _054180_, _054181_);
  and g_092270_(_054170_, _054181_, _054183_);
  or g_092271_(_054052_, _054175_, _054184_);
  and g_092272_(_054158_, _054164_, _054185_);
  or g_092273_(_054157_, _054165_, _054186_);
  and g_092274_(_054124_, _054186_, _054187_);
  or g_092275_(_054125_, _054185_, _054188_);
  and g_092276_(_054100_, _054188_, _054189_);
  or g_092277_(_054101_, _054187_, _054190_);
  and g_092278_(_054128_, _054189_, _054191_);
  or g_092279_(_054126_, _054190_, _054192_);
  and g_092280_(_054057_, _054060_, _054194_);
  not g_092281_(_054194_, _054195_);
  and g_092282_(_054090_, _054092_, _054196_);
  or g_092283_(_054089_, _054091_, _054197_);
  and g_092284_(_054065_, _054196_, _054198_);
  or g_092285_(_054066_, _054197_, _054199_);
  and g_092286_(_054195_, _054199_, _054200_);
  or g_092287_(_054194_, _054198_, _054201_);
  and g_092288_(_054192_, _054200_, _054202_);
  or g_092289_(_054191_, _054201_, _054203_);
  and g_092290_(_054184_, _054202_, _054205_);
  or g_092291_(_054183_, _054203_, _054206_);
  and g_092292_(_054941_, _054037_, _054207_);
  or g_092293_(out[544], _054038_, _054208_);
  and g_092294_(_054025_, _054208_, _054209_);
  or g_092295_(_054024_, _054207_, _054210_);
  and g_092296_(_054177_, _054209_, _054211_);
  or g_092297_(_054178_, _054210_, _054212_);
  and g_092298_(_054044_, _054211_, _054213_);
  or g_092299_(_054045_, _054212_, _054214_);
  and g_092300_(_054170_, _054213_, _054216_);
  or g_092301_(_054172_, _054214_, _054217_);
  and g_092302_(_054206_, _054217_, _054218_);
  or g_092303_(_054205_, _054216_, _054219_);
  and g_092304_(_054001_, _054219_, _054220_);
  or g_092305_(_054002_, _054218_, _054221_);
  and g_092306_(_054053_, _054218_, _054222_);
  or g_092307_(_054054_, _054219_, _054223_);
  and g_092308_(_054221_, _054223_, _054224_);
  or g_092309_(_054220_, _054222_, _054225_);
  xor g_092310_(out[564], _022318_, _054227_);
  xor g_092311_(_055051_, _022318_, _054228_);
  and g_092312_(_054129_, _054218_, _054229_);
  or g_092313_(_054130_, _054219_, _054230_);
  and g_092314_(_054136_, _054219_, _054231_);
  or g_092315_(_054135_, _054218_, _054232_);
  and g_092316_(_054230_, _054232_, _054233_);
  or g_092317_(_054229_, _054231_, _054234_);
  and g_092318_(_054227_, _054233_, _054235_);
  or g_092319_(_054228_, _054234_, _054236_);
  xor g_092320_(out[565], _022329_, _054238_);
  xor g_092321_(_055040_, _022329_, _054239_);
  and g_092322_(_054145_, _054218_, _054240_);
  or g_092323_(_054144_, _054219_, _054241_);
  and g_092324_(_054152_, _054219_, _054242_);
  or g_092325_(_054151_, _054218_, _054243_);
  and g_092326_(_054241_, _054243_, _054244_);
  or g_092327_(_054240_, _054242_, _054245_);
  and g_092328_(_054238_, _054245_, _054246_);
  or g_092329_(_054239_, _054244_, _054247_);
  and g_092330_(_054236_, _054247_, _054249_);
  or g_092331_(_054235_, _054246_, _054250_);
  xor g_092332_(out[563], _022296_, _054251_);
  not g_092333_(_054251_, _054252_);
  or g_092334_(_054022_, _054218_, _054253_);
  or g_092335_(_054015_, _054219_, _054254_);
  and g_092336_(_054253_, _054254_, _054255_);
  not g_092337_(_054255_, _054256_);
  and g_092338_(_054251_, _054256_, _054257_);
  or g_092339_(_054252_, _054255_, _054258_);
  or g_092340_(out[561], out[562], _054260_);
  xor g_092341_(out[561], out[562], _054261_);
  xor g_092342_(_055062_, out[562], _054262_);
  and g_092343_(_054005_, _054218_, _054263_);
  or g_092344_(_054004_, _054219_, _054264_);
  and g_092345_(_054012_, _054219_, _054265_);
  or g_092346_(_054011_, _054218_, _054266_);
  and g_092347_(_054264_, _054266_, _054267_);
  or g_092348_(_054263_, _054265_, _054268_);
  and g_092349_(_054262_, _054267_, _054269_);
  or g_092350_(_054261_, _054268_, _054271_);
  and g_092351_(_054258_, _054271_, _054272_);
  or g_092352_(_054257_, _054269_, _054273_);
  and g_092353_(_054252_, _054255_, _054274_);
  or g_092354_(_054251_, _054256_, _054275_);
  and g_092355_(_054261_, _054268_, _054276_);
  or g_092356_(_054262_, _054267_, _054277_);
  and g_092357_(_054275_, _054277_, _054278_);
  or g_092358_(_054274_, _054276_, _054279_);
  and g_092359_(_054272_, _054278_, _054280_);
  or g_092360_(_054273_, _054279_, _054282_);
  or g_092361_(_054930_, _054219_, _054283_);
  or g_092362_(_054030_, _054218_, _054284_);
  and g_092363_(_054283_, _054284_, _054285_);
  and g_092364_(out[561], _054285_, _054286_);
  not g_092365_(_054286_, _054287_);
  and g_092366_(_054038_, _054219_, _054288_);
  or g_092367_(_054037_, _054218_, _054289_);
  and g_092368_(_054941_, _054218_, _054290_);
  or g_092369_(out[544], _054219_, _054291_);
  and g_092370_(_054289_, _054291_, _054293_);
  or g_092371_(_054288_, _054290_, _054294_);
  and g_092372_(out[560], _054294_, _054295_);
  or g_092373_(_055073_, _054293_, _054296_);
  xor g_092374_(out[561], _054285_, _054297_);
  xor g_092375_(_055062_, _054285_, _054298_);
  and g_092376_(_054296_, _054297_, _054299_);
  or g_092377_(_054295_, _054298_, _054300_);
  and g_092378_(_054287_, _054300_, _054301_);
  or g_092379_(_054286_, _054299_, _054302_);
  and g_092380_(_054280_, _054302_, _054304_);
  or g_092381_(_054282_, _054301_, _054305_);
  and g_092382_(_054273_, _054275_, _054306_);
  or g_092383_(_054272_, _054274_, _054307_);
  and g_092384_(_054305_, _054307_, _054308_);
  or g_092385_(_054304_, _054306_, _054309_);
  and g_092386_(_054228_, _054234_, _054310_);
  or g_092387_(_054227_, _054233_, _054311_);
  and g_092388_(_054309_, _054311_, _054312_);
  or g_092389_(_054308_, _054310_, _054313_);
  and g_092390_(_054249_, _054313_, _054315_);
  or g_092391_(_054250_, _054312_, _054316_);
  and g_092392_(_022274_, _022417_, _054317_);
  or g_092393_(_022285_, _022406_, _054318_);
  xor g_092394_(out[570], _022384_, _054319_);
  xor g_092395_(_055128_, _022384_, _054320_);
  and g_092396_(_054224_, _054319_, _054321_);
  or g_092397_(_054225_, _054320_, _054322_);
  and g_092398_(_054318_, _054322_, _054323_);
  or g_092399_(_054317_, _054321_, _054324_);
  and g_092400_(_054225_, _054320_, _054326_);
  or g_092401_(_054224_, _054319_, _054327_);
  and g_092402_(_054075_, _054218_, _054328_);
  or g_092403_(_054074_, _054219_, _054329_);
  and g_092404_(_054073_, _054219_, _054330_);
  or g_092405_(_054071_, _054218_, _054331_);
  and g_092406_(_054329_, _054331_, _054332_);
  or g_092407_(_054328_, _054330_, _054333_);
  xor g_092408_(out[569], _022373_, _054334_);
  xor g_092409_(_055117_, _022373_, _054335_);
  and g_092410_(_054332_, _054335_, _054337_);
  or g_092411_(_054333_, _054334_, _054338_);
  and g_092412_(_022285_, _022406_, _054339_);
  or g_092413_(_022274_, _022417_, _054340_);
  and g_092414_(_054333_, _054334_, _054341_);
  or g_092415_(_054332_, _054335_, _054342_);
  xor g_092416_(out[568], _022362_, _054343_);
  xor g_092417_(_055106_, _022362_, _054344_);
  and g_092418_(_054078_, _054218_, _054345_);
  or g_092419_(_054079_, _054219_, _054346_);
  and g_092420_(_054086_, _054219_, _054348_);
  or g_092421_(_054085_, _054218_, _054349_);
  and g_092422_(_054346_, _054349_, _054350_);
  or g_092423_(_054345_, _054348_, _054351_);
  and g_092424_(_054343_, _054350_, _054352_);
  or g_092425_(_054344_, _054351_, _054353_);
  and g_092426_(_054342_, _054353_, _054354_);
  or g_092427_(_054341_, _054352_, _054355_);
  and g_092428_(_054344_, _054351_, _054356_);
  or g_092429_(_054343_, _054350_, _054357_);
  and g_092430_(_054338_, _054354_, _054359_);
  or g_092431_(_054337_, _054355_, _054360_);
  and g_092432_(_054327_, _054340_, _054361_);
  or g_092433_(_054326_, _054339_, _054362_);
  and g_092434_(_054323_, _054361_, _054363_);
  or g_092435_(_054324_, _054362_, _054364_);
  and g_092436_(_054357_, _054363_, _054365_);
  or g_092437_(_054356_, _054364_, _054366_);
  and g_092438_(_054359_, _054365_, _054367_);
  or g_092439_(_054360_, _054366_, _054368_);
  xor g_092440_(out[567], _022351_, _054370_);
  xor g_092441_(_055018_, _022351_, _054371_);
  or g_092442_(_054114_, _054219_, _054372_);
  or g_092443_(_054120_, _054218_, _054373_);
  and g_092444_(_054372_, _054373_, _054374_);
  not g_092445_(_054374_, _054375_);
  and g_092446_(_054371_, _054375_, _054376_);
  or g_092447_(_054370_, _054374_, _054377_);
  xor g_092448_(out[566], _022340_, _054378_);
  not g_092449_(_054378_, _054379_);
  or g_092450_(_054102_, _054219_, _054381_);
  or g_092451_(_054109_, _054218_, _054382_);
  and g_092452_(_054381_, _054382_, _054383_);
  not g_092453_(_054383_, _054384_);
  and g_092454_(_054379_, _054383_, _054385_);
  or g_092455_(_054378_, _054384_, _054386_);
  and g_092456_(_054377_, _054386_, _054387_);
  or g_092457_(_054376_, _054385_, _054388_);
  and g_092458_(_054239_, _054244_, _054389_);
  and g_092459_(_054370_, _054374_, _054390_);
  or g_092460_(_054371_, _054375_, _054392_);
  and g_092461_(_054378_, _054384_, _054393_);
  or g_092462_(_054390_, _054393_, _054394_);
  or g_092463_(_054389_, _054394_, _054395_);
  or g_092464_(_054388_, _054395_, _054396_);
  not g_092465_(_054396_, _054397_);
  and g_092466_(_054367_, _054397_, _054398_);
  or g_092467_(_054368_, _054396_, _054399_);
  and g_092468_(_054316_, _054398_, _054400_);
  or g_092469_(_054315_, _054399_, _054401_);
  and g_092470_(_054338_, _054355_, _054403_);
  or g_092471_(_054337_, _054354_, _054404_);
  and g_092472_(_054363_, _054403_, _054405_);
  or g_092473_(_054364_, _054404_, _054406_);
  and g_092474_(_054324_, _054340_, _054407_);
  or g_092475_(_054323_, _054339_, _054408_);
  and g_092476_(_054406_, _054408_, _054409_);
  or g_092477_(_054405_, _054407_, _054410_);
  and g_092478_(_054388_, _054392_, _054411_);
  or g_092479_(_054387_, _054390_, _054412_);
  and g_092480_(_054367_, _054411_, _054414_);
  or g_092481_(_054368_, _054412_, _054415_);
  and g_092482_(_054409_, _054415_, _054416_);
  or g_092483_(_054410_, _054414_, _054417_);
  and g_092484_(_054401_, _054416_, _054418_);
  or g_092485_(_054400_, _054417_, _054419_);
  and g_092486_(_055073_, _054293_, _054420_);
  or g_092487_(out[560], _054294_, _054421_);
  and g_092488_(_054311_, _054421_, _054422_);
  or g_092489_(_054310_, _054420_, _054423_);
  and g_092490_(_054249_, _054422_, _054425_);
  or g_092491_(_054250_, _054423_, _054426_);
  and g_092492_(_054280_, _054425_, _054427_);
  or g_092493_(_054282_, _054426_, _054428_);
  and g_092494_(_054299_, _054427_, _054429_);
  or g_092495_(_054300_, _054428_, _054430_);
  and g_092496_(_054398_, _054429_, _054431_);
  or g_092497_(_054399_, _054430_, _054432_);
  and g_092498_(_054419_, _054432_, _054433_);
  or g_092499_(_054418_, _054431_, _054434_);
  and g_092500_(_054225_, _054434_, _054436_);
  or g_092501_(_054224_, _054433_, _054437_);
  and g_092502_(_054319_, _054433_, _054438_);
  or g_092503_(_054320_, _054434_, _054439_);
  and g_092504_(_054437_, _054439_, _054440_);
  or g_092505_(_054436_, _054438_, _054441_);
  xor g_092506_(out[586], _022538_, _054442_);
  not g_092507_(_054442_, _054443_);
  and g_092508_(_054440_, _054442_, _054444_);
  or g_092509_(_054441_, _054443_, _054445_);
  and g_092510_(_022428_, _022571_, _054447_);
  or g_092511_(_022439_, _022560_, _054448_);
  and g_092512_(_054445_, _054448_, _054449_);
  or g_092513_(_054444_, _054447_, _054450_);
  and g_092514_(_054335_, _054433_, _054451_);
  or g_092515_(_054334_, _054434_, _054452_);
  and g_092516_(_054333_, _054434_, _054453_);
  or g_092517_(_054332_, _054433_, _054454_);
  and g_092518_(_054452_, _054454_, _054455_);
  or g_092519_(_054451_, _054453_, _054456_);
  xor g_092520_(out[585], _022527_, _054458_);
  not g_092521_(_054458_, _054459_);
  and g_092522_(_054455_, _054459_, _054460_);
  or g_092523_(_054456_, _054458_, _054461_);
  and g_092524_(_054441_, _054443_, _054462_);
  or g_092525_(_054440_, _054442_, _054463_);
  and g_092526_(_022439_, _022560_, _054464_);
  or g_092527_(_022428_, _022571_, _054465_);
  and g_092528_(_054463_, _054465_, _054466_);
  or g_092529_(_054462_, _054464_, _054467_);
  and g_092530_(_054461_, _054466_, _054469_);
  or g_092531_(_054460_, _054467_, _054470_);
  and g_092532_(_054449_, _054469_, _054471_);
  or g_092533_(_054450_, _054470_, _054472_);
  xor g_092534_(out[584], _022516_, _054473_);
  xor g_092535_(_055238_, _022516_, _054474_);
  and g_092536_(_054343_, _054433_, _054475_);
  or g_092537_(_054344_, _054434_, _054476_);
  and g_092538_(_054351_, _054434_, _054477_);
  or g_092539_(_054350_, _054433_, _054478_);
  and g_092540_(_054476_, _054478_, _054480_);
  or g_092541_(_054475_, _054477_, _054481_);
  and g_092542_(_054474_, _054481_, _054482_);
  not g_092543_(_054482_, _054483_);
  and g_092544_(_054456_, _054458_, _054484_);
  or g_092545_(_054455_, _054459_, _054485_);
  and g_092546_(_054473_, _054480_, _054486_);
  or g_092547_(_054474_, _054481_, _054487_);
  and g_092548_(_054485_, _054487_, _054488_);
  or g_092549_(_054484_, _054486_, _054489_);
  and g_092550_(_054483_, _054488_, _054491_);
  or g_092551_(_054482_, _054489_, _054492_);
  and g_092552_(_054471_, _054491_, _054493_);
  or g_092553_(_054472_, _054492_, _054494_);
  xor g_092554_(out[582], _022494_, _054495_);
  not g_092555_(_054495_, _054496_);
  or g_092556_(_054378_, _054434_, _054497_);
  or g_092557_(_054383_, _054433_, _054498_);
  and g_092558_(_054497_, _054498_, _054499_);
  not g_092559_(_054499_, _054500_);
  and g_092560_(_054496_, _054499_, _054502_);
  or g_092561_(_054495_, _054500_, _054503_);
  xor g_092562_(out[583], _022505_, _054504_);
  xor g_092563_(_055150_, _022505_, _054505_);
  or g_092564_(_054371_, _054434_, _054506_);
  or g_092565_(_054374_, _054433_, _054507_);
  and g_092566_(_054506_, _054507_, _054508_);
  not g_092567_(_054508_, _054509_);
  and g_092568_(_054505_, _054509_, _054510_);
  or g_092569_(_054504_, _054508_, _054511_);
  and g_092570_(_054503_, _054511_, _054513_);
  or g_092571_(_054502_, _054510_, _054514_);
  and g_092572_(_054504_, _054508_, _054515_);
  or g_092573_(_054505_, _054509_, _054516_);
  and g_092574_(_054495_, _054500_, _054517_);
  or g_092575_(_054496_, _054499_, _054518_);
  and g_092576_(_054516_, _054518_, _054519_);
  or g_092577_(_054515_, _054517_, _054520_);
  and g_092578_(_054513_, _054519_, _054521_);
  or g_092579_(_054514_, _054520_, _054522_);
  xor g_092580_(out[581], _022483_, _054524_);
  not g_092581_(_054524_, _054525_);
  and g_092582_(_054239_, _054433_, _054526_);
  or g_092583_(_054238_, _054434_, _054527_);
  and g_092584_(_054245_, _054434_, _054528_);
  or g_092585_(_054244_, _054433_, _054529_);
  and g_092586_(_054527_, _054529_, _054530_);
  or g_092587_(_054526_, _054528_, _054531_);
  and g_092588_(_054524_, _054531_, _054532_);
  or g_092589_(_054525_, _054530_, _054533_);
  xor g_092590_(out[580], _022472_, _054535_);
  xor g_092591_(_055183_, _022472_, _054536_);
  and g_092592_(_054227_, _054433_, _054537_);
  or g_092593_(_054228_, _054434_, _054538_);
  and g_092594_(_054234_, _054434_, _054539_);
  or g_092595_(_054233_, _054433_, _054540_);
  and g_092596_(_054538_, _054540_, _054541_);
  or g_092597_(_054537_, _054539_, _054542_);
  and g_092598_(_054535_, _054541_, _054543_);
  or g_092599_(_054536_, _054542_, _054544_);
  and g_092600_(_054533_, _054544_, _054546_);
  or g_092601_(_054532_, _054543_, _054547_);
  and g_092602_(_054525_, _054530_, _054548_);
  or g_092603_(_054524_, _054531_, _054549_);
  and g_092604_(_054536_, _054542_, _054550_);
  not g_092605_(_054550_, _054551_);
  and g_092606_(_054549_, _054551_, _054552_);
  or g_092607_(_054548_, _054550_, _054553_);
  and g_092608_(_054546_, _054552_, _054554_);
  or g_092609_(_054547_, _054553_, _054555_);
  and g_092610_(_054521_, _054554_, _054557_);
  or g_092611_(_054522_, _054555_, _054558_);
  and g_092612_(_054493_, _054557_, _054559_);
  or g_092613_(_054494_, _054558_, _054560_);
  xor g_092614_(out[579], _022450_, _054561_);
  not g_092615_(_054561_, _054562_);
  or g_092616_(_054255_, _054433_, _054563_);
  or g_092617_(_054251_, _054434_, _054564_);
  and g_092618_(_054563_, _054564_, _054565_);
  not g_092619_(_054565_, _054566_);
  and g_092620_(_054562_, _054565_, _054568_);
  or g_092621_(_054561_, _054566_, _054569_);
  or g_092622_(out[577], out[578], _054570_);
  xor g_092623_(out[577], out[578], _054571_);
  xor g_092624_(_055194_, out[578], _054572_);
  and g_092625_(_054268_, _054434_, _054573_);
  and g_092626_(_054262_, _054433_, _054574_);
  or g_092627_(_054573_, _054574_, _054575_);
  or g_092628_(_054571_, _054575_, _054576_);
  not g_092629_(_054576_, _054577_);
  and g_092630_(_054561_, _054566_, _054579_);
  or g_092631_(_054562_, _054565_, _054580_);
  and g_092632_(_054576_, _054580_, _054581_);
  or g_092633_(_054577_, _054579_, _054582_);
  or g_092634_(_055062_, _054434_, _054583_);
  or g_092635_(_054285_, _054433_, _054584_);
  and g_092636_(_054583_, _054584_, _054585_);
  and g_092637_(out[577], _054585_, _054586_);
  not g_092638_(_054586_, _054587_);
  and g_092639_(_054294_, _054434_, _054588_);
  or g_092640_(_054293_, _054433_, _054590_);
  and g_092641_(_055073_, _054433_, _054591_);
  or g_092642_(out[560], _054434_, _054592_);
  and g_092643_(_054590_, _054592_, _054593_);
  or g_092644_(_054588_, _054591_, _054594_);
  and g_092645_(out[576], _054594_, _054595_);
  or g_092646_(_055205_, _054593_, _054596_);
  xor g_092647_(out[577], _054585_, _054597_);
  xor g_092648_(_055194_, _054585_, _054598_);
  and g_092649_(_054596_, _054597_, _054599_);
  or g_092650_(_054595_, _054598_, _054601_);
  and g_092651_(_054587_, _054601_, _054602_);
  or g_092652_(_054586_, _054599_, _054603_);
  xor g_092653_(_054572_, _054575_, _054604_);
  or g_092654_(_054602_, _054604_, _054605_);
  and g_092655_(_054581_, _054605_, _054606_);
  or g_092656_(_054568_, _054579_, _054607_);
  or g_092657_(_054604_, _054607_, _054608_);
  not g_092658_(_054608_, _054609_);
  and g_092659_(_054603_, _054609_, _054610_);
  and g_092660_(_054569_, _054582_, _054612_);
  or g_092661_(_054610_, _054612_, _054613_);
  or g_092662_(_054568_, _054606_, _054614_);
  and g_092663_(_054559_, _054613_, _054615_);
  or g_092664_(_054560_, _054614_, _054616_);
  and g_092665_(_054514_, _054516_, _054617_);
  or g_092666_(_054513_, _054515_, _054618_);
  and g_092667_(_054547_, _054549_, _054619_);
  or g_092668_(_054546_, _054548_, _054620_);
  and g_092669_(_054521_, _054619_, _054621_);
  or g_092670_(_054522_, _054620_, _054623_);
  and g_092671_(_054618_, _054623_, _054624_);
  or g_092672_(_054617_, _054621_, _054625_);
  and g_092673_(_054493_, _054625_, _054626_);
  or g_092674_(_054494_, _054624_, _054627_);
  or g_092675_(_054472_, _054488_, _054628_);
  not g_092676_(_054628_, _054629_);
  and g_092677_(_054450_, _054465_, _054630_);
  or g_092678_(_054449_, _054464_, _054631_);
  and g_092679_(_054628_, _054631_, _054632_);
  or g_092680_(_054629_, _054630_, _054634_);
  and g_092681_(_054627_, _054632_, _054635_);
  or g_092682_(_054626_, _054634_, _054636_);
  and g_092683_(_054616_, _054635_, _054637_);
  or g_092684_(_054615_, _054636_, _054638_);
  and g_092685_(_055205_, _054593_, _054639_);
  or g_092686_(out[576], _054594_, _054640_);
  and g_092687_(_054599_, _054640_, _054641_);
  or g_092688_(_054601_, _054639_, _054642_);
  and g_092689_(_054559_, _054641_, _054643_);
  or g_092690_(_054560_, _054642_, _054645_);
  and g_092691_(_054609_, _054643_, _054646_);
  or g_092692_(_054608_, _054645_, _054647_);
  and g_092693_(_054638_, _054647_, _054648_);
  or g_092694_(_054637_, _054646_, _054649_);
  and g_092695_(_054441_, _054649_, _054650_);
  or g_092696_(_054440_, _054648_, _054651_);
  and g_092697_(_054442_, _054648_, _054652_);
  or g_092698_(_054443_, _054649_, _054653_);
  and g_092699_(_054651_, _054653_, _054654_);
  or g_092700_(_054650_, _054652_, _054656_);
  and g_092701_(_022582_, _022725_, _054657_);
  or g_092702_(_022593_, _022714_, _054658_);
  xor g_092703_(out[602], _022692_, _054659_);
  xor g_092704_(_055392_, _022692_, _054660_);
  and g_092705_(_054654_, _054659_, _054661_);
  or g_092706_(_054656_, _054660_, _054662_);
  and g_092707_(_054658_, _054662_, _054663_);
  or g_092708_(_054657_, _054661_, _054664_);
  and g_092709_(_022593_, _022714_, _054665_);
  or g_092710_(_022582_, _022725_, _054667_);
  and g_092711_(_054656_, _054660_, _054668_);
  or g_092712_(_054654_, _054659_, _054669_);
  and g_092713_(_054667_, _054669_, _054670_);
  or g_092714_(_054665_, _054668_, _054671_);
  or g_092715_(_054458_, _054649_, _054672_);
  not g_092716_(_054672_, _054673_);
  and g_092717_(_054456_, _054649_, _054674_);
  not g_092718_(_054674_, _054675_);
  and g_092719_(_054672_, _054675_, _054676_);
  or g_092720_(_054673_, _054674_, _054678_);
  xor g_092721_(out[601], _022681_, _054679_);
  xor g_092722_(_055381_, _022681_, _054680_);
  and g_092723_(_054676_, _054680_, _054681_);
  or g_092724_(_054678_, _054679_, _054682_);
  and g_092725_(_054670_, _054682_, _054683_);
  or g_092726_(_054671_, _054681_, _054684_);
  and g_092727_(_054663_, _054683_, _054685_);
  or g_092728_(_054664_, _054684_, _054686_);
  xor g_092729_(out[600], _022670_, _054687_);
  xor g_092730_(_055370_, _022670_, _054689_);
  or g_092731_(_054474_, _054649_, _054690_);
  not g_092732_(_054690_, _054691_);
  and g_092733_(_054481_, _054649_, _054692_);
  not g_092734_(_054692_, _054693_);
  and g_092735_(_054690_, _054693_, _054694_);
  or g_092736_(_054691_, _054692_, _054695_);
  and g_092737_(_054687_, _054694_, _054696_);
  or g_092738_(_054689_, _054695_, _054697_);
  and g_092739_(_054678_, _054679_, _054698_);
  or g_092740_(_054676_, _054680_, _054700_);
  and g_092741_(_054697_, _054700_, _054701_);
  or g_092742_(_054696_, _054698_, _054702_);
  and g_092743_(_054689_, _054695_, _054703_);
  or g_092744_(_054687_, _054694_, _054704_);
  and g_092745_(_054701_, _054704_, _054705_);
  or g_092746_(_054702_, _054703_, _054706_);
  and g_092747_(_054685_, _054705_, _054707_);
  or g_092748_(_054686_, _054706_, _054708_);
  xor g_092749_(out[598], _022648_, _054709_);
  not g_092750_(_054709_, _054711_);
  or g_092751_(_054495_, _054649_, _054712_);
  or g_092752_(_054499_, _054648_, _054713_);
  and g_092753_(_054712_, _054713_, _054714_);
  not g_092754_(_054714_, _054715_);
  or g_092755_(_054709_, _054715_, _054716_);
  xor g_092756_(_054711_, _054714_, _054717_);
  xor g_092757_(_054709_, _054714_, _054718_);
  xor g_092758_(out[599], _022659_, _054719_);
  not g_092759_(_054719_, _054720_);
  or g_092760_(_054505_, _054649_, _054722_);
  or g_092761_(_054508_, _054648_, _054723_);
  and g_092762_(_054722_, _054723_, _054724_);
  not g_092763_(_054724_, _054725_);
  and g_092764_(_054719_, _054724_, _054726_);
  xor g_092765_(out[597], _022637_, _054727_);
  xor g_092766_(_055304_, _022637_, _054728_);
  or g_092767_(_054524_, _054649_, _054729_);
  not g_092768_(_054729_, _054730_);
  and g_092769_(_054531_, _054649_, _054731_);
  not g_092770_(_054731_, _054733_);
  and g_092771_(_054729_, _054733_, _054734_);
  or g_092772_(_054730_, _054731_, _054735_);
  and g_092773_(_054728_, _054734_, _054736_);
  or g_092774_(_054727_, _054735_, _054737_);
  or g_092775_(_054719_, _054724_, _054738_);
  xor g_092776_(_054719_, _054724_, _054739_);
  xor g_092777_(_054720_, _054724_, _054740_);
  and g_092778_(_054717_, _054739_, _054741_);
  or g_092779_(_054718_, _054740_, _054742_);
  and g_092780_(_054737_, _054741_, _054744_);
  or g_092781_(_054736_, _054742_, _054745_);
  and g_092782_(_054727_, _054735_, _054746_);
  or g_092783_(_054728_, _054734_, _054747_);
  xor g_092784_(out[596], _022626_, _054748_);
  xor g_092785_(_055315_, _022626_, _054749_);
  or g_092786_(_054536_, _054649_, _054750_);
  not g_092787_(_054750_, _054751_);
  and g_092788_(_054542_, _054649_, _054752_);
  not g_092789_(_054752_, _054753_);
  and g_092790_(_054750_, _054753_, _054755_);
  or g_092791_(_054751_, _054752_, _054756_);
  and g_092792_(_054748_, _054755_, _054757_);
  or g_092793_(_054749_, _054756_, _054758_);
  and g_092794_(_054747_, _054758_, _054759_);
  or g_092795_(_054746_, _054757_, _054760_);
  and g_092796_(_054744_, _054760_, _054761_);
  or g_092797_(_054745_, _054759_, _054762_);
  and g_092798_(_054716_, _054738_, _054763_);
  or g_092799_(_054726_, _054763_, _054764_);
  not g_092800_(_054764_, _054766_);
  and g_092801_(_054762_, _054764_, _054767_);
  or g_092802_(_054761_, _054766_, _054768_);
  and g_092803_(_054707_, _054768_, _054769_);
  or g_092804_(_054708_, _054767_, _054770_);
  and g_092805_(_054749_, _054756_, _054771_);
  or g_092806_(_054748_, _054755_, _054772_);
  and g_092807_(_054759_, _054772_, _054773_);
  or g_092808_(_054760_, _054771_, _054774_);
  and g_092809_(_054744_, _054773_, _054775_);
  or g_092810_(_054745_, _054774_, _054777_);
  and g_092811_(_054707_, _054775_, _054778_);
  or g_092812_(_054708_, _054777_, _054779_);
  xor g_092813_(out[595], _022604_, _054780_);
  xor g_092814_(_055359_, _022604_, _054781_);
  or g_092815_(_054565_, _054648_, _054782_);
  or g_092816_(_054561_, _054649_, _054783_);
  and g_092817_(_054782_, _054783_, _054784_);
  not g_092818_(_054784_, _054785_);
  or g_092819_(_054781_, _054784_, _054786_);
  and g_092820_(_054781_, _054784_, _054788_);
  xor g_092821_(_054781_, _054784_, _054789_);
  xor g_092822_(_054780_, _054784_, _054790_);
  or g_092823_(out[593], out[594], _054791_);
  xor g_092824_(out[593], out[594], _054792_);
  xor g_092825_(_055326_, out[594], _054793_);
  and g_092826_(_054575_, _054649_, _054794_);
  and g_092827_(_054572_, _054648_, _054795_);
  or g_092828_(_054794_, _054795_, _054796_);
  or g_092829_(_054792_, _054796_, _054797_);
  xor g_092830_(_054792_, _054796_, _054799_);
  xor g_092831_(_054793_, _054796_, _054800_);
  and g_092832_(_054789_, _054799_, _054801_);
  or g_092833_(_054790_, _054800_, _054802_);
  or g_092834_(_055194_, _054649_, _054803_);
  or g_092835_(_054585_, _054648_, _054804_);
  and g_092836_(_054803_, _054804_, _054805_);
  and g_092837_(out[593], _054805_, _054806_);
  and g_092838_(_054801_, _054806_, _054807_);
  not g_092839_(_054807_, _054808_);
  and g_092840_(_054786_, _054797_, _054810_);
  or g_092841_(_054788_, _054810_, _054811_);
  not g_092842_(_054811_, _054812_);
  and g_092843_(_054594_, _054649_, _054813_);
  not g_092844_(_054813_, _054814_);
  or g_092845_(out[576], _054649_, _054815_);
  not g_092846_(_054815_, _054816_);
  and g_092847_(_054814_, _054815_, _054817_);
  or g_092848_(_054813_, _054816_, _054818_);
  and g_092849_(out[592], _054818_, _054819_);
  or g_092850_(_055337_, _054817_, _054821_);
  xor g_092851_(out[593], _054805_, _054822_);
  xor g_092852_(_055326_, _054805_, _054823_);
  and g_092853_(_054821_, _054822_, _054824_);
  or g_092854_(_054819_, _054823_, _054825_);
  and g_092855_(_054801_, _054824_, _054826_);
  or g_092856_(_054802_, _054825_, _054827_);
  and g_092857_(_054808_, _054811_, _054828_);
  or g_092858_(_054807_, _054812_, _054829_);
  and g_092859_(_054827_, _054828_, _054830_);
  or g_092860_(_054826_, _054829_, _054832_);
  and g_092861_(_054778_, _054832_, _054833_);
  or g_092862_(_054779_, _054830_, _054834_);
  and g_092863_(_054664_, _054667_, _054835_);
  or g_092864_(_054663_, _054665_, _054836_);
  and g_092865_(_054685_, _054702_, _054837_);
  or g_092866_(_054686_, _054701_, _054838_);
  and g_092867_(_054770_, _054838_, _054839_);
  or g_092868_(_054769_, _054837_, _054840_);
  and g_092869_(_054834_, _054839_, _054841_);
  or g_092870_(_054833_, _054840_, _054843_);
  and g_092871_(_054836_, _054841_, _054844_);
  or g_092872_(_054835_, _054843_, _054845_);
  or g_092873_(out[592], _054818_, _054846_);
  and g_092874_(_054826_, _054846_, _054847_);
  and g_092875_(_054778_, _054847_, _054848_);
  not g_092876_(_054848_, _054849_);
  and g_092877_(_054845_, _054849_, _054850_);
  or g_092878_(_054844_, _054848_, _054851_);
  and g_092879_(_054656_, _054851_, _054852_);
  or g_092880_(_054654_, _054850_, _054854_);
  and g_092881_(_054659_, _054850_, _054855_);
  or g_092882_(_054660_, _054851_, _054856_);
  and g_092883_(_054854_, _054856_, _054857_);
  or g_092884_(_054852_, _054855_, _054858_);
  and g_092885_(_053998_, _054858_, _054859_);
  or g_092886_(_053997_, _054857_, _054860_);
  and g_092887_(_053997_, _054857_, _054861_);
  or g_092888_(_053998_, _054858_, _054862_);
  and g_092889_(_054680_, _054850_, _054863_);
  or g_092890_(_054679_, _054851_, _054865_);
  and g_092891_(_054678_, _054851_, _054866_);
  or g_092892_(_054676_, _054850_, _054867_);
  and g_092893_(_054865_, _054867_, _054868_);
  or g_092894_(_054863_, _054866_, _054869_);
  xor g_092895_(out[617], _022835_, _054870_);
  xor g_092896_(_055513_, _022835_, _054871_);
  and g_092897_(_054868_, _054871_, _054872_);
  or g_092898_(_054869_, _054870_, _054873_);
  and g_092899_(_022736_, _022879_, _054874_);
  or g_092900_(_022747_, _022868_, _054876_);
  and g_092901_(_022747_, _022868_, _054877_);
  or g_092902_(_022736_, _022879_, _054878_);
  and g_092903_(_054869_, _054870_, _054879_);
  or g_092904_(_054868_, _054871_, _054880_);
  xor g_092905_(out[616], _022824_, _054881_);
  xor g_092906_(_055502_, _022824_, _054882_);
  and g_092907_(_054687_, _054850_, _054883_);
  or g_092908_(_054689_, _054851_, _054884_);
  and g_092909_(_054695_, _054851_, _054885_);
  or g_092910_(_054694_, _054850_, _054887_);
  and g_092911_(_054884_, _054887_, _054888_);
  or g_092912_(_054883_, _054885_, _054889_);
  and g_092913_(_054881_, _054888_, _054890_);
  or g_092914_(_054882_, _054889_, _054891_);
  and g_092915_(_054880_, _054891_, _054892_);
  or g_092916_(_054879_, _054890_, _054893_);
  and g_092917_(_054882_, _054889_, _054894_);
  or g_092918_(_054881_, _054888_, _054895_);
  and g_092919_(_054873_, _054892_, _054896_);
  or g_092920_(_054872_, _054893_, _054898_);
  and g_092921_(_054860_, _054876_, _054899_);
  or g_092922_(_054859_, _054874_, _054900_);
  and g_092923_(_054862_, _054878_, _054901_);
  or g_092924_(_054861_, _054877_, _054902_);
  and g_092925_(_054899_, _054901_, _054903_);
  or g_092926_(_054900_, _054902_, _054904_);
  and g_092927_(_054895_, _054903_, _054905_);
  or g_092928_(_054894_, _054904_, _054906_);
  and g_092929_(_054896_, _054905_, _054907_);
  or g_092930_(_054898_, _054906_, _054909_);
  xor g_092931_(out[614], _022802_, _054910_);
  xor g_092932_(_055425_, _022802_, _054911_);
  and g_092933_(_054711_, _054850_, _054912_);
  or g_092934_(_054709_, _054851_, _054913_);
  and g_092935_(_054715_, _054851_, _054914_);
  or g_092936_(_054714_, _054850_, _054915_);
  and g_092937_(_054913_, _054915_, _054916_);
  or g_092938_(_054912_, _054914_, _054917_);
  and g_092939_(_054911_, _054916_, _054918_);
  or g_092940_(_054910_, _054917_, _054920_);
  xor g_092941_(out[615], _022813_, _054921_);
  xor g_092942_(_055414_, _022813_, _054922_);
  and g_092943_(_054719_, _054850_, _054923_);
  or g_092944_(_054720_, _054851_, _054924_);
  and g_092945_(_054725_, _054851_, _054925_);
  or g_092946_(_054724_, _054850_, _054926_);
  and g_092947_(_054924_, _054926_, _054927_);
  or g_092948_(_054923_, _054925_, _054928_);
  and g_092949_(_054922_, _054928_, _054929_);
  or g_092950_(_054921_, _054927_, _054931_);
  and g_092951_(_054920_, _054931_, _054932_);
  or g_092952_(_054918_, _054929_, _054933_);
  and g_092953_(_054921_, _054927_, _054934_);
  or g_092954_(_054922_, _054928_, _054935_);
  and g_092955_(_054910_, _054917_, _054936_);
  or g_092956_(_054911_, _054916_, _054937_);
  and g_092957_(_054935_, _054937_, _054938_);
  or g_092958_(_054934_, _054936_, _054939_);
  and g_092959_(_054932_, _054938_, _054940_);
  or g_092960_(_054933_, _054939_, _054942_);
  xor g_092961_(out[613], _022791_, _054943_);
  and g_092962_(_054728_, _054850_, _054944_);
  or g_092963_(_054727_, _054851_, _054945_);
  and g_092964_(_054735_, _054851_, _054946_);
  or g_092965_(_054734_, _054850_, _054947_);
  and g_092966_(_054945_, _054947_, _054948_);
  or g_092967_(_054944_, _054946_, _054949_);
  and g_092968_(_054943_, _054949_, _054950_);
  xor g_092969_(out[612], _022780_, _054951_);
  xor g_092970_(_055447_, _022780_, _054953_);
  or g_092971_(_054749_, _054851_, _054954_);
  or g_092972_(_054755_, _054850_, _054955_);
  and g_092973_(_054954_, _054955_, _054956_);
  or g_092974_(_054943_, _054949_, _054957_);
  and g_092975_(_054951_, _054956_, _054958_);
  xor g_092976_(_054943_, _054949_, _054959_);
  xor g_092977_(_054943_, _054948_, _054960_);
  xor g_092978_(_054951_, _054956_, _054961_);
  xor g_092979_(_054953_, _054956_, _054962_);
  and g_092980_(_054940_, _054961_, _054964_);
  or g_092981_(_054942_, _054962_, _054965_);
  and g_092982_(_054959_, _054964_, _054966_);
  or g_092983_(_054960_, _054965_, _054967_);
  and g_092984_(_054785_, _054851_, _054968_);
  or g_092985_(_054784_, _054850_, _054969_);
  and g_092986_(_054781_, _054850_, _054970_);
  or g_092987_(_054780_, _054851_, _054971_);
  and g_092988_(_054969_, _054971_, _054972_);
  or g_092989_(_054968_, _054970_, _054973_);
  and g_092990_(_053994_, _054973_, _054975_);
  or g_092991_(_053996_, _054972_, _054976_);
  or g_092992_(out[609], out[610], _054977_);
  xor g_092993_(out[609], out[610], _054978_);
  xor g_092994_(_055458_, out[610], _054979_);
  and g_092995_(_054796_, _054851_, _054980_);
  not g_092996_(_054980_, _054981_);
  and g_092997_(_054793_, _054850_, _054982_);
  or g_092998_(_054792_, _054851_, _054983_);
  and g_092999_(_054981_, _054983_, _054984_);
  or g_093000_(_054980_, _054982_, _054986_);
  and g_093001_(_054979_, _054984_, _054987_);
  or g_093002_(_054978_, _054986_, _054988_);
  and g_093003_(_053996_, _054972_, _054989_);
  or g_093004_(_053994_, _054973_, _054990_);
  and g_093005_(_054976_, _054990_, _054991_);
  or g_093006_(_054975_, _054989_, _054992_);
  xor g_093007_(_054979_, _054984_, _054993_);
  xor g_093008_(_054978_, _054984_, _054994_);
  and g_093009_(_054991_, _054993_, _054995_);
  or g_093010_(_054992_, _054994_, _054997_);
  or g_093011_(_055326_, _054851_, _054998_);
  or g_093012_(_054805_, _054850_, _054999_);
  and g_093013_(_054998_, _054999_, _055000_);
  and g_093014_(out[609], _055000_, _055001_);
  not g_093015_(_055001_, _055002_);
  and g_093016_(_054818_, _054851_, _055003_);
  or g_093017_(_054817_, _054850_, _055004_);
  and g_093018_(_055337_, _054850_, _055005_);
  or g_093019_(out[592], _054851_, _055006_);
  and g_093020_(_055004_, _055006_, _055008_);
  or g_093021_(_055003_, _055005_, _055009_);
  and g_093022_(out[608], _055009_, _055010_);
  or g_093023_(_055469_, _055008_, _055011_);
  xor g_093024_(out[609], _055000_, _055012_);
  xor g_093025_(_055458_, _055000_, _055013_);
  and g_093026_(_055011_, _055012_, _055014_);
  or g_093027_(_055010_, _055013_, _055015_);
  and g_093028_(_055002_, _055015_, _055016_);
  or g_093029_(_055001_, _055014_, _055017_);
  and g_093030_(_054995_, _055017_, _055019_);
  or g_093031_(_054997_, _055016_, _055020_);
  and g_093032_(_054987_, _054990_, _055021_);
  or g_093033_(_054988_, _054989_, _055022_);
  and g_093034_(_054976_, _055022_, _055023_);
  or g_093035_(_054975_, _055021_, _055024_);
  and g_093036_(_055020_, _055023_, _055025_);
  or g_093037_(_055019_, _055024_, _055026_);
  and g_093038_(_054966_, _055026_, _055027_);
  or g_093039_(_054967_, _055025_, _055028_);
  or g_093040_(_054950_, _054958_, _055030_);
  and g_093041_(_054957_, _055030_, _055031_);
  and g_093042_(_054940_, _055031_, _055032_);
  not g_093043_(_055032_, _055033_);
  and g_093044_(_054933_, _054935_, _055034_);
  or g_093045_(_054932_, _054934_, _055035_);
  and g_093046_(_055033_, _055035_, _055036_);
  or g_093047_(_055032_, _055034_, _055037_);
  and g_093048_(_055028_, _055036_, _055038_);
  or g_093049_(_055027_, _055037_, _055039_);
  and g_093050_(_054907_, _055039_, _055041_);
  or g_093051_(_054909_, _055038_, _055042_);
  and g_093052_(_054873_, _054893_, _055043_);
  or g_093053_(_054872_, _054892_, _055044_);
  and g_093054_(_054903_, _055043_, _055045_);
  or g_093055_(_054904_, _055044_, _055046_);
  and g_093056_(_054861_, _054878_, _055047_);
  or g_093057_(_054862_, _054877_, _055048_);
  and g_093058_(_054876_, _055048_, _055049_);
  or g_093059_(_054874_, _055047_, _055050_);
  and g_093060_(_055046_, _055049_, _055052_);
  or g_093061_(_055045_, _055050_, _055053_);
  and g_093062_(_055042_, _055052_, _055054_);
  or g_093063_(_055041_, _055053_, _055055_);
  and g_093064_(_055469_, _055008_, _055056_);
  or g_093065_(out[608], _055009_, _055057_);
  and g_093066_(_055014_, _055057_, _055058_);
  or g_093067_(_055015_, _055056_, _055059_);
  and g_093068_(_054995_, _055058_, _055060_);
  or g_093069_(_054997_, _055059_, _055061_);
  and g_093070_(_054907_, _055060_, _055063_);
  or g_093071_(_054909_, _055061_, _055064_);
  and g_093072_(_054966_, _055063_, _055065_);
  or g_093073_(_054967_, _055064_, _055066_);
  and g_093074_(_055055_, _055066_, _055067_);
  or g_093075_(_055054_, _055065_, _055068_);
  or g_093076_(_053994_, _055068_, _055069_);
  or g_093077_(_054972_, _055067_, _055070_);
  and g_093078_(_055069_, _055070_, _055071_);
  xor g_093079_(out[628], _022934_, _055072_);
  and g_093080_(_054953_, _055067_, _055074_);
  and g_093081_(_054956_, _055068_, _055075_);
  or g_093082_(_055074_, _055075_, _055076_);
  and g_093083_(_055072_, _055076_, _055077_);
  not g_093084_(_055077_, _055078_);
  xor g_093085_(_055568_, _022945_, _055079_);
  or g_093086_(_054948_, _055067_, _055080_);
  or g_093087_(_054943_, _055068_, _055081_);
  and g_093088_(_055080_, _055081_, _055082_);
  or g_093089_(_055079_, _055082_, _055083_);
  not g_093090_(_055083_, _055085_);
  and g_093091_(_055078_, _055083_, _055086_);
  or g_093092_(_055077_, _055085_, _055087_);
  xor g_093093_(_055623_, _022912_, _055088_);
  or g_093094_(_055071_, _055088_, _055089_);
  or g_093095_(out[625], out[626], _055090_);
  xor g_093096_(out[625], out[626], _055091_);
  xor g_093097_(_055590_, out[626], _055092_);
  and g_093098_(_054986_, _055068_, _055093_);
  and g_093099_(_054979_, _055067_, _055094_);
  or g_093100_(_055093_, _055094_, _055096_);
  not g_093101_(_055096_, _055097_);
  or g_093102_(_055091_, _055096_, _055098_);
  and g_093103_(_055089_, _055098_, _055099_);
  and g_093104_(_055071_, _055088_, _055100_);
  xor g_093105_(_055071_, _055088_, _055101_);
  xor g_093106_(_055091_, _055096_, _055102_);
  and g_093107_(_055101_, _055102_, _055103_);
  or g_093108_(_055458_, _055068_, _055104_);
  or g_093109_(_055000_, _055067_, _055105_);
  and g_093110_(_055104_, _055105_, _055107_);
  and g_093111_(out[625], _055107_, _055108_);
  or g_093112_(_055008_, _055067_, _055109_);
  or g_093113_(out[608], _055068_, _055110_);
  and g_093114_(_055109_, _055110_, _055111_);
  not g_093115_(_055111_, _055112_);
  or g_093116_(_055601_, _055111_, _055113_);
  xor g_093117_(out[625], _055107_, _055114_);
  and g_093118_(_055113_, _055114_, _055115_);
  or g_093119_(_055108_, _055115_, _055116_);
  and g_093120_(_055103_, _055116_, _055118_);
  or g_093121_(_055099_, _055100_, _055119_);
  not g_093122_(_055119_, _055120_);
  or g_093123_(_055118_, _055120_, _055121_);
  or g_093124_(_055072_, _055076_, _055122_);
  and g_093125_(_055121_, _055122_, _055123_);
  or g_093126_(_055087_, _055123_, _055124_);
  and g_093127_(_022890_, _023033_, _055125_);
  or g_093128_(_022901_, _023022_, _055126_);
  and g_093129_(_053997_, _055067_, _055127_);
  not g_093130_(_055127_, _055129_);
  and g_093131_(_054858_, _055068_, _055130_);
  or g_093132_(_054857_, _055067_, _055131_);
  and g_093133_(_055129_, _055131_, _055132_);
  or g_093134_(_055127_, _055130_, _055133_);
  xor g_093135_(out[634], _023000_, _055134_);
  not g_093136_(_055134_, _055135_);
  and g_093137_(_055132_, _055134_, _055136_);
  or g_093138_(_055133_, _055135_, _055137_);
  and g_093139_(_055126_, _055137_, _055138_);
  or g_093140_(_055125_, _055136_, _055140_);
  or g_093141_(_055132_, _055134_, _055141_);
  or g_093142_(_054868_, _055067_, _055142_);
  or g_093143_(_054870_, _055068_, _055143_);
  and g_093144_(_055142_, _055143_, _055144_);
  not g_093145_(_055144_, _055145_);
  xor g_093146_(out[633], _022989_, _055146_);
  xor g_093147_(_055645_, _022989_, _055147_);
  and g_093148_(_055144_, _055147_, _055148_);
  or g_093149_(_055145_, _055146_, _055149_);
  or g_093150_(_022890_, _023033_, _055151_);
  or g_093151_(_055144_, _055147_, _055152_);
  not g_093152_(_055152_, _055153_);
  xor g_093153_(out[632], _022978_, _055154_);
  or g_093154_(_054888_, _055067_, _055155_);
  or g_093155_(_054882_, _055068_, _055156_);
  and g_093156_(_055155_, _055156_, _055157_);
  and g_093157_(_055154_, _055157_, _055158_);
  not g_093158_(_055158_, _055159_);
  and g_093159_(_055152_, _055159_, _055160_);
  or g_093160_(_055153_, _055158_, _055162_);
  or g_093161_(_055154_, _055157_, _055163_);
  not g_093162_(_055163_, _055164_);
  and g_093163_(_055149_, _055160_, _055165_);
  or g_093164_(_055148_, _055162_, _055166_);
  and g_093165_(_055141_, _055151_, _055167_);
  not g_093166_(_055167_, _055168_);
  and g_093167_(_055138_, _055167_, _055169_);
  or g_093168_(_055140_, _055168_, _055170_);
  and g_093169_(_055163_, _055169_, _055171_);
  or g_093170_(_055164_, _055170_, _055173_);
  and g_093171_(_055165_, _055171_, _055174_);
  or g_093172_(_055166_, _055173_, _055175_);
  xor g_093173_(out[631], _022967_, _055176_);
  xor g_093174_(_055546_, _022967_, _055177_);
  and g_093175_(_054928_, _055068_, _055178_);
  or g_093176_(_054927_, _055067_, _055179_);
  and g_093177_(_054921_, _055067_, _055180_);
  or g_093178_(_054922_, _055068_, _055181_);
  and g_093179_(_055179_, _055181_, _055182_);
  or g_093180_(_055178_, _055180_, _055184_);
  and g_093181_(_055177_, _055184_, _055185_);
  or g_093182_(_055177_, _055184_, _055186_);
  xor g_093183_(_055176_, _055182_, _055187_);
  xor g_093184_(_055177_, _055182_, _055188_);
  xor g_093185_(out[630], _022956_, _055189_);
  not g_093186_(_055189_, _055190_);
  and g_093187_(_054917_, _055068_, _055191_);
  or g_093188_(_054916_, _055067_, _055192_);
  and g_093189_(_054911_, _055067_, _055193_);
  or g_093190_(_054910_, _055068_, _055195_);
  and g_093191_(_055192_, _055195_, _055196_);
  or g_093192_(_055191_, _055193_, _055197_);
  and g_093193_(_055190_, _055196_, _055198_);
  and g_093194_(_055079_, _055082_, _055199_);
  xor g_093195_(_055189_, _055196_, _055200_);
  or g_093196_(_055199_, _055200_, _055201_);
  not g_093197_(_055201_, _055202_);
  and g_093198_(_055187_, _055202_, _055203_);
  or g_093199_(_055188_, _055201_, _055204_);
  or g_093200_(_055175_, _055204_, _055206_);
  and g_093201_(_055162_, _055169_, _055207_);
  and g_093202_(_055149_, _055207_, _055208_);
  and g_093203_(_055140_, _055151_, _055209_);
  or g_093204_(_055208_, _055209_, _055210_);
  and g_093205_(_055186_, _055198_, _055211_);
  and g_093206_(_055124_, _055203_, _055212_);
  or g_093207_(_055211_, _055212_, _055213_);
  or g_093208_(_055185_, _055213_, _055214_);
  and g_093209_(_055174_, _055214_, _055215_);
  or g_093210_(_055210_, _055215_, _055217_);
  or g_093211_(out[624], _055112_, _055218_);
  and g_093212_(_055122_, _055218_, _055219_);
  and g_093213_(_055086_, _055115_, _055220_);
  and g_093214_(_055103_, _055219_, _055221_);
  and g_093215_(_055220_, _055221_, _055222_);
  not g_093216_(_055222_, _055223_);
  or g_093217_(_055206_, _055223_, _055224_);
  and g_093218_(_055217_, _055224_, _055225_);
  not g_093219_(_055225_, _055226_);
  or g_093220_(_055071_, _055225_, _055228_);
  and g_093221_(_055088_, _055225_, _055229_);
  not g_093222_(_055229_, _055230_);
  and g_093223_(_055228_, _055230_, _055231_);
  not g_093224_(_055231_, _055232_);
  and g_093225_(_023044_, _023187_, _055233_);
  or g_093226_(_023055_, _023176_, _055234_);
  or g_093227_(_055132_, _055225_, _055235_);
  not g_093228_(_055235_, _055236_);
  and g_093229_(_055134_, _055225_, _055237_);
  not g_093230_(_055237_, _055239_);
  and g_093231_(_055235_, _055239_, _055240_);
  or g_093232_(_055236_, _055237_, _055241_);
  xor g_093233_(out[650], _023154_, _055242_);
  xor g_093234_(_055788_, _023154_, _055243_);
  and g_093235_(_055240_, _055242_, _055244_);
  or g_093236_(_055241_, _055243_, _055245_);
  and g_093237_(_055234_, _055245_, _055246_);
  or g_093238_(_055233_, _055244_, _055247_);
  and g_093239_(_055241_, _055243_, _055248_);
  or g_093240_(_055240_, _055242_, _055250_);
  and g_093241_(_023055_, _023176_, _055251_);
  or g_093242_(_023044_, _023187_, _055252_);
  and g_093243_(_055250_, _055252_, _055253_);
  or g_093244_(_055248_, _055251_, _055254_);
  and g_093245_(_055246_, _055253_, _055255_);
  or g_093246_(_055247_, _055254_, _055256_);
  or g_093247_(_055146_, _055226_, _055257_);
  or g_093248_(_055144_, _055225_, _055258_);
  and g_093249_(_055257_, _055258_, _055259_);
  not g_093250_(_055259_, _055261_);
  xor g_093251_(out[649], _023143_, _055262_);
  xor g_093252_(_055777_, _023143_, _055263_);
  and g_093253_(_055261_, _055262_, _055264_);
  or g_093254_(_055259_, _055263_, _055265_);
  xor g_093255_(out[648], _023132_, _055266_);
  and g_093256_(_055154_, _055225_, _055267_);
  not g_093257_(_055267_, _055268_);
  or g_093258_(_055157_, _055225_, _055269_);
  and g_093259_(_055268_, _055269_, _055270_);
  and g_093260_(_055266_, _055270_, _055272_);
  not g_093261_(_055272_, _055273_);
  and g_093262_(_055265_, _055273_, _055274_);
  or g_093263_(_055264_, _055272_, _055275_);
  or g_093264_(_055266_, _055270_, _055276_);
  not g_093265_(_055276_, _055277_);
  and g_093266_(_055259_, _055263_, _055278_);
  or g_093267_(_055261_, _055262_, _055279_);
  and g_093268_(_055276_, _055279_, _055280_);
  or g_093269_(_055277_, _055278_, _055281_);
  and g_093270_(_055274_, _055280_, _055283_);
  or g_093271_(_055275_, _055281_, _055284_);
  and g_093272_(_055255_, _055283_, _055285_);
  or g_093273_(_055256_, _055284_, _055286_);
  xor g_093274_(out[646], _023110_, _055287_);
  not g_093275_(_055287_, _055288_);
  and g_093276_(_055196_, _055226_, _055289_);
  or g_093277_(_055197_, _055225_, _055290_);
  and g_093278_(_055189_, _055225_, _055291_);
  not g_093279_(_055291_, _055292_);
  or g_093280_(_055289_, _055291_, _055294_);
  and g_093281_(_055290_, _055292_, _055295_);
  or g_093282_(_055287_, _055295_, _055296_);
  xor g_093283_(out[647], _023121_, _055297_);
  not g_093284_(_055297_, _055298_);
  and g_093285_(_055176_, _055225_, _055299_);
  not g_093286_(_055299_, _055300_);
  and g_093287_(_055184_, _055226_, _055301_);
  or g_093288_(_055182_, _055225_, _055302_);
  and g_093289_(_055300_, _055302_, _055303_);
  or g_093290_(_055299_, _055301_, _055305_);
  or g_093291_(_055297_, _055303_, _055306_);
  and g_093292_(_055296_, _055306_, _055307_);
  and g_093293_(_055297_, _055303_, _055308_);
  or g_093294_(_055298_, _055305_, _055309_);
  or g_093295_(_055288_, _055294_, _055310_);
  and g_093296_(_055309_, _055310_, _055311_);
  xor g_093297_(_055287_, _055294_, _055312_);
  xor g_093298_(_055298_, _055303_, _055313_);
  and g_093299_(_055307_, _055311_, _055314_);
  or g_093300_(_055312_, _055313_, _055316_);
  xor g_093301_(out[645], _023099_, _055317_);
  xor g_093302_(_055700_, _023099_, _055318_);
  and g_093303_(_055079_, _055225_, _055319_);
  not g_093304_(_055319_, _055320_);
  or g_093305_(_055082_, _055225_, _055321_);
  not g_093306_(_055321_, _055322_);
  and g_093307_(_055320_, _055321_, _055323_);
  or g_093308_(_055319_, _055322_, _055324_);
  and g_093309_(_055317_, _055324_, _055325_);
  or g_093310_(_055318_, _055323_, _055327_);
  xor g_093311_(out[644], _023088_, _055328_);
  xor g_093312_(_055711_, _023088_, _055329_);
  or g_093313_(_055076_, _055225_, _055330_);
  not g_093314_(_055330_, _055331_);
  and g_093315_(_055072_, _055225_, _055332_);
  not g_093316_(_055332_, _055333_);
  and g_093317_(_055330_, _055333_, _055334_);
  or g_093318_(_055331_, _055332_, _055335_);
  and g_093319_(_055328_, _055334_, _055336_);
  or g_093320_(_055329_, _055335_, _055338_);
  and g_093321_(_055327_, _055338_, _055339_);
  or g_093322_(_055325_, _055336_, _055340_);
  and g_093323_(_055318_, _055323_, _055341_);
  or g_093324_(_055317_, _055324_, _055342_);
  and g_093325_(_055329_, _055335_, _055343_);
  or g_093326_(_055328_, _055334_, _055344_);
  and g_093327_(_055342_, _055344_, _055345_);
  or g_093328_(_055341_, _055343_, _055346_);
  and g_093329_(_055339_, _055345_, _055347_);
  or g_093330_(_055340_, _055346_, _055349_);
  and g_093331_(_055314_, _055347_, _055350_);
  or g_093332_(_055316_, _055349_, _055351_);
  and g_093333_(_055285_, _055350_, _055352_);
  or g_093334_(_055286_, _055351_, _055353_);
  xor g_093335_(out[643], _023066_, _055354_);
  and g_093336_(_055232_, _055354_, _055355_);
  or g_093337_(out[641], out[642], _055356_);
  xor g_093338_(out[641], out[642], _055357_);
  xor g_093339_(_055722_, out[642], _055358_);
  or g_093340_(_055091_, _055226_, _055360_);
  or g_093341_(_055097_, _055225_, _055361_);
  and g_093342_(_055360_, _055361_, _055362_);
  and g_093343_(_055358_, _055362_, _055363_);
  or g_093344_(_055355_, _055363_, _055364_);
  or g_093345_(_055232_, _055354_, _055365_);
  xor g_093346_(_055232_, _055354_, _055366_);
  xor g_093347_(_055231_, _055354_, _055367_);
  xor g_093348_(_055358_, _055362_, _055368_);
  xor g_093349_(_055357_, _055362_, _055369_);
  and g_093350_(_055366_, _055368_, _055371_);
  or g_093351_(_055367_, _055369_, _055372_);
  or g_093352_(_055590_, _055226_, _055373_);
  or g_093353_(_055107_, _055225_, _055374_);
  and g_093354_(_055373_, _055374_, _055375_);
  and g_093355_(out[641], _055375_, _055376_);
  or g_093356_(_055111_, _055225_, _055377_);
  or g_093357_(out[624], _055226_, _055378_);
  and g_093358_(_055377_, _055378_, _055379_);
  not g_093359_(_055379_, _055380_);
  and g_093360_(out[640], _055380_, _055382_);
  or g_093361_(_055733_, _055379_, _055383_);
  xor g_093362_(out[641], _055375_, _055384_);
  xor g_093363_(_055722_, _055375_, _055385_);
  and g_093364_(_055383_, _055384_, _055386_);
  or g_093365_(_055382_, _055385_, _055387_);
  or g_093366_(_055376_, _055386_, _055388_);
  and g_093367_(_055371_, _055388_, _055389_);
  and g_093368_(_055364_, _055365_, _055390_);
  or g_093369_(_055389_, _055390_, _055391_);
  and g_093370_(_055352_, _055391_, _055393_);
  not g_093371_(_055393_, _055394_);
  or g_093372_(_055307_, _055308_, _055395_);
  not g_093373_(_055395_, _055396_);
  and g_093374_(_055340_, _055342_, _055397_);
  or g_093375_(_055316_, _055339_, _055398_);
  and g_093376_(_055314_, _055397_, _055399_);
  or g_093377_(_055341_, _055398_, _055400_);
  and g_093378_(_055395_, _055400_, _055401_);
  or g_093379_(_055396_, _055399_, _055402_);
  and g_093380_(_055285_, _055402_, _055404_);
  or g_093381_(_055286_, _055401_, _055405_);
  and g_093382_(_055247_, _055252_, _055406_);
  or g_093383_(_055246_, _055251_, _055407_);
  and g_093384_(_055255_, _055275_, _055408_);
  or g_093385_(_055256_, _055274_, _055409_);
  and g_093386_(_055279_, _055408_, _055410_);
  or g_093387_(_055278_, _055409_, _055411_);
  and g_093388_(_055407_, _055411_, _055412_);
  or g_093389_(_055406_, _055410_, _055413_);
  and g_093390_(_055405_, _055412_, _055415_);
  or g_093391_(_055404_, _055413_, _055416_);
  and g_093392_(_055394_, _055415_, _055417_);
  or g_093393_(_055393_, _055416_, _055418_);
  and g_093394_(_055733_, _055379_, _055419_);
  or g_093395_(out[640], _055380_, _055420_);
  and g_093396_(_055371_, _055420_, _055421_);
  or g_093397_(_055372_, _055419_, _055422_);
  and g_093398_(_055386_, _055421_, _055423_);
  or g_093399_(_055387_, _055422_, _055424_);
  and g_093400_(_055352_, _055423_, _055426_);
  or g_093401_(_055353_, _055424_, _055427_);
  and g_093402_(_055418_, _055427_, _055428_);
  or g_093403_(_055417_, _055426_, _055429_);
  or g_093404_(_055231_, _055428_, _055430_);
  or g_093405_(_055354_, _055429_, _055431_);
  and g_093406_(_055430_, _055431_, _055432_);
  not g_093407_(_055432_, _055433_);
  and g_093408_(_053992_, _055433_, _055434_);
  or g_093409_(_053993_, _055432_, _055435_);
  or g_093410_(out[657], out[658], _055437_);
  xor g_093411_(out[657], out[658], _055438_);
  xor g_093412_(_055854_, out[658], _055439_);
  or g_093413_(_055357_, _055429_, _055440_);
  or g_093414_(_055362_, _055428_, _055441_);
  and g_093415_(_055440_, _055441_, _055442_);
  not g_093416_(_055442_, _055443_);
  and g_093417_(_055439_, _055442_, _055444_);
  or g_093418_(_055438_, _055443_, _055445_);
  and g_093419_(_055435_, _055445_, _055446_);
  or g_093420_(_055434_, _055444_, _055448_);
  and g_093421_(_053993_, _055432_, _055449_);
  or g_093422_(_053992_, _055433_, _055450_);
  and g_093423_(_055438_, _055443_, _055451_);
  or g_093424_(_055439_, _055442_, _055452_);
  and g_093425_(_055450_, _055452_, _055453_);
  or g_093426_(_055449_, _055451_, _055454_);
  and g_093427_(_055446_, _055453_, _055455_);
  or g_093428_(_055448_, _055454_, _055456_);
  or g_093429_(_055722_, _055429_, _055457_);
  or g_093430_(_055375_, _055428_, _055459_);
  and g_093431_(_055457_, _055459_, _055460_);
  and g_093432_(out[657], _055460_, _055461_);
  not g_093433_(_055461_, _055462_);
  or g_093434_(_055379_, _055428_, _055463_);
  not g_093435_(_055463_, _055464_);
  and g_093436_(_055733_, _055428_, _055465_);
  not g_093437_(_055465_, _055466_);
  and g_093438_(_055463_, _055466_, _055467_);
  or g_093439_(_055464_, _055465_, _055468_);
  and g_093440_(out[656], _055468_, _055470_);
  or g_093441_(_055865_, _055467_, _055471_);
  xor g_093442_(out[657], _055460_, _055472_);
  xor g_093443_(_055854_, _055460_, _055473_);
  and g_093444_(_055471_, _055472_, _055474_);
  or g_093445_(_055470_, _055473_, _055475_);
  and g_093446_(_055462_, _055475_, _055476_);
  or g_093447_(_055461_, _055474_, _055477_);
  and g_093448_(_055455_, _055477_, _055478_);
  or g_093449_(_055456_, _055476_, _055479_);
  and g_093450_(_055448_, _055450_, _055481_);
  or g_093451_(_055446_, _055449_, _055482_);
  and g_093452_(_055479_, _055482_, _055483_);
  or g_093453_(_055478_, _055481_, _055484_);
  and g_093454_(_055241_, _055429_, _055485_);
  or g_093455_(_055240_, _055428_, _055486_);
  and g_093456_(_055242_, _055428_, _055487_);
  or g_093457_(_055243_, _055429_, _055488_);
  and g_093458_(_055486_, _055488_, _055489_);
  or g_093459_(_055485_, _055487_, _055490_);
  or g_093460_(_053990_, _055489_, _055492_);
  not g_093461_(_055492_, _055493_);
  and g_093462_(_053990_, _055489_, _055494_);
  or g_093463_(_053991_, _055490_, _055495_);
  and g_093464_(_023198_, _023330_, _055496_);
  or g_093465_(_023198_, _023330_, _055497_);
  xor g_093466_(_023198_, _023330_, _055498_);
  xor g_093467_(_023209_, _023330_, _055499_);
  and g_093468_(_055495_, _055498_, _055500_);
  or g_093469_(_055494_, _055499_, _055501_);
  and g_093470_(_055492_, _055500_, _055503_);
  or g_093471_(_055493_, _055501_, _055504_);
  xor g_093472_(out[665], _023297_, _055505_);
  xor g_093473_(_055909_, _023297_, _055506_);
  and g_093474_(_055263_, _055428_, _055507_);
  not g_093475_(_055507_, _055508_);
  or g_093476_(_055259_, _055428_, _055509_);
  not g_093477_(_055509_, _055510_);
  and g_093478_(_055508_, _055509_, _055511_);
  or g_093479_(_055507_, _055510_, _055512_);
  and g_093480_(_055505_, _055512_, _055514_);
  or g_093481_(_055506_, _055511_, _055515_);
  xor g_093482_(out[664], _023286_, _055516_);
  not g_093483_(_055516_, _055517_);
  and g_093484_(_055266_, _055428_, _055518_);
  not g_093485_(_055518_, _055519_);
  or g_093486_(_055270_, _055428_, _055520_);
  not g_093487_(_055520_, _055521_);
  and g_093488_(_055519_, _055520_, _055522_);
  or g_093489_(_055518_, _055521_, _055523_);
  and g_093490_(_055516_, _055522_, _055525_);
  or g_093491_(_055517_, _055523_, _055526_);
  and g_093492_(_055515_, _055526_, _055527_);
  or g_093493_(_055514_, _055525_, _055528_);
  and g_093494_(_055506_, _055511_, _055529_);
  or g_093495_(_055505_, _055512_, _055530_);
  and g_093496_(_055517_, _055523_, _055531_);
  or g_093497_(_055516_, _055522_, _055532_);
  and g_093498_(_055530_, _055532_, _055533_);
  or g_093499_(_055529_, _055531_, _055534_);
  and g_093500_(_055527_, _055533_, _055536_);
  or g_093501_(_055528_, _055534_, _055537_);
  and g_093502_(_055503_, _055536_, _055538_);
  or g_093503_(_055504_, _055537_, _055539_);
  xor g_093504_(out[661], _023253_, _055540_);
  xor g_093505_(_055832_, _023253_, _055541_);
  and g_093506_(_055318_, _055428_, _055542_);
  or g_093507_(_055317_, _055429_, _055543_);
  and g_093508_(_055324_, _055429_, _055544_);
  or g_093509_(_055323_, _055428_, _055545_);
  and g_093510_(_055543_, _055545_, _055547_);
  or g_093511_(_055542_, _055544_, _055548_);
  and g_093512_(_055540_, _055548_, _055549_);
  or g_093513_(_055541_, _055547_, _055550_);
  and g_093514_(_055541_, _055547_, _055551_);
  or g_093515_(_055540_, _055548_, _055552_);
  xor g_093516_(out[662], _023264_, _055553_);
  xor g_093517_(_055821_, _023264_, _055554_);
  and g_093518_(_055288_, _055428_, _055555_);
  or g_093519_(_055287_, _055429_, _055556_);
  and g_093520_(_055295_, _055429_, _055558_);
  or g_093521_(_055294_, _055428_, _055559_);
  and g_093522_(_055556_, _055559_, _055560_);
  or g_093523_(_055555_, _055558_, _055561_);
  or g_093524_(_055554_, _055560_, _055562_);
  not g_093525_(_055562_, _055563_);
  xor g_093526_(out[660], _023242_, _055564_);
  not g_093527_(_055564_, _055565_);
  and g_093528_(_055328_, _055428_, _055566_);
  not g_093529_(_055566_, _055567_);
  or g_093530_(_055334_, _055428_, _055569_);
  not g_093531_(_055569_, _055570_);
  and g_093532_(_055567_, _055569_, _055571_);
  or g_093533_(_055566_, _055570_, _055572_);
  and g_093534_(_055565_, _055572_, _055573_);
  or g_093535_(_055564_, _055571_, _055574_);
  and g_093536_(_055554_, _055560_, _055575_);
  or g_093537_(_055553_, _055561_, _055576_);
  xor g_093538_(out[663], _023275_, _055577_);
  not g_093539_(_055577_, _055578_);
  and g_093540_(_055297_, _055428_, _055580_);
  or g_093541_(_055298_, _055429_, _055581_);
  and g_093542_(_055305_, _055429_, _055582_);
  or g_093543_(_055303_, _055428_, _055583_);
  and g_093544_(_055581_, _055583_, _055584_);
  or g_093545_(_055580_, _055582_, _055585_);
  and g_093546_(_055578_, _055585_, _055586_);
  or g_093547_(_055577_, _055584_, _055587_);
  and g_093548_(_055576_, _055587_, _055588_);
  or g_093549_(_055575_, _055586_, _055589_);
  and g_093550_(_055577_, _055584_, _055591_);
  not g_093551_(_055591_, _055592_);
  and g_093552_(_055564_, _055571_, _055593_);
  or g_093553_(_055565_, _055572_, _055594_);
  and g_093554_(_055550_, _055574_, _055595_);
  or g_093555_(_055549_, _055573_, _055596_);
  and g_093556_(_055552_, _055595_, _055597_);
  or g_093557_(_055551_, _055596_, _055598_);
  and g_093558_(_055594_, _055597_, _055599_);
  or g_093559_(_055593_, _055598_, _055600_);
  and g_093560_(_055562_, _055588_, _055602_);
  or g_093561_(_055563_, _055589_, _055603_);
  and g_093562_(_055592_, _055602_, _055604_);
  or g_093563_(_055591_, _055603_, _055605_);
  and g_093564_(_055599_, _055604_, _055606_);
  or g_093565_(_055600_, _055605_, _055607_);
  and g_093566_(_055538_, _055606_, _055608_);
  and g_093567_(_055484_, _055608_, _055609_);
  or g_093568_(_055504_, _055527_, _055610_);
  or g_093569_(_055529_, _055610_, _055611_);
  and g_093570_(_055494_, _055497_, _055613_);
  or g_093571_(_055496_, _055613_, _055614_);
  not g_093572_(_055614_, _055615_);
  and g_093573_(_055611_, _055615_, _055616_);
  not g_093574_(_055616_, _055617_);
  and g_093575_(_055550_, _055594_, _055618_);
  or g_093576_(_055549_, _055593_, _055619_);
  and g_093577_(_055552_, _055562_, _055620_);
  or g_093578_(_055551_, _055563_, _055621_);
  and g_093579_(_055619_, _055620_, _055622_);
  or g_093580_(_055618_, _055621_, _055624_);
  and g_093581_(_055588_, _055624_, _055625_);
  or g_093582_(_055589_, _055622_, _055626_);
  and g_093583_(_055592_, _055626_, _055627_);
  or g_093584_(_055591_, _055625_, _055628_);
  and g_093585_(_055538_, _055627_, _055629_);
  or g_093586_(_055617_, _055629_, _055630_);
  or g_093587_(_055483_, _055607_, _055631_);
  and g_093588_(_055628_, _055631_, _055632_);
  or g_093589_(_055539_, _055632_, _055633_);
  and g_093590_(_055616_, _055633_, _055635_);
  or g_093591_(_055609_, _055630_, _055636_);
  or g_093592_(out[656], _055468_, _055637_);
  and g_093593_(_055474_, _055637_, _055638_);
  and g_093594_(_055608_, _055638_, _055639_);
  not g_093595_(_055639_, _055640_);
  and g_093596_(_055455_, _055639_, _055641_);
  or g_093597_(_055456_, _055640_, _055642_);
  and g_093598_(_055636_, _055642_, _055643_);
  or g_093599_(_055635_, _055641_, _055644_);
  and g_093600_(_053990_, _055643_, _055646_);
  or g_093601_(_053991_, _055644_, _055647_);
  or g_093602_(_055489_, _055643_, _055648_);
  not g_093603_(_055648_, _055649_);
  and g_093604_(_055647_, _055648_, _055650_);
  or g_093605_(_055646_, _055649_, _055651_);
  xor g_093606_(out[679], _023418_, _055652_);
  not g_093607_(_055652_, _055653_);
  or g_093608_(_055584_, _055643_, _055654_);
  or g_093609_(_055578_, _055644_, _055655_);
  and g_093610_(_055654_, _055655_, _055657_);
  and g_093611_(_055652_, _055657_, _055658_);
  or g_093612_(_055652_, _055657_, _055659_);
  xor g_093613_(_055653_, _055657_, _055660_);
  xor g_093614_(out[677], _023396_, _055661_);
  xor g_093615_(_055964_, _023396_, _055662_);
  or g_093616_(_055547_, _055643_, _055663_);
  or g_093617_(_055540_, _055644_, _055664_);
  and g_093618_(_055663_, _055664_, _055665_);
  not g_093619_(_055665_, _055666_);
  and g_093620_(_055662_, _055665_, _055668_);
  xor g_093621_(out[678], _023407_, _055669_);
  or g_093622_(_055560_, _055643_, _055670_);
  not g_093623_(_055670_, _055671_);
  and g_093624_(_055554_, _055643_, _055672_);
  not g_093625_(_055672_, _055673_);
  and g_093626_(_055670_, _055673_, _055674_);
  or g_093627_(_055671_, _055672_, _055675_);
  or g_093628_(_055669_, _055675_, _055676_);
  xor g_093629_(_055669_, _055674_, _055677_);
  or g_093630_(_055660_, _055677_, _055679_);
  or g_093631_(_055668_, _055679_, _055680_);
  or g_093632_(_023341_, _023473_, _055681_);
  not g_093633_(_055681_, _055682_);
  xor g_093634_(out[682], _023451_, _055683_);
  xor g_093635_(_000087_, _023451_, _055684_);
  and g_093636_(_055650_, _055683_, _055685_);
  or g_093637_(_055651_, _055684_, _055686_);
  and g_093638_(_055681_, _055686_, _055687_);
  or g_093639_(_055682_, _055685_, _055688_);
  and g_093640_(_055651_, _055684_, _055690_);
  and g_093641_(_023341_, _023473_, _055691_);
  or g_093642_(_055688_, _055691_, _055692_);
  or g_093643_(_055690_, _055692_, _055693_);
  or g_093644_(_055511_, _055643_, _055694_);
  not g_093645_(_055694_, _055695_);
  and g_093646_(_055506_, _055643_, _055696_);
  not g_093647_(_055696_, _055697_);
  and g_093648_(_055694_, _055697_, _055698_);
  or g_093649_(_055695_, _055696_, _055699_);
  xor g_093650_(out[681], _023440_, _055701_);
  xor g_093651_(_000076_, _023440_, _055702_);
  and g_093652_(_055699_, _055701_, _055703_);
  or g_093653_(_055698_, _055702_, _055704_);
  xor g_093654_(out[680], _023429_, _055705_);
  not g_093655_(_055705_, _055706_);
  or g_093656_(_055522_, _055643_, _055707_);
  not g_093657_(_055707_, _055708_);
  and g_093658_(_055516_, _055643_, _055709_);
  not g_093659_(_055709_, _055710_);
  and g_093660_(_055707_, _055710_, _055712_);
  or g_093661_(_055708_, _055709_, _055713_);
  and g_093662_(_055705_, _055712_, _055714_);
  or g_093663_(_055706_, _055713_, _055715_);
  and g_093664_(_055704_, _055715_, _055716_);
  or g_093665_(_055703_, _055714_, _055717_);
  and g_093666_(_055706_, _055713_, _055718_);
  and g_093667_(_055698_, _055702_, _055719_);
  or g_093668_(_055718_, _055719_, _055720_);
  or g_093669_(_055717_, _055720_, _055721_);
  or g_093670_(_055693_, _055721_, _055723_);
  and g_093671_(_055661_, _055666_, _055724_);
  or g_093672_(_055662_, _055665_, _055725_);
  xor g_093673_(out[676], _023385_, _055726_);
  not g_093674_(_055726_, _055727_);
  and g_093675_(_055564_, _055643_, _055728_);
  and g_093676_(_055572_, _055644_, _055729_);
  or g_093677_(_055728_, _055729_, _055730_);
  not g_093678_(_055730_, _055731_);
  and g_093679_(_055726_, _055731_, _055732_);
  or g_093680_(_055727_, _055730_, _055734_);
  and g_093681_(_055725_, _055734_, _055735_);
  or g_093682_(_055724_, _055732_, _055736_);
  and g_093683_(_055727_, _055730_, _055737_);
  or g_093684_(_055736_, _055737_, _055738_);
  or g_093685_(_055680_, _055738_, _055739_);
  or g_093686_(_055723_, _055739_, _055740_);
  or g_093687_(out[673], out[674], _055741_);
  xor g_093688_(_000021_, out[674], _055742_);
  not g_093689_(_055742_, _055743_);
  and g_093690_(_055443_, _055644_, _055745_);
  and g_093691_(_055439_, _055643_, _055746_);
  or g_093692_(_055745_, _055746_, _055747_);
  or g_093693_(_055743_, _055747_, _055748_);
  xor g_093694_(out[675], _023363_, _055749_);
  xor g_093695_(_000054_, _023363_, _055750_);
  or g_093696_(_055432_, _055643_, _055751_);
  or g_093697_(_053992_, _055644_, _055752_);
  and g_093698_(_055751_, _055752_, _055753_);
  not g_093699_(_055753_, _055754_);
  or g_093700_(_055750_, _055753_, _055756_);
  and g_093701_(_055748_, _055756_, _055757_);
  and g_093702_(_055750_, _055753_, _055758_);
  xor g_093703_(_055749_, _055753_, _055759_);
  xor g_093704_(_055742_, _055747_, _055760_);
  or g_093705_(_055740_, _055759_, _055761_);
  or g_093706_(_055760_, _055761_, _055762_);
  and g_093707_(out[657], _055643_, _055763_);
  or g_093708_(_055460_, _055643_, _055764_);
  not g_093709_(_055764_, _055765_);
  or g_093710_(_055763_, _055765_, _055767_);
  or g_093711_(_000021_, _055767_, _055768_);
  or g_093712_(_055762_, _055768_, _055769_);
  or g_093713_(_055680_, _055735_, _055770_);
  and g_093714_(_055659_, _055676_, _055771_);
  or g_093715_(_055658_, _055771_, _055772_);
  and g_093716_(_055770_, _055772_, _055773_);
  or g_093717_(_055723_, _055773_, _055774_);
  or g_093718_(_055757_, _055758_, _055775_);
  or g_093719_(_055740_, _055775_, _055776_);
  or g_093720_(_055687_, _055691_, _055778_);
  or g_093721_(_055716_, _055719_, _055779_);
  or g_093722_(_055693_, _055779_, _055780_);
  and g_093723_(_055778_, _055780_, _055781_);
  and g_093724_(_055776_, _055781_, _055782_);
  and g_093725_(_055774_, _055782_, _055783_);
  and g_093726_(_055769_, _055783_, _055784_);
  and g_093727_(_055468_, _055644_, _055785_);
  and g_093728_(_055865_, _055643_, _055786_);
  or g_093729_(_055785_, _055786_, _055787_);
  not g_093730_(_055787_, _055789_);
  and g_093731_(out[672], _055787_, _055790_);
  xor g_093732_(out[673], _055767_, _055791_);
  or g_093733_(_055790_, _055791_, _055792_);
  or g_093734_(_055762_, _055792_, _055793_);
  or g_093735_(out[672], _055787_, _055794_);
  or g_093736_(_055793_, _055794_, _055795_);
  and g_093737_(_055784_, _055795_, _055796_);
  not g_093738_(_055796_, _055797_);
  or g_093739_(_055650_, _055797_, _055798_);
  or g_093740_(_055684_, _055796_, _055800_);
  and g_093741_(_055798_, _055800_, _055801_);
  not g_093742_(_055801_, _055802_);
  xor g_093743_(out[698], _023605_, _055803_);
  and g_093744_(_055801_, _055803_, _055804_);
  and g_093745_(_023495_, _023638_, _055805_);
  or g_093746_(_023495_, _023638_, _055806_);
  xor g_093747_(_023506_, _023627_, _055807_);
  xor g_093748_(_023506_, _023638_, _055808_);
  xor g_093749_(_055801_, _055803_, _055809_);
  xor g_093750_(_055802_, _055803_, _055811_);
  and g_093751_(_055807_, _055809_, _055812_);
  or g_093752_(_055808_, _055811_, _055813_);
  or g_093753_(_055701_, _055796_, _055814_);
  not g_093754_(_055814_, _055815_);
  and g_093755_(_055699_, _055796_, _055816_);
  or g_093756_(_055698_, _055797_, _055817_);
  and g_093757_(_055814_, _055817_, _055818_);
  or g_093758_(_055815_, _055816_, _055819_);
  xor g_093759_(out[697], _023594_, _055820_);
  xor g_093760_(_000208_, _023594_, _055822_);
  and g_093761_(_055818_, _055822_, _055823_);
  or g_093762_(_055819_, _055820_, _055824_);
  xor g_093763_(out[696], _023583_, _055825_);
  not g_093764_(_055825_, _055826_);
  and g_093765_(_055705_, _055797_, _055827_);
  or g_093766_(_055706_, _055796_, _055828_);
  and g_093767_(_055713_, _055796_, _055829_);
  not g_093768_(_055829_, _055830_);
  and g_093769_(_055828_, _055830_, _055831_);
  or g_093770_(_055827_, _055829_, _055833_);
  and g_093771_(_055826_, _055833_, _055834_);
  or g_093772_(_055825_, _055831_, _055835_);
  and g_093773_(_055824_, _055835_, _055836_);
  or g_093774_(_055823_, _055834_, _055837_);
  and g_093775_(_055819_, _055820_, _055838_);
  or g_093776_(_055818_, _055822_, _055839_);
  and g_093777_(_055825_, _055831_, _055840_);
  or g_093778_(_055826_, _055833_, _055841_);
  and g_093779_(_055839_, _055841_, _055842_);
  or g_093780_(_055838_, _055840_, _055844_);
  and g_093781_(_055836_, _055842_, _055845_);
  or g_093782_(_055837_, _055844_, _055846_);
  and g_093783_(_055812_, _055845_, _055847_);
  or g_093784_(_055813_, _055846_, _055848_);
  xor g_093785_(out[694], _023561_, _055849_);
  xor g_093786_(_000120_, _023561_, _055850_);
  or g_093787_(_055669_, _055796_, _055851_);
  not g_093788_(_055851_, _055852_);
  and g_093789_(_055675_, _055796_, _055853_);
  or g_093790_(_055674_, _055797_, _055855_);
  and g_093791_(_055851_, _055855_, _055856_);
  or g_093792_(_055852_, _055853_, _055857_);
  and g_093793_(_055849_, _055857_, _055858_);
  or g_093794_(_055850_, _055856_, _055859_);
  xor g_093795_(out[693], _023550_, _055860_);
  xor g_093796_(_000131_, _023550_, _055861_);
  or g_093797_(_055661_, _055796_, _055862_);
  not g_093798_(_055862_, _055863_);
  and g_093799_(_055666_, _055796_, _055864_);
  or g_093800_(_055665_, _055797_, _055866_);
  and g_093801_(_055862_, _055866_, _055867_);
  or g_093802_(_055863_, _055864_, _055868_);
  and g_093803_(_055861_, _055867_, _055869_);
  or g_093804_(_055860_, _055868_, _055870_);
  and g_093805_(_055859_, _055870_, _055871_);
  or g_093806_(_055858_, _055869_, _055872_);
  xor g_093807_(out[695], _023572_, _055873_);
  xor g_093808_(_000109_, _023572_, _055874_);
  and g_093809_(_055657_, _055796_, _055875_);
  not g_093810_(_055875_, _055877_);
  or g_093811_(_055652_, _055796_, _055878_);
  not g_093812_(_055878_, _055879_);
  or g_093813_(_055875_, _055879_, _055880_);
  and g_093814_(_055877_, _055878_, _055881_);
  and g_093815_(_055873_, _055880_, _055882_);
  or g_093816_(_055874_, _055881_, _055883_);
  xor g_093817_(out[692], _023539_, _055884_);
  not g_093818_(_055884_, _055885_);
  and g_093819_(_055730_, _055796_, _055886_);
  not g_093820_(_055886_, _055888_);
  and g_093821_(_055726_, _055797_, _055889_);
  or g_093822_(_055727_, _055796_, _055890_);
  and g_093823_(_055888_, _055890_, _055891_);
  or g_093824_(_055886_, _055889_, _055892_);
  and g_093825_(_055885_, _055892_, _055893_);
  or g_093826_(_055884_, _055891_, _055894_);
  and g_093827_(_055883_, _055894_, _055895_);
  or g_093828_(_055882_, _055893_, _055896_);
  and g_093829_(_055871_, _055895_, _055897_);
  or g_093830_(_055872_, _055896_, _055899_);
  and g_093831_(_055850_, _055856_, _055900_);
  or g_093832_(_055849_, _055857_, _055901_);
  and g_093833_(_055874_, _055881_, _055902_);
  or g_093834_(_055873_, _055880_, _055903_);
  and g_093835_(_055901_, _055903_, _055904_);
  or g_093836_(_055900_, _055902_, _055905_);
  and g_093837_(_055860_, _055868_, _055906_);
  or g_093838_(_055861_, _055867_, _055907_);
  and g_093839_(_055884_, _055891_, _055908_);
  or g_093840_(_055885_, _055892_, _055910_);
  and g_093841_(_055907_, _055910_, _055911_);
  or g_093842_(_055906_, _055908_, _055912_);
  and g_093843_(_055904_, _055911_, _055913_);
  or g_093844_(_055905_, _055912_, _055914_);
  and g_093845_(_055897_, _055913_, _055915_);
  or g_093846_(_055899_, _055914_, _055916_);
  and g_093847_(_055847_, _055915_, _055917_);
  or g_093848_(_055848_, _055916_, _055918_);
  xor g_093849_(out[691], _023517_, _055919_);
  xor g_093850_(_000186_, _023517_, _055921_);
  and g_093851_(_055754_, _055796_, _055922_);
  or g_093852_(_055753_, _055797_, _055923_);
  or g_093853_(_055749_, _055796_, _055924_);
  not g_093854_(_055924_, _055925_);
  and g_093855_(_055923_, _055924_, _055926_);
  or g_093856_(_055922_, _055925_, _055927_);
  and g_093857_(_055919_, _055927_, _055928_);
  or g_093858_(out[689], out[690], _055929_);
  xor g_093859_(out[689], out[690], _055930_);
  xor g_093860_(_000153_, out[690], _055932_);
  and g_093861_(_055747_, _055796_, _055933_);
  not g_093862_(_055933_, _055934_);
  or g_093863_(_055743_, _055796_, _055935_);
  and g_093864_(_055934_, _055935_, _055936_);
  and g_093865_(_055932_, _055936_, _055937_);
  or g_093866_(_055928_, _055937_, _055938_);
  or g_093867_(_055919_, _055927_, _055939_);
  xor g_093868_(_055921_, _055926_, _055940_);
  xor g_093869_(_055919_, _055926_, _055941_);
  xor g_093870_(_055932_, _055936_, _055943_);
  xor g_093871_(_055930_, _055936_, _055944_);
  and g_093872_(_055940_, _055943_, _055945_);
  or g_093873_(_055941_, _055944_, _055946_);
  or g_093874_(_000021_, _055796_, _055947_);
  and g_093875_(_055767_, _055796_, _055948_);
  not g_093876_(_055948_, _055949_);
  and g_093877_(_055947_, _055949_, _055950_);
  and g_093878_(out[689], _055950_, _055951_);
  not g_093879_(_055951_, _055952_);
  and g_093880_(out[672], _055797_, _055954_);
  or g_093881_(_000032_, _055784_, _055955_);
  and g_093882_(_055789_, _055796_, _055956_);
  or g_093883_(_055787_, _055797_, _055957_);
  and g_093884_(_055955_, _055957_, _055958_);
  or g_093885_(_055954_, _055956_, _055959_);
  and g_093886_(out[688], _055958_, _055960_);
  or g_093887_(_000164_, _055959_, _055961_);
  xor g_093888_(out[689], _055950_, _055962_);
  xor g_093889_(_000153_, _055950_, _055963_);
  and g_093890_(_055961_, _055962_, _000000_);
  or g_093891_(_055960_, _055963_, _000001_);
  and g_093892_(_055952_, _000001_, _000002_);
  or g_093893_(_055951_, _000000_, _000003_);
  and g_093894_(_055945_, _000003_, _000004_);
  or g_093895_(_055946_, _000002_, _000005_);
  and g_093896_(_055938_, _055939_, _000006_);
  not g_093897_(_000006_, _000007_);
  and g_093898_(_000005_, _000007_, _000008_);
  or g_093899_(_000004_, _000006_, _000009_);
  and g_093900_(_055917_, _000009_, _000011_);
  or g_093901_(_055918_, _000008_, _000012_);
  or g_093902_(_055872_, _055911_, _000013_);
  and g_093903_(_055904_, _000013_, _000014_);
  or g_093904_(_055848_, _055882_, _000015_);
  or g_093905_(_000014_, _000015_, _000016_);
  not g_093906_(_000016_, _000017_);
  or g_093907_(_055823_, _055842_, _000018_);
  and g_093908_(_055812_, _055844_, _000019_);
  and g_093909_(_055824_, _000019_, _000020_);
  or g_093910_(_055813_, _000018_, _000022_);
  or g_093911_(_055804_, _055805_, _000023_);
  and g_093912_(_055806_, _000023_, _000024_);
  not g_093913_(_000024_, _000025_);
  and g_093914_(_000022_, _000025_, _000026_);
  or g_093915_(_000020_, _000024_, _000027_);
  and g_093916_(_000012_, _000026_, _000028_);
  or g_093917_(_000011_, _000027_, _000029_);
  and g_093918_(_000016_, _000028_, _000030_);
  or g_093919_(_000017_, _000029_, _000031_);
  or g_093920_(out[688], _055958_, _000033_);
  and g_093921_(_055945_, _000033_, _000034_);
  and g_093922_(_000000_, _000034_, _000035_);
  and g_093923_(_055917_, _000035_, _000036_);
  not g_093924_(_000036_, _000037_);
  and g_093925_(_000031_, _000037_, _000038_);
  or g_093926_(_000030_, _000036_, _000039_);
  or g_093927_(_055801_, _000038_, _000040_);
  not g_093928_(_000040_, _000041_);
  and g_093929_(_055803_, _000038_, _000042_);
  not g_093930_(_000042_, _000044_);
  and g_093931_(_000040_, _000044_, _000045_);
  or g_093932_(_000041_, _000042_, _000046_);
  and g_093933_(_053988_, _000045_, _000047_);
  or g_093934_(_053989_, _000047_, _000048_);
  not g_093935_(_000048_, _000049_);
  or g_093936_(_023649_, _023792_, _000050_);
  or g_093937_(_053988_, _000045_, _000051_);
  and g_093938_(_000050_, _000051_, _000052_);
  and g_093939_(_000049_, _000052_, _000053_);
  xor g_093940_(out[712], _023737_, _000055_);
  or g_093941_(_055826_, _000039_, _000056_);
  or g_093942_(_055831_, _000038_, _000057_);
  and g_093943_(_000056_, _000057_, _000058_);
  and g_093944_(_000055_, _000058_, _000059_);
  and g_093945_(_055822_, _000038_, _000060_);
  and g_093946_(_055819_, _000039_, _000061_);
  or g_093947_(_000060_, _000061_, _000062_);
  xor g_093948_(out[713], _023748_, _000063_);
  and g_093949_(_000062_, _000063_, _000064_);
  or g_093950_(_000062_, _000063_, _000066_);
  xor g_093951_(_000055_, _000058_, _000067_);
  xor g_093952_(_000062_, _000063_, _000068_);
  and g_093953_(_000053_, _000068_, _000069_);
  and g_093954_(_000067_, _000069_, _000070_);
  not g_093955_(_000070_, _000071_);
  xor g_093956_(out[710], _023715_, _000072_);
  xor g_093957_(_000252_, _023715_, _000073_);
  and g_093958_(_055850_, _000038_, _000074_);
  not g_093959_(_000074_, _000075_);
  and g_093960_(_055857_, _000039_, _000077_);
  or g_093961_(_055856_, _000038_, _000078_);
  and g_093962_(_000075_, _000078_, _000079_);
  or g_093963_(_000074_, _000077_, _000080_);
  and g_093964_(_000073_, _000079_, _000081_);
  or g_093965_(_000072_, _000080_, _000082_);
  xor g_093966_(out[711], _023726_, _000083_);
  xor g_093967_(_000241_, _023726_, _000084_);
  and g_093968_(_055873_, _000038_, _000085_);
  or g_093969_(_055874_, _000039_, _000086_);
  or g_093970_(_055880_, _000038_, _000088_);
  not g_093971_(_000088_, _000089_);
  and g_093972_(_000086_, _000088_, _000090_);
  or g_093973_(_000085_, _000089_, _000091_);
  and g_093974_(_000084_, _000091_, _000092_);
  or g_093975_(_000083_, _000090_, _000093_);
  and g_093976_(_000082_, _000093_, _000094_);
  or g_093977_(_000081_, _000092_, _000095_);
  or g_093978_(_000073_, _000079_, _000096_);
  or g_093979_(_000084_, _000091_, _000097_);
  and g_093980_(_000096_, _000097_, _000099_);
  not g_093981_(_000099_, _000100_);
  and g_093982_(_000094_, _000099_, _000101_);
  or g_093983_(_000095_, _000100_, _000102_);
  xor g_093984_(out[708], _023693_, _000103_);
  and g_093985_(_055884_, _000038_, _000104_);
  not g_093986_(_000104_, _000105_);
  or g_093987_(_055891_, _000038_, _000106_);
  not g_093988_(_000106_, _000107_);
  and g_093989_(_000105_, _000106_, _000108_);
  or g_093990_(_000104_, _000107_, _000110_);
  and g_093991_(_000103_, _000108_, _000111_);
  xor g_093992_(out[709], _023704_, _000112_);
  and g_093993_(_055861_, _000038_, _000113_);
  not g_093994_(_000113_, _000114_);
  or g_093995_(_055867_, _000038_, _000115_);
  not g_093996_(_000115_, _000116_);
  and g_093997_(_000114_, _000115_, _000117_);
  or g_093998_(_000113_, _000116_, _000118_);
  and g_093999_(_000112_, _000118_, _000119_);
  or g_094000_(_000111_, _000119_, _000121_);
  not g_094001_(_000121_, _000122_);
  or g_094002_(_000112_, _000118_, _000123_);
  or g_094003_(_000103_, _000108_, _000124_);
  and g_094004_(_000123_, _000124_, _000125_);
  not g_094005_(_000125_, _000126_);
  and g_094006_(_000122_, _000125_, _000127_);
  or g_094007_(_000121_, _000126_, _000128_);
  and g_094008_(_000101_, _000127_, _000129_);
  or g_094009_(_000102_, _000128_, _000130_);
  xor g_094010_(out[707], _023671_, _000132_);
  or g_094011_(_055926_, _000038_, _000133_);
  not g_094012_(_000133_, _000134_);
  and g_094013_(_055921_, _000038_, _000135_);
  not g_094014_(_000135_, _000136_);
  and g_094015_(_000133_, _000136_, _000137_);
  or g_094016_(_000134_, _000135_, _000138_);
  or g_094017_(_000132_, _000138_, _000139_);
  or g_094018_(out[705], out[706], _000140_);
  xor g_094019_(out[705], out[706], _000141_);
  xor g_094020_(_000285_, out[706], _000143_);
  or g_094021_(_055930_, _000039_, _000144_);
  or g_094022_(_055936_, _000038_, _000145_);
  and g_094023_(_000144_, _000145_, _000146_);
  and g_094024_(_000143_, _000146_, _000147_);
  and g_094025_(_000132_, _000138_, _000148_);
  xor g_094026_(_000132_, _000138_, _000149_);
  xor g_094027_(_000143_, _000146_, _000150_);
  and g_094028_(_000149_, _000150_, _000151_);
  or g_094029_(_000153_, _000039_, _000152_);
  or g_094030_(_055950_, _000038_, _000154_);
  and g_094031_(_000152_, _000154_, _000155_);
  and g_094032_(out[705], _000155_, _000156_);
  and g_094033_(out[688], _000038_, _000157_);
  not g_094034_(_000157_, _000158_);
  and g_094035_(_055959_, _000039_, _000159_);
  or g_094036_(_055958_, _000038_, _000160_);
  or g_094037_(_000157_, _000159_, _000161_);
  and g_094038_(_000158_, _000160_, _000162_);
  and g_094039_(out[704], _000162_, _000163_);
  or g_094040_(_000296_, _000161_, _000165_);
  xor g_094041_(out[705], _000155_, _000166_);
  xor g_094042_(_000285_, _000155_, _000167_);
  and g_094043_(_000165_, _000166_, _000168_);
  or g_094044_(_000163_, _000167_, _000169_);
  or g_094045_(_000156_, _000168_, _000170_);
  and g_094046_(_000151_, _000170_, _000171_);
  or g_094047_(_000147_, _000148_, _000172_);
  and g_094048_(_000139_, _000172_, _000173_);
  or g_094049_(_000171_, _000173_, _000174_);
  and g_094050_(_000129_, _000174_, _000176_);
  and g_094051_(_000095_, _000097_, _000177_);
  and g_094052_(_000121_, _000123_, _000178_);
  and g_094053_(_000101_, _000178_, _000179_);
  or g_094054_(_000177_, _000179_, _000180_);
  or g_094055_(_000176_, _000180_, _000181_);
  and g_094056_(_000070_, _000181_, _000182_);
  and g_094057_(_000048_, _000050_, _000183_);
  and g_094058_(_000059_, _000066_, _000184_);
  or g_094059_(_000064_, _000184_, _000185_);
  and g_094060_(_000053_, _000185_, _000187_);
  or g_094061_(_000183_, _000187_, _000188_);
  or g_094062_(_000182_, _000188_, _000189_);
  or g_094063_(out[704], _000162_, _000190_);
  and g_094064_(_000151_, _000190_, _000191_);
  not g_094065_(_000191_, _000192_);
  or g_094066_(_000169_, _000192_, _000193_);
  or g_094067_(_000130_, _000193_, _000194_);
  or g_094068_(_000071_, _000194_, _000195_);
  and g_094069_(_000189_, _000195_, _000196_);
  not g_094070_(_000196_, _000198_);
  and g_094071_(_053988_, _000196_, _000199_);
  not g_094072_(_000199_, _000200_);
  and g_094073_(_000046_, _000198_, _000201_);
  or g_094074_(_000045_, _000196_, _000202_);
  and g_094075_(_000200_, _000202_, _000203_);
  or g_094076_(_000199_, _000201_, _000204_);
  and g_094077_(_053983_, _000203_, _000205_);
  or g_094078_(_053985_, _000204_, _000206_);
  and g_094079_(_053987_, _000206_, _000207_);
  or g_094080_(_053986_, _000205_, _000209_);
  or g_094081_(_023803_, _023946_, _000210_);
  or g_094082_(_053983_, _000203_, _000211_);
  and g_094083_(_000210_, _000211_, _000212_);
  or g_094084_(_000062_, _000196_, _000213_);
  not g_094085_(_000213_, _000214_);
  and g_094086_(_000063_, _000196_, _000215_);
  or g_094087_(_000214_, _000215_, _000216_);
  not g_094088_(_000216_, _000217_);
  xor g_094089_(out[729], _023902_, _000218_);
  xor g_094090_(_000472_, _023902_, _000220_);
  or g_094091_(_000217_, _000218_, _000221_);
  xor g_094092_(out[728], _023891_, _000222_);
  or g_094093_(_000058_, _000196_, _000223_);
  and g_094094_(_000055_, _000196_, _000224_);
  not g_094095_(_000224_, _000225_);
  and g_094096_(_000223_, _000225_, _000226_);
  or g_094097_(_000222_, _000226_, _000227_);
  or g_094098_(_000216_, _000220_, _000228_);
  not g_094099_(_000228_, _000229_);
  and g_094100_(_000222_, _000226_, _000231_);
  not g_094101_(_000231_, _000232_);
  and g_094102_(_000228_, _000232_, _000233_);
  or g_094103_(_000229_, _000231_, _000234_);
  and g_094104_(_000221_, _000233_, _000235_);
  and g_094105_(_000207_, _000212_, _000236_);
  and g_094106_(_000227_, _000236_, _000237_);
  and g_094107_(_000235_, _000237_, _000238_);
  or g_094108_(out[721], out[722], _000239_);
  xor g_094109_(out[721], out[722], _000240_);
  xor g_094110_(_000417_, out[722], _000242_);
  or g_094111_(_000146_, _000196_, _000243_);
  or g_094112_(_000141_, _000198_, _000244_);
  and g_094113_(_000243_, _000244_, _000245_);
  and g_094114_(_000242_, _000245_, _000246_);
  xor g_094115_(out[723], _023825_, _000247_);
  or g_094116_(_000137_, _000196_, _000248_);
  or g_094117_(_000132_, _000198_, _000249_);
  and g_094118_(_000248_, _000249_, _000250_);
  not g_094119_(_000250_, _000251_);
  and g_094120_(_000247_, _000251_, _000253_);
  or g_094121_(_000246_, _000253_, _000254_);
  or g_094122_(_000285_, _000198_, _000255_);
  or g_094123_(_000155_, _000196_, _000256_);
  and g_094124_(_000255_, _000256_, _000257_);
  and g_094125_(out[721], _000257_, _000258_);
  and g_094126_(out[704], _000196_, _000259_);
  not g_094127_(_000259_, _000260_);
  or g_094128_(_000162_, _000196_, _000261_);
  not g_094129_(_000261_, _000262_);
  or g_094130_(_000259_, _000262_, _000264_);
  and g_094131_(_000260_, _000261_, _000265_);
  or g_094132_(_000428_, _000264_, _000266_);
  xor g_094133_(out[721], _000257_, _000267_);
  and g_094134_(_000266_, _000267_, _000268_);
  or g_094135_(_000258_, _000268_, _000269_);
  xor g_094136_(_000242_, _000245_, _000270_);
  xor g_094137_(out[726], _023869_, _000271_);
  or g_094138_(_000079_, _000196_, _000272_);
  not g_094139_(_000272_, _000273_);
  and g_094140_(_000073_, _000196_, _000275_);
  or g_094141_(_000072_, _000198_, _000276_);
  and g_094142_(_000272_, _000276_, _000277_);
  or g_094143_(_000273_, _000275_, _000278_);
  or g_094144_(_000271_, _000278_, _000279_);
  xor g_094145_(out[727], _023880_, _000280_);
  xor g_094146_(_000373_, _023880_, _000281_);
  or g_094147_(_000090_, _000196_, _000282_);
  or g_094148_(_000084_, _000198_, _000283_);
  and g_094149_(_000282_, _000283_, _000284_);
  or g_094150_(_000280_, _000284_, _000286_);
  and g_094151_(_000279_, _000286_, _000287_);
  and g_094152_(_000280_, _000284_, _000288_);
  xor g_094153_(_000271_, _000278_, _000289_);
  xor g_094154_(_000271_, _000277_, _000290_);
  xor g_094155_(_000280_, _000284_, _000291_);
  xor g_094156_(_000281_, _000284_, _000292_);
  and g_094157_(_000289_, _000291_, _000293_);
  or g_094158_(_000290_, _000292_, _000294_);
  xor g_094159_(out[724], _023847_, _000295_);
  not g_094160_(_000295_, _000297_);
  and g_094161_(_000110_, _000198_, _000298_);
  or g_094162_(_000108_, _000196_, _000299_);
  and g_094163_(_000103_, _000196_, _000300_);
  not g_094164_(_000300_, _000301_);
  and g_094165_(_000299_, _000301_, _000302_);
  or g_094166_(_000298_, _000300_, _000303_);
  or g_094167_(_000297_, _000303_, _000304_);
  xor g_094168_(_000395_, _023858_, _000305_);
  or g_094169_(_000117_, _000196_, _000306_);
  or g_094170_(_000112_, _000198_, _000308_);
  and g_094171_(_000306_, _000308_, _000309_);
  or g_094172_(_000305_, _000309_, _000310_);
  and g_094173_(_000304_, _000310_, _000311_);
  and g_094174_(_000305_, _000309_, _000312_);
  xor g_094175_(_000295_, _000302_, _000313_);
  xor g_094176_(_000305_, _000309_, _000314_);
  and g_094177_(_000293_, _000314_, _000315_);
  and g_094178_(_000313_, _000315_, _000316_);
  or g_094179_(_000247_, _000251_, _000317_);
  xor g_094180_(_000247_, _000251_, _000319_);
  and g_094181_(_000270_, _000319_, _000320_);
  and g_094182_(_000269_, _000320_, _000321_);
  and g_094183_(_000254_, _000317_, _000322_);
  or g_094184_(_000321_, _000322_, _000323_);
  and g_094185_(_000316_, _000323_, _000324_);
  or g_094186_(_000294_, _000311_, _000325_);
  or g_094187_(_000312_, _000325_, _000326_);
  or g_094188_(_000287_, _000288_, _000327_);
  and g_094189_(_000326_, _000327_, _000328_);
  not g_094190_(_000328_, _000330_);
  or g_094191_(_000324_, _000330_, _000331_);
  and g_094192_(_000238_, _000331_, _000332_);
  and g_094193_(_000209_, _000210_, _000333_);
  and g_094194_(_000234_, _000236_, _000334_);
  and g_094195_(_000221_, _000334_, _000335_);
  or g_094196_(_000333_, _000335_, _000336_);
  or g_094197_(_000332_, _000336_, _000337_);
  or g_094198_(out[720], _000265_, _000338_);
  and g_094199_(_000268_, _000338_, _000339_);
  and g_094200_(_000320_, _000339_, _000341_);
  and g_094201_(_000316_, _000341_, _000342_);
  and g_094202_(_000238_, _000342_, _000343_);
  not g_094203_(_000343_, _000344_);
  and g_094204_(_000337_, _000344_, _000345_);
  not g_094205_(_000345_, _000346_);
  and g_094206_(_053983_, _000345_, _000347_);
  not g_094207_(_000347_, _000348_);
  and g_094208_(_000204_, _000346_, _000349_);
  or g_094209_(_000203_, _000345_, _000350_);
  and g_094210_(_000348_, _000350_, _000352_);
  or g_094211_(_000347_, _000349_, _000353_);
  xor g_094212_(out[739], _023979_, _000354_);
  xor g_094213_(_000582_, _023979_, _000355_);
  or g_094214_(_000247_, _000346_, _000356_);
  or g_094215_(_000250_, _000345_, _000357_);
  and g_094216_(_000356_, _000357_, _000358_);
  not g_094217_(_000358_, _000359_);
  and g_094218_(_000354_, _000359_, _000360_);
  or g_094219_(out[737], out[738], _000361_);
  xor g_094220_(_000549_, out[738], _000363_);
  or g_094221_(_000245_, _000345_, _000364_);
  or g_094222_(_000240_, _000346_, _000365_);
  and g_094223_(_000364_, _000365_, _000366_);
  and g_094224_(_000363_, _000366_, _000367_);
  or g_094225_(_000360_, _000367_, _000368_);
  or g_094226_(_000354_, _000359_, _000369_);
  xor g_094227_(_000355_, _000358_, _000370_);
  xor g_094228_(_000363_, _000366_, _000371_);
  and g_094229_(_000370_, _000371_, _000372_);
  or g_094230_(_000417_, _000346_, _000374_);
  or g_094231_(_000257_, _000345_, _000375_);
  and g_094232_(_000374_, _000375_, _000376_);
  and g_094233_(out[737], _000376_, _000377_);
  and g_094234_(_000265_, _000346_, _000378_);
  and g_094235_(_000428_, _000345_, _000379_);
  or g_094236_(_000378_, _000379_, _000380_);
  and g_094237_(out[736], _000380_, _000381_);
  not g_094238_(_000381_, _000382_);
  xor g_094239_(out[737], _000376_, _000383_);
  xor g_094240_(_000549_, _000376_, _000385_);
  and g_094241_(_000382_, _000383_, _000386_);
  or g_094242_(_000381_, _000385_, _000387_);
  or g_094243_(_000377_, _000386_, _000388_);
  and g_094244_(_000372_, _000388_, _000389_);
  and g_094245_(_000368_, _000369_, _000390_);
  or g_094246_(_000389_, _000390_, _000391_);
  not g_094247_(_000391_, _000392_);
  and g_094248_(_023957_, _024100_, _000393_);
  or g_094249_(_023968_, _024089_, _000394_);
  xor g_094250_(out[746], _024067_, _000396_);
  xor g_094251_(_000615_, _024067_, _000397_);
  and g_094252_(_000352_, _000396_, _000398_);
  or g_094253_(_000353_, _000397_, _000399_);
  and g_094254_(_000394_, _000399_, _000400_);
  or g_094255_(_000393_, _000398_, _000401_);
  and g_094256_(_000353_, _000397_, _000402_);
  or g_094257_(_000352_, _000396_, _000403_);
  or g_094258_(_000216_, _000345_, _000404_);
  or g_094259_(_000218_, _000346_, _000405_);
  and g_094260_(_000404_, _000405_, _000407_);
  not g_094261_(_000407_, _000408_);
  xor g_094262_(out[745], _024056_, _000409_);
  xor g_094263_(_000604_, _024056_, _000410_);
  and g_094264_(_000407_, _000410_, _000411_);
  or g_094265_(_000408_, _000409_, _000412_);
  and g_094266_(_023968_, _024089_, _000413_);
  or g_094267_(_023957_, _024100_, _000414_);
  xor g_094268_(out[744], _024045_, _000415_);
  or g_094269_(_000226_, _000345_, _000416_);
  and g_094270_(_000222_, _000345_, _000418_);
  not g_094271_(_000418_, _000419_);
  and g_094272_(_000416_, _000419_, _000420_);
  and g_094273_(_000415_, _000420_, _000421_);
  not g_094274_(_000421_, _000422_);
  or g_094275_(_000407_, _000410_, _000423_);
  not g_094276_(_000423_, _000424_);
  and g_094277_(_000422_, _000423_, _000425_);
  or g_094278_(_000421_, _000424_, _000426_);
  or g_094279_(_000415_, _000420_, _000427_);
  not g_094280_(_000427_, _000429_);
  and g_094281_(_000412_, _000425_, _000430_);
  or g_094282_(_000411_, _000426_, _000431_);
  and g_094283_(_000403_, _000414_, _000432_);
  or g_094284_(_000402_, _000413_, _000433_);
  and g_094285_(_000400_, _000432_, _000434_);
  or g_094286_(_000401_, _000433_, _000435_);
  and g_094287_(_000427_, _000434_, _000436_);
  or g_094288_(_000429_, _000435_, _000437_);
  and g_094289_(_000430_, _000436_, _000438_);
  or g_094290_(_000431_, _000437_, _000440_);
  xor g_094291_(out[743], _024034_, _000441_);
  not g_094292_(_000441_, _000442_);
  and g_094293_(_000284_, _000346_, _000443_);
  and g_094294_(_000281_, _000345_, _000444_);
  or g_094295_(_000443_, _000444_, _000445_);
  or g_094296_(_000441_, _000445_, _000446_);
  xor g_094297_(out[742], _024023_, _000447_);
  not g_094298_(_000447_, _000448_);
  or g_094299_(_000277_, _000345_, _000449_);
  or g_094300_(_000271_, _000346_, _000451_);
  and g_094301_(_000449_, _000451_, _000452_);
  not g_094302_(_000452_, _000453_);
  or g_094303_(_000447_, _000453_, _000454_);
  and g_094304_(_000446_, _000454_, _000455_);
  and g_094305_(_000441_, _000445_, _000456_);
  xor g_094306_(_000448_, _000452_, _000457_);
  xor g_094307_(_000447_, _000452_, _000458_);
  xor g_094308_(_000441_, _000445_, _000459_);
  xor g_094309_(_000442_, _000445_, _000460_);
  and g_094310_(_000457_, _000459_, _000462_);
  or g_094311_(_000458_, _000460_, _000463_);
  xor g_094312_(out[740], _024001_, _000464_);
  or g_094313_(_000297_, _000346_, _000465_);
  or g_094314_(_000302_, _000345_, _000466_);
  and g_094315_(_000465_, _000466_, _000467_);
  and g_094316_(_000464_, _000467_, _000468_);
  not g_094317_(_000468_, _000469_);
  xor g_094318_(out[741], _024012_, _000470_);
  xor g_094319_(_000527_, _024012_, _000471_);
  or g_094320_(_000309_, _000345_, _000473_);
  not g_094321_(_000473_, _000474_);
  and g_094322_(_000305_, _000345_, _000475_);
  not g_094323_(_000475_, _000476_);
  and g_094324_(_000473_, _000476_, _000477_);
  or g_094325_(_000474_, _000475_, _000478_);
  and g_094326_(_000470_, _000478_, _000479_);
  or g_094327_(_000471_, _000477_, _000480_);
  and g_094328_(_000469_, _000480_, _000481_);
  or g_094329_(_000468_, _000479_, _000482_);
  and g_094330_(_000471_, _000477_, _000484_);
  or g_094331_(_000470_, _000478_, _000485_);
  or g_094332_(_000464_, _000467_, _000486_);
  and g_094333_(_000485_, _000486_, _000487_);
  not g_094334_(_000487_, _000488_);
  and g_094335_(_000481_, _000487_, _000489_);
  or g_094336_(_000482_, _000488_, _000490_);
  and g_094337_(_000462_, _000489_, _000491_);
  or g_094338_(_000463_, _000490_, _000492_);
  and g_094339_(_000438_, _000491_, _000493_);
  or g_094340_(_000440_, _000492_, _000495_);
  and g_094341_(_000391_, _000493_, _000496_);
  or g_094342_(_000392_, _000495_, _000497_);
  or g_094343_(_000455_, _000456_, _000498_);
  not g_094344_(_000498_, _000499_);
  and g_094345_(_000462_, _000482_, _000500_);
  or g_094346_(_000463_, _000481_, _000501_);
  and g_094347_(_000485_, _000500_, _000502_);
  or g_094348_(_000484_, _000501_, _000503_);
  and g_094349_(_000498_, _000503_, _000504_);
  or g_094350_(_000499_, _000502_, _000506_);
  and g_094351_(_000438_, _000506_, _000507_);
  or g_094352_(_000440_, _000504_, _000508_);
  and g_094353_(_000426_, _000434_, _000509_);
  or g_094354_(_000425_, _000435_, _000510_);
  and g_094355_(_000412_, _000509_, _000511_);
  or g_094356_(_000411_, _000510_, _000512_);
  and g_094357_(_000401_, _000414_, _000513_);
  or g_094358_(_000400_, _000413_, _000514_);
  and g_094359_(_000512_, _000514_, _000515_);
  or g_094360_(_000511_, _000513_, _000517_);
  and g_094361_(_000508_, _000515_, _000518_);
  or g_094362_(_000507_, _000517_, _000519_);
  and g_094363_(_000497_, _000518_, _000520_);
  or g_094364_(_000496_, _000519_, _000521_);
  or g_094365_(out[736], _000380_, _000522_);
  and g_094366_(_000372_, _000522_, _000523_);
  not g_094367_(_000523_, _000524_);
  and g_094368_(_000386_, _000523_, _000525_);
  or g_094369_(_000387_, _000524_, _000526_);
  and g_094370_(_000493_, _000525_, _000528_);
  or g_094371_(_000495_, _000526_, _000529_);
  and g_094372_(_000521_, _000529_, _000530_);
  or g_094373_(_000520_, _000528_, _000531_);
  and g_094374_(_000353_, _000531_, _000532_);
  or g_094375_(_000352_, _000530_, _000533_);
  and g_094376_(_000396_, _000530_, _000534_);
  or g_094377_(_000397_, _000531_, _000535_);
  and g_094378_(_000533_, _000535_, _000536_);
  or g_094379_(_000532_, _000534_, _000537_);
  and g_094380_(_024111_, _024254_, _000539_);
  or g_094381_(_024122_, _024243_, _000540_);
  xor g_094382_(out[762], _024221_, _000541_);
  xor g_094383_(_000747_, _024221_, _000542_);
  and g_094384_(_000536_, _000541_, _000543_);
  or g_094385_(_000537_, _000542_, _000544_);
  and g_094386_(_000540_, _000544_, _000545_);
  or g_094387_(_000539_, _000543_, _000546_);
  and g_094388_(_000537_, _000542_, _000547_);
  or g_094389_(_000536_, _000541_, _000548_);
  and g_094390_(_024122_, _024243_, _000550_);
  or g_094391_(_024111_, _024254_, _000551_);
  and g_094392_(_000548_, _000551_, _000552_);
  or g_094393_(_000547_, _000550_, _000553_);
  and g_094394_(_000545_, _000552_, _000554_);
  or g_094395_(_000546_, _000553_, _000555_);
  and g_094396_(_000410_, _000530_, _000556_);
  not g_094397_(_000556_, _000557_);
  or g_094398_(_000407_, _000530_, _000558_);
  not g_094399_(_000558_, _000559_);
  and g_094400_(_000557_, _000558_, _000561_);
  or g_094401_(_000556_, _000559_, _000562_);
  xor g_094402_(out[761], _024210_, _000563_);
  not g_094403_(_000563_, _000564_);
  and g_094404_(_000562_, _000563_, _000565_);
  or g_094405_(_000561_, _000564_, _000566_);
  xor g_094406_(out[760], _024199_, _000567_);
  xor g_094407_(_000725_, _024199_, _000568_);
  and g_094408_(_000415_, _000530_, _000569_);
  not g_094409_(_000569_, _000570_);
  or g_094410_(_000420_, _000530_, _000572_);
  not g_094411_(_000572_, _000573_);
  and g_094412_(_000570_, _000572_, _000574_);
  or g_094413_(_000569_, _000573_, _000575_);
  and g_094414_(_000567_, _000574_, _000576_);
  or g_094415_(_000568_, _000575_, _000577_);
  and g_094416_(_000566_, _000577_, _000578_);
  or g_094417_(_000565_, _000576_, _000579_);
  and g_094418_(_000568_, _000575_, _000580_);
  or g_094419_(_000567_, _000574_, _000581_);
  and g_094420_(_000561_, _000564_, _000583_);
  or g_094421_(_000562_, _000563_, _000584_);
  and g_094422_(_000581_, _000584_, _000585_);
  or g_094423_(_000580_, _000583_, _000586_);
  and g_094424_(_000578_, _000585_, _000587_);
  or g_094425_(_000579_, _000586_, _000588_);
  and g_094426_(_000554_, _000587_, _000589_);
  or g_094427_(_000555_, _000588_, _000590_);
  xor g_094428_(out[758], _024177_, _000591_);
  not g_094429_(_000591_, _000592_);
  and g_094430_(_000448_, _000530_, _000594_);
  not g_094431_(_000594_, _000595_);
  or g_094432_(_000452_, _000530_, _000596_);
  not g_094433_(_000596_, _000597_);
  and g_094434_(_000595_, _000596_, _000598_);
  or g_094435_(_000594_, _000597_, _000599_);
  and g_094436_(_000592_, _000598_, _000600_);
  xor g_094437_(out[759], _024188_, _000601_);
  xor g_094438_(_000637_, _024188_, _000602_);
  and g_094439_(_000441_, _000530_, _000603_);
  or g_094440_(_000445_, _000530_, _000605_);
  not g_094441_(_000605_, _000606_);
  or g_094442_(_000603_, _000606_, _000607_);
  and g_094443_(_000602_, _000607_, _000608_);
  or g_094444_(_000600_, _000608_, _000609_);
  or g_094445_(_000602_, _000607_, _000610_);
  xor g_094446_(_000602_, _000607_, _000611_);
  xor g_094447_(_000601_, _000607_, _000612_);
  xor g_094448_(_000592_, _000598_, _000613_);
  xor g_094449_(_000591_, _000598_, _000614_);
  and g_094450_(_000611_, _000613_, _000616_);
  or g_094451_(_000612_, _000614_, _000617_);
  xor g_094452_(out[757], _024166_, _000618_);
  not g_094453_(_000618_, _000619_);
  and g_094454_(_000471_, _000530_, _000620_);
  and g_094455_(_000478_, _000531_, _000621_);
  or g_094456_(_000620_, _000621_, _000622_);
  or g_094457_(_000618_, _000622_, _000623_);
  xor g_094458_(out[756], _024155_, _000624_);
  xor g_094459_(_000670_, _024155_, _000625_);
  and g_094460_(_000464_, _000530_, _000627_);
  not g_094461_(_000627_, _000628_);
  or g_094462_(_000467_, _000530_, _000629_);
  not g_094463_(_000629_, _000630_);
  and g_094464_(_000628_, _000629_, _000631_);
  or g_094465_(_000627_, _000630_, _000632_);
  and g_094466_(_000624_, _000631_, _000633_);
  or g_094467_(_000625_, _000632_, _000634_);
  and g_094468_(_000618_, _000622_, _000635_);
  and g_094469_(_000625_, _000632_, _000636_);
  not g_094470_(_000636_, _000638_);
  xor g_094471_(_000618_, _000622_, _000639_);
  xor g_094472_(_000619_, _000622_, _000640_);
  and g_094473_(_000634_, _000639_, _000641_);
  or g_094474_(_000633_, _000640_, _000642_);
  and g_094475_(_000638_, _000641_, _000643_);
  or g_094476_(_000636_, _000642_, _000644_);
  and g_094477_(_000616_, _000643_, _000645_);
  or g_094478_(_000617_, _000644_, _000646_);
  and g_094479_(_000589_, _000645_, _000647_);
  or g_094480_(_000590_, _000646_, _000649_);
  or g_094481_(out[753], out[754], _000650_);
  xor g_094482_(out[753], out[754], _000651_);
  xor g_094483_(_000681_, out[754], _000652_);
  and g_094484_(_000363_, _000530_, _000653_);
  or g_094485_(_000366_, _000530_, _000654_);
  not g_094486_(_000654_, _000655_);
  or g_094487_(_000653_, _000655_, _000656_);
  not g_094488_(_000656_, _000657_);
  and g_094489_(_000652_, _000657_, _000658_);
  xor g_094490_(_000652_, _000656_, _000660_);
  xor g_094491_(out[755], _024133_, _000661_);
  and g_094492_(_000359_, _000531_, _000662_);
  and g_094493_(_000355_, _000530_, _000663_);
  or g_094494_(_000662_, _000663_, _000664_);
  not g_094495_(_000664_, _000665_);
  or g_094496_(_000661_, _000664_, _000666_);
  and g_094497_(_000661_, _000664_, _000667_);
  xor g_094498_(_000661_, _000665_, _000668_);
  or g_094499_(_000660_, _000668_, _000669_);
  or g_094500_(_000649_, _000669_, _000671_);
  not g_094501_(_000671_, _000672_);
  and g_094502_(out[737], _000530_, _000673_);
  or g_094503_(_000376_, _000530_, _000674_);
  not g_094504_(_000674_, _000675_);
  or g_094505_(_000673_, _000675_, _000676_);
  not g_094506_(_000676_, _000677_);
  and g_094507_(out[753], _000677_, _000678_);
  or g_094508_(_000681_, _000676_, _000679_);
  and g_094509_(_000672_, _000678_, _000680_);
  or g_094510_(_000671_, _000679_, _000682_);
  and g_094511_(_000609_, _000610_, _000683_);
  or g_094512_(_000633_, _000635_, _000684_);
  and g_094513_(_000616_, _000684_, _000685_);
  and g_094514_(_000623_, _000685_, _000686_);
  or g_094515_(_000683_, _000686_, _000687_);
  not g_094516_(_000687_, _000688_);
  and g_094517_(_000589_, _000687_, _000689_);
  or g_094518_(_000590_, _000688_, _000690_);
  or g_094519_(_000658_, _000667_, _000691_);
  and g_094520_(_000666_, _000691_, _000693_);
  not g_094521_(_000693_, _000694_);
  and g_094522_(_000647_, _000693_, _000695_);
  or g_094523_(_000649_, _000694_, _000696_);
  and g_094524_(_000554_, _000579_, _000697_);
  or g_094525_(_000555_, _000578_, _000698_);
  and g_094526_(_000584_, _000697_, _000699_);
  or g_094527_(_000583_, _000698_, _000700_);
  and g_094528_(_000546_, _000551_, _000701_);
  or g_094529_(_000545_, _000550_, _000702_);
  and g_094530_(_000700_, _000702_, _000704_);
  or g_094531_(_000699_, _000701_, _000705_);
  and g_094532_(_000696_, _000704_, _000706_);
  or g_094533_(_000695_, _000705_, _000707_);
  and g_094534_(_000690_, _000706_, _000708_);
  or g_094535_(_000689_, _000707_, _000709_);
  and g_094536_(_000682_, _000708_, _000710_);
  or g_094537_(_000680_, _000709_, _000711_);
  and g_094538_(_000380_, _000531_, _000712_);
  and g_094539_(_000560_, _000530_, _000713_);
  or g_094540_(_000712_, _000713_, _000715_);
  not g_094541_(_000715_, _000716_);
  and g_094542_(out[752], _000715_, _000717_);
  xor g_094543_(out[753], _000676_, _000718_);
  or g_094544_(_000717_, _000718_, _000719_);
  or g_094545_(_000671_, _000719_, _000720_);
  or g_094546_(out[752], _000715_, _000721_);
  or g_094547_(_000720_, _000721_, _000722_);
  not g_094548_(_000722_, _000723_);
  and g_094549_(_000710_, _000722_, _000724_);
  or g_094550_(_000711_, _000723_, _000726_);
  and g_094551_(_000537_, _000724_, _000727_);
  or g_094552_(_000536_, _000726_, _000728_);
  or g_094553_(_000542_, _000724_, _000729_);
  not g_094554_(_000729_, _000730_);
  and g_094555_(_000728_, _000729_, _000731_);
  or g_094556_(_000727_, _000730_, _000732_);
  xor g_094557_(out[775], _024342_, _000733_);
  xor g_094558_(_000769_, _024342_, _000734_);
  and g_094559_(_000607_, _000724_, _000735_);
  and g_094560_(_000601_, _000726_, _000737_);
  or g_094561_(_000735_, _000737_, _000738_);
  not g_094562_(_000738_, _000739_);
  and g_094563_(_000733_, _000739_, _000740_);
  or g_094564_(_000733_, _000739_, _000741_);
  xor g_094565_(_000734_, _000738_, _000742_);
  xor g_094566_(_000733_, _000738_, _000743_);
  xor g_094567_(out[773], _024320_, _000744_);
  and g_094568_(_000619_, _000726_, _000745_);
  and g_094569_(_000622_, _000724_, _000746_);
  or g_094570_(_000745_, _000746_, _000748_);
  or g_094571_(_000744_, _000748_, _000749_);
  xor g_094572_(out[774], _024331_, _000750_);
  and g_094573_(_000592_, _000726_, _000751_);
  and g_094574_(_000599_, _000724_, _000752_);
  or g_094575_(_000751_, _000752_, _000753_);
  or g_094576_(_000750_, _000753_, _000754_);
  xor g_094577_(_000750_, _000753_, _000755_);
  and g_094578_(_000749_, _000755_, _000756_);
  not g_094579_(_000756_, _000757_);
  and g_094580_(_000742_, _000756_, _000759_);
  or g_094581_(_000743_, _000757_, _000760_);
  and g_094582_(_024265_, _024408_, _000761_);
  or g_094583_(_024276_, _024397_, _000762_);
  xor g_094584_(out[778], _024375_, _000763_);
  xor g_094585_(_000879_, _024375_, _000764_);
  and g_094586_(_000731_, _000763_, _000765_);
  or g_094587_(_000732_, _000764_, _000766_);
  and g_094588_(_000762_, _000766_, _000767_);
  or g_094589_(_000761_, _000765_, _000768_);
  and g_094590_(_000732_, _000764_, _000770_);
  not g_094591_(_000770_, _000771_);
  and g_094592_(_024276_, _024397_, _000772_);
  or g_094593_(_024265_, _024408_, _000773_);
  and g_094594_(_000767_, _000773_, _000774_);
  or g_094595_(_000768_, _000772_, _000775_);
  and g_094596_(_000771_, _000774_, _000776_);
  or g_094597_(_000770_, _000775_, _000777_);
  or g_094598_(_000563_, _000724_, _000778_);
  not g_094599_(_000778_, _000779_);
  and g_094600_(_000562_, _000724_, _000781_);
  not g_094601_(_000781_, _000782_);
  and g_094602_(_000778_, _000782_, _000783_);
  or g_094603_(_000779_, _000781_, _000784_);
  xor g_094604_(out[777], _024364_, _000785_);
  not g_094605_(_000785_, _000786_);
  and g_094606_(_000784_, _000785_, _000787_);
  not g_094607_(_000787_, _000788_);
  xor g_094608_(out[776], _024353_, _000789_);
  xor g_094609_(_000857_, _024353_, _000790_);
  or g_094610_(_000568_, _000724_, _000792_);
  not g_094611_(_000792_, _000793_);
  and g_094612_(_000575_, _000724_, _000794_);
  not g_094613_(_000794_, _000795_);
  and g_094614_(_000792_, _000795_, _000796_);
  or g_094615_(_000793_, _000794_, _000797_);
  and g_094616_(_000789_, _000796_, _000798_);
  or g_094617_(_000790_, _000797_, _000799_);
  and g_094618_(_000788_, _000799_, _000800_);
  or g_094619_(_000787_, _000798_, _000801_);
  and g_094620_(_000783_, _000786_, _000803_);
  or g_094621_(_000784_, _000785_, _000804_);
  and g_094622_(_000790_, _000797_, _000805_);
  not g_094623_(_000805_, _000806_);
  and g_094624_(_000804_, _000806_, _000807_);
  or g_094625_(_000803_, _000805_, _000808_);
  and g_094626_(_000800_, _000807_, _000809_);
  or g_094627_(_000801_, _000808_, _000810_);
  and g_094628_(_000776_, _000809_, _000811_);
  or g_094629_(_000777_, _000810_, _000812_);
  xor g_094630_(_000802_, _024309_, _000814_);
  and g_094631_(_000632_, _000724_, _000815_);
  and g_094632_(_000624_, _000726_, _000816_);
  or g_094633_(_000815_, _000816_, _000817_);
  and g_094634_(_000814_, _000817_, _000818_);
  and g_094635_(_000744_, _000748_, _000819_);
  or g_094636_(_000814_, _000817_, _000820_);
  not g_094637_(_000820_, _000821_);
  or g_094638_(_000819_, _000821_, _000822_);
  or g_094639_(_000818_, _000822_, _000823_);
  or g_094640_(_000760_, _000823_, _000825_);
  or g_094641_(_000812_, _000825_, _000826_);
  or g_094642_(out[769], out[770], _000827_);
  xor g_094643_(out[769], out[770], _000828_);
  xor g_094644_(_000813_, out[770], _000829_);
  and g_094645_(_000652_, _000726_, _000830_);
  and g_094646_(_000656_, _000724_, _000831_);
  or g_094647_(_000830_, _000831_, _000832_);
  not g_094648_(_000832_, _000833_);
  xor g_094649_(out[771], _024287_, _000834_);
  and g_094650_(_000664_, _000724_, _000836_);
  not g_094651_(_000836_, _000837_);
  or g_094652_(_000661_, _000724_, _000838_);
  not g_094653_(_000838_, _000839_);
  and g_094654_(_000837_, _000838_, _000840_);
  or g_094655_(_000836_, _000839_, _000841_);
  or g_094656_(_000834_, _000841_, _000842_);
  and g_094657_(_000829_, _000833_, _000843_);
  and g_094658_(_000834_, _000841_, _000844_);
  or g_094659_(_000843_, _000844_, _000845_);
  xor g_094660_(_000834_, _000840_, _000847_);
  xor g_094661_(_000829_, _000832_, _000848_);
  or g_094662_(_000826_, _000847_, _000849_);
  or g_094663_(_000848_, _000849_, _000850_);
  or g_094664_(_000677_, _000726_, _000851_);
  or g_094665_(_000681_, _000724_, _000852_);
  and g_094666_(_000851_, _000852_, _000853_);
  and g_094667_(out[769], _000853_, _000854_);
  not g_094668_(_000854_, _000855_);
  or g_094669_(_000850_, _000855_, _000856_);
  and g_094670_(_000759_, _000822_, _000858_);
  and g_094671_(_000741_, _000754_, _000859_);
  or g_094672_(_000740_, _000859_, _000860_);
  not g_094673_(_000860_, _000861_);
  or g_094674_(_000858_, _000861_, _000862_);
  and g_094675_(_000811_, _000862_, _000863_);
  not g_094676_(_000863_, _000864_);
  and g_094677_(_000842_, _000845_, _000865_);
  not g_094678_(_000865_, _000866_);
  or g_094679_(_000826_, _000866_, _000867_);
  or g_094680_(_000777_, _000800_, _000869_);
  or g_094681_(_000803_, _000869_, _000870_);
  or g_094682_(_000767_, _000772_, _000871_);
  and g_094683_(_000870_, _000871_, _000872_);
  and g_094684_(_000867_, _000872_, _000873_);
  and g_094685_(_000864_, _000873_, _000874_);
  and g_094686_(_000856_, _000874_, _000875_);
  or g_094687_(_000692_, _000710_, _000876_);
  not g_094688_(_000876_, _000877_);
  and g_094689_(_000716_, _000724_, _000878_);
  or g_094690_(_000877_, _000878_, _000880_);
  not g_094691_(_000880_, _000881_);
  and g_094692_(out[768], _000881_, _000882_);
  xor g_094693_(_000813_, _000853_, _000883_);
  or g_094694_(_000882_, _000883_, _000884_);
  or g_094695_(_000850_, _000884_, _000885_);
  or g_094696_(out[768], _000881_, _000886_);
  or g_094697_(_000885_, _000886_, _000887_);
  and g_094698_(_000875_, _000887_, _000888_);
  not g_094699_(_000888_, _000889_);
  and g_094700_(_000732_, _000888_, _000891_);
  not g_094701_(_000891_, _000892_);
  or g_094702_(_000764_, _000888_, _000893_);
  not g_094703_(_000893_, _000894_);
  and g_094704_(_000892_, _000893_, _000895_);
  or g_094705_(_000891_, _000894_, _000896_);
  and g_094706_(_053982_, _000896_, _000897_);
  or g_094707_(_053981_, _000895_, _000898_);
  or g_094708_(_000785_, _000888_, _000899_);
  or g_094709_(_000783_, _000889_, _000900_);
  and g_094710_(_000899_, _000900_, _000902_);
  xor g_094711_(_001000_, _024518_, _000903_);
  and g_094712_(_000902_, _000903_, _000904_);
  not g_094713_(_000904_, _000905_);
  and g_094714_(_000898_, _000905_, _000906_);
  or g_094715_(_000897_, _000904_, _000907_);
  and g_094716_(_024430_, _024551_, _000908_);
  or g_094717_(_024419_, _024562_, _000909_);
  xor g_094718_(out[792], _024507_, _000910_);
  or g_094719_(_000790_, _000888_, _000911_);
  or g_094720_(_000796_, _000889_, _000913_);
  and g_094721_(_000911_, _000913_, _000914_);
  or g_094722_(_000910_, _000914_, _000915_);
  not g_094723_(_000915_, _000916_);
  and g_094724_(_000909_, _000915_, _000917_);
  or g_094725_(_000908_, _000916_, _000918_);
  and g_094726_(_000906_, _000917_, _000919_);
  or g_094727_(_000907_, _000918_, _000920_);
  and g_094728_(_024419_, _024562_, _000921_);
  or g_094729_(_024430_, _024551_, _000922_);
  and g_094730_(_053981_, _000895_, _000924_);
  or g_094731_(_053982_, _000896_, _000925_);
  and g_094732_(_000922_, _000925_, _000926_);
  or g_094733_(_000921_, _000924_, _000927_);
  and g_094734_(_000910_, _000914_, _000928_);
  not g_094735_(_000928_, _000929_);
  or g_094736_(_000902_, _000903_, _000930_);
  not g_094737_(_000930_, _000931_);
  and g_094738_(_000929_, _000930_, _000932_);
  or g_094739_(_000928_, _000931_, _000933_);
  and g_094740_(_000926_, _000932_, _000935_);
  or g_094741_(_000927_, _000933_, _000936_);
  and g_094742_(_000919_, _000935_, _000937_);
  or g_094743_(_000920_, _000936_, _000938_);
  xor g_094744_(out[790], _024485_, _000939_);
  xor g_094745_(_000912_, _024485_, _000940_);
  or g_094746_(_000750_, _000888_, _000941_);
  not g_094747_(_000941_, _000942_);
  and g_094748_(_000753_, _000888_, _000943_);
  not g_094749_(_000943_, _000944_);
  and g_094750_(_000941_, _000944_, _000946_);
  or g_094751_(_000942_, _000943_, _000947_);
  and g_094752_(_000940_, _000946_, _000948_);
  or g_094753_(_000939_, _000947_, _000949_);
  xor g_094754_(out[791], _024496_, _000950_);
  not g_094755_(_000950_, _000951_);
  or g_094756_(_000734_, _000888_, _000952_);
  not g_094757_(_000952_, _000953_);
  and g_094758_(_000738_, _000888_, _000954_);
  not g_094759_(_000954_, _000955_);
  and g_094760_(_000952_, _000955_, _000957_);
  or g_094761_(_000953_, _000954_, _000958_);
  and g_094762_(_000951_, _000958_, _000959_);
  or g_094763_(_000950_, _000957_, _000960_);
  and g_094764_(_000949_, _000960_, _000961_);
  or g_094765_(_000948_, _000959_, _000962_);
  and g_094766_(_000950_, _000957_, _000963_);
  not g_094767_(_000963_, _000964_);
  or g_094768_(_000940_, _000946_, _000965_);
  not g_094769_(_000965_, _000966_);
  and g_094770_(_000961_, _000965_, _000968_);
  or g_094771_(_000962_, _000966_, _000969_);
  and g_094772_(_000964_, _000968_, _000970_);
  or g_094773_(_000963_, _000969_, _000971_);
  xor g_094774_(out[788], _024463_, _000972_);
  and g_094775_(_000817_, _000888_, _000973_);
  not g_094776_(_000973_, _000974_);
  or g_094777_(_000814_, _000888_, _000975_);
  and g_094778_(_000974_, _000975_, _000976_);
  and g_094779_(_000972_, _000976_, _000977_);
  not g_094780_(_000977_, _000979_);
  xor g_094781_(out[789], _024474_, _000980_);
  xor g_094782_(_000923_, _024474_, _000981_);
  or g_094783_(_000744_, _000888_, _000982_);
  and g_094784_(_000748_, _000888_, _000983_);
  not g_094785_(_000983_, _000984_);
  and g_094786_(_000982_, _000984_, _000985_);
  not g_094787_(_000985_, _000986_);
  or g_094788_(_000981_, _000985_, _000987_);
  not g_094789_(_000987_, _000988_);
  and g_094790_(_000979_, _000987_, _000990_);
  or g_094791_(_000977_, _000988_, _000991_);
  and g_094792_(_000981_, _000985_, _000992_);
  or g_094793_(_000980_, _000986_, _000993_);
  or g_094794_(_000972_, _000976_, _000994_);
  not g_094795_(_000994_, _000995_);
  and g_094796_(_000993_, _000994_, _000996_);
  or g_094797_(_000992_, _000995_, _000997_);
  and g_094798_(_000990_, _000996_, _000998_);
  or g_094799_(_000991_, _000997_, _000999_);
  and g_094800_(_000970_, _000998_, _001001_);
  or g_094801_(_000971_, _000999_, _001002_);
  xor g_094802_(out[787], _024441_, _001003_);
  xor g_094803_(_000978_, _024441_, _001004_);
  or g_094804_(_000840_, _000889_, _001005_);
  or g_094805_(_000834_, _000888_, _001006_);
  and g_094806_(_001005_, _001006_, _001007_);
  or g_094807_(_001004_, _001007_, _001008_);
  or g_094808_(out[785], out[786], _001009_);
  xor g_094809_(out[785], out[786], _001010_);
  xor g_094810_(_000945_, out[786], _001012_);
  or g_094811_(_000828_, _000888_, _001013_);
  or g_094812_(_000833_, _000889_, _001014_);
  and g_094813_(_001013_, _001014_, _001015_);
  not g_094814_(_001015_, _001016_);
  or g_094815_(_001010_, _001016_, _001017_);
  and g_094816_(_001004_, _001007_, _001018_);
  xor g_094817_(_001004_, _001007_, _001019_);
  xor g_094818_(_001003_, _001007_, _001020_);
  xor g_094819_(_001012_, _001015_, _001021_);
  xor g_094820_(_001010_, _001015_, _001023_);
  and g_094821_(_001019_, _001021_, _001024_);
  or g_094822_(_001020_, _001023_, _001025_);
  or g_094823_(_000853_, _000889_, _001026_);
  or g_094824_(_000813_, _000888_, _001027_);
  and g_094825_(_001026_, _001027_, _001028_);
  and g_094826_(out[785], _001028_, _001029_);
  not g_094827_(_001029_, _001030_);
  or g_094828_(_000824_, _000875_, _001031_);
  not g_094829_(_001031_, _001032_);
  and g_094830_(_000880_, _000888_, _001034_);
  not g_094831_(_001034_, _001035_);
  and g_094832_(_001031_, _001035_, _001036_);
  or g_094833_(_001032_, _001034_, _001037_);
  and g_094834_(out[784], _001036_, _001038_);
  or g_094835_(_000956_, _001037_, _001039_);
  xor g_094836_(out[785], _001028_, _001040_);
  xor g_094837_(_000945_, _001028_, _001041_);
  and g_094838_(_001039_, _001040_, _001042_);
  or g_094839_(_001038_, _001041_, _001043_);
  and g_094840_(_001030_, _001043_, _001045_);
  or g_094841_(_001029_, _001042_, _001046_);
  and g_094842_(_001024_, _001046_, _001047_);
  or g_094843_(_001025_, _001045_, _001048_);
  or g_094844_(_001017_, _001018_, _001049_);
  and g_094845_(_001008_, _001049_, _001050_);
  not g_094846_(_001050_, _001051_);
  and g_094847_(_001048_, _001050_, _001052_);
  or g_094848_(_001047_, _001051_, _001053_);
  and g_094849_(_001001_, _001053_, _001054_);
  or g_094850_(_001002_, _001052_, _001056_);
  or g_094851_(_000961_, _000963_, _001057_);
  not g_094852_(_001057_, _001058_);
  and g_094853_(_000991_, _000993_, _001059_);
  or g_094854_(_000990_, _000992_, _001060_);
  and g_094855_(_000970_, _001059_, _001061_);
  or g_094856_(_000971_, _001060_, _001062_);
  and g_094857_(_001057_, _001062_, _001063_);
  or g_094858_(_001058_, _001061_, _001064_);
  and g_094859_(_001056_, _001063_, _001065_);
  or g_094860_(_001054_, _001064_, _001067_);
  and g_094861_(_000937_, _001067_, _001068_);
  or g_094862_(_000938_, _001065_, _001069_);
  and g_094863_(_000906_, _000933_, _001070_);
  or g_094864_(_000907_, _000932_, _001071_);
  and g_094865_(_000926_, _001071_, _001072_);
  or g_094866_(_000927_, _001070_, _001073_);
  and g_094867_(_000909_, _001073_, _001074_);
  or g_094868_(_000908_, _001072_, _001075_);
  and g_094869_(_001069_, _001075_, _001076_);
  or g_094870_(_001068_, _001074_, _001078_);
  or g_094871_(out[784], _001036_, _001079_);
  not g_094872_(_001079_, _001080_);
  or g_094873_(_001043_, _001080_, _001081_);
  not g_094874_(_001081_, _001082_);
  and g_094875_(_001024_, _001082_, _001083_);
  or g_094876_(_001025_, _001081_, _001084_);
  and g_094877_(_000937_, _001083_, _001085_);
  or g_094878_(_000938_, _001084_, _001086_);
  and g_094879_(_001001_, _001085_, _001087_);
  or g_094880_(_001002_, _001086_, _001089_);
  and g_094881_(_001078_, _001089_, _001090_);
  or g_094882_(_001076_, _001087_, _001091_);
  and g_094883_(_053981_, _001090_, _001092_);
  or g_094884_(_053982_, _001091_, _001093_);
  and g_094885_(_000896_, _001091_, _001094_);
  or g_094886_(_000895_, _001090_, _001095_);
  and g_094887_(_001093_, _001095_, _001096_);
  or g_094888_(_001092_, _001094_, _001097_);
  and g_094889_(_000956_, _001090_, _001098_);
  and g_094890_(_001036_, _001091_, _001100_);
  or g_094891_(_001098_, _001100_, _001101_);
  or g_094892_(out[800], _001101_, _001102_);
  not g_094893_(_001102_, _001103_);
  and g_094894_(_024573_, _024716_, _001104_);
  or g_094895_(_024584_, _024705_, _001105_);
  xor g_094896_(out[810], _024683_, _001106_);
  xor g_094897_(_001143_, _024683_, _001107_);
  and g_094898_(_001096_, _001106_, _001108_);
  or g_094899_(_001097_, _001107_, _001109_);
  and g_094900_(_001105_, _001109_, _001111_);
  or g_094901_(_001104_, _001108_, _001112_);
  and g_094902_(_024584_, _024705_, _001113_);
  or g_094903_(_024573_, _024716_, _001114_);
  xor g_094904_(_001121_, _024661_, _001115_);
  or g_094905_(_000914_, _001090_, _001116_);
  not g_094906_(_001116_, _001117_);
  and g_094907_(_000910_, _001090_, _001118_);
  or g_094908_(_001117_, _001118_, _001119_);
  and g_094909_(_001115_, _001119_, _001120_);
  not g_094910_(_001120_, _001122_);
  and g_094911_(_001097_, _001107_, _001123_);
  or g_094912_(_001096_, _001106_, _001124_);
  or g_094913_(_000902_, _001090_, _001125_);
  not g_094914_(_001125_, _001126_);
  and g_094915_(_000903_, _001090_, _001127_);
  not g_094916_(_001127_, _001128_);
  and g_094917_(_001125_, _001128_, _001129_);
  or g_094918_(_001126_, _001127_, _001130_);
  xor g_094919_(out[809], _024672_, _001131_);
  not g_094920_(_001131_, _001133_);
  and g_094921_(_001129_, _001133_, _001134_);
  or g_094922_(_001130_, _001131_, _001135_);
  and g_094923_(_001124_, _001135_, _001136_);
  or g_094924_(_001123_, _001134_, _001137_);
  or g_094925_(_001115_, _001119_, _001138_);
  not g_094926_(_001138_, _001139_);
  and g_094927_(_001130_, _001131_, _001140_);
  not g_094928_(_001140_, _001141_);
  and g_094929_(_001138_, _001141_, _001142_);
  or g_094930_(_001139_, _001140_, _001144_);
  and g_094931_(_001111_, _001114_, _001145_);
  or g_094932_(_001112_, _001113_, _001146_);
  and g_094933_(_001136_, _001145_, _001147_);
  or g_094934_(_001137_, _001146_, _001148_);
  and g_094935_(_001122_, _001147_, _001149_);
  or g_094936_(_001120_, _001148_, _001150_);
  and g_094937_(_001142_, _001149_, _001151_);
  or g_094938_(_001144_, _001150_, _001152_);
  xor g_094939_(out[806], _024639_, _001153_);
  and g_094940_(_000947_, _001091_, _001155_);
  and g_094941_(_000940_, _001090_, _001156_);
  or g_094942_(_001155_, _001156_, _001157_);
  or g_094943_(_001153_, _001157_, _001158_);
  not g_094944_(_001158_, _001159_);
  xor g_094945_(out[807], _024650_, _001160_);
  xor g_094946_(_001033_, _024650_, _001161_);
  and g_094947_(_000958_, _001091_, _001162_);
  and g_094948_(_000950_, _001090_, _001163_);
  or g_094949_(_001162_, _001163_, _001164_);
  not g_094950_(_001164_, _001166_);
  and g_094951_(_001161_, _001164_, _001167_);
  not g_094952_(_001167_, _001168_);
  and g_094953_(_001158_, _001168_, _001169_);
  or g_094954_(_001159_, _001167_, _001170_);
  and g_094955_(_001160_, _001166_, _001171_);
  or g_094956_(_001161_, _001164_, _001172_);
  xor g_094957_(_001066_, _024617_, _001173_);
  and g_094958_(_000972_, _001090_, _001174_);
  or g_094959_(_000976_, _001090_, _001175_);
  not g_094960_(_001175_, _001177_);
  or g_094961_(_001174_, _001177_, _001178_);
  and g_094962_(_001173_, _001178_, _001179_);
  not g_094963_(_001179_, _001180_);
  and g_094964_(_001172_, _001180_, _001181_);
  or g_094965_(_001171_, _001179_, _001182_);
  and g_094966_(_001169_, _001181_, _001183_);
  or g_094967_(_001170_, _001182_, _001184_);
  xor g_094968_(out[805], _024628_, _001185_);
  and g_094969_(_000986_, _001091_, _001186_);
  and g_094970_(_000981_, _001090_, _001188_);
  or g_094971_(_001186_, _001188_, _001189_);
  and g_094972_(_001185_, _001189_, _001190_);
  not g_094973_(_001190_, _001191_);
  or g_094974_(_001173_, _001178_, _001192_);
  not g_094975_(_001192_, _001193_);
  and g_094976_(_001191_, _001192_, _001194_);
  or g_094977_(_001190_, _001193_, _001195_);
  or g_094978_(_001185_, _001189_, _001196_);
  not g_094979_(_001196_, _001197_);
  and g_094980_(_001153_, _001157_, _001199_);
  not g_094981_(_001199_, _001200_);
  and g_094982_(_001196_, _001200_, _001201_);
  or g_094983_(_001197_, _001199_, _001202_);
  and g_094984_(_001194_, _001201_, _001203_);
  or g_094985_(_001195_, _001202_, _001204_);
  and g_094986_(_001183_, _001203_, _001205_);
  or g_094987_(_001184_, _001204_, _001206_);
  and g_094988_(_001151_, _001205_, _001207_);
  or g_094989_(_001152_, _001206_, _001208_);
  or g_094990_(out[801], out[802], _001210_);
  xor g_094991_(out[801], out[802], _001211_);
  xor g_094992_(_001077_, out[802], _001212_);
  or g_094993_(_001015_, _001090_, _001213_);
  not g_094994_(_001213_, _001214_);
  and g_094995_(_001012_, _001090_, _001215_);
  not g_094996_(_001215_, _001216_);
  and g_094997_(_001213_, _001216_, _001217_);
  or g_094998_(_001214_, _001215_, _001218_);
  and g_094999_(_001212_, _001217_, _001219_);
  xor g_095000_(out[803], _024595_, _001221_);
  xor g_095001_(_001110_, _024595_, _001222_);
  and g_095002_(_001004_, _001090_, _001223_);
  not g_095003_(_001223_, _001224_);
  or g_095004_(_001007_, _001090_, _001225_);
  not g_095005_(_001225_, _001226_);
  and g_095006_(_001224_, _001225_, _001227_);
  or g_095007_(_001223_, _001226_, _001228_);
  and g_095008_(_001221_, _001228_, _001229_);
  or g_095009_(_001219_, _001229_, _001230_);
  and g_095010_(_001211_, _001218_, _001232_);
  and g_095011_(_001222_, _001227_, _001233_);
  or g_095012_(_001221_, _001228_, _001234_);
  or g_095013_(_001232_, _001233_, _001235_);
  xor g_095014_(_001212_, _001217_, _001236_);
  xor g_095015_(_001222_, _001227_, _001237_);
  and g_095016_(_001236_, _001237_, _001238_);
  or g_095017_(_001230_, _001235_, _001239_);
  and g_095018_(out[785], _001090_, _001240_);
  not g_095019_(_001240_, _001241_);
  or g_095020_(_001028_, _001090_, _001243_);
  not g_095021_(_001243_, _001244_);
  and g_095022_(_001241_, _001243_, _001245_);
  or g_095023_(_001240_, _001244_, _001246_);
  and g_095024_(out[801], _001245_, _001247_);
  and g_095025_(out[800], _001101_, _001248_);
  not g_095026_(_001248_, _001249_);
  xor g_095027_(out[801], _001245_, _001250_);
  xor g_095028_(_001077_, _001245_, _001251_);
  and g_095029_(_001249_, _001250_, _001252_);
  or g_095030_(_001248_, _001251_, _001254_);
  and g_095031_(_001238_, _001252_, _001255_);
  or g_095032_(_001239_, _001254_, _001256_);
  and g_095033_(_001207_, _001255_, _001257_);
  or g_095034_(_001208_, _001256_, _001258_);
  and g_095035_(_001102_, _001257_, _001259_);
  or g_095036_(_001103_, _001258_, _001260_);
  and g_095037_(_001136_, _001144_, _001261_);
  or g_095038_(_001112_, _001261_, _001262_);
  and g_095039_(_001114_, _001262_, _001263_);
  not g_095040_(_001263_, _001265_);
  and g_095041_(_001195_, _001201_, _001266_);
  or g_095042_(_001170_, _001266_, _001267_);
  and g_095043_(_001172_, _001267_, _001268_);
  and g_095044_(_001151_, _001268_, _001269_);
  not g_095045_(_001269_, _001270_);
  and g_095046_(_001230_, _001234_, _001271_);
  and g_095047_(_001238_, _001247_, _001272_);
  or g_095048_(_001271_, _001272_, _001273_);
  not g_095049_(_001273_, _001274_);
  and g_095050_(_001256_, _001274_, _001276_);
  or g_095051_(_001255_, _001273_, _001277_);
  and g_095052_(_001207_, _001277_, _001278_);
  or g_095053_(_001208_, _001276_, _001279_);
  and g_095054_(_001265_, _001279_, _001280_);
  or g_095055_(_001263_, _001278_, _001281_);
  and g_095056_(_001270_, _001280_, _001282_);
  or g_095057_(_001269_, _001281_, _001283_);
  and g_095058_(_001260_, _001283_, _001284_);
  or g_095059_(_001259_, _001282_, _001285_);
  and g_095060_(_001097_, _001285_, _001287_);
  or g_095061_(_001096_, _001284_, _001288_);
  and g_095062_(_001106_, _001284_, _001289_);
  or g_095063_(_001107_, _001285_, _001290_);
  and g_095064_(_001288_, _001290_, _001291_);
  or g_095065_(_001287_, _001289_, _001292_);
  xor g_095066_(out[820], _024771_, _001293_);
  not g_095067_(_001293_, _001294_);
  or g_095068_(_001173_, _001285_, _001295_);
  and g_095069_(_001178_, _001285_, _001296_);
  not g_095070_(_001296_, _001298_);
  and g_095071_(_001295_, _001298_, _001299_);
  not g_095072_(_001299_, _001300_);
  and g_095073_(_001293_, _001299_, _001301_);
  not g_095074_(_001301_, _001302_);
  xor g_095075_(out[821], _024782_, _001303_);
  xor g_095076_(_001187_, _024782_, _001304_);
  or g_095077_(_001185_, _001285_, _001305_);
  not g_095078_(_001305_, _001306_);
  and g_095079_(_001189_, _001285_, _001307_);
  not g_095080_(_001307_, _001309_);
  and g_095081_(_001305_, _001309_, _001310_);
  or g_095082_(_001306_, _001307_, _001311_);
  and g_095083_(_001303_, _001311_, _001312_);
  or g_095084_(_001304_, _001310_, _001313_);
  and g_095085_(_001302_, _001313_, _001314_);
  or g_095086_(_001301_, _001312_, _001315_);
  and g_095087_(_001101_, _001285_, _001316_);
  not g_095088_(_001316_, _001317_);
  or g_095089_(out[800], _001285_, _001318_);
  not g_095090_(_001318_, _001320_);
  and g_095091_(_001317_, _001318_, _001321_);
  or g_095092_(_001316_, _001320_, _001322_);
  and g_095093_(out[816], _001322_, _001323_);
  or g_095094_(_001220_, _001321_, _001324_);
  or g_095095_(_001077_, _001285_, _001325_);
  not g_095096_(_001325_, _001326_);
  and g_095097_(_001246_, _001285_, _001327_);
  or g_095098_(_001245_, _001284_, _001328_);
  and g_095099_(_001325_, _001328_, _001329_);
  or g_095100_(_001326_, _001327_, _001331_);
  and g_095101_(out[817], _001329_, _001332_);
  or g_095102_(_001209_, _001331_, _001333_);
  xor g_095103_(out[817], _001329_, _001334_);
  xor g_095104_(_001209_, _001329_, _001335_);
  and g_095105_(_001324_, _001334_, _001336_);
  or g_095106_(_001323_, _001335_, _001337_);
  or g_095107_(out[817], out[818], _001338_);
  xor g_095108_(out[817], out[818], _001339_);
  xor g_095109_(_001209_, out[818], _001340_);
  and g_095110_(_001218_, _001285_, _001342_);
  or g_095111_(_001217_, _001284_, _001343_);
  and g_095112_(_001212_, _001284_, _001344_);
  or g_095113_(_001211_, _001285_, _001345_);
  and g_095114_(_001343_, _001345_, _001346_);
  or g_095115_(_001342_, _001344_, _001347_);
  xor g_095116_(out[819], _024749_, _001348_);
  xor g_095117_(_001242_, _024749_, _001349_);
  and g_095118_(_001228_, _001285_, _001350_);
  or g_095119_(_001227_, _001284_, _001351_);
  and g_095120_(_001222_, _001284_, _001353_);
  or g_095121_(_001221_, _001285_, _001354_);
  and g_095122_(_001351_, _001354_, _001355_);
  or g_095123_(_001350_, _001353_, _001356_);
  and g_095124_(_001349_, _001355_, _001357_);
  or g_095125_(_001348_, _001356_, _001358_);
  and g_095126_(_001340_, _001346_, _001359_);
  or g_095127_(_001339_, _001347_, _001360_);
  xor g_095128_(_001340_, _001346_, _001361_);
  xor g_095129_(_001339_, _001346_, _001362_);
  and g_095130_(_001358_, _001361_, _001364_);
  or g_095131_(_001357_, _001362_, _001365_);
  and g_095132_(_001336_, _001364_, _001366_);
  or g_095133_(_001337_, _001365_, _001367_);
  and g_095134_(_001348_, _001356_, _001368_);
  or g_095135_(_001349_, _001355_, _001369_);
  and g_095136_(_001360_, _001369_, _001370_);
  or g_095137_(_001359_, _001368_, _001371_);
  and g_095138_(_001358_, _001371_, _001372_);
  or g_095139_(_001357_, _001370_, _001373_);
  and g_095140_(_001332_, _001364_, _001375_);
  or g_095141_(_001333_, _001365_, _001376_);
  and g_095142_(_001373_, _001376_, _001377_);
  or g_095143_(_001372_, _001375_, _001378_);
  and g_095144_(_001367_, _001377_, _001379_);
  or g_095145_(_001366_, _001378_, _001380_);
  and g_095146_(_001294_, _001300_, _001381_);
  or g_095147_(_001293_, _001299_, _001382_);
  and g_095148_(_001380_, _001382_, _001383_);
  or g_095149_(_001379_, _001381_, _001384_);
  and g_095150_(_001314_, _001384_, _001386_);
  or g_095151_(_001315_, _001383_, _001387_);
  and g_095152_(_024727_, _024870_, _001388_);
  or g_095153_(_024738_, _024859_, _001389_);
  xor g_095154_(out[826], _024837_, _001390_);
  xor g_095155_(_001275_, _024837_, _001391_);
  and g_095156_(_001291_, _001390_, _001392_);
  or g_095157_(_001292_, _001391_, _001393_);
  and g_095158_(_001389_, _001393_, _001394_);
  or g_095159_(_001388_, _001392_, _001395_);
  and g_095160_(_024738_, _024859_, _001397_);
  or g_095161_(_024727_, _024870_, _001398_);
  and g_095162_(_001292_, _001391_, _001399_);
  or g_095163_(_001291_, _001390_, _001400_);
  and g_095164_(_001398_, _001400_, _001401_);
  or g_095165_(_001397_, _001399_, _001402_);
  and g_095166_(_001394_, _001401_, _001403_);
  or g_095167_(_001395_, _001402_, _001404_);
  or g_095168_(_001131_, _001285_, _001405_);
  not g_095169_(_001405_, _001406_);
  and g_095170_(_001130_, _001285_, _001408_);
  not g_095171_(_001408_, _001409_);
  and g_095172_(_001405_, _001409_, _001410_);
  or g_095173_(_001406_, _001408_, _001411_);
  xor g_095174_(out[825], _024826_, _001412_);
  xor g_095175_(_001264_, _024826_, _001413_);
  and g_095176_(_001411_, _001412_, _001414_);
  or g_095177_(_001410_, _001413_, _001415_);
  xor g_095178_(out[824], _024815_, _001416_);
  not g_095179_(_001416_, _001417_);
  or g_095180_(_001115_, _001285_, _001419_);
  not g_095181_(_001419_, _001420_);
  and g_095182_(_001119_, _001285_, _001421_);
  not g_095183_(_001421_, _001422_);
  and g_095184_(_001419_, _001422_, _001423_);
  or g_095185_(_001420_, _001421_, _001424_);
  and g_095186_(_001416_, _001423_, _001425_);
  or g_095187_(_001417_, _001424_, _001426_);
  and g_095188_(_001415_, _001426_, _001427_);
  or g_095189_(_001414_, _001425_, _001428_);
  and g_095190_(_001410_, _001413_, _001430_);
  not g_095191_(_001430_, _001431_);
  or g_095192_(_001416_, _001423_, _001432_);
  not g_095193_(_001432_, _001433_);
  and g_095194_(_001427_, _001431_, _001434_);
  or g_095195_(_001428_, _001430_, _001435_);
  and g_095196_(_001403_, _001434_, _001436_);
  or g_095197_(_001404_, _001435_, _001437_);
  and g_095198_(_001432_, _001436_, _001438_);
  or g_095199_(_001433_, _001437_, _001439_);
  xor g_095200_(_001176_, _024793_, _001441_);
  or g_095201_(_001153_, _001285_, _001442_);
  and g_095202_(_001157_, _001285_, _001443_);
  not g_095203_(_001443_, _001444_);
  and g_095204_(_001442_, _001444_, _001445_);
  and g_095205_(_001441_, _001445_, _001446_);
  not g_095206_(_001446_, _001447_);
  xor g_095207_(out[823], _024804_, _001448_);
  not g_095208_(_001448_, _001449_);
  or g_095209_(_001161_, _001285_, _001450_);
  or g_095210_(_001166_, _001284_, _001452_);
  and g_095211_(_001450_, _001452_, _001453_);
  not g_095212_(_001453_, _001454_);
  or g_095213_(_001448_, _001453_, _001455_);
  not g_095214_(_001455_, _001456_);
  and g_095215_(_001447_, _001455_, _001457_);
  or g_095216_(_001446_, _001456_, _001458_);
  and g_095217_(_001304_, _001310_, _001459_);
  or g_095218_(_001303_, _001311_, _001460_);
  and g_095219_(_001448_, _001453_, _001461_);
  or g_095220_(_001449_, _001454_, _001463_);
  or g_095221_(_001441_, _001445_, _001464_);
  not g_095222_(_001464_, _001465_);
  and g_095223_(_001460_, _001463_, _001466_);
  or g_095224_(_001459_, _001461_, _001467_);
  and g_095225_(_001464_, _001466_, _001468_);
  or g_095226_(_001458_, _001465_, _001469_);
  and g_095227_(_001457_, _001468_, _001470_);
  or g_095228_(_001467_, _001469_, _001471_);
  and g_095229_(_001438_, _001470_, _001472_);
  or g_095230_(_001439_, _001471_, _001474_);
  and g_095231_(_001387_, _001472_, _001475_);
  or g_095232_(_001386_, _001474_, _001476_);
  and g_095233_(_001395_, _001398_, _001477_);
  or g_095234_(_001394_, _001397_, _001478_);
  and g_095235_(_001403_, _001428_, _001479_);
  or g_095236_(_001404_, _001427_, _001480_);
  and g_095237_(_001431_, _001479_, _001481_);
  or g_095238_(_001430_, _001480_, _001482_);
  and g_095239_(_001478_, _001482_, _001483_);
  or g_095240_(_001477_, _001481_, _001485_);
  and g_095241_(_001458_, _001463_, _001486_);
  or g_095242_(_001457_, _001461_, _001487_);
  and g_095243_(_001438_, _001486_, _001488_);
  or g_095244_(_001439_, _001487_, _001489_);
  and g_095245_(_001483_, _001489_, _001490_);
  or g_095246_(_001485_, _001488_, _001491_);
  and g_095247_(_001476_, _001490_, _001492_);
  or g_095248_(_001475_, _001491_, _001493_);
  or g_095249_(out[816], _001322_, _001494_);
  and g_095250_(_001369_, _001494_, _001496_);
  and g_095251_(_001382_, _001496_, _001497_);
  not g_095252_(_001497_, _001498_);
  and g_095253_(_001314_, _001497_, _001499_);
  or g_095254_(_001315_, _001498_, _001500_);
  and g_095255_(_001366_, _001499_, _001501_);
  or g_095256_(_001367_, _001500_, _001502_);
  and g_095257_(_001472_, _001501_, _001503_);
  or g_095258_(_001474_, _001502_, _001504_);
  and g_095259_(_001493_, _001504_, _001505_);
  or g_095260_(_001492_, _001503_, _001507_);
  and g_095261_(_001292_, _001507_, _001508_);
  or g_095262_(_001291_, _001505_, _001509_);
  and g_095263_(_001390_, _001505_, _001510_);
  or g_095264_(_001391_, _001507_, _001511_);
  and g_095265_(_001509_, _001511_, _001512_);
  or g_095266_(_001508_, _001510_, _001513_);
  or g_095267_(out[833], out[834], _001514_);
  xor g_095268_(out[833], out[834], _001515_);
  xor g_095269_(_001341_, out[834], _001516_);
  or g_095270_(_001346_, _001505_, _001518_);
  or g_095271_(_001339_, _001507_, _001519_);
  and g_095272_(_001518_, _001519_, _001520_);
  not g_095273_(_001520_, _001521_);
  and g_095274_(_001516_, _001520_, _001522_);
  or g_095275_(_001515_, _001521_, _001523_);
  xor g_095276_(out[835], _024903_, _001524_);
  xor g_095277_(_001374_, _024903_, _001525_);
  and g_095278_(_001356_, _001507_, _001526_);
  or g_095279_(_001355_, _001505_, _001527_);
  and g_095280_(_001349_, _001505_, _001529_);
  or g_095281_(_001348_, _001507_, _001530_);
  and g_095282_(_001527_, _001530_, _001531_);
  or g_095283_(_001526_, _001529_, _001532_);
  or g_095284_(_001525_, _001531_, _001533_);
  not g_095285_(_001533_, _001534_);
  and g_095286_(_001523_, _001533_, _001535_);
  or g_095287_(_001522_, _001534_, _001536_);
  or g_095288_(_001209_, _001507_, _001537_);
  or g_095289_(_001329_, _001505_, _001538_);
  and g_095290_(_001537_, _001538_, _001540_);
  and g_095291_(out[833], _001540_, _001541_);
  not g_095292_(_001541_, _001542_);
  and g_095293_(out[816], _001505_, _001543_);
  not g_095294_(_001543_, _001544_);
  and g_095295_(_001321_, _001507_, _001545_);
  or g_095296_(_001322_, _001505_, _001546_);
  or g_095297_(_001543_, _001545_, _001547_);
  and g_095298_(_001544_, _001546_, _001548_);
  and g_095299_(out[832], _001548_, _001549_);
  or g_095300_(_001352_, _001547_, _001551_);
  xor g_095301_(out[833], _001540_, _001552_);
  xor g_095302_(_001341_, _001540_, _001553_);
  and g_095303_(_001551_, _001552_, _001554_);
  or g_095304_(_001549_, _001553_, _001555_);
  and g_095305_(_001542_, _001555_, _001556_);
  or g_095306_(_001541_, _001554_, _001557_);
  xor g_095307_(_001516_, _001520_, _001558_);
  xor g_095308_(_001515_, _001520_, _001559_);
  and g_095309_(_001557_, _001558_, _001560_);
  or g_095310_(_001556_, _001559_, _001562_);
  and g_095311_(_001535_, _001562_, _001563_);
  or g_095312_(_001536_, _001560_, _001564_);
  and g_095313_(_024881_, _025024_, _001565_);
  or g_095314_(_024892_, _025013_, _001566_);
  xor g_095315_(out[842], _024991_, _001567_);
  not g_095316_(_001567_, _001568_);
  and g_095317_(_001512_, _001567_, _001569_);
  or g_095318_(_001513_, _001568_, _001570_);
  and g_095319_(_001566_, _001570_, _001571_);
  or g_095320_(_001565_, _001569_, _001573_);
  and g_095321_(_024892_, _025013_, _001574_);
  or g_095322_(_024881_, _025024_, _001575_);
  and g_095323_(_001513_, _001568_, _001576_);
  or g_095324_(_001512_, _001567_, _001577_);
  and g_095325_(_001575_, _001577_, _001578_);
  or g_095326_(_001574_, _001576_, _001579_);
  and g_095327_(_001413_, _001505_, _001580_);
  not g_095328_(_001580_, _001581_);
  or g_095329_(_001410_, _001505_, _001582_);
  not g_095330_(_001582_, _001584_);
  and g_095331_(_001581_, _001582_, _001585_);
  or g_095332_(_001580_, _001584_, _001586_);
  xor g_095333_(out[841], _024980_, _001587_);
  xor g_095334_(_001396_, _024980_, _001588_);
  and g_095335_(_001585_, _001588_, _001589_);
  not g_095336_(_001589_, _001590_);
  or g_095337_(_001579_, _001589_, _001591_);
  or g_095338_(_001573_, _001591_, _001592_);
  xor g_095339_(out[840], _024969_, _001593_);
  not g_095340_(_001593_, _001595_);
  and g_095341_(_001416_, _001505_, _001596_);
  not g_095342_(_001596_, _001597_);
  or g_095343_(_001423_, _001505_, _001598_);
  not g_095344_(_001598_, _001599_);
  and g_095345_(_001597_, _001598_, _001600_);
  or g_095346_(_001596_, _001599_, _001601_);
  or g_095347_(_001593_, _001600_, _001602_);
  not g_095348_(_001602_, _001603_);
  and g_095349_(_001586_, _001587_, _001604_);
  or g_095350_(_001585_, _001588_, _001606_);
  and g_095351_(_001593_, _001600_, _001607_);
  or g_095352_(_001595_, _001601_, _001608_);
  and g_095353_(_001606_, _001608_, _001609_);
  or g_095354_(_001604_, _001607_, _001610_);
  or g_095355_(_001603_, _001610_, _001611_);
  and g_095356_(_001590_, _001609_, _001612_);
  and g_095357_(_001571_, _001578_, _001613_);
  and g_095358_(_001602_, _001613_, _001614_);
  and g_095359_(_001612_, _001614_, _001615_);
  or g_095360_(_001592_, _001611_, _001617_);
  xor g_095361_(out[838], _024947_, _001618_);
  not g_095362_(_001618_, _001619_);
  and g_095363_(_001441_, _001505_, _001620_);
  not g_095364_(_001620_, _001621_);
  or g_095365_(_001445_, _001505_, _001622_);
  not g_095366_(_001622_, _001623_);
  and g_095367_(_001621_, _001622_, _001624_);
  or g_095368_(_001620_, _001623_, _001625_);
  or g_095369_(_001618_, _001625_, _001626_);
  xor g_095370_(out[839], _024958_, _001628_);
  not g_095371_(_001628_, _001629_);
  and g_095372_(_001448_, _001505_, _001630_);
  not g_095373_(_001630_, _001631_);
  or g_095374_(_001453_, _001505_, _001632_);
  not g_095375_(_001632_, _001633_);
  and g_095376_(_001631_, _001632_, _001634_);
  or g_095377_(_001630_, _001633_, _001635_);
  or g_095378_(_001628_, _001634_, _001636_);
  and g_095379_(_001626_, _001636_, _001637_);
  and g_095380_(_001628_, _001634_, _001639_);
  or g_095381_(_001629_, _001635_, _001640_);
  or g_095382_(_001619_, _001624_, _001641_);
  and g_095383_(_001640_, _001641_, _001642_);
  xor g_095384_(_001618_, _001624_, _001643_);
  xor g_095385_(_001629_, _001634_, _001644_);
  and g_095386_(_001637_, _001642_, _001645_);
  or g_095387_(_001643_, _001644_, _001646_);
  xor g_095388_(out[837], _024936_, _001647_);
  xor g_095389_(_001319_, _024936_, _001648_);
  and g_095390_(_001304_, _001505_, _001650_);
  or g_095391_(_001303_, _001507_, _001651_);
  and g_095392_(_001311_, _001507_, _001652_);
  or g_095393_(_001310_, _001505_, _001653_);
  and g_095394_(_001651_, _001653_, _001654_);
  or g_095395_(_001650_, _001652_, _001655_);
  or g_095396_(_001648_, _001654_, _001656_);
  not g_095397_(_001656_, _001657_);
  xor g_095398_(out[836], _024925_, _001658_);
  not g_095399_(_001658_, _001659_);
  and g_095400_(_001293_, _001505_, _001661_);
  not g_095401_(_001661_, _001662_);
  or g_095402_(_001299_, _001505_, _001663_);
  not g_095403_(_001663_, _001664_);
  and g_095404_(_001662_, _001663_, _001665_);
  or g_095405_(_001661_, _001664_, _001666_);
  and g_095406_(_001658_, _001665_, _001667_);
  or g_095407_(_001659_, _001666_, _001668_);
  and g_095408_(_001656_, _001668_, _001669_);
  or g_095409_(_001657_, _001667_, _001670_);
  and g_095410_(_001659_, _001666_, _001672_);
  or g_095411_(_001658_, _001665_, _001673_);
  and g_095412_(_001648_, _001654_, _001674_);
  or g_095413_(_001647_, _001655_, _001675_);
  and g_095414_(_001525_, _001531_, _001676_);
  or g_095415_(_001524_, _001532_, _001677_);
  and g_095416_(_001675_, _001677_, _001678_);
  or g_095417_(_001674_, _001676_, _001679_);
  and g_095418_(_001673_, _001678_, _001680_);
  or g_095419_(_001672_, _001679_, _001681_);
  and g_095420_(_001669_, _001680_, _001683_);
  or g_095421_(_001670_, _001681_, _001684_);
  and g_095422_(_001645_, _001683_, _001685_);
  or g_095423_(_001646_, _001684_, _001686_);
  and g_095424_(_001615_, _001685_, _001687_);
  or g_095425_(_001617_, _001686_, _001688_);
  and g_095426_(_001564_, _001687_, _001689_);
  or g_095427_(_001563_, _001688_, _001690_);
  and g_095428_(_001645_, _001670_, _001691_);
  not g_095429_(_001691_, _001692_);
  and g_095430_(_001675_, _001691_, _001694_);
  or g_095431_(_001674_, _001692_, _001695_);
  or g_095432_(_001637_, _001639_, _001696_);
  not g_095433_(_001696_, _001697_);
  and g_095434_(_001695_, _001696_, _001698_);
  or g_095435_(_001694_, _001697_, _001699_);
  and g_095436_(_001615_, _001699_, _001700_);
  or g_095437_(_001617_, _001698_, _001701_);
  and g_095438_(_001573_, _001575_, _001702_);
  not g_095439_(_001702_, _001703_);
  and g_095440_(_001610_, _001613_, _001705_);
  and g_095441_(_001590_, _001705_, _001706_);
  or g_095442_(_001592_, _001609_, _001707_);
  and g_095443_(_001690_, _001707_, _001708_);
  or g_095444_(_001689_, _001706_, _001709_);
  and g_095445_(_001701_, _001708_, _001710_);
  or g_095446_(_001700_, _001709_, _001711_);
  and g_095447_(_001703_, _001710_, _001712_);
  or g_095448_(_001702_, _001711_, _001713_);
  or g_095449_(out[832], _001548_, _001714_);
  and g_095450_(_001533_, _001714_, _001716_);
  not g_095451_(_001716_, _001717_);
  or g_095452_(_001559_, _001717_, _001718_);
  or g_095453_(_001555_, _001718_, _001719_);
  not g_095454_(_001719_, _001720_);
  and g_095455_(_001687_, _001720_, _001721_);
  or g_095456_(_001688_, _001719_, _001722_);
  and g_095457_(_001713_, _001722_, _001723_);
  or g_095458_(_001712_, _001721_, _001724_);
  or g_095459_(_001512_, _001723_, _001725_);
  not g_095460_(_001725_, _001727_);
  and g_095461_(_001567_, _001723_, _001728_);
  not g_095462_(_001728_, _001729_);
  and g_095463_(_001725_, _001729_, _001730_);
  or g_095464_(_001727_, _001728_, _001731_);
  and g_095465_(_025035_, _025178_, _001732_);
  or g_095466_(_025046_, _025167_, _001733_);
  xor g_095467_(out[858], _025145_, _001734_);
  not g_095468_(_001734_, _001735_);
  and g_095469_(_001730_, _001734_, _001736_);
  or g_095470_(_001731_, _001735_, _001738_);
  and g_095471_(_001733_, _001738_, _001739_);
  or g_095472_(_001732_, _001736_, _001740_);
  or g_095473_(_001730_, _001734_, _001741_);
  or g_095474_(_025035_, _025178_, _001742_);
  and g_095475_(_001741_, _001742_, _001743_);
  not g_095476_(_001743_, _001744_);
  and g_095477_(_001739_, _001743_, _001745_);
  or g_095478_(_001740_, _001744_, _001746_);
  or g_095479_(_001587_, _001724_, _001747_);
  or g_095480_(_001585_, _001723_, _001749_);
  and g_095481_(_001747_, _001749_, _001750_);
  not g_095482_(_001750_, _001751_);
  xor g_095483_(out[857], _025134_, _001752_);
  xor g_095484_(_001528_, _025134_, _001753_);
  or g_095485_(_001750_, _001753_, _001754_);
  not g_095486_(_001754_, _001755_);
  xor g_095487_(out[856], _025123_, _001756_);
  or g_095488_(_001595_, _001724_, _001757_);
  or g_095489_(_001600_, _001723_, _001758_);
  and g_095490_(_001757_, _001758_, _001760_);
  and g_095491_(_001756_, _001760_, _001761_);
  not g_095492_(_001761_, _001762_);
  and g_095493_(_001754_, _001762_, _001763_);
  or g_095494_(_001755_, _001761_, _001764_);
  or g_095495_(_001756_, _001760_, _001765_);
  not g_095496_(_001765_, _001766_);
  and g_095497_(_001750_, _001753_, _001767_);
  or g_095498_(_001751_, _001752_, _001768_);
  and g_095499_(_001765_, _001768_, _001769_);
  or g_095500_(_001766_, _001767_, _001771_);
  and g_095501_(_001763_, _001769_, _001772_);
  or g_095502_(_001764_, _001771_, _001773_);
  and g_095503_(_001745_, _001772_, _001774_);
  or g_095504_(_001746_, _001773_, _001775_);
  xor g_095505_(out[854], _025101_, _001776_);
  xor g_095506_(_001440_, _025101_, _001777_);
  and g_095507_(_001619_, _001723_, _001778_);
  or g_095508_(_001618_, _001724_, _001779_);
  and g_095509_(_001625_, _001724_, _001780_);
  or g_095510_(_001624_, _001723_, _001782_);
  and g_095511_(_001779_, _001782_, _001783_);
  or g_095512_(_001778_, _001780_, _001784_);
  and g_095513_(_001777_, _001783_, _001785_);
  or g_095514_(_001776_, _001784_, _001786_);
  xor g_095515_(out[855], _025112_, _001787_);
  xor g_095516_(_001429_, _025112_, _001788_);
  and g_095517_(_001628_, _001723_, _001789_);
  or g_095518_(_001629_, _001724_, _001790_);
  and g_095519_(_001635_, _001724_, _001791_);
  or g_095520_(_001634_, _001723_, _001793_);
  and g_095521_(_001790_, _001793_, _001794_);
  or g_095522_(_001789_, _001791_, _001795_);
  and g_095523_(_001788_, _001795_, _001796_);
  or g_095524_(_001787_, _001794_, _001797_);
  and g_095525_(_001786_, _001797_, _001798_);
  or g_095526_(_001785_, _001796_, _001799_);
  and g_095527_(_001787_, _001794_, _001800_);
  not g_095528_(_001800_, _001801_);
  and g_095529_(_001776_, _001784_, _001802_);
  or g_095530_(_001777_, _001783_, _001804_);
  or g_095531_(_001800_, _001802_, _001805_);
  and g_095532_(_001798_, _001801_, _001806_);
  and g_095533_(_001804_, _001806_, _001807_);
  or g_095534_(_001799_, _001805_, _001808_);
  xor g_095535_(out[852], _025079_, _001809_);
  or g_095536_(_001659_, _001724_, _001810_);
  or g_095537_(_001665_, _001723_, _001811_);
  and g_095538_(_001810_, _001811_, _001812_);
  and g_095539_(_001809_, _001812_, _001813_);
  not g_095540_(_001813_, _001815_);
  or g_095541_(_001809_, _001812_, _001816_);
  xor g_095542_(out[853], _025090_, _001817_);
  xor g_095543_(_001451_, _025090_, _001818_);
  or g_095544_(_001647_, _001724_, _001819_);
  or g_095545_(_001654_, _001723_, _001820_);
  and g_095546_(_001819_, _001820_, _001821_);
  not g_095547_(_001821_, _001822_);
  and g_095548_(_001818_, _001821_, _001823_);
  or g_095549_(_001817_, _001822_, _001824_);
  and g_095550_(_001817_, _001822_, _001826_);
  or g_095551_(_001818_, _001821_, _001827_);
  and g_095552_(_001816_, _001827_, _001828_);
  and g_095553_(_001824_, _001828_, _001829_);
  and g_095554_(_001815_, _001829_, _001830_);
  and g_095555_(_001807_, _001830_, _001831_);
  not g_095556_(_001831_, _001832_);
  and g_095557_(_001774_, _001831_, _001833_);
  or g_095558_(_001775_, _001832_, _001834_);
  xor g_095559_(out[851], _025057_, _001835_);
  xor g_095560_(_001506_, _025057_, _001837_);
  or g_095561_(_001531_, _001723_, _001838_);
  or g_095562_(_001524_, _001724_, _001839_);
  and g_095563_(_001838_, _001839_, _001840_);
  not g_095564_(_001840_, _001841_);
  and g_095565_(_001835_, _001841_, _001842_);
  or g_095566_(_001837_, _001840_, _001843_);
  or g_095567_(out[849], out[850], _001844_);
  xor g_095568_(out[849], out[850], _001845_);
  xor g_095569_(_001473_, out[850], _001846_);
  or g_095570_(_001520_, _001723_, _001848_);
  or g_095571_(_001515_, _001724_, _001849_);
  and g_095572_(_001848_, _001849_, _001850_);
  and g_095573_(_001846_, _001850_, _001851_);
  not g_095574_(_001851_, _001852_);
  and g_095575_(_001843_, _001852_, _001853_);
  or g_095576_(_001846_, _001850_, _001854_);
  and g_095577_(_001837_, _001840_, _001855_);
  or g_095578_(_001835_, _001841_, _001856_);
  and g_095579_(_001854_, _001856_, _001857_);
  xor g_095580_(_001845_, _001850_, _001859_);
  or g_095581_(_001842_, _001855_, _001860_);
  and g_095582_(_001853_, _001857_, _001861_);
  or g_095583_(_001859_, _001860_, _001862_);
  or g_095584_(_001341_, _001724_, _001863_);
  or g_095585_(_001540_, _001723_, _001864_);
  and g_095586_(_001863_, _001864_, _001865_);
  and g_095587_(out[849], _001865_, _001866_);
  not g_095588_(_001866_, _001867_);
  and g_095589_(_001548_, _001724_, _001868_);
  and g_095590_(_001352_, _001723_, _001870_);
  or g_095591_(_001868_, _001870_, _001871_);
  and g_095592_(out[848], _001871_, _001872_);
  not g_095593_(_001872_, _001873_);
  xor g_095594_(out[849], _001865_, _001874_);
  xor g_095595_(_001473_, _001865_, _001875_);
  and g_095596_(_001873_, _001874_, _001876_);
  or g_095597_(_001872_, _001875_, _001877_);
  and g_095598_(_001867_, _001877_, _001878_);
  or g_095599_(_001866_, _001876_, _001879_);
  and g_095600_(_001861_, _001879_, _001881_);
  or g_095601_(_001862_, _001878_, _001882_);
  and g_095602_(_001851_, _001856_, _001883_);
  or g_095603_(_001853_, _001855_, _001884_);
  or g_095604_(_001842_, _001883_, _001885_);
  and g_095605_(_001882_, _001884_, _001886_);
  or g_095606_(_001881_, _001885_, _001887_);
  and g_095607_(_001833_, _001887_, _001888_);
  or g_095608_(_001834_, _001886_, _001889_);
  or g_095609_(_001798_, _001800_, _001890_);
  not g_095610_(_001890_, _001892_);
  and g_095611_(_001815_, _001827_, _001893_);
  or g_095612_(_001813_, _001826_, _001894_);
  and g_095613_(_001824_, _001894_, _001895_);
  or g_095614_(_001808_, _001893_, _001896_);
  and g_095615_(_001807_, _001895_, _001897_);
  or g_095616_(_001823_, _001896_, _001898_);
  and g_095617_(_001890_, _001898_, _001899_);
  or g_095618_(_001892_, _001897_, _001900_);
  and g_095619_(_001774_, _001900_, _001901_);
  or g_095620_(_001775_, _001899_, _001903_);
  and g_095621_(_001740_, _001742_, _001904_);
  not g_095622_(_001904_, _001905_);
  or g_095623_(_001763_, _001767_, _001906_);
  and g_095624_(_001745_, _001764_, _001907_);
  and g_095625_(_001768_, _001907_, _001908_);
  or g_095626_(_001746_, _001906_, _001909_);
  and g_095627_(_001905_, _001909_, _001910_);
  or g_095628_(_001904_, _001908_, _001911_);
  and g_095629_(_001903_, _001910_, _001912_);
  or g_095630_(_001901_, _001911_, _001914_);
  and g_095631_(_001889_, _001912_, _001915_);
  or g_095632_(_001888_, _001914_, _001916_);
  or g_095633_(out[848], _001871_, _001917_);
  and g_095634_(_001861_, _001917_, _001918_);
  not g_095635_(_001918_, _001919_);
  and g_095636_(_001876_, _001918_, _001920_);
  or g_095637_(_001877_, _001919_, _001921_);
  and g_095638_(_001833_, _001920_, _001922_);
  or g_095639_(_001834_, _001921_, _001923_);
  and g_095640_(_001916_, _001923_, _001925_);
  or g_095641_(_001915_, _001922_, _001926_);
  or g_095642_(_001730_, _001925_, _001927_);
  or g_095643_(_001735_, _001926_, _001928_);
  and g_095644_(_001927_, _001928_, _001929_);
  and g_095645_(_053979_, _001929_, _001930_);
  or g_095646_(_053980_, _001930_, _001931_);
  not g_095647_(_001931_, _001932_);
  xor g_095648_(out[873], _025288_, _001933_);
  and g_095649_(_001753_, _001925_, _001934_);
  and g_095650_(_001751_, _001926_, _001936_);
  or g_095651_(_001934_, _001936_, _001937_);
  or g_095652_(_001933_, _001937_, _001938_);
  or g_095653_(_025189_, _025321_, _001939_);
  or g_095654_(_053979_, _001929_, _001940_);
  and g_095655_(_001939_, _001940_, _001941_);
  and g_095656_(_001938_, _001941_, _001942_);
  and g_095657_(_001932_, _001942_, _001943_);
  and g_095658_(_001933_, _001937_, _001944_);
  and g_095659_(_001756_, _001925_, _001945_);
  not g_095660_(_001945_, _001947_);
  or g_095661_(_001760_, _001925_, _001948_);
  and g_095662_(_001947_, _001948_, _001949_);
  xor g_095663_(out[872], _025277_, _001950_);
  and g_095664_(_001949_, _001950_, _001951_);
  or g_095665_(_001944_, _001951_, _001952_);
  not g_095666_(_001952_, _001953_);
  or g_095667_(_001949_, _001950_, _001954_);
  and g_095668_(_001953_, _001954_, _001955_);
  and g_095669_(_001943_, _001955_, _001956_);
  xor g_095670_(out[870], _025255_, _001958_);
  xor g_095671_(_001572_, _025255_, _001959_);
  and g_095672_(_001777_, _001925_, _001960_);
  not g_095673_(_001960_, _001961_);
  and g_095674_(_001784_, _001926_, _001962_);
  or g_095675_(_001783_, _001925_, _001963_);
  and g_095676_(_001961_, _001963_, _001964_);
  or g_095677_(_001960_, _001962_, _001965_);
  and g_095678_(_001959_, _001964_, _001966_);
  or g_095679_(_001958_, _001965_, _001967_);
  xor g_095680_(out[871], _025266_, _001969_);
  xor g_095681_(_001561_, _025266_, _001970_);
  and g_095682_(_001787_, _001925_, _001971_);
  or g_095683_(_001788_, _001926_, _001972_);
  or g_095684_(_001794_, _001925_, _001973_);
  not g_095685_(_001973_, _001974_);
  and g_095686_(_001972_, _001973_, _001975_);
  or g_095687_(_001971_, _001974_, _001976_);
  and g_095688_(_001970_, _001976_, _001977_);
  or g_095689_(_001969_, _001975_, _001978_);
  and g_095690_(_001967_, _001978_, _001980_);
  or g_095691_(_001966_, _001977_, _001981_);
  or g_095692_(_001970_, _001976_, _001982_);
  or g_095693_(_001959_, _001964_, _001983_);
  and g_095694_(_001980_, _001983_, _001984_);
  and g_095695_(_001982_, _001984_, _001985_);
  xor g_095696_(out[868], _025233_, _001986_);
  and g_095697_(_001809_, _001925_, _001987_);
  not g_095698_(_001987_, _001988_);
  or g_095699_(_001812_, _001925_, _001989_);
  and g_095700_(_001988_, _001989_, _001991_);
  and g_095701_(_001986_, _001991_, _001992_);
  xor g_095702_(out[869], _025244_, _001993_);
  and g_095703_(_001818_, _001925_, _001994_);
  not g_095704_(_001994_, _001995_);
  or g_095705_(_001821_, _001925_, _001996_);
  not g_095706_(_001996_, _001997_);
  and g_095707_(_001995_, _001996_, _001998_);
  or g_095708_(_001994_, _001997_, _001999_);
  and g_095709_(_001993_, _001999_, _002000_);
  or g_095710_(_001992_, _002000_, _002002_);
  not g_095711_(_002002_, _002003_);
  or g_095712_(_001993_, _001999_, _002004_);
  or g_095713_(_001986_, _001991_, _002005_);
  and g_095714_(_002004_, _002005_, _002006_);
  and g_095715_(_002003_, _002006_, _002007_);
  and g_095716_(_001985_, _002007_, _002008_);
  xor g_095717_(out[867], _025211_, _002009_);
  and g_095718_(_001841_, _001926_, _002010_);
  and g_095719_(_001837_, _001925_, _002011_);
  or g_095720_(_002010_, _002011_, _002013_);
  or g_095721_(_002009_, _002013_, _002014_);
  and g_095722_(_002009_, _002013_, _002015_);
  or g_095723_(out[865], out[866], _002016_);
  xor g_095724_(_001605_, out[866], _002017_);
  or g_095725_(_001845_, _001926_, _002018_);
  or g_095726_(_001850_, _001925_, _002019_);
  and g_095727_(_002018_, _002019_, _002020_);
  and g_095728_(_002017_, _002020_, _002021_);
  or g_095729_(_002015_, _002021_, _002022_);
  and g_095730_(_002014_, _002022_, _002024_);
  xor g_095731_(_002009_, _002013_, _002025_);
  xor g_095732_(_002017_, _002020_, _002026_);
  and g_095733_(_002025_, _002026_, _002027_);
  or g_095734_(_001473_, _001926_, _002028_);
  or g_095735_(_001865_, _001925_, _002029_);
  and g_095736_(_002028_, _002029_, _002030_);
  and g_095737_(out[865], _002030_, _002031_);
  and g_095738_(_002027_, _002031_, _002032_);
  or g_095739_(_002024_, _002032_, _002033_);
  and g_095740_(_002008_, _002033_, _002035_);
  and g_095741_(_001871_, _001926_, _002036_);
  and g_095742_(_001484_, _001925_, _002037_);
  or g_095743_(_002036_, _002037_, _002038_);
  and g_095744_(out[864], _002038_, _002039_);
  not g_095745_(_002039_, _002040_);
  xor g_095746_(out[865], _002030_, _002041_);
  and g_095747_(_002040_, _002041_, _002042_);
  and g_095748_(_002027_, _002042_, _002043_);
  and g_095749_(_002008_, _002043_, _002044_);
  and g_095750_(_002002_, _002004_, _002046_);
  and g_095751_(_001985_, _002046_, _002047_);
  and g_095752_(_001981_, _001982_, _002048_);
  or g_095753_(_002047_, _002048_, _002049_);
  or g_095754_(_002035_, _002049_, _002050_);
  or g_095755_(_002044_, _002050_, _002051_);
  and g_095756_(_001956_, _002051_, _002052_);
  and g_095757_(_001943_, _001952_, _002053_);
  and g_095758_(_001931_, _001939_, _002054_);
  or g_095759_(_002053_, _002054_, _002055_);
  or g_095760_(_002052_, _002055_, _002057_);
  or g_095761_(out[864], _002038_, _002058_);
  and g_095762_(_001956_, _002058_, _002059_);
  and g_095763_(_002044_, _002059_, _002060_);
  not g_095764_(_002060_, _002061_);
  and g_095765_(_002057_, _002061_, _002062_);
  not g_095766_(_002062_, _002063_);
  and g_095767_(_053979_, _002062_, _002064_);
  not g_095768_(_002064_, _002065_);
  or g_095769_(_001929_, _002062_, _002066_);
  and g_095770_(_002065_, _002066_, _002068_);
  xor g_095771_(_001770_, _025365_, _002069_);
  and g_095772_(_002009_, _002062_, _002070_);
  or g_095773_(_002013_, _002062_, _002071_);
  not g_095774_(_002071_, _002072_);
  or g_095775_(_002070_, _002072_, _002073_);
  or g_095776_(_002069_, _002073_, _002074_);
  or g_095777_(out[881], out[882], _002075_);
  xor g_095778_(out[881], out[882], _002076_);
  xor g_095779_(_001737_, out[882], _002077_);
  or g_095780_(_002020_, _002062_, _002079_);
  and g_095781_(_002017_, _002062_, _002080_);
  not g_095782_(_002080_, _002081_);
  and g_095783_(_002079_, _002081_, _002082_);
  and g_095784_(_002077_, _002082_, _002083_);
  not g_095785_(_002083_, _002084_);
  and g_095786_(_002069_, _002073_, _002085_);
  xor g_095787_(_002077_, _002082_, _002086_);
  xor g_095788_(_002069_, _002073_, _002087_);
  and g_095789_(_002086_, _002087_, _002088_);
  or g_095790_(_001605_, _002063_, _002090_);
  or g_095791_(_002030_, _002062_, _002091_);
  and g_095792_(_002090_, _002091_, _002092_);
  and g_095793_(out[881], _002092_, _002093_);
  and g_095794_(out[864], _002062_, _002094_);
  not g_095795_(_002094_, _002095_);
  or g_095796_(_002038_, _002062_, _002096_);
  not g_095797_(_002096_, _002097_);
  or g_095798_(_002094_, _002097_, _002098_);
  and g_095799_(_002095_, _002096_, _002099_);
  and g_095800_(out[880], _002099_, _002101_);
  or g_095801_(_001748_, _002098_, _002102_);
  xor g_095802_(out[881], _002092_, _002103_);
  xor g_095803_(_001737_, _002092_, _002104_);
  and g_095804_(_002102_, _002103_, _002105_);
  or g_095805_(_002101_, _002104_, _002106_);
  or g_095806_(_002093_, _002105_, _002107_);
  and g_095807_(_002088_, _002107_, _002108_);
  or g_095808_(_002084_, _002085_, _002109_);
  and g_095809_(_002074_, _002109_, _002110_);
  not g_095810_(_002110_, _002112_);
  or g_095811_(_002108_, _002112_, _002113_);
  and g_095812_(_025343_, _025486_, _002114_);
  or g_095813_(_025354_, _025475_, _002115_);
  xor g_095814_(out[890], _025453_, _002116_);
  and g_095815_(_002068_, _002116_, _002117_);
  not g_095816_(_002117_, _002118_);
  and g_095817_(_002115_, _002118_, _002119_);
  or g_095818_(_002114_, _002117_, _002120_);
  xor g_095819_(out[889], _025442_, _002121_);
  xor g_095820_(_001792_, _025442_, _002123_);
  or g_095821_(_001937_, _002062_, _002124_);
  not g_095822_(_002124_, _002125_);
  and g_095823_(_001933_, _002062_, _002126_);
  or g_095824_(_002125_, _002126_, _002127_);
  not g_095825_(_002127_, _002128_);
  and g_095826_(_002123_, _002127_, _002129_);
  or g_095827_(_002121_, _002128_, _002130_);
  or g_095828_(_025343_, _025486_, _002131_);
  or g_095829_(_002068_, _002116_, _002132_);
  and g_095830_(_002131_, _002132_, _002134_);
  or g_095831_(_002123_, _002127_, _002135_);
  not g_095832_(_002135_, _002136_);
  xor g_095833_(out[888], _025431_, _002137_);
  or g_095834_(_001949_, _002062_, _002138_);
  and g_095835_(_001950_, _002062_, _002139_);
  not g_095836_(_002139_, _002140_);
  and g_095837_(_002138_, _002140_, _002141_);
  and g_095838_(_002137_, _002141_, _002142_);
  not g_095839_(_002142_, _002143_);
  and g_095840_(_002135_, _002143_, _002145_);
  or g_095841_(_002136_, _002142_, _002146_);
  or g_095842_(_002137_, _002141_, _002147_);
  and g_095843_(_002130_, _002145_, _002148_);
  or g_095844_(_002129_, _002146_, _002149_);
  and g_095845_(_002119_, _002134_, _002150_);
  and g_095846_(_002147_, _002150_, _002151_);
  not g_095847_(_002151_, _002152_);
  and g_095848_(_002148_, _002151_, _002153_);
  or g_095849_(_002149_, _002152_, _002154_);
  xor g_095850_(out[886], _025409_, _002156_);
  xor g_095851_(_001704_, _025409_, _002157_);
  or g_095852_(_001964_, _002062_, _002158_);
  not g_095853_(_002158_, _002159_);
  and g_095854_(_001959_, _002062_, _002160_);
  or g_095855_(_001958_, _002063_, _002161_);
  and g_095856_(_002158_, _002161_, _002162_);
  or g_095857_(_002159_, _002160_, _002163_);
  and g_095858_(_002156_, _002163_, _002164_);
  or g_095859_(_002157_, _002162_, _002165_);
  xor g_095860_(_001715_, _025398_, _002167_);
  or g_095861_(_001998_, _002062_, _002168_);
  or g_095862_(_001993_, _002063_, _002169_);
  and g_095863_(_002168_, _002169_, _002170_);
  and g_095864_(_002167_, _002170_, _002171_);
  not g_095865_(_002171_, _002172_);
  and g_095866_(_002165_, _002172_, _002173_);
  or g_095867_(_002164_, _002171_, _002174_);
  xor g_095868_(out[887], _025420_, _002175_);
  xor g_095869_(_001693_, _025420_, _002176_);
  and g_095870_(_001976_, _002063_, _002178_);
  or g_095871_(_001975_, _002062_, _002179_);
  and g_095872_(_001969_, _002062_, _002180_);
  or g_095873_(_001970_, _002063_, _002181_);
  and g_095874_(_002179_, _002181_, _002182_);
  or g_095875_(_002178_, _002180_, _002183_);
  and g_095876_(_002175_, _002182_, _002184_);
  or g_095877_(_002176_, _002183_, _002185_);
  xor g_095878_(out[884], _025387_, _002186_);
  and g_095879_(_001986_, _002062_, _002187_);
  not g_095880_(_002187_, _002189_);
  or g_095881_(_001991_, _002062_, _002190_);
  and g_095882_(_002189_, _002190_, _002191_);
  or g_095883_(_002186_, _002191_, _002192_);
  not g_095884_(_002192_, _002193_);
  or g_095885_(_002184_, _002193_, _002194_);
  or g_095886_(_002174_, _002194_, _002195_);
  and g_095887_(_002186_, _002191_, _002196_);
  not g_095888_(_002196_, _002197_);
  or g_095889_(_002167_, _002170_, _002198_);
  not g_095890_(_002198_, _002200_);
  or g_095891_(_002196_, _002200_, _002201_);
  and g_095892_(_002157_, _002162_, _002202_);
  or g_095893_(_002156_, _002163_, _002203_);
  and g_095894_(_002176_, _002183_, _002204_);
  or g_095895_(_002175_, _002182_, _002205_);
  and g_095896_(_002203_, _002205_, _002206_);
  or g_095897_(_002202_, _002204_, _002207_);
  or g_095898_(_002201_, _002207_, _002208_);
  and g_095899_(_002185_, _002206_, _002209_);
  and g_095900_(_002173_, _002209_, _002211_);
  and g_095901_(_002192_, _002198_, _002212_);
  and g_095902_(_002197_, _002212_, _002213_);
  and g_095903_(_002211_, _002213_, _002214_);
  or g_095904_(_002195_, _002208_, _002215_);
  or g_095905_(_002154_, _002215_, _002216_);
  and g_095906_(_002173_, _002201_, _002217_);
  or g_095907_(_002207_, _002217_, _002218_);
  and g_095908_(_002185_, _002218_, _002219_);
  and g_095909_(_002120_, _002131_, _002220_);
  and g_095910_(_002130_, _002146_, _002222_);
  and g_095911_(_002150_, _002222_, _002223_);
  and g_095912_(_002113_, _002214_, _002224_);
  or g_095913_(_002219_, _002224_, _002225_);
  and g_095914_(_002153_, _002225_, _002226_);
  or g_095915_(_002223_, _002226_, _002227_);
  or g_095916_(_002220_, _002227_, _002228_);
  or g_095917_(out[880], _002099_, _002229_);
  and g_095918_(_002088_, _002229_, _002230_);
  not g_095919_(_002230_, _002231_);
  or g_095920_(_002106_, _002231_, _002233_);
  or g_095921_(_002216_, _002233_, _002234_);
  and g_095922_(_002228_, _002234_, _002235_);
  not g_095923_(_002235_, _002236_);
  or g_095924_(_002068_, _002235_, _002237_);
  not g_095925_(_002237_, _002238_);
  and g_095926_(_002116_, _002235_, _002239_);
  or g_095927_(_002238_, _002239_, _002240_);
  and g_095928_(_025497_, _025640_, _002241_);
  or g_095929_(_025508_, _025629_, _002242_);
  xor g_095930_(_001935_, _025607_, _002244_);
  or g_095931_(_002240_, _002244_, _002245_);
  not g_095932_(_002245_, _002246_);
  and g_095933_(_002242_, _002245_, _002247_);
  or g_095934_(_002241_, _002246_, _002248_);
  or g_095935_(_025497_, _025640_, _002249_);
  and g_095936_(_002240_, _002244_, _002250_);
  not g_095937_(_002250_, _002251_);
  and g_095938_(_002247_, _002251_, _002252_);
  and g_095939_(_002249_, _002252_, _002253_);
  and g_095940_(_002123_, _002235_, _002255_);
  and g_095941_(_002128_, _002236_, _002256_);
  or g_095942_(_002255_, _002256_, _002257_);
  xor g_095943_(out[905], _025596_, _002258_);
  not g_095944_(_002258_, _002259_);
  and g_095945_(_002257_, _002258_, _002260_);
  not g_095946_(_002260_, _002261_);
  xor g_095947_(_001913_, _025585_, _002262_);
  and g_095948_(_002137_, _002235_, _002263_);
  or g_095949_(_002141_, _002235_, _002264_);
  not g_095950_(_002264_, _002266_);
  or g_095951_(_002263_, _002266_, _002267_);
  or g_095952_(_002262_, _002267_, _002268_);
  not g_095953_(_002268_, _002269_);
  and g_095954_(_002261_, _002268_, _002270_);
  or g_095955_(_002260_, _002269_, _002271_);
  and g_095956_(_002262_, _002267_, _002272_);
  not g_095957_(_002272_, _002273_);
  or g_095958_(_002257_, _002258_, _002274_);
  and g_095959_(_002273_, _002274_, _002275_);
  and g_095960_(_002270_, _002275_, _002277_);
  and g_095961_(_002253_, _002277_, _002278_);
  xor g_095962_(out[901], _025552_, _002279_);
  xor g_095963_(_001847_, _025552_, _002280_);
  and g_095964_(_002167_, _002235_, _002281_);
  not g_095965_(_002281_, _002282_);
  or g_095966_(_002170_, _002235_, _002283_);
  not g_095967_(_002283_, _002284_);
  and g_095968_(_002282_, _002283_, _002285_);
  or g_095969_(_002281_, _002284_, _002286_);
  or g_095970_(_002279_, _002286_, _002288_);
  and g_095971_(_002278_, _002288_, _002289_);
  not g_095972_(_002289_, _002290_);
  xor g_095973_(out[902], _025563_, _002291_);
  not g_095974_(_002291_, _002292_);
  and g_095975_(_002162_, _002236_, _002293_);
  or g_095976_(_002163_, _002235_, _002294_);
  and g_095977_(_002156_, _002235_, _002295_);
  not g_095978_(_002295_, _002296_);
  or g_095979_(_002293_, _002295_, _002297_);
  and g_095980_(_002294_, _002296_, _002299_);
  and g_095981_(_002292_, _002297_, _002300_);
  xor g_095982_(out[903], _025574_, _002301_);
  not g_095983_(_002301_, _002302_);
  and g_095984_(_002175_, _002235_, _002303_);
  not g_095985_(_002303_, _002304_);
  and g_095986_(_002183_, _002236_, _002305_);
  or g_095987_(_002182_, _002235_, _002306_);
  and g_095988_(_002304_, _002306_, _002307_);
  or g_095989_(_002303_, _002305_, _002308_);
  and g_095990_(_002302_, _002308_, _002310_);
  or g_095991_(_002300_, _002310_, _002311_);
  and g_095992_(_002291_, _002299_, _002312_);
  and g_095993_(_002301_, _002307_, _002313_);
  or g_095994_(_002302_, _002308_, _002314_);
  or g_095995_(_002312_, _002313_, _002315_);
  xor g_095996_(_002292_, _002297_, _002316_);
  xor g_095997_(_002301_, _002307_, _002317_);
  and g_095998_(_002316_, _002317_, _002318_);
  or g_095999_(_002311_, _002315_, _002319_);
  xor g_096000_(out[900], _025541_, _002321_);
  xor g_096001_(_001858_, _025541_, _002322_);
  and g_096002_(_002186_, _002235_, _002323_);
  not g_096003_(_002323_, _002324_);
  or g_096004_(_002191_, _002235_, _002325_);
  not g_096005_(_002325_, _002326_);
  and g_096006_(_002324_, _002325_, _002327_);
  or g_096007_(_002323_, _002326_, _002328_);
  and g_096008_(_002322_, _002328_, _002329_);
  or g_096009_(_002321_, _002327_, _002330_);
  or g_096010_(out[897], out[898], _002332_);
  xor g_096011_(out[897], out[898], _002333_);
  xor g_096012_(_001869_, out[898], _002334_);
  or g_096013_(_002082_, _002235_, _002335_);
  not g_096014_(_002335_, _002336_);
  and g_096015_(_002077_, _002235_, _002337_);
  or g_096016_(_002336_, _002337_, _002338_);
  not g_096017_(_002338_, _002339_);
  and g_096018_(_002333_, _002338_, _002340_);
  xor g_096019_(out[899], _025519_, _002341_);
  xor g_096020_(_001902_, _025519_, _002343_);
  or g_096021_(_002073_, _002235_, _002344_);
  not g_096022_(_002344_, _002345_);
  and g_096023_(_002069_, _002235_, _002346_);
  or g_096024_(_002345_, _002346_, _002347_);
  not g_096025_(_002347_, _002348_);
  and g_096026_(_002343_, _002348_, _002349_);
  or g_096027_(_002341_, _002347_, _002350_);
  or g_096028_(_002340_, _002349_, _002351_);
  or g_096029_(_002329_, _002351_, _002352_);
  and g_096030_(_002321_, _002327_, _002354_);
  or g_096031_(_002322_, _002328_, _002355_);
  and g_096032_(_002279_, _002286_, _002356_);
  or g_096033_(_002280_, _002285_, _002357_);
  and g_096034_(_002355_, _002357_, _002358_);
  or g_096035_(_002354_, _002356_, _002359_);
  and g_096036_(_002334_, _002339_, _002360_);
  and g_096037_(_002341_, _002347_, _002361_);
  or g_096038_(_002360_, _002361_, _002362_);
  or g_096039_(_002359_, _002362_, _002363_);
  or g_096040_(_002352_, _002363_, _002365_);
  xor g_096041_(_002341_, _002347_, _002366_);
  and g_096042_(_002318_, _002358_, _002367_);
  and g_096043_(_002330_, _002367_, _002368_);
  xor g_096044_(_002333_, _002338_, _002369_);
  and g_096045_(_002366_, _002368_, _002370_);
  and g_096046_(_002369_, _002370_, _002371_);
  or g_096047_(_002319_, _002365_, _002372_);
  and g_096048_(out[881], _002235_, _002373_);
  not g_096049_(_002373_, _002374_);
  or g_096050_(_002092_, _002235_, _002376_);
  not g_096051_(_002376_, _002377_);
  and g_096052_(_002374_, _002376_, _002378_);
  or g_096053_(_002373_, _002377_, _002379_);
  and g_096054_(out[897], _002378_, _002380_);
  or g_096055_(_001869_, _002379_, _002381_);
  and g_096056_(_002099_, _002236_, _002382_);
  and g_096057_(_001748_, _002235_, _002383_);
  or g_096058_(_002382_, _002383_, _002384_);
  and g_096059_(out[896], _002384_, _002385_);
  not g_096060_(_002385_, _002387_);
  xor g_096061_(out[897], _002378_, _002388_);
  xor g_096062_(_001869_, _002378_, _002389_);
  and g_096063_(_002387_, _002388_, _002390_);
  or g_096064_(_002385_, _002389_, _002391_);
  and g_096065_(_002381_, _002391_, _002392_);
  or g_096066_(_002380_, _002390_, _002393_);
  and g_096067_(_002371_, _002393_, _002394_);
  or g_096068_(_002372_, _002392_, _002395_);
  and g_096069_(_002330_, _002350_, _002396_);
  and g_096070_(_002362_, _002396_, _002398_);
  or g_096071_(_002359_, _002398_, _002399_);
  not g_096072_(_002399_, _002400_);
  and g_096073_(_002318_, _002399_, _002401_);
  or g_096074_(_002319_, _002400_, _002402_);
  and g_096075_(_002371_, _002390_, _002403_);
  or g_096076_(_002372_, _002391_, _002404_);
  and g_096077_(_002395_, _002402_, _002405_);
  or g_096078_(_002394_, _002401_, _002406_);
  and g_096079_(_002289_, _002406_, _002407_);
  or g_096080_(_002290_, _002405_, _002409_);
  and g_096081_(_002311_, _002314_, _002410_);
  and g_096082_(_002278_, _002410_, _002411_);
  and g_096083_(_002248_, _002249_, _002412_);
  and g_096084_(_002271_, _002274_, _002413_);
  and g_096085_(_002253_, _002413_, _002414_);
  or g_096086_(_002412_, _002414_, _002415_);
  or g_096087_(_002411_, _002415_, _002416_);
  not g_096088_(_002416_, _002417_);
  and g_096089_(_002409_, _002417_, _002418_);
  or g_096090_(_002407_, _002416_, _002420_);
  or g_096091_(out[896], _002384_, _002421_);
  and g_096092_(_002289_, _002421_, _002422_);
  not g_096093_(_002422_, _002423_);
  and g_096094_(_002403_, _002422_, _002424_);
  or g_096095_(_002404_, _002423_, _002425_);
  and g_096096_(_002420_, _002425_, _002426_);
  or g_096097_(_002418_, _002424_, _002427_);
  and g_096098_(_002240_, _002427_, _002428_);
  not g_096099_(_002428_, _002429_);
  or g_096100_(_002244_, _002427_, _002431_);
  not g_096101_(_002431_, _002432_);
  and g_096102_(_002429_, _002431_, _002433_);
  or g_096103_(_002428_, _002432_, _002434_);
  and g_096104_(_053978_, _002434_, _002435_);
  xor g_096105_(out[919], _025728_, _002436_);
  xor g_096106_(_001957_, _025728_, _002437_);
  and g_096107_(_002308_, _002427_, _002438_);
  or g_096108_(_002307_, _002426_, _002439_);
  and g_096109_(_002301_, _002426_, _002440_);
  or g_096110_(_002302_, _002427_, _002442_);
  and g_096111_(_002439_, _002442_, _002443_);
  or g_096112_(_002438_, _002440_, _002444_);
  and g_096113_(_002436_, _002443_, _002445_);
  xor g_096114_(_002045_, _025739_, _002446_);
  and g_096115_(_002267_, _002427_, _002447_);
  or g_096116_(_002262_, _002427_, _002448_);
  not g_096117_(_002448_, _002449_);
  or g_096118_(_002447_, _002449_, _002450_);
  and g_096119_(_002446_, _002450_, _002451_);
  or g_096120_(_002445_, _002451_, _002453_);
  and g_096121_(_025651_, _025794_, _002454_);
  or g_096122_(_025662_, _025783_, _002455_);
  and g_096123_(_053977_, _002433_, _002456_);
  or g_096124_(_053978_, _002434_, _002457_);
  and g_096125_(_002455_, _002457_, _002458_);
  or g_096126_(_002454_, _002456_, _002459_);
  xor g_096127_(out[921], _025750_, _002460_);
  not g_096128_(_002460_, _002461_);
  and g_096129_(_002257_, _002427_, _002462_);
  and g_096130_(_002259_, _002426_, _002464_);
  or g_096131_(_002462_, _002464_, _002465_);
  not g_096132_(_002465_, _002466_);
  and g_096133_(_002460_, _002465_, _002467_);
  not g_096134_(_002467_, _002468_);
  or g_096135_(_002446_, _002450_, _002469_);
  not g_096136_(_002469_, _002470_);
  and g_096137_(_002468_, _002469_, _002471_);
  or g_096138_(_002467_, _002470_, _002472_);
  and g_096139_(_025662_, _025783_, _002473_);
  and g_096140_(_002461_, _002466_, _002475_);
  or g_096141_(_002435_, _002473_, _002476_);
  or g_096142_(_002459_, _002476_, _002477_);
  or g_096143_(_002453_, _002475_, _002478_);
  or g_096144_(_002472_, _002478_, _002479_);
  or g_096145_(_002477_, _002479_, _002480_);
  xor g_096146_(out[916], _025695_, _002481_);
  not g_096147_(_002481_, _002482_);
  and g_096148_(_002328_, _002427_, _002483_);
  and g_096149_(_002321_, _002426_, _002484_);
  or g_096150_(_002483_, _002484_, _002486_);
  or g_096151_(_002482_, _002486_, _002487_);
  xor g_096152_(out[917], _025706_, _002488_);
  xor g_096153_(_001979_, _025706_, _002489_);
  and g_096154_(_002286_, _002427_, _002490_);
  or g_096155_(_002285_, _002426_, _002491_);
  and g_096156_(_002280_, _002426_, _002492_);
  or g_096157_(_002279_, _002427_, _002493_);
  and g_096158_(_002491_, _002493_, _002494_);
  or g_096159_(_002490_, _002492_, _002495_);
  and g_096160_(_002488_, _002495_, _002497_);
  or g_096161_(_002489_, _002494_, _002498_);
  and g_096162_(_002437_, _002444_, _002499_);
  or g_096163_(_002436_, _002443_, _002500_);
  xor g_096164_(out[918], _025717_, _002501_);
  xor g_096165_(_001968_, _025717_, _002502_);
  and g_096166_(_002299_, _002427_, _002503_);
  or g_096167_(_002297_, _002426_, _002504_);
  and g_096168_(_002292_, _002426_, _002505_);
  or g_096169_(_002291_, _002427_, _002506_);
  and g_096170_(_002504_, _002506_, _002508_);
  or g_096171_(_002503_, _002505_, _002509_);
  and g_096172_(_002501_, _002509_, _002510_);
  or g_096173_(_002499_, _002510_, _002511_);
  and g_096174_(_002489_, _002494_, _002512_);
  and g_096175_(_002502_, _002508_, _002513_);
  or g_096176_(_002501_, _002509_, _002514_);
  xor g_096177_(_002481_, _002486_, _002515_);
  or g_096178_(_002512_, _002515_, _002516_);
  or g_096179_(_002497_, _002513_, _002517_);
  or g_096180_(_002511_, _002517_, _002519_);
  or g_096181_(_002516_, _002519_, _002520_);
  or g_096182_(_002480_, _002520_, _002521_);
  not g_096183_(_002521_, _002522_);
  xor g_096184_(out[915], _025673_, _002523_);
  and g_096185_(_002347_, _002427_, _002524_);
  and g_096186_(_002343_, _002426_, _002525_);
  or g_096187_(_002524_, _002525_, _002526_);
  and g_096188_(_002523_, _002526_, _002527_);
  or g_096189_(out[913], out[914], _002528_);
  xor g_096190_(out[913], out[914], _002530_);
  xor g_096191_(_002001_, out[914], _002531_);
  and g_096192_(_002338_, _002427_, _002532_);
  and g_096193_(_002334_, _002426_, _002533_);
  or g_096194_(_002532_, _002533_, _002534_);
  and g_096195_(_002530_, _002534_, _002535_);
  or g_096196_(_002530_, _002534_, _002536_);
  not g_096197_(_002536_, _002537_);
  or g_096198_(_002523_, _002526_, _002538_);
  xor g_096199_(_002523_, _002526_, _002539_);
  and g_096200_(_002536_, _002539_, _002541_);
  not g_096201_(_002541_, _002542_);
  xor g_096202_(_002530_, _002534_, _002543_);
  and g_096203_(_002539_, _002543_, _002544_);
  or g_096204_(_002535_, _002542_, _002545_);
  or g_096205_(_001869_, _002427_, _002546_);
  or g_096206_(_002378_, _002426_, _002547_);
  and g_096207_(_002546_, _002547_, _002548_);
  and g_096208_(out[913], _002548_, _002549_);
  and g_096209_(_002384_, _002427_, _002550_);
  and g_096210_(_001880_, _002426_, _002552_);
  or g_096211_(_002550_, _002552_, _002553_);
  and g_096212_(out[912], _002553_, _002554_);
  not g_096213_(_002554_, _002555_);
  xor g_096214_(out[913], _002548_, _002556_);
  xor g_096215_(_002001_, _002548_, _002557_);
  and g_096216_(_002555_, _002556_, _002558_);
  or g_096217_(_002554_, _002557_, _002559_);
  and g_096218_(_002544_, _002558_, _002560_);
  or g_096219_(_002545_, _002559_, _002561_);
  and g_096220_(_002544_, _002549_, _002563_);
  and g_096221_(_002537_, _002538_, _002564_);
  or g_096222_(_002527_, _002564_, _002565_);
  or g_096223_(_002563_, _002565_, _002566_);
  not g_096224_(_002566_, _002567_);
  and g_096225_(_002561_, _002567_, _002568_);
  or g_096226_(_002560_, _002566_, _002569_);
  and g_096227_(_002522_, _002569_, _002570_);
  or g_096228_(_002521_, _002568_, _002571_);
  and g_096229_(_002487_, _002498_, _002572_);
  or g_096230_(_002511_, _002572_, _002574_);
  or g_096231_(_002512_, _002574_, _002575_);
  and g_096232_(_002500_, _002514_, _002576_);
  and g_096233_(_002575_, _002576_, _002577_);
  or g_096234_(_002480_, _002577_, _002578_);
  or g_096235_(_002435_, _002475_, _002579_);
  or g_096236_(_002471_, _002579_, _002580_);
  and g_096237_(_002458_, _002580_, _002581_);
  or g_096238_(_002473_, _002581_, _002582_);
  and g_096239_(_002578_, _002582_, _002583_);
  not g_096240_(_002583_, _002585_);
  and g_096241_(_002571_, _002583_, _002586_);
  or g_096242_(_002570_, _002585_, _002587_);
  or g_096243_(out[912], _002553_, _002588_);
  not g_096244_(_002588_, _002589_);
  and g_096245_(_002560_, _002588_, _002590_);
  or g_096246_(_002561_, _002589_, _002591_);
  and g_096247_(_002522_, _002590_, _002592_);
  or g_096248_(_002521_, _002591_, _002593_);
  and g_096249_(_002587_, _002593_, _002594_);
  or g_096250_(_002586_, _002592_, _002596_);
  and g_096251_(_053977_, _002594_, _002597_);
  or g_096252_(_053978_, _002596_, _002598_);
  and g_096253_(_002434_, _002596_, _002599_);
  or g_096254_(_002433_, _002594_, _002600_);
  and g_096255_(_002598_, _002600_, _002601_);
  or g_096256_(_002597_, _002599_, _002602_);
  and g_096257_(_053975_, _002601_, _002603_);
  or g_096258_(_053976_, _002602_, _002604_);
  and g_096259_(_053974_, _002604_, _002605_);
  or g_096260_(_053972_, _002603_, _002607_);
  and g_096261_(_053976_, _002602_, _002608_);
  not g_096262_(_002608_, _002609_);
  and g_096263_(_025805_, _025948_, _002610_);
  or g_096264_(_025816_, _025937_, _002611_);
  or g_096265_(_002608_, _002610_, _002612_);
  and g_096266_(_002605_, _002611_, _002613_);
  and g_096267_(_002609_, _002613_, _002614_);
  or g_096268_(_002607_, _002612_, _002615_);
  and g_096269_(_002465_, _002596_, _002616_);
  not g_096270_(_002616_, _002618_);
  or g_096271_(_002460_, _002596_, _002619_);
  not g_096272_(_002619_, _002620_);
  and g_096273_(_002618_, _002619_, _002621_);
  or g_096274_(_002616_, _002620_, _002622_);
  and g_096275_(_053970_, _002622_, _002623_);
  or g_096276_(_053971_, _002621_, _002624_);
  and g_096277_(_002450_, _002596_, _002625_);
  not g_096278_(_002625_, _002626_);
  or g_096279_(_002446_, _002596_, _002627_);
  not g_096280_(_002627_, _002629_);
  and g_096281_(_002626_, _002627_, _002630_);
  or g_096282_(_002625_, _002629_, _002631_);
  xor g_096283_(out[936], _025893_, _002632_);
  not g_096284_(_002632_, _002633_);
  and g_096285_(_002630_, _002632_, _002634_);
  or g_096286_(_002631_, _002633_, _002635_);
  and g_096287_(_002624_, _002635_, _002636_);
  or g_096288_(_002623_, _002634_, _002637_);
  and g_096289_(_053971_, _002621_, _002638_);
  or g_096290_(_053970_, _002622_, _002640_);
  and g_096291_(_002631_, _002633_, _002641_);
  or g_096292_(_002630_, _002632_, _002642_);
  and g_096293_(_002640_, _002642_, _002643_);
  or g_096294_(_002638_, _002641_, _002644_);
  and g_096295_(_002636_, _002643_, _002645_);
  or g_096296_(_002637_, _002644_, _002646_);
  and g_096297_(_002614_, _002645_, _002647_);
  or g_096298_(_002615_, _002646_, _002648_);
  xor g_096299_(out[933], _025860_, _002649_);
  xor g_096300_(_002089_, _025860_, _002651_);
  and g_096301_(_002495_, _002596_, _002652_);
  or g_096302_(_002494_, _002594_, _002653_);
  and g_096303_(_002489_, _002594_, _002654_);
  or g_096304_(_002488_, _002596_, _002655_);
  and g_096305_(_002653_, _002655_, _002656_);
  or g_096306_(_002652_, _002654_, _002657_);
  and g_096307_(_002651_, _002656_, _002658_);
  not g_096308_(_002658_, _002659_);
  xor g_096309_(_002100_, _025849_, _002660_);
  and g_096310_(_002481_, _002594_, _002662_);
  and g_096311_(_002486_, _002596_, _002663_);
  or g_096312_(_002662_, _002663_, _002664_);
  and g_096313_(_002660_, _002664_, _002665_);
  or g_096314_(_002658_, _002665_, _002666_);
  not g_096315_(_002666_, _002667_);
  xor g_096316_(out[935], _025882_, _002668_);
  not g_096317_(_002668_, _002669_);
  and g_096318_(_002444_, _002596_, _002670_);
  not g_096319_(_002670_, _002671_);
  and g_096320_(_002436_, _002594_, _002673_);
  or g_096321_(_002437_, _002596_, _002674_);
  and g_096322_(_002671_, _002674_, _002675_);
  or g_096323_(_002670_, _002673_, _002676_);
  and g_096324_(_002668_, _002675_, _002677_);
  or g_096325_(_002669_, _002676_, _002678_);
  xor g_096326_(out[934], _025871_, _002679_);
  not g_096327_(_002679_, _002680_);
  or g_096328_(_002508_, _002594_, _002681_);
  or g_096329_(_002501_, _002596_, _002682_);
  and g_096330_(_002681_, _002682_, _002684_);
  or g_096331_(_002680_, _002684_, _002685_);
  not g_096332_(_002685_, _002686_);
  and g_096333_(_002678_, _002685_, _002687_);
  or g_096334_(_002677_, _002686_, _002688_);
  and g_096335_(_002667_, _002687_, _002689_);
  or g_096336_(_002666_, _002688_, _002690_);
  and g_096337_(_002680_, _002684_, _002691_);
  and g_096338_(_002669_, _002676_, _002692_);
  or g_096339_(_002691_, _002692_, _002693_);
  not g_096340_(_002693_, _002695_);
  and g_096341_(_002649_, _002657_, _002696_);
  not g_096342_(_002696_, _002697_);
  or g_096343_(_002660_, _002664_, _002698_);
  not g_096344_(_002698_, _002699_);
  and g_096345_(_002697_, _002698_, _002700_);
  or g_096346_(_002696_, _002699_, _002701_);
  and g_096347_(_002695_, _002700_, _002702_);
  or g_096348_(_002693_, _002701_, _002703_);
  and g_096349_(_002689_, _002702_, _002704_);
  or g_096350_(_002690_, _002703_, _002706_);
  and g_096351_(_002647_, _002704_, _002707_);
  or g_096352_(_002648_, _002706_, _002708_);
  xor g_096353_(out[931], _025827_, _002709_);
  xor g_096354_(_002144_, _025827_, _002710_);
  and g_096355_(_002526_, _002596_, _002711_);
  not g_096356_(_002711_, _002712_);
  or g_096357_(_002523_, _002596_, _002713_);
  not g_096358_(_002713_, _002714_);
  and g_096359_(_002712_, _002713_, _002715_);
  or g_096360_(_002711_, _002714_, _002717_);
  and g_096361_(_002709_, _002717_, _002718_);
  or g_096362_(out[929], out[930], _002719_);
  xor g_096363_(out[929], out[930], _002720_);
  xor g_096364_(_002111_, out[930], _002721_);
  or g_096365_(_002530_, _002596_, _002722_);
  and g_096366_(_002534_, _002596_, _002723_);
  not g_096367_(_002723_, _002724_);
  and g_096368_(_002722_, _002724_, _002725_);
  and g_096369_(_002721_, _002725_, _002726_);
  or g_096370_(_002718_, _002726_, _002728_);
  or g_096371_(_002709_, _002717_, _002729_);
  xor g_096372_(_002710_, _002715_, _002730_);
  xor g_096373_(_002721_, _002725_, _002731_);
  and g_096374_(_002730_, _002731_, _002732_);
  not g_096375_(_002732_, _002733_);
  or g_096376_(_002001_, _002596_, _002734_);
  or g_096377_(_002548_, _002594_, _002735_);
  and g_096378_(_002734_, _002735_, _002736_);
  and g_096379_(out[929], _002736_, _002737_);
  not g_096380_(_002737_, _002739_);
  and g_096381_(_002553_, _002596_, _002740_);
  not g_096382_(_002740_, _002741_);
  or g_096383_(out[912], _002596_, _002742_);
  not g_096384_(_002742_, _002743_);
  and g_096385_(_002741_, _002742_, _002744_);
  or g_096386_(_002740_, _002743_, _002745_);
  and g_096387_(out[928], _002745_, _002746_);
  or g_096388_(_002122_, _002744_, _002747_);
  xor g_096389_(out[929], _002736_, _002748_);
  xor g_096390_(_002111_, _002736_, _002750_);
  and g_096391_(_002747_, _002748_, _002751_);
  or g_096392_(_002746_, _002750_, _002752_);
  and g_096393_(_002739_, _002752_, _002753_);
  or g_096394_(_002737_, _002751_, _002754_);
  and g_096395_(_002732_, _002754_, _002755_);
  or g_096396_(_002733_, _002753_, _002756_);
  and g_096397_(_002728_, _002729_, _002757_);
  not g_096398_(_002757_, _002758_);
  and g_096399_(_002756_, _002758_, _002759_);
  or g_096400_(_002755_, _002757_, _002761_);
  and g_096401_(_002707_, _002761_, _002762_);
  or g_096402_(_002708_, _002759_, _002763_);
  and g_096403_(_002659_, _002685_, _002764_);
  and g_096404_(_002701_, _002764_, _002765_);
  or g_096405_(_002693_, _002765_, _002766_);
  and g_096406_(_002647_, _002766_, _002767_);
  not g_096407_(_002767_, _002768_);
  and g_096408_(_002678_, _002767_, _002769_);
  or g_096409_(_002677_, _002768_, _002770_);
  or g_096410_(_002605_, _002610_, _002772_);
  not g_096411_(_002772_, _002773_);
  and g_096412_(_002637_, _002640_, _002774_);
  or g_096413_(_002636_, _002638_, _002775_);
  and g_096414_(_002614_, _002774_, _002776_);
  or g_096415_(_002615_, _002775_, _002777_);
  and g_096416_(_002772_, _002777_, _002778_);
  or g_096417_(_002773_, _002776_, _002779_);
  and g_096418_(_002763_, _002778_, _002780_);
  or g_096419_(_002762_, _002779_, _002781_);
  and g_096420_(_002770_, _002780_, _002783_);
  or g_096421_(_002769_, _002781_, _002784_);
  and g_096422_(_002122_, _002744_, _002785_);
  or g_096423_(_002733_, _002785_, _002786_);
  or g_096424_(_002752_, _002786_, _002787_);
  or g_096425_(_002708_, _002787_, _002788_);
  not g_096426_(_002788_, _002789_);
  and g_096427_(_002784_, _002788_, _002790_);
  or g_096428_(_002783_, _002789_, _002791_);
  or g_096429_(_053970_, _002791_, _002792_);
  or g_096430_(_002621_, _002790_, _002794_);
  and g_096431_(_002792_, _002794_, _002795_);
  not g_096432_(_002795_, _002796_);
  and g_096433_(_025970_, _026080_, _002797_);
  or g_096434_(_025959_, _026091_, _002798_);
  xor g_096435_(out[954], _026058_, _002799_);
  not g_096436_(_002799_, _002800_);
  and g_096437_(_002602_, _002791_, _002801_);
  and g_096438_(_053975_, _002790_, _002802_);
  or g_096439_(_002801_, _002802_, _002803_);
  not g_096440_(_002803_, _002805_);
  and g_096441_(_002799_, _002805_, _002806_);
  or g_096442_(_002800_, _002803_, _002807_);
  and g_096443_(_002798_, _002807_, _002808_);
  or g_096444_(_002797_, _002806_, _002809_);
  and g_096445_(_025959_, _026091_, _002810_);
  or g_096446_(_025970_, _026080_, _002811_);
  and g_096447_(_002800_, _002803_, _002812_);
  or g_096448_(_002799_, _002805_, _002813_);
  or g_096449_(_002810_, _002812_, _002814_);
  and g_096450_(_002808_, _002813_, _002816_);
  and g_096451_(_002811_, _002816_, _002817_);
  or g_096452_(_002809_, _002814_, _002818_);
  xor g_096453_(out[953], _026047_, _002819_);
  not g_096454_(_002819_, _002820_);
  and g_096455_(_002796_, _002819_, _002821_);
  or g_096456_(_002795_, _002820_, _002822_);
  and g_096457_(_002632_, _002790_, _002823_);
  not g_096458_(_002823_, _002824_);
  or g_096459_(_002630_, _002790_, _002825_);
  not g_096460_(_002825_, _002827_);
  and g_096461_(_002824_, _002825_, _002828_);
  or g_096462_(_002823_, _002827_, _002829_);
  xor g_096463_(out[952], _026036_, _002830_);
  xor g_096464_(_002265_, _026036_, _002831_);
  and g_096465_(_002828_, _002830_, _002832_);
  or g_096466_(_002829_, _002831_, _002833_);
  and g_096467_(_002822_, _002833_, _002834_);
  or g_096468_(_002821_, _002832_, _002835_);
  and g_096469_(_002795_, _002820_, _002836_);
  or g_096470_(_002796_, _002819_, _002838_);
  and g_096471_(_002829_, _002831_, _002839_);
  or g_096472_(_002828_, _002830_, _002840_);
  and g_096473_(_002838_, _002840_, _002841_);
  or g_096474_(_002836_, _002839_, _002842_);
  and g_096475_(_002834_, _002841_, _002843_);
  or g_096476_(_002835_, _002842_, _002844_);
  and g_096477_(_002817_, _002843_, _002845_);
  or g_096478_(_002818_, _002844_, _002846_);
  xor g_096479_(out[951], _026025_, _002847_);
  xor g_096480_(_002188_, _026025_, _002849_);
  and g_096481_(_002668_, _002790_, _002850_);
  not g_096482_(_002850_, _002851_);
  or g_096483_(_002675_, _002790_, _002852_);
  not g_096484_(_002852_, _002853_);
  and g_096485_(_002851_, _002852_, _002854_);
  or g_096486_(_002850_, _002853_, _002855_);
  and g_096487_(_002849_, _002855_, _002856_);
  or g_096488_(_002847_, _002854_, _002857_);
  xor g_096489_(out[950], _026014_, _002858_);
  not g_096490_(_002858_, _002860_);
  or g_096491_(_002679_, _002791_, _002861_);
  or g_096492_(_002684_, _002790_, _002862_);
  and g_096493_(_002861_, _002862_, _002863_);
  not g_096494_(_002863_, _002864_);
  and g_096495_(_002860_, _002863_, _002865_);
  or g_096496_(_002858_, _002864_, _002866_);
  and g_096497_(_002857_, _002866_, _002867_);
  or g_096498_(_002856_, _002865_, _002868_);
  and g_096499_(_002858_, _002864_, _002869_);
  and g_096500_(_002847_, _002854_, _002871_);
  or g_096501_(_002849_, _002855_, _002872_);
  or g_096502_(_002869_, _002871_, _002873_);
  or g_096503_(_002868_, _002873_, _002874_);
  not g_096504_(_002874_, _002875_);
  xor g_096505_(out[949], _026003_, _002876_);
  xor g_096506_(_002210_, _026003_, _002877_);
  and g_096507_(_002651_, _002790_, _002878_);
  not g_096508_(_002878_, _002879_);
  or g_096509_(_002656_, _002790_, _002880_);
  not g_096510_(_002880_, _002882_);
  and g_096511_(_002879_, _002880_, _002883_);
  or g_096512_(_002878_, _002882_, _002884_);
  and g_096513_(_002877_, _002883_, _002885_);
  or g_096514_(_002876_, _002884_, _002886_);
  and g_096515_(_002876_, _002884_, _002887_);
  or g_096516_(_002877_, _002883_, _002888_);
  or g_096517_(_002885_, _002887_, _002889_);
  xor g_096518_(out[948], _025992_, _002890_);
  not g_096519_(_002890_, _002891_);
  and g_096520_(_002660_, _002790_, _002893_);
  not g_096521_(_002893_, _002894_);
  or g_096522_(_002664_, _002790_, _002895_);
  and g_096523_(_002894_, _002895_, _002896_);
  not g_096524_(_002896_, _002897_);
  and g_096525_(_002890_, _002897_, _002898_);
  or g_096526_(_002891_, _002896_, _002899_);
  xor g_096527_(_002890_, _002896_, _002900_);
  or g_096528_(_002889_, _002900_, _002901_);
  not g_096529_(_002901_, _002902_);
  or g_096530_(out[945], out[946], _002904_);
  xor g_096531_(out[945], out[946], _002905_);
  xor g_096532_(_054336_, out[946], _002906_);
  or g_096533_(_002725_, _002790_, _002907_);
  or g_096534_(_002720_, _002791_, _002908_);
  and g_096535_(_002907_, _002908_, _002909_);
  and g_096536_(_002906_, _002909_, _002910_);
  not g_096537_(_002910_, _002911_);
  xor g_096538_(out[947], _025981_, _002912_);
  not g_096539_(_002912_, _002913_);
  and g_096540_(_002717_, _002791_, _002915_);
  or g_096541_(_002715_, _002790_, _002916_);
  and g_096542_(_002710_, _002790_, _002917_);
  or g_096543_(_002709_, _002791_, _002918_);
  and g_096544_(_002916_, _002918_, _002919_);
  or g_096545_(_002915_, _002917_, _002920_);
  and g_096546_(_002913_, _002919_, _002921_);
  or g_096547_(_002912_, _002920_, _002922_);
  xor g_096548_(_002906_, _002909_, _002923_);
  xor g_096549_(_002905_, _002909_, _002924_);
  and g_096550_(_002922_, _002923_, _002926_);
  or g_096551_(_002921_, _002924_, _002927_);
  or g_096552_(_002913_, _002919_, _002928_);
  not g_096553_(_002928_, _002929_);
  and g_096554_(out[929], _002790_, _002930_);
  or g_096555_(_002736_, _002790_, _002931_);
  not g_096556_(_002931_, _002932_);
  or g_096557_(_002930_, _002932_, _002933_);
  or g_096558_(_054336_, _002933_, _002934_);
  or g_096559_(_002744_, _002790_, _002935_);
  or g_096560_(out[928], _002791_, _002937_);
  and g_096561_(_002935_, _002937_, _002938_);
  not g_096562_(_002938_, _002939_);
  and g_096563_(out[944], _002939_, _002940_);
  or g_096564_(_002232_, _002938_, _002941_);
  xor g_096565_(_054336_, _002933_, _002942_);
  xor g_096566_(out[945], _002933_, _002943_);
  and g_096567_(_002926_, _002928_, _002944_);
  or g_096568_(_002927_, _002929_, _002945_);
  and g_096569_(_002941_, _002942_, _002946_);
  or g_096570_(_002940_, _002943_, _002948_);
  and g_096571_(_002944_, _002946_, _002949_);
  or g_096572_(_002945_, _002948_, _002950_);
  and g_096573_(_002911_, _002928_, _002951_);
  or g_096574_(_002910_, _002929_, _002952_);
  and g_096575_(_002922_, _002952_, _002953_);
  or g_096576_(_002921_, _002951_, _002954_);
  and g_096577_(_002950_, _002954_, _002955_);
  or g_096578_(_002949_, _002953_, _002956_);
  or g_096579_(_002927_, _002934_, _002957_);
  not g_096580_(_002957_, _002959_);
  and g_096581_(_002955_, _002957_, _002960_);
  or g_096582_(_002956_, _002959_, _002961_);
  and g_096583_(_002902_, _002961_, _002962_);
  or g_096584_(_002901_, _002960_, _002963_);
  and g_096585_(_002886_, _002898_, _002964_);
  or g_096586_(_002885_, _002899_, _002965_);
  or g_096587_(_002887_, _002964_, _002966_);
  and g_096588_(_002888_, _002965_, _002967_);
  and g_096589_(_002963_, _002967_, _002968_);
  or g_096590_(_002962_, _002966_, _002970_);
  and g_096591_(_002875_, _002970_, _002971_);
  or g_096592_(_002874_, _002968_, _002972_);
  and g_096593_(_002868_, _002872_, _002973_);
  or g_096594_(_002867_, _002871_, _002974_);
  and g_096595_(_002972_, _002974_, _002975_);
  or g_096596_(_002971_, _002973_, _002976_);
  and g_096597_(_002845_, _002976_, _002977_);
  or g_096598_(_002846_, _002975_, _002978_);
  and g_096599_(_002809_, _002811_, _002979_);
  or g_096600_(_002808_, _002810_, _002981_);
  and g_096601_(_002835_, _002838_, _002982_);
  or g_096602_(_002834_, _002836_, _002983_);
  and g_096603_(_002817_, _002982_, _002984_);
  or g_096604_(_002818_, _002983_, _002985_);
  and g_096605_(_002981_, _002985_, _002986_);
  or g_096606_(_002979_, _002984_, _002987_);
  and g_096607_(_002978_, _002986_, _002988_);
  or g_096608_(_002977_, _002987_, _002989_);
  and g_096609_(_002232_, _002938_, _002990_);
  or g_096610_(_002874_, _002901_, _002992_);
  or g_096611_(_002990_, _002992_, _002993_);
  or g_096612_(_002950_, _002993_, _002994_);
  not g_096613_(_002994_, _002995_);
  and g_096614_(_002845_, _002995_, _002996_);
  or g_096615_(_002846_, _002994_, _002997_);
  and g_096616_(_002989_, _002997_, _002998_);
  or g_096617_(_002988_, _002996_, _002999_);
  or g_096618_(_002795_, _002998_, _003000_);
  or g_096619_(_002819_, _002999_, _003001_);
  and g_096620_(_003000_, _003001_, _003003_);
  or g_096621_(_053897_, _053965_, _003004_);
  or g_096622_(_053892_, _053966_, _003005_);
  and g_096623_(_003004_, _003005_, _003006_);
  or g_096624_(_002919_, _002998_, _003007_);
  or g_096625_(_002912_, _002999_, _003008_);
  and g_096626_(_003007_, _003008_, _003009_);
  and g_096627_(out[465], _053965_, _003010_);
  and g_096628_(_053876_, _053966_, _003011_);
  or g_096629_(_003010_, _003011_, _003012_);
  and g_096630_(out[945], _002998_, _003014_);
  and g_096631_(_002933_, _002999_, _003015_);
  or g_096632_(_003014_, _003015_, _003016_);
  xor g_096633_(_003012_, _003016_, _003017_);
  and g_096634_(_053838_, _053965_, _003018_);
  not g_096635_(_003018_, _003019_);
  and g_096636_(_053845_, _053966_, _003020_);
  or g_096637_(_053844_, _053965_, _003021_);
  and g_096638_(_003019_, _003021_, _003022_);
  or g_096639_(_003018_, _003020_, _003023_);
  and g_096640_(_002876_, _002998_, _003025_);
  or g_096641_(_002877_, _002999_, _003026_);
  and g_096642_(_002883_, _002999_, _003027_);
  not g_096643_(_003027_, _003028_);
  and g_096644_(_003026_, _003028_, _003029_);
  or g_096645_(_003025_, _003027_, _003030_);
  or g_096646_(_053914_, _053965_, _003031_);
  or g_096647_(out[464], _053966_, _003032_);
  and g_096648_(_003031_, _003032_, _003033_);
  or g_096649_(_002938_, _002998_, _003034_);
  or g_096650_(out[944], _002999_, _003036_);
  and g_096651_(_003034_, _003036_, _003037_);
  xor g_096652_(_003033_, _003037_, _003038_);
  and g_096653_(_053774_, _053965_, _003039_);
  or g_096654_(_053776_, _053966_, _003040_);
  and g_096655_(_053773_, _053966_, _003041_);
  or g_096656_(_053772_, _053965_, _003042_);
  and g_096657_(_003040_, _003042_, _003043_);
  or g_096658_(_003039_, _003041_, _003044_);
  and g_096659_(_002830_, _002998_, _003045_);
  or g_096660_(_002831_, _002999_, _003047_);
  and g_096661_(_002829_, _002999_, _003048_);
  or g_096662_(_002828_, _002998_, _003049_);
  and g_096663_(_003047_, _003049_, _003050_);
  or g_096664_(_003045_, _003048_, _003051_);
  and g_096665_(_003043_, _003051_, _003052_);
  and g_096666_(_003044_, _003050_, _003053_);
  or g_096667_(_053881_, _053966_, _003054_);
  or g_096668_(_053886_, _053965_, _003055_);
  and g_096669_(_003054_, _003055_, _003056_);
  and g_096670_(_002905_, _002998_, _003058_);
  and g_096671_(_002909_, _002999_, _003059_);
  or g_096672_(_003058_, _003059_, _003060_);
  or g_096673_(_053827_, _053966_, _003061_);
  or g_096674_(_053833_, _053965_, _003062_);
  and g_096675_(_003061_, _003062_, _003063_);
  or g_096676_(_002891_, _002999_, _003064_);
  or g_096677_(_002897_, _002998_, _003065_);
  and g_096678_(_003064_, _003065_, _003066_);
  and g_096679_(_053816_, _053965_, _003067_);
  or g_096680_(_053817_, _053966_, _003069_);
  and g_096681_(_053824_, _053966_, _003070_);
  or g_096682_(_053823_, _053965_, _003071_);
  and g_096683_(_003069_, _003071_, _003072_);
  or g_096684_(_003067_, _003070_, _003073_);
  and g_096685_(_002847_, _002998_, _003074_);
  or g_096686_(_002849_, _002999_, _003075_);
  and g_096687_(_002855_, _002999_, _003076_);
  or g_096688_(_002854_, _002998_, _003077_);
  and g_096689_(_003075_, _003077_, _003078_);
  or g_096690_(_003074_, _003076_, _003080_);
  and g_096691_(_003072_, _003080_, _003081_);
  or g_096692_(_053811_, _053966_, _003082_);
  or g_096693_(_053815_, _053965_, _003083_);
  and g_096694_(_003082_, _003083_, _003084_);
  or g_096695_(_002863_, _002998_, _003085_);
  or g_096696_(_002858_, _002999_, _003086_);
  and g_096697_(_003085_, _003086_, _003087_);
  and g_096698_(_003073_, _003078_, _003088_);
  or g_096699_(_053760_, _053965_, _003089_);
  or g_096700_(_026157_, _053966_, _003091_);
  and g_096701_(_003089_, _003091_, _003092_);
  or g_096702_(_002805_, _002998_, _003093_);
  or g_096703_(_002800_, _002999_, _003094_);
  and g_096704_(_003093_, _003094_, _003095_);
  or g_096705_(_026113_, _003052_, _003096_);
  or g_096706_(_003053_, _003081_, _003097_);
  or g_096707_(_003096_, _003097_, _003098_);
  and g_096708_(_003022_, _003029_, _003099_);
  and g_096709_(_003023_, _003030_, _003100_);
  or g_096710_(_003088_, _003100_, _003102_);
  or g_096711_(_003099_, _003102_, _003103_);
  or g_096712_(_003098_, _003103_, _003104_);
  xor g_096713_(_003084_, _003087_, _003105_);
  or g_096714_(_003038_, _003105_, _003106_);
  xor g_096715_(_003056_, _003060_, _003107_);
  or g_096716_(_003017_, _003107_, _003108_);
  or g_096717_(_003106_, _003108_, _003109_);
  xor g_096718_(_053969_, _003003_, _003110_);
  xor g_096719_(_003006_, _003009_, _003111_);
  or g_096720_(_003110_, _003111_, _003113_);
  xor g_096721_(_003063_, _003066_, _003114_);
  xor g_096722_(_003092_, _003095_, _003115_);
  or g_096723_(_003114_, _003115_, _003116_);
  or g_096724_(_003113_, _003116_, _003117_);
  or g_096725_(_003109_, _003117_, _003118_);
  or g_096726_(_003104_, _003118_, _003119_);
  not g_096727_(_003119_, _003120_);
  or g_096728_(out[467], _053880_, _003121_);
  not g_096729_(_003121_, _003122_);
  and g_096730_(out[468], _003121_, _003124_);
  or g_096731_(_054292_, _003122_, _003125_);
  and g_096732_(out[469], _003124_, _003126_);
  and g_096733_(out[470], _003126_, _003127_);
  or g_096734_(out[471], _003127_, _003128_);
  xor g_096735_(out[471], _003127_, _003129_);
  xor g_096736_(_054237_, _003127_, _003130_);
  and g_096737_(out[472], _003128_, _003131_);
  or g_096738_(out[473], _003131_, _003132_);
  or g_096739_(out[474], _003132_, _003133_);
  xor g_096740_(out[474], _003132_, _003135_);
  not g_096741_(_003135_, _003136_);
  or g_096742_(out[419], _053270_, _003137_);
  not g_096743_(_003137_, _003138_);
  and g_096744_(out[420], _003137_, _003139_);
  or g_096745_(_053995_, _003138_, _003140_);
  and g_096746_(out[421], _003139_, _003141_);
  and g_096747_(out[422], _003141_, _003142_);
  or g_096748_(out[423], _003142_, _003143_);
  and g_096749_(out[424], _003143_, _003144_);
  or g_096750_(out[425], _003144_, _003146_);
  not g_096751_(_003146_, _003147_);
  or g_096752_(out[426], _003146_, _003148_);
  xor g_096753_(out[426], _003146_, _003149_);
  xor g_096754_(_004751_, _003146_, _003150_);
  or g_096755_(out[3], _005851_, _003151_);
  and g_096756_(out[4], _003151_, _003152_);
  not g_096757_(_003152_, _003153_);
  and g_096758_(out[5], _003152_, _003154_);
  and g_096759_(out[6], _003154_, _003155_);
  or g_096760_(out[7], _003155_, _003157_);
  and g_096761_(out[8], _003157_, _003158_);
  or g_096762_(out[9], _003158_, _003159_);
  or g_096763_(out[10], _003159_, _003160_);
  xor g_096764_(out[11], _003160_, _003161_);
  xor g_096765_(_002298_, _003160_, _003162_);
  or g_096766_(out[19], _005818_, _003163_);
  and g_096767_(out[20], _003163_, _003164_);
  not g_096768_(_003164_, _003165_);
  and g_096769_(out[21], _003164_, _003166_);
  and g_096770_(out[22], _003166_, _003168_);
  or g_096771_(out[23], _003168_, _003169_);
  and g_096772_(out[24], _003169_, _003170_);
  or g_096773_(out[25], _003170_, _003171_);
  or g_096774_(out[26], _003171_, _003172_);
  xor g_096775_(out[27], _003172_, _003173_);
  xor g_096776_(_002430_, _003172_, _003174_);
  and g_096777_(_003161_, _003173_, _003175_);
  or g_096778_(_003162_, _003174_, _003176_);
  or g_096779_(out[35], _007831_, _003177_);
  not g_096780_(_003177_, _003179_);
  and g_096781_(out[36], _003177_, _003180_);
  or g_096782_(_002606_, _003179_, _003181_);
  and g_096783_(out[37], _003180_, _003182_);
  and g_096784_(out[38], _003182_, _003183_);
  or g_096785_(out[39], _003183_, _003184_);
  and g_096786_(out[40], _003184_, _003185_);
  or g_096787_(out[41], _003185_, _003186_);
  not g_096788_(_003186_, _003187_);
  or g_096789_(out[42], _003186_, _003188_);
  xor g_096790_(out[43], _003188_, _003190_);
  xor g_096791_(_002562_, _003188_, _003191_);
  and g_096792_(_003175_, _003190_, _003192_);
  or g_096793_(_003176_, _003191_, _003193_);
  or g_096794_(out[51], _010823_, _003194_);
  not g_096795_(_003194_, _003195_);
  and g_096796_(out[52], _003194_, _003196_);
  or g_096797_(_002738_, _003195_, _003197_);
  and g_096798_(out[53], _003196_, _003198_);
  and g_096799_(out[54], _003198_, _003199_);
  or g_096800_(out[55], _003199_, _003201_);
  and g_096801_(out[56], _003201_, _003202_);
  or g_096802_(out[57], _003202_, _003203_);
  not g_096803_(_003203_, _003204_);
  or g_096804_(out[58], _003203_, _003205_);
  xor g_096805_(out[59], _003205_, _003206_);
  xor g_096806_(_002694_, _003205_, _003207_);
  and g_096807_(_003192_, _003206_, _003208_);
  or g_096808_(_003193_, _003207_, _003209_);
  or g_096809_(out[67], _026608_, _003210_);
  not g_096810_(_003210_, _003212_);
  and g_096811_(out[68], _003210_, _003213_);
  or g_096812_(_002870_, _003212_, _003214_);
  and g_096813_(out[69], _003213_, _003215_);
  and g_096814_(out[70], _003215_, _003216_);
  or g_096815_(out[71], _003216_, _003217_);
  and g_096816_(out[72], _003217_, _003218_);
  or g_096817_(out[73], _003218_, _003219_);
  not g_096818_(_003219_, _003220_);
  or g_096819_(out[74], _003219_, _003221_);
  xor g_096820_(out[75], _003221_, _003223_);
  xor g_096821_(_002826_, _003221_, _003224_);
  and g_096822_(_003208_, _003223_, _003225_);
  or g_096823_(_003209_, _003224_, _003226_);
  or g_096824_(out[83], _026575_, _003227_);
  not g_096825_(_003227_, _003228_);
  and g_096826_(out[84], _003227_, _003229_);
  or g_096827_(_003002_, _003228_, _003230_);
  and g_096828_(out[85], _003229_, _003231_);
  and g_096829_(out[86], _003231_, _003232_);
  or g_096830_(out[87], _003232_, _003234_);
  and g_096831_(out[88], _003234_, _003235_);
  or g_096832_(out[89], _003235_, _003236_);
  not g_096833_(_003236_, _003237_);
  or g_096834_(out[90], _003236_, _003238_);
  xor g_096835_(out[91], _003238_, _003239_);
  xor g_096836_(_002958_, _003238_, _003240_);
  and g_096837_(_003225_, _003239_, _003241_);
  or g_096838_(_003226_, _003240_, _003242_);
  or g_096839_(out[99], _031195_, _003243_);
  not g_096840_(_003243_, _003245_);
  and g_096841_(out[100], _003243_, _003246_);
  or g_096842_(_003134_, _003245_, _003247_);
  and g_096843_(out[101], _003246_, _003248_);
  and g_096844_(out[102], _003248_, _003249_);
  or g_096845_(out[103], _003249_, _003250_);
  and g_096846_(out[104], _003250_, _003251_);
  or g_096847_(out[105], _003251_, _003252_);
  not g_096848_(_003252_, _003253_);
  or g_096849_(out[106], _003252_, _003254_);
  xor g_096850_(out[107], _003254_, _003256_);
  xor g_096851_(_003090_, _003254_, _003257_);
  and g_096852_(_003241_, _003256_, _003258_);
  or g_096853_(_003242_, _003257_, _003259_);
  or g_096854_(out[115], _034110_, _003260_);
  not g_096855_(_003260_, _003261_);
  and g_096856_(out[116], _003260_, _003262_);
  or g_096857_(_003266_, _003261_, _003263_);
  and g_096858_(out[117], _003262_, _003264_);
  and g_096859_(out[118], _003264_, _003265_);
  or g_096860_(out[119], _003265_, _003267_);
  and g_096861_(out[120], _003267_, _003268_);
  or g_096862_(out[121], _003268_, _003269_);
  not g_096863_(_003269_, _003270_);
  or g_096864_(out[122], _003269_, _003271_);
  xor g_096865_(out[123], _003271_, _003272_);
  xor g_096866_(_003222_, _003271_, _003273_);
  and g_096867_(_003258_, _003272_, _003274_);
  or g_096868_(_003259_, _003273_, _003275_);
  or g_096869_(out[131], _036178_, _003276_);
  not g_096870_(_003276_, _003278_);
  and g_096871_(out[132], _003276_, _003279_);
  or g_096872_(_003398_, _003278_, _003280_);
  and g_096873_(out[133], _003279_, _003281_);
  and g_096874_(out[134], _003281_, _003282_);
  or g_096875_(out[135], _003282_, _003283_);
  and g_096876_(out[136], _003283_, _003284_);
  or g_096877_(out[137], _003284_, _003285_);
  not g_096878_(_003285_, _003286_);
  or g_096879_(out[138], _003285_, _003287_);
  xor g_096880_(out[139], _003287_, _003289_);
  xor g_096881_(_003354_, _003287_, _003290_);
  and g_096882_(_003274_, _003289_, _003291_);
  or g_096883_(_003275_, _003290_, _003292_);
  or g_096884_(out[147], _038455_, _003293_);
  not g_096885_(_003293_, _003294_);
  and g_096886_(out[148], _003293_, _003295_);
  or g_096887_(_003530_, _003294_, _003296_);
  and g_096888_(out[149], _003295_, _003297_);
  and g_096889_(out[150], _003297_, _003298_);
  or g_096890_(out[151], _003298_, _003300_);
  and g_096891_(out[152], _003300_, _003301_);
  or g_096892_(out[153], _003301_, _003302_);
  not g_096893_(_003302_, _003303_);
  or g_096894_(out[154], _003302_, _003304_);
  xor g_096895_(out[155], _003304_, _003305_);
  xor g_096896_(_003486_, _003304_, _003306_);
  and g_096897_(_003291_, _003305_, _003307_);
  or g_096898_(_003292_, _003306_, _003308_);
  or g_096899_(out[163], _040556_, _003309_);
  not g_096900_(_003309_, _003311_);
  and g_096901_(out[164], _003309_, _003312_);
  or g_096902_(_003662_, _003311_, _003313_);
  and g_096903_(out[165], _003312_, _003314_);
  and g_096904_(out[166], _003314_, _003315_);
  or g_096905_(out[167], _003315_, _003316_);
  and g_096906_(out[168], _003316_, _003317_);
  or g_096907_(out[169], _003317_, _003318_);
  or g_096908_(out[170], _003318_, _003319_);
  xor g_096909_(out[171], _003319_, _003320_);
  xor g_096910_(_003618_, _003319_, _003322_);
  and g_096911_(_003307_, _003320_, _003323_);
  or g_096912_(_003308_, _003322_, _003324_);
  or g_096913_(out[179], _042679_, _003325_);
  not g_096914_(_003325_, _003326_);
  and g_096915_(out[180], _003325_, _003327_);
  or g_096916_(_003794_, _003326_, _003328_);
  and g_096917_(out[181], _003327_, _003329_);
  and g_096918_(out[182], _003329_, _003330_);
  or g_096919_(out[183], _003330_, _003331_);
  and g_096920_(out[184], _003331_, _003333_);
  or g_096921_(out[185], _003333_, _003334_);
  not g_096922_(_003334_, _003335_);
  or g_096923_(out[186], _003334_, _003336_);
  xor g_096924_(out[187], _003336_, _003337_);
  xor g_096925_(_003750_, _003336_, _003338_);
  and g_096926_(_003323_, _003337_, _003339_);
  or g_096927_(_003324_, _003338_, _003340_);
  or g_096928_(out[195], _044516_, _003341_);
  not g_096929_(_003341_, _003342_);
  and g_096930_(out[196], _003341_, _003344_);
  or g_096931_(_003926_, _003342_, _003345_);
  and g_096932_(out[197], _003344_, _003346_);
  and g_096933_(out[198], _003346_, _003347_);
  or g_096934_(out[199], _003347_, _003348_);
  and g_096935_(out[200], _003348_, _003349_);
  or g_096936_(out[201], _003349_, _003350_);
  not g_096937_(_003350_, _003351_);
  or g_096938_(out[202], _003350_, _003352_);
  xor g_096939_(out[203], _003352_, _003353_);
  not g_096940_(_003353_, _003355_);
  and g_096941_(_003339_, _003353_, _003356_);
  or g_096942_(_003340_, _003355_, _003357_);
  or g_096943_(out[211], _046870_, _003358_);
  and g_096944_(out[212], _003358_, _003359_);
  and g_096945_(out[213], _003359_, _003360_);
  and g_096946_(out[214], _003360_, _003361_);
  or g_096947_(out[215], _003361_, _003362_);
  and g_096948_(out[216], _003362_, _003363_);
  or g_096949_(out[217], _003363_, _003364_);
  not g_096950_(_003364_, _003366_);
  or g_096951_(out[218], _003364_, _003367_);
  xor g_096952_(out[219], _003367_, _003368_);
  xor g_096953_(_003992_, _003367_, _003369_);
  and g_096954_(_003356_, _003368_, _003370_);
  or g_096955_(_003357_, _003369_, _003371_);
  or g_096956_(out[227], _047805_, _003372_);
  not g_096957_(_003372_, _003373_);
  and g_096958_(out[228], _003372_, _003374_);
  or g_096959_(_004168_, _003373_, _003375_);
  and g_096960_(out[229], _003374_, _003377_);
  and g_096961_(out[230], _003377_, _003378_);
  or g_096962_(out[231], _003378_, _003379_);
  and g_096963_(out[232], _003379_, _003380_);
  or g_096964_(out[233], _003380_, _003381_);
  not g_096965_(_003381_, _003382_);
  or g_096966_(out[234], _003381_, _003383_);
  xor g_096967_(out[235], _003383_, _003384_);
  xor g_096968_(_004124_, _003383_, _003385_);
  and g_096969_(_003370_, _003384_, _003386_);
  or g_096970_(_003371_, _003385_, _003388_);
  or g_096971_(out[243], _050467_, _003389_);
  and g_096972_(out[244], _003389_, _003390_);
  and g_096973_(out[245], _003390_, _003391_);
  and g_096974_(out[246], _003391_, _003392_);
  or g_096975_(out[247], _003392_, _003393_);
  and g_096976_(out[248], _003393_, _003394_);
  or g_096977_(out[249], _003394_, _003395_);
  not g_096978_(_003395_, _003396_);
  or g_096979_(out[250], _003395_, _003397_);
  xor g_096980_(out[251], _003397_, _003399_);
  xor g_096981_(_004245_, _003397_, _003400_);
  and g_096982_(_003386_, _003399_, _003401_);
  or g_096983_(_003388_, _003400_, _003402_);
  or g_096984_(out[259], _051425_, _003403_);
  and g_096985_(out[260], _003403_, _003404_);
  and g_096986_(out[261], _003404_, _003405_);
  and g_096987_(out[262], _003405_, _003406_);
  or g_096988_(out[263], _003406_, _003407_);
  and g_096989_(out[264], _003407_, _003408_);
  or g_096990_(out[265], _003408_, _003410_);
  not g_096991_(_003410_, _003411_);
  or g_096992_(out[266], _003410_, _003412_);
  xor g_096993_(out[267], _003412_, _003413_);
  xor g_096994_(_004366_, _003412_, _003414_);
  and g_096995_(_003401_, _003413_, _003415_);
  or g_096996_(_003402_, _003414_, _003416_);
  or g_096997_(out[275], _051640_, _003417_);
  not g_096998_(_003417_, _003418_);
  and g_096999_(out[276], _003417_, _003419_);
  or g_097000_(_053104_, _003418_, _003421_);
  and g_097001_(out[277], _003419_, _003422_);
  and g_097002_(out[278], _003422_, _003423_);
  or g_097003_(out[279], _003423_, _003424_);
  and g_097004_(out[280], _003424_, _003425_);
  or g_097005_(out[281], _003425_, _003426_);
  not g_097006_(_003426_, _003427_);
  or g_097007_(out[282], _003426_, _003428_);
  xor g_097008_(out[283], _003428_, _003429_);
  xor g_097009_(_004432_, _003428_, _003430_);
  and g_097010_(_003415_, _003429_, _003432_);
  or g_097011_(_003416_, _003430_, _003433_);
  or g_097012_(out[291], _051815_, _003434_);
  not g_097013_(_003434_, _003435_);
  and g_097014_(out[292], _003434_, _003436_);
  or g_097015_(_053203_, _003435_, _003437_);
  and g_097016_(out[293], _003436_, _003438_);
  and g_097017_(out[294], _003438_, _003439_);
  or g_097018_(out[295], _003439_, _003440_);
  and g_097019_(out[296], _003440_, _003441_);
  or g_097020_(out[297], _003441_, _003443_);
  or g_097021_(out[298], _003443_, _003444_);
  xor g_097022_(out[299], _003444_, _003445_);
  xor g_097023_(_004465_, _003444_, _003446_);
  and g_097024_(_003432_, _003445_, _003447_);
  or g_097025_(_003433_, _003446_, _003448_);
  or g_097026_(out[307], _051956_, _003449_);
  and g_097027_(out[308], _003449_, _003450_);
  and g_097028_(out[309], _003450_, _003451_);
  and g_097029_(out[310], _003451_, _003452_);
  or g_097030_(out[311], _003452_, _003454_);
  and g_097031_(out[312], _003454_, _003455_);
  or g_097032_(out[313], _003455_, _003456_);
  or g_097033_(out[314], _003456_, _003457_);
  xor g_097034_(out[315], _003457_, _003458_);
  xor g_097035_(_004498_, _003457_, _003459_);
  and g_097036_(_003447_, _003458_, _003460_);
  or g_097037_(_003448_, _003459_, _003461_);
  or g_097038_(out[323], _052166_, _003462_);
  not g_097039_(_003462_, _003463_);
  and g_097040_(out[324], _003462_, _003465_);
  or g_097041_(_053401_, _003463_, _003466_);
  and g_097042_(out[325], _003465_, _003467_);
  and g_097043_(out[326], _003467_, _003468_);
  or g_097044_(out[327], _003468_, _003469_);
  and g_097045_(out[328], _003469_, _003470_);
  or g_097046_(out[329], _003470_, _003471_);
  not g_097047_(_003471_, _003472_);
  or g_097048_(out[330], _003471_, _003473_);
  xor g_097049_(out[331], _003473_, _003474_);
  xor g_097050_(_004531_, _003473_, _003476_);
  and g_097051_(_003460_, _003474_, _003477_);
  or g_097052_(_003461_, _003476_, _003478_);
  or g_097053_(out[339], _052353_, _003479_);
  not g_097054_(_003479_, _003480_);
  and g_097055_(out[340], _003479_, _003481_);
  or g_097056_(_053500_, _003480_, _003482_);
  and g_097057_(out[341], _003481_, _003483_);
  and g_097058_(out[342], _003483_, _003484_);
  or g_097059_(out[343], _003484_, _003485_);
  and g_097060_(out[344], _003485_, _003487_);
  or g_097061_(out[345], _003487_, _003488_);
  not g_097062_(_003488_, _003489_);
  or g_097063_(out[346], _003488_, _003490_);
  xor g_097064_(out[347], _003490_, _003491_);
  xor g_097065_(_004564_, _003490_, _003492_);
  and g_097066_(_003477_, _003491_, _003493_);
  or g_097067_(_003478_, _003492_, _003494_);
  or g_097068_(out[355], _052547_, _003495_);
  not g_097069_(_003495_, _003496_);
  and g_097070_(out[356], _003495_, _003498_);
  or g_097071_(_053599_, _003496_, _003499_);
  and g_097072_(out[357], _003498_, _003500_);
  and g_097073_(out[358], _003500_, _003501_);
  or g_097074_(out[359], _003501_, _003502_);
  and g_097075_(out[360], _003502_, _003503_);
  or g_097076_(out[361], _003503_, _003504_);
  or g_097077_(out[362], _003504_, _003505_);
  xor g_097078_(out[363], _003505_, _003506_);
  xor g_097079_(_004597_, _003505_, _003507_);
  and g_097080_(_003493_, _003506_, _003509_);
  or g_097081_(_003494_, _003507_, _003510_);
  or g_097082_(out[371], _052741_, _003511_);
  not g_097083_(_003511_, _003512_);
  and g_097084_(out[372], _003511_, _003513_);
  or g_097085_(_053698_, _003512_, _003514_);
  and g_097086_(out[373], _003513_, _003515_);
  and g_097087_(out[374], _003515_, _003516_);
  or g_097088_(out[375], _003516_, _003517_);
  and g_097089_(out[376], _003517_, _003518_);
  or g_097090_(out[377], _003518_, _003520_);
  not g_097091_(_003520_, _003521_);
  or g_097092_(out[378], _003520_, _003522_);
  xor g_097093_(out[379], _003522_, _003523_);
  xor g_097094_(_004630_, _003522_, _003524_);
  and g_097095_(_003509_, _003523_, _003525_);
  or g_097096_(_003510_, _003524_, _003526_);
  or g_097097_(out[387], _052921_, _003527_);
  not g_097098_(_003527_, _003528_);
  and g_097099_(out[388], _003527_, _003529_);
  or g_097100_(_053797_, _003528_, _003531_);
  and g_097101_(out[389], _003529_, _003532_);
  and g_097102_(out[390], _003532_, _003533_);
  or g_097103_(out[391], _003533_, _003534_);
  and g_097104_(out[392], _003534_, _003535_);
  or g_097105_(out[393], _003535_, _003536_);
  or g_097106_(out[394], _003536_, _003537_);
  xor g_097107_(out[395], _003537_, _003538_);
  not g_097108_(_003538_, _003539_);
  and g_097109_(_003525_, _003538_, _003540_);
  or g_097110_(_003526_, _003539_, _003542_);
  or g_097111_(out[403], _053009_, _003543_);
  not g_097112_(_003543_, _003544_);
  and g_097113_(out[404], _003543_, _003545_);
  or g_097114_(_053896_, _003544_, _003546_);
  and g_097115_(out[405], _003545_, _003547_);
  and g_097116_(out[406], _003547_, _003548_);
  or g_097117_(out[407], _003548_, _003549_);
  and g_097118_(out[408], _003549_, _003550_);
  or g_097119_(out[409], _003550_, _003551_);
  or g_097120_(out[410], _003551_, _003553_);
  xor g_097121_(out[411], _003553_, _003554_);
  xor g_097122_(_004696_, _003553_, _003555_);
  and g_097123_(_003540_, _003554_, _003556_);
  or g_097124_(_003542_, _003555_, _003557_);
  xor g_097125_(out[427], _003148_, _003558_);
  xor g_097126_(_004729_, _003148_, _003559_);
  and g_097127_(_003556_, _003559_, _003560_);
  or g_097128_(_003557_, _003558_, _003561_);
  xor g_097129_(out[250], _003395_, _003562_);
  xor g_097130_(_004355_, _003395_, _003564_);
  xor g_097131_(out[106], _003252_, _003565_);
  xor g_097132_(_003211_, _003252_, _003566_);
  and g_097133_(_003161_, _003174_, _003567_);
  or g_097134_(_003162_, _003173_, _003568_);
  xor g_097135_(out[10], _003159_, _003569_);
  xor g_097136_(_002419_, _003159_, _003570_);
  xor g_097137_(out[26], _003171_, _003571_);
  not g_097138_(_003571_, _003572_);
  and g_097139_(_003570_, _003571_, _003573_);
  or g_097140_(_003569_, _003572_, _003575_);
  and g_097141_(_003568_, _003575_, _003576_);
  or g_097142_(_003567_, _003573_, _003577_);
  and g_097143_(_003162_, _003173_, _003578_);
  or g_097144_(_003161_, _003174_, _003579_);
  and g_097145_(_003569_, _003572_, _003580_);
  or g_097146_(_003570_, _003571_, _003581_);
  and g_097147_(_003579_, _003581_, _003582_);
  or g_097148_(_003578_, _003580_, _003583_);
  and g_097149_(_003576_, _003582_, _003584_);
  or g_097150_(_003577_, _003583_, _003586_);
  and g_097151_(out[9], _003158_, _003587_);
  xor g_097152_(out[9], _003158_, _003588_);
  xor g_097153_(_002408_, _003158_, _003589_);
  and g_097154_(out[25], _003170_, _003590_);
  xor g_097155_(out[25], _003170_, _003591_);
  xor g_097156_(_002540_, _003170_, _003592_);
  and g_097157_(_003588_, _003592_, _003593_);
  or g_097158_(_003589_, _003591_, _003594_);
  and g_097159_(_003589_, _003591_, _003595_);
  or g_097160_(_003588_, _003592_, _003597_);
  and g_097161_(_003594_, _003597_, _003598_);
  or g_097162_(_003593_, _003595_, _003599_);
  xor g_097163_(out[8], _003157_, _003600_);
  xor g_097164_(_002397_, _003157_, _003601_);
  xor g_097165_(out[24], _003169_, _003602_);
  xor g_097166_(_002529_, _003169_, _003603_);
  and g_097167_(_003600_, _003603_, _003604_);
  or g_097168_(_003601_, _003602_, _003605_);
  xor g_097169_(_003601_, _003602_, _003606_);
  xor g_097170_(_003600_, _003602_, _003608_);
  and g_097171_(_003598_, _003606_, _003609_);
  or g_097172_(_003599_, _003608_, _003610_);
  and g_097173_(_003584_, _003609_, _003611_);
  or g_097174_(_003586_, _003610_, _003612_);
  xor g_097175_(out[7], _003155_, _003613_);
  xor g_097176_(_002309_, _003155_, _003614_);
  xor g_097177_(out[23], _003168_, _003615_);
  xor g_097178_(_002441_, _003168_, _003616_);
  and g_097179_(_003614_, _003615_, _003617_);
  or g_097180_(_003613_, _003616_, _003619_);
  xor g_097181_(out[6], _003154_, _003620_);
  xor g_097182_(_002320_, _003154_, _003621_);
  xor g_097183_(out[22], _003166_, _003622_);
  xor g_097184_(_002452_, _003166_, _003623_);
  and g_097185_(_003620_, _003623_, _003624_);
  or g_097186_(_003621_, _003622_, _003625_);
  and g_097187_(_003619_, _003625_, _003626_);
  or g_097188_(_003617_, _003624_, _003627_);
  and g_097189_(_003621_, _003622_, _003628_);
  or g_097190_(_003620_, _003623_, _003630_);
  and g_097191_(_003613_, _003616_, _003631_);
  or g_097192_(_003614_, _003615_, _003632_);
  and g_097193_(_003630_, _003632_, _003633_);
  or g_097194_(_003628_, _003631_, _003634_);
  and g_097195_(_003626_, _003633_, _003635_);
  or g_097196_(_003627_, _003634_, _003636_);
  or g_097197_(_005301_, _005851_, _003637_);
  not g_097198_(_003637_, _003638_);
  and g_097199_(_003153_, _003637_, _003639_);
  or g_097200_(_003152_, _003638_, _003641_);
  or g_097201_(_005466_, _005818_, _003642_);
  not g_097202_(_003642_, _003643_);
  and g_097203_(_003165_, _003642_, _003644_);
  or g_097204_(_003164_, _003643_, _003645_);
  and g_097205_(_003639_, _003645_, _003646_);
  or g_097206_(_003641_, _003644_, _003647_);
  xor g_097207_(out[5], _003152_, _003648_);
  xor g_097208_(_002331_, _003152_, _003649_);
  xor g_097209_(out[21], _003164_, _003650_);
  xor g_097210_(_002463_, _003164_, _003652_);
  and g_097211_(_003648_, _003652_, _003653_);
  or g_097212_(_003649_, _003650_, _003654_);
  and g_097213_(_003647_, _003654_, _003655_);
  or g_097214_(_003646_, _003653_, _003656_);
  and g_097215_(_003649_, _003650_, _003657_);
  or g_097216_(_003648_, _003652_, _003658_);
  and g_097217_(_003641_, _003644_, _003659_);
  or g_097218_(_003639_, _003645_, _003660_);
  and g_097219_(_003658_, _003660_, _003661_);
  or g_097220_(_003657_, _003659_, _003663_);
  and g_097221_(_003655_, _003661_, _003664_);
  or g_097222_(_003656_, _003663_, _003665_);
  and g_097223_(_003635_, _003664_, _003666_);
  or g_097224_(_003636_, _003665_, _003667_);
  and g_097225_(_006313_, _003666_, _003668_);
  or g_097226_(_006324_, _003667_, _003669_);
  and g_097227_(_003611_, _003668_, _003670_);
  or g_097228_(_003612_, _003669_, _003671_);
  xor g_097229_(out[3], _005851_, _003672_);
  xor g_097230_(out[19], _005818_, _003674_);
  xor g_097231_(_002518_, _005818_, _003675_);
  and g_097232_(_003672_, _003675_, _003676_);
  or g_097233_(_003672_, _003675_, _003677_);
  and g_097234_(_005906_, _003677_, _003678_);
  or g_097235_(_003676_, _003678_, _003679_);
  and g_097236_(_006126_, _003679_, _003680_);
  not g_097237_(_003680_, _003681_);
  and g_097238_(_003666_, _003681_, _003682_);
  or g_097239_(_003667_, _003680_, _003683_);
  and g_097240_(_003656_, _003658_, _003685_);
  or g_097241_(_003655_, _003657_, _003686_);
  and g_097242_(_003635_, _003685_, _003687_);
  or g_097243_(_003636_, _003686_, _003688_);
  and g_097244_(_003627_, _003632_, _003689_);
  or g_097245_(_003626_, _003631_, _003690_);
  and g_097246_(_003688_, _003690_, _003691_);
  or g_097247_(_003687_, _003689_, _003692_);
  and g_097248_(_003683_, _003691_, _003693_);
  or g_097249_(_003682_, _003692_, _003694_);
  and g_097250_(_003611_, _003694_, _003696_);
  or g_097251_(_003612_, _003693_, _003697_);
  and g_097252_(_003598_, _003604_, _003698_);
  or g_097253_(_003599_, _003605_, _003699_);
  and g_097254_(_003597_, _003699_, _003700_);
  or g_097255_(_003595_, _003698_, _003701_);
  and g_097256_(_003584_, _003701_, _003702_);
  or g_097257_(_003586_, _003700_, _003703_);
  and g_097258_(_003577_, _003579_, _003704_);
  or g_097259_(_003576_, _003578_, _003705_);
  and g_097260_(_003703_, _003705_, _003707_);
  or g_097261_(_003702_, _003704_, _003708_);
  and g_097262_(_003697_, _003707_, _003709_);
  or g_097263_(_003696_, _003708_, _003710_);
  and g_097264_(_003671_, _003710_, _003711_);
  or g_097265_(_003670_, _003709_, _003712_);
  and g_097266_(_005862_, _003712_, _003713_);
  and g_097267_(_005829_, _003711_, _003714_);
  or g_097268_(_003713_, _003714_, _003715_);
  not g_097269_(_003715_, _003716_);
  and g_097270_(out[41], _003185_, _003718_);
  xor g_097271_(out[41], _003185_, _003719_);
  or g_097272_(_003187_, _003718_, _003720_);
  and g_097273_(_003588_, _003712_, _003721_);
  or g_097274_(_003589_, _003711_, _003722_);
  and g_097275_(_003591_, _003711_, _003723_);
  or g_097276_(_003592_, _003712_, _003724_);
  and g_097277_(_003722_, _003724_, _003725_);
  or g_097278_(_003721_, _003723_, _003726_);
  and g_097279_(_003719_, _003725_, _003727_);
  or g_097280_(_003720_, _003726_, _003729_);
  xor g_097281_(out[40], _003184_, _003730_);
  xor g_097282_(_002661_, _003184_, _003731_);
  or g_097283_(_003602_, _003712_, _003732_);
  not g_097284_(_003732_, _003733_);
  and g_097285_(_003601_, _003712_, _003734_);
  or g_097286_(_003600_, _003711_, _003735_);
  and g_097287_(_003732_, _003735_, _003736_);
  or g_097288_(_003733_, _003734_, _003737_);
  and g_097289_(_003731_, _003736_, _003738_);
  or g_097290_(_003730_, _003737_, _003740_);
  and g_097291_(_003729_, _003740_, _003741_);
  or g_097292_(_003727_, _003738_, _003742_);
  and g_097293_(_003720_, _003726_, _003743_);
  or g_097294_(_003719_, _003725_, _003744_);
  and g_097295_(_003730_, _003737_, _003745_);
  or g_097296_(_003731_, _003736_, _003746_);
  and g_097297_(_003744_, _003746_, _003747_);
  or g_097298_(_003743_, _003745_, _003748_);
  and g_097299_(_003741_, _003747_, _003749_);
  or g_097300_(_003742_, _003748_, _003751_);
  and g_097301_(_003175_, _003191_, _003752_);
  or g_097302_(_003176_, _003190_, _003753_);
  and g_097303_(_003569_, _003712_, _003754_);
  or g_097304_(_003570_, _003711_, _003755_);
  and g_097305_(_003571_, _003711_, _003756_);
  or g_097306_(_003572_, _003712_, _003757_);
  and g_097307_(_003755_, _003757_, _003758_);
  or g_097308_(_003754_, _003756_, _003759_);
  xor g_097309_(out[42], _003186_, _003760_);
  xor g_097310_(_002683_, _003186_, _003762_);
  and g_097311_(_003758_, _003760_, _003763_);
  or g_097312_(_003759_, _003762_, _003764_);
  and g_097313_(_003753_, _003764_, _003765_);
  or g_097314_(_003752_, _003763_, _003766_);
  and g_097315_(_003176_, _003190_, _003767_);
  or g_097316_(_003175_, _003191_, _003768_);
  and g_097317_(_003759_, _003762_, _003769_);
  or g_097318_(_003758_, _003760_, _003770_);
  and g_097319_(_003768_, _003770_, _003771_);
  or g_097320_(_003767_, _003769_, _003773_);
  and g_097321_(_003765_, _003771_, _003774_);
  or g_097322_(_003766_, _003773_, _003775_);
  and g_097323_(_003749_, _003774_, _003776_);
  or g_097324_(_003751_, _003775_, _003777_);
  and g_097325_(_007842_, _003716_, _003778_);
  or g_097326_(_007853_, _003715_, _003779_);
  xor g_097327_(out[35], _007831_, _003780_);
  xor g_097328_(_002650_, _007831_, _003781_);
  and g_097329_(_003672_, _003712_, _003782_);
  not g_097330_(_003782_, _003784_);
  and g_097331_(_003674_, _003711_, _003785_);
  or g_097332_(_003675_, _003712_, _003786_);
  and g_097333_(_003784_, _003786_, _003787_);
  or g_097334_(_003782_, _003785_, _003788_);
  and g_097335_(_003780_, _003787_, _003789_);
  or g_097336_(_003781_, _003788_, _003790_);
  and g_097337_(_003779_, _003790_, _003791_);
  or g_097338_(_003778_, _003789_, _003792_);
  or g_097339_(_002485_, _003712_, _003793_);
  or g_097340_(_002353_, _003711_, _003795_);
  and g_097341_(_003793_, _003795_, _003796_);
  and g_097342_(out[33], _003796_, _003797_);
  not g_097343_(_003797_, _003798_);
  and g_097344_(_002364_, _003712_, _003799_);
  or g_097345_(out[0], _003711_, _003800_);
  and g_097346_(_002496_, _003711_, _003801_);
  or g_097347_(out[16], _003712_, _003802_);
  and g_097348_(_003800_, _003802_, _003803_);
  or g_097349_(_003799_, _003801_, _003804_);
  and g_097350_(out[32], _003804_, _003806_);
  or g_097351_(_002628_, _003803_, _003807_);
  xor g_097352_(out[33], _003796_, _003808_);
  xor g_097353_(_002617_, _003796_, _003809_);
  and g_097354_(_003807_, _003808_, _003810_);
  or g_097355_(_003806_, _003809_, _003811_);
  and g_097356_(_003798_, _003811_, _003812_);
  or g_097357_(_003797_, _003810_, _003813_);
  xor g_097358_(_007853_, _003715_, _003814_);
  xor g_097359_(_007842_, _003715_, _003815_);
  and g_097360_(_003813_, _003814_, _003817_);
  or g_097361_(_003812_, _003815_, _003818_);
  and g_097362_(_003791_, _003818_, _003819_);
  or g_097363_(_003792_, _003817_, _003820_);
  xor g_097364_(out[38], _003182_, _003821_);
  xor g_097365_(_002584_, _003182_, _003822_);
  and g_097366_(_003621_, _003712_, _003823_);
  or g_097367_(_003620_, _003711_, _003824_);
  and g_097368_(_003623_, _003711_, _003825_);
  or g_097369_(_003622_, _003712_, _003826_);
  and g_097370_(_003824_, _003826_, _003828_);
  or g_097371_(_003823_, _003825_, _003829_);
  and g_097372_(_003822_, _003828_, _003830_);
  or g_097373_(_003821_, _003829_, _003831_);
  xor g_097374_(out[39], _003183_, _003832_);
  xor g_097375_(_002573_, _003183_, _003833_);
  and g_097376_(_003613_, _003712_, _003834_);
  or g_097377_(_003614_, _003711_, _003835_);
  and g_097378_(_003615_, _003711_, _003836_);
  or g_097379_(_003616_, _003712_, _003837_);
  and g_097380_(_003835_, _003837_, _003839_);
  or g_097381_(_003834_, _003836_, _003840_);
  and g_097382_(_003832_, _003839_, _003841_);
  or g_097383_(_003833_, _003840_, _003842_);
  and g_097384_(_003831_, _003842_, _003843_);
  or g_097385_(_003830_, _003841_, _003844_);
  and g_097386_(_003821_, _003829_, _003845_);
  or g_097387_(_003822_, _003828_, _003846_);
  and g_097388_(_003833_, _003840_, _003847_);
  or g_097389_(_003832_, _003839_, _003848_);
  and g_097390_(_003846_, _003848_, _003850_);
  or g_097391_(_003845_, _003847_, _003851_);
  and g_097392_(_003843_, _003850_, _003852_);
  or g_097393_(_003844_, _003851_, _003853_);
  xor g_097394_(out[37], _003180_, _003854_);
  xor g_097395_(_002595_, _003180_, _003855_);
  and g_097396_(_003652_, _003711_, _003856_);
  or g_097397_(_003650_, _003712_, _003857_);
  and g_097398_(_003649_, _003712_, _003858_);
  or g_097399_(_003648_, _003711_, _003859_);
  and g_097400_(_003857_, _003859_, _003861_);
  or g_097401_(_003856_, _003858_, _003862_);
  and g_097402_(_003855_, _003861_, _003863_);
  or g_097403_(_003854_, _003862_, _003864_);
  or g_097404_(_005147_, _007831_, _003865_);
  not g_097405_(_003865_, _003866_);
  and g_097406_(_003181_, _003865_, _003867_);
  or g_097407_(_003180_, _003866_, _003868_);
  and g_097408_(_003641_, _003712_, _003869_);
  or g_097409_(_003639_, _003711_, _003870_);
  and g_097410_(_003645_, _003711_, _003872_);
  or g_097411_(_003644_, _003712_, _003873_);
  and g_097412_(_003870_, _003873_, _003874_);
  or g_097413_(_003869_, _003872_, _003875_);
  and g_097414_(_003868_, _003874_, _003876_);
  or g_097415_(_003867_, _003875_, _003877_);
  and g_097416_(_003864_, _003877_, _003878_);
  or g_097417_(_003863_, _003876_, _003879_);
  and g_097418_(_003854_, _003862_, _003880_);
  or g_097419_(_003855_, _003861_, _003881_);
  and g_097420_(_003867_, _003875_, _003883_);
  or g_097421_(_003868_, _003874_, _003884_);
  and g_097422_(_003881_, _003884_, _003885_);
  or g_097423_(_003880_, _003883_, _003886_);
  and g_097424_(_003878_, _003885_, _003887_);
  or g_097425_(_003879_, _003886_, _003888_);
  and g_097426_(_003852_, _003887_, _003889_);
  or g_097427_(_003853_, _003888_, _003890_);
  and g_097428_(_003781_, _003788_, _003891_);
  or g_097429_(_003780_, _003787_, _003892_);
  and g_097430_(_003889_, _003892_, _003894_);
  or g_097431_(_003890_, _003891_, _003895_);
  or g_097432_(_003815_, _003891_, _003896_);
  and g_097433_(_003820_, _003894_, _003897_);
  or g_097434_(_003819_, _003895_, _003898_);
  and g_097435_(_003879_, _003881_, _003899_);
  or g_097436_(_003878_, _003880_, _003900_);
  and g_097437_(_003852_, _003899_, _003901_);
  or g_097438_(_003853_, _003900_, _003902_);
  and g_097439_(_003844_, _003848_, _003903_);
  not g_097440_(_003903_, _003905_);
  and g_097441_(_003902_, _003905_, _003906_);
  or g_097442_(_003901_, _003903_, _003907_);
  and g_097443_(_003898_, _003906_, _003908_);
  or g_097444_(_003897_, _003907_, _003909_);
  and g_097445_(_003776_, _003909_, _003910_);
  or g_097446_(_003777_, _003908_, _003911_);
  and g_097447_(_003766_, _003768_, _003912_);
  or g_097448_(_003765_, _003767_, _003913_);
  and g_097449_(_003742_, _003771_, _003914_);
  or g_097450_(_003741_, _003773_, _003916_);
  and g_097451_(_003744_, _003914_, _003917_);
  or g_097452_(_003743_, _003916_, _003918_);
  and g_097453_(_003913_, _003918_, _003919_);
  or g_097454_(_003912_, _003917_, _003920_);
  and g_097455_(_003911_, _003919_, _003921_);
  or g_097456_(_003910_, _003920_, _003922_);
  and g_097457_(_002628_, _003803_, _003923_);
  or g_097458_(_003789_, _003923_, _003924_);
  or g_097459_(_003811_, _003924_, _003925_);
  or g_097460_(_003896_, _003925_, _003927_);
  or g_097461_(_003890_, _003927_, _003928_);
  not g_097462_(_003928_, _003929_);
  and g_097463_(_003776_, _003929_, _003930_);
  or g_097464_(_003777_, _003928_, _003931_);
  and g_097465_(_003922_, _003931_, _003932_);
  or g_097466_(_003921_, _003930_, _003933_);
  and g_097467_(_003715_, _003933_, _003934_);
  and g_097468_(_007842_, _003932_, _003935_);
  or g_097469_(_003934_, _003935_, _003936_);
  not g_097470_(_003936_, _003938_);
  and g_097471_(_003192_, _003207_, _003939_);
  or g_097472_(_003193_, _003206_, _003940_);
  and g_097473_(_003759_, _003933_, _003941_);
  or g_097474_(_003758_, _003932_, _003942_);
  and g_097475_(_003760_, _003932_, _003943_);
  or g_097476_(_003762_, _003933_, _003944_);
  and g_097477_(_003942_, _003944_, _003945_);
  or g_097478_(_003941_, _003943_, _003946_);
  xor g_097479_(out[58], _003203_, _003947_);
  xor g_097480_(_002815_, _003203_, _003949_);
  and g_097481_(_003945_, _003947_, _003950_);
  or g_097482_(_003946_, _003949_, _003951_);
  and g_097483_(_003940_, _003951_, _003952_);
  or g_097484_(_003939_, _003950_, _003953_);
  and g_097485_(_003193_, _003206_, _003954_);
  or g_097486_(_003192_, _003207_, _003955_);
  and g_097487_(_003946_, _003949_, _003956_);
  or g_097488_(_003945_, _003947_, _003957_);
  and g_097489_(_003955_, _003957_, _003958_);
  or g_097490_(_003954_, _003956_, _003960_);
  and g_097491_(_003952_, _003958_, _003961_);
  or g_097492_(_003953_, _003960_, _003962_);
  and g_097493_(_003720_, _003932_, _003963_);
  or g_097494_(_003719_, _003933_, _003964_);
  and g_097495_(_003725_, _003933_, _003965_);
  or g_097496_(_003726_, _003932_, _003966_);
  and g_097497_(_003964_, _003966_, _003967_);
  or g_097498_(_003963_, _003965_, _003968_);
  and g_097499_(out[57], _003202_, _003969_);
  xor g_097500_(out[57], _003202_, _003971_);
  or g_097501_(_003204_, _003969_, _003972_);
  and g_097502_(_003968_, _003971_, _003973_);
  or g_097503_(_003967_, _003972_, _003974_);
  xor g_097504_(out[56], _003201_, _003975_);
  xor g_097505_(_002793_, _003201_, _003976_);
  and g_097506_(_003731_, _003932_, _003977_);
  or g_097507_(_003730_, _003933_, _003978_);
  and g_097508_(_003737_, _003933_, _003979_);
  or g_097509_(_003736_, _003932_, _003980_);
  and g_097510_(_003978_, _003980_, _003982_);
  or g_097511_(_003977_, _003979_, _003983_);
  and g_097512_(_003976_, _003982_, _003984_);
  or g_097513_(_003975_, _003983_, _003985_);
  and g_097514_(_003974_, _003985_, _003986_);
  or g_097515_(_003973_, _003984_, _003987_);
  and g_097516_(_003967_, _003972_, _003988_);
  or g_097517_(_003968_, _003971_, _003989_);
  and g_097518_(_003975_, _003983_, _003990_);
  or g_097519_(_003976_, _003982_, _003991_);
  and g_097520_(_003989_, _003991_, _003993_);
  or g_097521_(_003988_, _003990_, _003994_);
  and g_097522_(_003986_, _003993_, _003995_);
  or g_097523_(_003987_, _003994_, _003996_);
  and g_097524_(_003961_, _003995_, _003997_);
  or g_097525_(_003962_, _003996_, _003998_);
  xor g_097526_(out[54], _003198_, _003999_);
  xor g_097527_(_002716_, _003198_, _004000_);
  or g_097528_(_003821_, _003933_, _004001_);
  or g_097529_(_003828_, _003932_, _004002_);
  and g_097530_(_004001_, _004002_, _004004_);
  and g_097531_(_004000_, _004004_, _004005_);
  xor g_097532_(_004000_, _004004_, _004006_);
  xor g_097533_(_003999_, _004004_, _004007_);
  xor g_097534_(out[55], _003199_, _004008_);
  xor g_097535_(_002705_, _003199_, _004009_);
  or g_097536_(_003833_, _003933_, _004010_);
  or g_097537_(_003839_, _003932_, _004011_);
  and g_097538_(_004010_, _004011_, _004012_);
  and g_097539_(_004008_, _004012_, _004013_);
  or g_097540_(_004008_, _004012_, _004015_);
  xor g_097541_(_004008_, _004012_, _004016_);
  xor g_097542_(_004009_, _004012_, _004017_);
  and g_097543_(_004006_, _004016_, _004018_);
  or g_097544_(_004007_, _004017_, _004019_);
  or g_097545_(_004993_, _010823_, _004020_);
  not g_097546_(_004020_, _004021_);
  and g_097547_(_003197_, _004020_, _004022_);
  or g_097548_(_003196_, _004021_, _004023_);
  and g_097549_(_003875_, _003933_, _004024_);
  or g_097550_(_003874_, _003932_, _004026_);
  and g_097551_(_003868_, _003932_, _004027_);
  or g_097552_(_003867_, _003933_, _004028_);
  and g_097553_(_004026_, _004028_, _004029_);
  or g_097554_(_004024_, _004027_, _004030_);
  and g_097555_(_004023_, _004029_, _004031_);
  or g_097556_(_004022_, _004030_, _004032_);
  xor g_097557_(out[53], _003196_, _004033_);
  xor g_097558_(_002727_, _003196_, _004034_);
  and g_097559_(_003855_, _003932_, _004035_);
  or g_097560_(_003854_, _003933_, _004037_);
  and g_097561_(_003862_, _003933_, _004038_);
  or g_097562_(_003861_, _003932_, _004039_);
  and g_097563_(_004037_, _004039_, _004040_);
  or g_097564_(_004035_, _004038_, _004041_);
  and g_097565_(_004034_, _004040_, _004042_);
  or g_097566_(_004033_, _004041_, _004043_);
  and g_097567_(_004032_, _004043_, _004044_);
  or g_097568_(_004031_, _004042_, _004045_);
  and g_097569_(_004033_, _004041_, _004046_);
  or g_097570_(_004034_, _004040_, _004048_);
  and g_097571_(_004022_, _004030_, _004049_);
  or g_097572_(_004023_, _004029_, _004050_);
  and g_097573_(_004048_, _004050_, _004051_);
  or g_097574_(_004046_, _004049_, _004052_);
  and g_097575_(_004044_, _004051_, _004053_);
  or g_097576_(_004045_, _004052_, _004054_);
  and g_097577_(_004018_, _004053_, _004055_);
  or g_097578_(_004019_, _004054_, _004056_);
  and g_097579_(_003997_, _004055_, _004057_);
  or g_097580_(_003998_, _004056_, _004059_);
  xor g_097581_(out[51], _010823_, _004060_);
  xor g_097582_(_002782_, _010823_, _004061_);
  and g_097583_(_003780_, _003932_, _004062_);
  or g_097584_(_003781_, _003933_, _004063_);
  and g_097585_(_003788_, _003933_, _004064_);
  or g_097586_(_003787_, _003932_, _004065_);
  and g_097587_(_004063_, _004065_, _004066_);
  or g_097588_(_004062_, _004064_, _004067_);
  and g_097589_(_004060_, _004066_, _004068_);
  or g_097590_(_004061_, _004067_, _004070_);
  and g_097591_(_004061_, _004067_, _004071_);
  or g_097592_(_004060_, _004066_, _004072_);
  and g_097593_(_010834_, _003938_, _004073_);
  or g_097594_(_010845_, _003936_, _004074_);
  and g_097595_(_004072_, _004073_, _004075_);
  or g_097596_(_004071_, _004074_, _004076_);
  and g_097597_(_004070_, _004076_, _004077_);
  or g_097598_(_004068_, _004075_, _004078_);
  or g_097599_(_002617_, _003933_, _004079_);
  or g_097600_(_003796_, _003932_, _004081_);
  and g_097601_(_004079_, _004081_, _004082_);
  and g_097602_(out[49], _004082_, _004083_);
  not g_097603_(_004083_, _004084_);
  and g_097604_(out[32], _003932_, _004085_);
  or g_097605_(_002628_, _003933_, _004086_);
  and g_097606_(_003803_, _003933_, _004087_);
  or g_097607_(_003804_, _003932_, _004088_);
  and g_097608_(_004086_, _004088_, _004089_);
  or g_097609_(_004085_, _004087_, _004090_);
  and g_097610_(out[48], _004089_, _004092_);
  or g_097611_(_002760_, _004090_, _004093_);
  xor g_097612_(out[49], _004082_, _004094_);
  xor g_097613_(_002749_, _004082_, _004095_);
  and g_097614_(_004093_, _004094_, _004096_);
  or g_097615_(_004092_, _004095_, _004097_);
  and g_097616_(_004084_, _004097_, _004098_);
  or g_097617_(_004083_, _004096_, _004099_);
  xor g_097618_(_010845_, _003936_, _004100_);
  xor g_097619_(_010834_, _003936_, _004101_);
  and g_097620_(_004072_, _004100_, _004103_);
  or g_097621_(_004071_, _004101_, _004104_);
  and g_097622_(_004099_, _004103_, _004105_);
  or g_097623_(_004098_, _004104_, _004106_);
  and g_097624_(_004077_, _004106_, _004107_);
  or g_097625_(_004078_, _004105_, _004108_);
  and g_097626_(_004057_, _004108_, _004109_);
  or g_097627_(_004059_, _004107_, _004110_);
  and g_097628_(_004018_, _004045_, _004111_);
  or g_097629_(_004019_, _004044_, _004112_);
  and g_097630_(_004048_, _004111_, _004114_);
  or g_097631_(_004046_, _004112_, _004115_);
  and g_097632_(_004005_, _004015_, _004116_);
  or g_097633_(_004013_, _004116_, _004117_);
  not g_097634_(_004117_, _004118_);
  and g_097635_(_004115_, _004118_, _004119_);
  or g_097636_(_004114_, _004117_, _004120_);
  and g_097637_(_003997_, _004120_, _004121_);
  or g_097638_(_003998_, _004119_, _004122_);
  and g_097639_(_003987_, _003989_, _004123_);
  or g_097640_(_003986_, _003988_, _004125_);
  and g_097641_(_003961_, _004123_, _004126_);
  or g_097642_(_003962_, _004125_, _004127_);
  and g_097643_(_003953_, _003955_, _004128_);
  or g_097644_(_003952_, _003954_, _004129_);
  and g_097645_(_004110_, _004129_, _004130_);
  or g_097646_(_004109_, _004128_, _004131_);
  and g_097647_(_004122_, _004127_, _004132_);
  or g_097648_(_004121_, _004126_, _004133_);
  and g_097649_(_004130_, _004132_, _004134_);
  or g_097650_(_004131_, _004133_, _004136_);
  and g_097651_(_002760_, _004090_, _004137_);
  or g_097652_(out[48], _004089_, _004138_);
  and g_097653_(_004070_, _004138_, _004139_);
  or g_097654_(_004068_, _004137_, _004140_);
  and g_097655_(_004096_, _004139_, _004141_);
  or g_097656_(_004097_, _004140_, _004142_);
  and g_097657_(_004103_, _004141_, _004143_);
  or g_097658_(_004104_, _004142_, _004144_);
  and g_097659_(_004057_, _004143_, _004145_);
  or g_097660_(_004059_, _004144_, _004147_);
  and g_097661_(_004136_, _004147_, _004148_);
  or g_097662_(_004134_, _004145_, _004149_);
  and g_097663_(_003936_, _004149_, _004150_);
  and g_097664_(_010834_, _004148_, _004151_);
  or g_097665_(_004150_, _004151_, _004152_);
  not g_097666_(_004152_, _004153_);
  and g_097667_(_003946_, _004149_, _004154_);
  or g_097668_(_003945_, _004148_, _004155_);
  and g_097669_(_003947_, _004148_, _004156_);
  or g_097670_(_003949_, _004149_, _004158_);
  and g_097671_(_004155_, _004158_, _004159_);
  or g_097672_(_004154_, _004156_, _004160_);
  xor g_097673_(out[74], _003219_, _004161_);
  xor g_097674_(_002947_, _003219_, _004162_);
  and g_097675_(_004159_, _004161_, _004163_);
  or g_097676_(_004160_, _004162_, _004164_);
  and g_097677_(_003208_, _003224_, _004165_);
  or g_097678_(_003209_, _003223_, _004166_);
  and g_097679_(_004164_, _004166_, _004167_);
  or g_097680_(_004163_, _004165_, _004169_);
  and g_097681_(_004160_, _004162_, _004170_);
  or g_097682_(_004159_, _004161_, _004171_);
  and g_097683_(_004167_, _004171_, _004172_);
  or g_097684_(_004169_, _004170_, _004173_);
  and g_097685_(_003209_, _003223_, _004174_);
  or g_097686_(_003208_, _003224_, _004175_);
  and g_097687_(_003968_, _004149_, _004176_);
  or g_097688_(_003967_, _004148_, _004177_);
  and g_097689_(_003972_, _004148_, _004178_);
  or g_097690_(_003971_, _004149_, _004180_);
  and g_097691_(_004177_, _004180_, _004181_);
  or g_097692_(_004176_, _004178_, _004182_);
  and g_097693_(out[73], _003218_, _004183_);
  xor g_097694_(out[73], _003218_, _004184_);
  or g_097695_(_003220_, _004183_, _004185_);
  and g_097696_(_004182_, _004184_, _004186_);
  or g_097697_(_004181_, _004185_, _004187_);
  and g_097698_(_004175_, _004187_, _004188_);
  or g_097699_(_004174_, _004186_, _004189_);
  xor g_097700_(out[72], _003217_, _004191_);
  xor g_097701_(_002925_, _003217_, _004192_);
  and g_097702_(_003976_, _004148_, _004193_);
  or g_097703_(_003975_, _004149_, _004194_);
  and g_097704_(_003983_, _004149_, _004195_);
  or g_097705_(_003982_, _004148_, _004196_);
  and g_097706_(_004194_, _004196_, _004197_);
  or g_097707_(_004193_, _004195_, _004198_);
  and g_097708_(_004192_, _004197_, _004199_);
  or g_097709_(_004191_, _004198_, _004200_);
  and g_097710_(_004181_, _004185_, _004202_);
  or g_097711_(_004182_, _004184_, _004203_);
  and g_097712_(_004200_, _004203_, _004204_);
  or g_097713_(_004199_, _004202_, _004205_);
  and g_097714_(_004191_, _004198_, _004206_);
  or g_097715_(_004192_, _004197_, _004207_);
  and g_097716_(_004204_, _004207_, _004208_);
  or g_097717_(_004205_, _004206_, _004209_);
  and g_097718_(_004188_, _004208_, _004210_);
  or g_097719_(_004189_, _004209_, _004211_);
  and g_097720_(_004172_, _004210_, _004213_);
  or g_097721_(_004173_, _004211_, _004214_);
  xor g_097722_(out[71], _003216_, _004215_);
  xor g_097723_(_002837_, _003216_, _004216_);
  or g_097724_(_004009_, _004149_, _004217_);
  or g_097725_(_004012_, _004148_, _004218_);
  and g_097726_(_004217_, _004218_, _004219_);
  and g_097727_(_004215_, _004219_, _004220_);
  xor g_097728_(out[70], _003215_, _004221_);
  xor g_097729_(_002848_, _003215_, _004222_);
  or g_097730_(_003999_, _004149_, _004224_);
  or g_097731_(_004004_, _004148_, _004225_);
  and g_097732_(_004224_, _004225_, _004226_);
  and g_097733_(_004222_, _004226_, _004227_);
  or g_097734_(_004215_, _004219_, _004228_);
  xor g_097735_(_004215_, _004219_, _004229_);
  xor g_097736_(_004216_, _004219_, _004230_);
  xor g_097737_(_004222_, _004226_, _004231_);
  xor g_097738_(_004221_, _004226_, _004232_);
  and g_097739_(_004229_, _004231_, _004233_);
  or g_097740_(_004230_, _004232_, _004235_);
  or g_097741_(_004861_, _026608_, _004236_);
  not g_097742_(_004236_, _004237_);
  and g_097743_(_003214_, _004236_, _004238_);
  or g_097744_(_003213_, _004237_, _004239_);
  and g_097745_(_004030_, _004149_, _004240_);
  or g_097746_(_004029_, _004148_, _004241_);
  and g_097747_(_004023_, _004148_, _004242_);
  or g_097748_(_004022_, _004149_, _004243_);
  and g_097749_(_004241_, _004243_, _004244_);
  or g_097750_(_004240_, _004242_, _004246_);
  and g_097751_(_004239_, _004244_, _004247_);
  or g_097752_(_004238_, _004246_, _004248_);
  xor g_097753_(out[69], _003213_, _004249_);
  xor g_097754_(_002859_, _003213_, _004250_);
  and g_097755_(_004034_, _004148_, _004251_);
  or g_097756_(_004033_, _004149_, _004252_);
  and g_097757_(_004041_, _004149_, _004253_);
  or g_097758_(_004040_, _004148_, _004254_);
  and g_097759_(_004252_, _004254_, _004255_);
  or g_097760_(_004251_, _004253_, _004257_);
  and g_097761_(_004250_, _004255_, _004258_);
  or g_097762_(_004249_, _004257_, _004259_);
  and g_097763_(_004248_, _004259_, _004260_);
  or g_097764_(_004247_, _004258_, _004261_);
  and g_097765_(_004249_, _004257_, _004262_);
  or g_097766_(_004250_, _004255_, _004263_);
  and g_097767_(_004238_, _004246_, _004264_);
  or g_097768_(_004239_, _004244_, _004265_);
  and g_097769_(_004263_, _004265_, _004266_);
  or g_097770_(_004262_, _004264_, _004268_);
  and g_097771_(_004260_, _004266_, _004269_);
  or g_097772_(_004261_, _004268_, _004270_);
  and g_097773_(_004233_, _004269_, _004271_);
  or g_097774_(_004235_, _004270_, _004272_);
  and g_097775_(_004213_, _004271_, _004273_);
  or g_097776_(_004214_, _004272_, _004274_);
  xor g_097777_(out[67], _026608_, _004275_);
  xor g_097778_(_002914_, _026608_, _004276_);
  and g_097779_(_004060_, _004148_, _004277_);
  not g_097780_(_004277_, _004279_);
  or g_097781_(_004066_, _004148_, _004280_);
  not g_097782_(_004280_, _004281_);
  and g_097783_(_004279_, _004280_, _004282_);
  or g_097784_(_004277_, _004281_, _004283_);
  and g_097785_(_004275_, _004282_, _004284_);
  or g_097786_(_004276_, _004283_, _004285_);
  or g_097787_(_026630_, _004152_, _004286_);
  not g_097788_(_004286_, _004287_);
  and g_097789_(_004285_, _004286_, _004288_);
  or g_097790_(_004284_, _004287_, _004290_);
  and g_097791_(_004276_, _004283_, _004291_);
  or g_097792_(_004275_, _004282_, _004292_);
  and g_097793_(_026630_, _004152_, _004293_);
  or g_097794_(_026619_, _004153_, _004294_);
  and g_097795_(_004292_, _004294_, _004295_);
  or g_097796_(_004291_, _004293_, _004296_);
  and g_097797_(_004288_, _004295_, _004297_);
  or g_097798_(_004290_, _004296_, _004298_);
  and g_097799_(out[49], _004148_, _004299_);
  not g_097800_(_004299_, _004301_);
  or g_097801_(_004082_, _004148_, _004302_);
  not g_097802_(_004302_, _004303_);
  and g_097803_(_004301_, _004302_, _004304_);
  or g_097804_(_004299_, _004303_, _004305_);
  and g_097805_(out[65], _004304_, _004306_);
  or g_097806_(_002881_, _004305_, _004307_);
  and g_097807_(out[48], _004148_, _004308_);
  not g_097808_(_004308_, _004309_);
  or g_097809_(_004089_, _004148_, _004310_);
  not g_097810_(_004310_, _004312_);
  and g_097811_(_004309_, _004310_, _004313_);
  or g_097812_(_004308_, _004312_, _004314_);
  and g_097813_(out[64], _004313_, _004315_);
  or g_097814_(_002892_, _004314_, _004316_);
  xor g_097815_(out[65], _004304_, _004317_);
  xor g_097816_(_002881_, _004304_, _004318_);
  and g_097817_(_004316_, _004317_, _004319_);
  or g_097818_(_004315_, _004318_, _004320_);
  and g_097819_(_004307_, _004320_, _004321_);
  or g_097820_(_004306_, _004319_, _004323_);
  and g_097821_(_004297_, _004323_, _004324_);
  or g_097822_(_004298_, _004321_, _004325_);
  and g_097823_(_004290_, _004292_, _004326_);
  or g_097824_(_004288_, _004291_, _004327_);
  and g_097825_(_004325_, _004327_, _004328_);
  or g_097826_(_004324_, _004326_, _004329_);
  and g_097827_(_004273_, _004329_, _004330_);
  or g_097828_(_004274_, _004328_, _004331_);
  and g_097829_(_004233_, _004261_, _004332_);
  or g_097830_(_004235_, _004260_, _004334_);
  and g_097831_(_004263_, _004332_, _004335_);
  or g_097832_(_004262_, _004334_, _004336_);
  and g_097833_(_004227_, _004228_, _004337_);
  or g_097834_(_004220_, _004337_, _004338_);
  not g_097835_(_004338_, _004339_);
  and g_097836_(_004336_, _004339_, _004340_);
  or g_097837_(_004335_, _004338_, _004341_);
  and g_097838_(_004213_, _004341_, _004342_);
  or g_097839_(_004214_, _004340_, _004343_);
  and g_097840_(_004199_, _004203_, _004345_);
  or g_097841_(_004200_, _004202_, _004346_);
  and g_097842_(_004187_, _004346_, _004347_);
  or g_097843_(_004186_, _004345_, _004348_);
  and g_097844_(_004172_, _004348_, _004349_);
  or g_097845_(_004173_, _004347_, _004350_);
  and g_097846_(_004167_, _004350_, _004351_);
  or g_097847_(_004169_, _004349_, _004352_);
  and g_097848_(_004175_, _004352_, _004353_);
  or g_097849_(_004174_, _004351_, _004354_);
  and g_097850_(_004343_, _004354_, _004356_);
  or g_097851_(_004342_, _004353_, _004357_);
  and g_097852_(_004331_, _004356_, _004358_);
  or g_097853_(_004330_, _004357_, _004359_);
  or g_097854_(out[64], _004313_, _004360_);
  and g_097855_(_004297_, _004360_, _004361_);
  not g_097856_(_004361_, _004362_);
  and g_097857_(_004319_, _004361_, _004363_);
  or g_097858_(_004320_, _004362_, _004364_);
  and g_097859_(_004273_, _004363_, _004365_);
  or g_097860_(_004274_, _004364_, _004367_);
  and g_097861_(_004359_, _004367_, _004368_);
  or g_097862_(_004358_, _004365_, _004369_);
  or g_097863_(_004153_, _004368_, _004370_);
  not g_097864_(_004370_, _004371_);
  and g_097865_(_026619_, _004368_, _004372_);
  not g_097866_(_004372_, _004373_);
  and g_097867_(_004370_, _004373_, _004374_);
  or g_097868_(_004371_, _004372_, _004375_);
  xor g_097869_(out[90], _003236_, _004376_);
  xor g_097870_(_003079_, _003236_, _004378_);
  and g_097871_(_004160_, _004369_, _004379_);
  or g_097872_(_004159_, _004368_, _004380_);
  and g_097873_(_004161_, _004368_, _004381_);
  or g_097874_(_004162_, _004369_, _004382_);
  and g_097875_(_004380_, _004382_, _004383_);
  or g_097876_(_004379_, _004381_, _004384_);
  and g_097877_(_004376_, _004383_, _004385_);
  or g_097878_(_004378_, _004384_, _004386_);
  and g_097879_(_003225_, _003240_, _004387_);
  or g_097880_(_003226_, _003239_, _004389_);
  and g_097881_(_004386_, _004389_, _004390_);
  or g_097882_(_004385_, _004387_, _004391_);
  and g_097883_(_004378_, _004384_, _004392_);
  or g_097884_(_004376_, _004383_, _004393_);
  and g_097885_(_003226_, _003239_, _004394_);
  or g_097886_(_003225_, _003240_, _004395_);
  and g_097887_(_004182_, _004369_, _004396_);
  or g_097888_(_004181_, _004368_, _004397_);
  and g_097889_(_004185_, _004368_, _004398_);
  not g_097890_(_004398_, _004400_);
  and g_097891_(_004397_, _004400_, _004401_);
  or g_097892_(_004396_, _004398_, _004402_);
  and g_097893_(out[89], _003235_, _004403_);
  xor g_097894_(out[89], _003235_, _004404_);
  or g_097895_(_003237_, _004403_, _004405_);
  and g_097896_(_004401_, _004405_, _004406_);
  or g_097897_(_004402_, _004404_, _004407_);
  xor g_097898_(out[88], _003234_, _004408_);
  xor g_097899_(_003057_, _003234_, _004409_);
  and g_097900_(_004192_, _004368_, _004411_);
  not g_097901_(_004411_, _004412_);
  or g_097902_(_004197_, _004368_, _004413_);
  not g_097903_(_004413_, _004414_);
  and g_097904_(_004412_, _004413_, _004415_);
  or g_097905_(_004411_, _004414_, _004416_);
  and g_097906_(_004408_, _004416_, _004417_);
  or g_097907_(_004409_, _004415_, _004418_);
  and g_097908_(_004402_, _004404_, _004419_);
  not g_097909_(_004419_, _004420_);
  and g_097910_(_004409_, _004415_, _004422_);
  or g_097911_(_004408_, _004416_, _004423_);
  and g_097912_(_004420_, _004423_, _004424_);
  or g_097913_(_004419_, _004422_, _004425_);
  and g_097914_(_004393_, _004395_, _004426_);
  or g_097915_(_004392_, _004394_, _004427_);
  and g_097916_(_004390_, _004426_, _004428_);
  or g_097917_(_004391_, _004427_, _004429_);
  and g_097918_(_004418_, _004420_, _004430_);
  or g_097919_(_004417_, _004419_, _004431_);
  and g_097920_(_004407_, _004423_, _004433_);
  or g_097921_(_004406_, _004422_, _004434_);
  and g_097922_(_004430_, _004433_, _004435_);
  or g_097923_(_004431_, _004434_, _004436_);
  and g_097924_(_004428_, _004435_, _004437_);
  or g_097925_(_004429_, _004436_, _004438_);
  xor g_097926_(out[86], _003231_, _004439_);
  not g_097927_(_004439_, _004440_);
  or g_097928_(_004221_, _004369_, _004441_);
  or g_097929_(_004226_, _004368_, _004442_);
  and g_097930_(_004441_, _004442_, _004444_);
  and g_097931_(_004440_, _004444_, _004445_);
  xor g_097932_(_004440_, _004444_, _004446_);
  xor g_097933_(_004439_, _004444_, _004447_);
  xor g_097934_(out[87], _003232_, _004448_);
  xor g_097935_(_002969_, _003232_, _004449_);
  or g_097936_(_004216_, _004369_, _004450_);
  or g_097937_(_004219_, _004368_, _004451_);
  and g_097938_(_004450_, _004451_, _004452_);
  or g_097939_(_004448_, _004452_, _004453_);
  and g_097940_(_004448_, _004452_, _004455_);
  xor g_097941_(_004448_, _004452_, _004456_);
  xor g_097942_(_004449_, _004452_, _004457_);
  and g_097943_(_004446_, _004456_, _004458_);
  or g_097944_(_004447_, _004457_, _004459_);
  or g_097945_(_011736_, _026575_, _004460_);
  not g_097946_(_004460_, _004461_);
  and g_097947_(_003230_, _004460_, _004462_);
  or g_097948_(_003229_, _004461_, _004463_);
  and g_097949_(_004246_, _004369_, _004464_);
  or g_097950_(_004244_, _004368_, _004466_);
  and g_097951_(_004239_, _004368_, _004467_);
  or g_097952_(_004238_, _004369_, _004468_);
  and g_097953_(_004466_, _004468_, _004469_);
  or g_097954_(_004464_, _004467_, _004470_);
  and g_097955_(_004463_, _004469_, _004471_);
  or g_097956_(_004462_, _004470_, _004472_);
  xor g_097957_(out[85], _003229_, _004473_);
  xor g_097958_(_002991_, _003229_, _004474_);
  and g_097959_(_004250_, _004368_, _004475_);
  or g_097960_(_004249_, _004369_, _004477_);
  and g_097961_(_004257_, _004369_, _004478_);
  or g_097962_(_004255_, _004368_, _004479_);
  and g_097963_(_004477_, _004479_, _004480_);
  or g_097964_(_004475_, _004478_, _004481_);
  and g_097965_(_004474_, _004480_, _004482_);
  or g_097966_(_004473_, _004481_, _004483_);
  and g_097967_(_004472_, _004483_, _004484_);
  or g_097968_(_004471_, _004482_, _004485_);
  and g_097969_(_004473_, _004481_, _004486_);
  or g_097970_(_004474_, _004480_, _004488_);
  and g_097971_(_004462_, _004470_, _004489_);
  or g_097972_(_004463_, _004469_, _004490_);
  and g_097973_(_004488_, _004490_, _004491_);
  or g_097974_(_004486_, _004489_, _004492_);
  and g_097975_(_004484_, _004491_, _004493_);
  or g_097976_(_004485_, _004492_, _004494_);
  and g_097977_(_004458_, _004493_, _004495_);
  or g_097978_(_004459_, _004494_, _004496_);
  and g_097979_(_004437_, _004495_, _004497_);
  or g_097980_(_004438_, _004496_, _004499_);
  xor g_097981_(out[83], _026575_, _004500_);
  xor g_097982_(_003046_, _026575_, _004501_);
  and g_097983_(_004275_, _004368_, _004502_);
  not g_097984_(_004502_, _004503_);
  or g_097985_(_004282_, _004368_, _004504_);
  not g_097986_(_004504_, _004505_);
  and g_097987_(_004503_, _004504_, _004506_);
  or g_097988_(_004502_, _004505_, _004507_);
  and g_097989_(_004500_, _004506_, _004508_);
  or g_097990_(_004501_, _004507_, _004510_);
  and g_097991_(_004501_, _004507_, _004511_);
  or g_097992_(_004500_, _004506_, _004512_);
  and g_097993_(_026586_, _004374_, _004513_);
  or g_097994_(_026597_, _004375_, _004514_);
  and g_097995_(_004512_, _004513_, _004515_);
  or g_097996_(_004511_, _004514_, _004516_);
  and g_097997_(_004510_, _004516_, _004517_);
  or g_097998_(_004508_, _004515_, _004518_);
  and g_097999_(out[65], _004368_, _004519_);
  not g_098000_(_004519_, _004521_);
  or g_098001_(_004304_, _004368_, _004522_);
  not g_098002_(_004522_, _004523_);
  and g_098003_(_004521_, _004522_, _004524_);
  or g_098004_(_004519_, _004523_, _004525_);
  and g_098005_(out[81], _004524_, _004526_);
  or g_098006_(_003013_, _004525_, _004527_);
  and g_098007_(out[64], _004368_, _004528_);
  not g_098008_(_004528_, _004529_);
  or g_098009_(_004313_, _004368_, _004530_);
  not g_098010_(_004530_, _004532_);
  and g_098011_(_004529_, _004530_, _004533_);
  or g_098012_(_004528_, _004532_, _004534_);
  and g_098013_(out[80], _004533_, _004535_);
  or g_098014_(_003024_, _004534_, _004536_);
  xor g_098015_(out[81], _004524_, _004537_);
  xor g_098016_(_003013_, _004524_, _004538_);
  and g_098017_(_004536_, _004537_, _004539_);
  or g_098018_(_004535_, _004538_, _004540_);
  and g_098019_(_004527_, _004540_, _004541_);
  or g_098020_(_004526_, _004539_, _004543_);
  xor g_098021_(_026586_, _004374_, _004544_);
  xor g_098022_(_026597_, _004374_, _004545_);
  and g_098023_(_004512_, _004544_, _004546_);
  or g_098024_(_004511_, _004545_, _004547_);
  and g_098025_(_004543_, _004546_, _004548_);
  or g_098026_(_004541_, _004547_, _004549_);
  and g_098027_(_004517_, _004549_, _004550_);
  or g_098028_(_004518_, _004548_, _004551_);
  and g_098029_(_004497_, _004551_, _004552_);
  or g_098030_(_004499_, _004550_, _004554_);
  and g_098031_(_004458_, _004485_, _004555_);
  or g_098032_(_004459_, _004484_, _004556_);
  and g_098033_(_004488_, _004555_, _004557_);
  or g_098034_(_004486_, _004556_, _004558_);
  and g_098035_(_004445_, _004453_, _004559_);
  or g_098036_(_004455_, _004559_, _004560_);
  not g_098037_(_004560_, _004561_);
  and g_098038_(_004558_, _004561_, _004562_);
  or g_098039_(_004557_, _004560_, _004563_);
  and g_098040_(_004437_, _004563_, _004565_);
  or g_098041_(_004438_, _004562_, _004566_);
  and g_098042_(_004425_, _004428_, _004567_);
  or g_098043_(_004424_, _004429_, _004568_);
  and g_098044_(_004407_, _004567_, _004569_);
  or g_098045_(_004406_, _004568_, _004570_);
  or g_098046_(_004390_, _004394_, _004571_);
  not g_098047_(_004571_, _004572_);
  and g_098048_(_004570_, _004571_, _004573_);
  or g_098049_(_004569_, _004572_, _004574_);
  and g_098050_(_004566_, _004573_, _004576_);
  or g_098051_(_004565_, _004574_, _004577_);
  and g_098052_(_004554_, _004576_, _004578_);
  or g_098053_(_004552_, _004577_, _004579_);
  and g_098054_(_003024_, _004534_, _004580_);
  or g_098055_(out[80], _004533_, _004581_);
  and g_098056_(_004510_, _004581_, _004582_);
  or g_098057_(_004508_, _004580_, _004583_);
  and g_098058_(_004539_, _004582_, _004584_);
  or g_098059_(_004540_, _004583_, _004585_);
  and g_098060_(_004546_, _004584_, _004587_);
  or g_098061_(_004547_, _004585_, _004588_);
  and g_098062_(_004497_, _004587_, _004589_);
  or g_098063_(_004499_, _004588_, _004590_);
  and g_098064_(_004579_, _004590_, _004591_);
  or g_098065_(_004578_, _004589_, _004592_);
  or g_098066_(_004374_, _004591_, _004593_);
  or g_098067_(_026597_, _004592_, _004594_);
  and g_098068_(_004593_, _004594_, _004595_);
  and g_098069_(_031206_, _004595_, _004596_);
  xor g_098070_(out[99], _031195_, _004598_);
  xor g_098071_(_003178_, _031195_, _004599_);
  and g_098072_(_004500_, _004591_, _004600_);
  or g_098073_(_004501_, _004592_, _004601_);
  and g_098074_(_004507_, _004592_, _004602_);
  or g_098075_(_004506_, _004591_, _004603_);
  and g_098076_(_004601_, _004603_, _004604_);
  or g_098077_(_004600_, _004602_, _004605_);
  and g_098078_(_004598_, _004604_, _004606_);
  or g_098079_(_004596_, _004606_, _004607_);
  or g_098080_(_003013_, _004592_, _004609_);
  or g_098081_(_004524_, _004591_, _004610_);
  and g_098082_(_004609_, _004610_, _004611_);
  and g_098083_(out[97], _004611_, _004612_);
  and g_098084_(out[80], _004591_, _004613_);
  or g_098085_(_003024_, _004592_, _004614_);
  and g_098086_(_004534_, _004592_, _004615_);
  or g_098087_(_004533_, _004591_, _004616_);
  and g_098088_(_004614_, _004616_, _004617_);
  or g_098089_(_004613_, _004615_, _004618_);
  and g_098090_(out[96], _004617_, _004620_);
  or g_098091_(_003156_, _004618_, _004621_);
  xor g_098092_(out[97], _004611_, _004622_);
  xor g_098093_(_003145_, _004611_, _004623_);
  and g_098094_(_004621_, _004622_, _004624_);
  or g_098095_(_004620_, _004623_, _004625_);
  or g_098096_(_004612_, _004624_, _004626_);
  xor g_098097_(_031206_, _004595_, _004627_);
  xor g_098098_(_031217_, _004595_, _004628_);
  and g_098099_(_004626_, _004627_, _004629_);
  or g_098100_(_004607_, _004629_, _004631_);
  not g_098101_(_004631_, _004632_);
  and g_098102_(_004384_, _004592_, _004633_);
  or g_098103_(_004383_, _004591_, _004634_);
  and g_098104_(_004376_, _004591_, _004635_);
  or g_098105_(_004378_, _004592_, _004636_);
  and g_098106_(_004634_, _004636_, _004637_);
  or g_098107_(_004633_, _004635_, _004638_);
  and g_098108_(_003565_, _004637_, _004639_);
  or g_098109_(_003566_, _004638_, _004640_);
  and g_098110_(_003241_, _003257_, _004642_);
  or g_098111_(_003242_, _003256_, _004643_);
  and g_098112_(_004640_, _004643_, _004644_);
  or g_098113_(_004639_, _004642_, _004645_);
  and g_098114_(_003566_, _004638_, _004646_);
  or g_098115_(_003565_, _004637_, _004647_);
  and g_098116_(_003242_, _003256_, _004648_);
  or g_098117_(_003241_, _003257_, _004649_);
  and g_098118_(out[105], _003251_, _004650_);
  xor g_098119_(out[105], _003251_, _004651_);
  or g_098120_(_003253_, _004650_, _004653_);
  and g_098121_(_004402_, _004592_, _004654_);
  or g_098122_(_004401_, _004591_, _004655_);
  and g_098123_(_004405_, _004591_, _004656_);
  or g_098124_(_004404_, _004592_, _004657_);
  and g_098125_(_004655_, _004657_, _004658_);
  or g_098126_(_004654_, _004656_, _004659_);
  and g_098127_(_004653_, _004658_, _004660_);
  or g_098128_(_004651_, _004659_, _004661_);
  xor g_098129_(out[104], _003250_, _004662_);
  xor g_098130_(_003189_, _003250_, _004664_);
  and g_098131_(_004409_, _004591_, _004665_);
  or g_098132_(_004408_, _004592_, _004666_);
  and g_098133_(_004416_, _004592_, _004667_);
  or g_098134_(_004415_, _004591_, _004668_);
  and g_098135_(_004666_, _004668_, _004669_);
  or g_098136_(_004665_, _004667_, _004670_);
  and g_098137_(_004662_, _004670_, _004671_);
  or g_098138_(_004664_, _004669_, _004672_);
  and g_098139_(_004651_, _004659_, _004673_);
  or g_098140_(_004653_, _004658_, _004675_);
  and g_098141_(_004672_, _004675_, _004676_);
  or g_098142_(_004671_, _004673_, _004677_);
  and g_098143_(_004664_, _004669_, _004678_);
  or g_098144_(_004662_, _004670_, _004679_);
  and g_098145_(_004644_, _004649_, _004680_);
  or g_098146_(_004645_, _004648_, _004681_);
  and g_098147_(_004647_, _004680_, _004682_);
  or g_098148_(_004646_, _004681_, _004683_);
  and g_098149_(_004661_, _004679_, _004684_);
  or g_098150_(_004660_, _004678_, _004686_);
  and g_098151_(_004676_, _004684_, _004687_);
  or g_098152_(_004677_, _004686_, _004688_);
  and g_098153_(_004682_, _004687_, _004689_);
  or g_098154_(_004683_, _004688_, _004690_);
  xor g_098155_(out[103], _003249_, _004691_);
  xor g_098156_(_003101_, _003249_, _004692_);
  or g_098157_(_004452_, _004591_, _004693_);
  or g_098158_(_004449_, _004592_, _004694_);
  and g_098159_(_004693_, _004694_, _004695_);
  and g_098160_(_004691_, _004695_, _004697_);
  or g_098161_(_004691_, _004695_, _004698_);
  xor g_098162_(_004691_, _004695_, _004699_);
  xor g_098163_(_004692_, _004695_, _004700_);
  xor g_098164_(out[102], _003248_, _004701_);
  xor g_098165_(_003112_, _003248_, _004702_);
  or g_098166_(_004444_, _004591_, _004703_);
  or g_098167_(_004439_, _004592_, _004704_);
  and g_098168_(_004703_, _004704_, _004705_);
  and g_098169_(_004702_, _004705_, _004706_);
  xor g_098170_(_004702_, _004705_, _004708_);
  xor g_098171_(_004701_, _004705_, _004709_);
  and g_098172_(_004699_, _004708_, _004710_);
  or g_098173_(_004700_, _004709_, _004711_);
  or g_098174_(_011890_, _031195_, _004712_);
  not g_098175_(_004712_, _004713_);
  and g_098176_(_003247_, _004712_, _004714_);
  or g_098177_(_003246_, _004713_, _004715_);
  and g_098178_(_004470_, _004592_, _004716_);
  or g_098179_(_004469_, _004591_, _004717_);
  and g_098180_(_004463_, _004591_, _004719_);
  or g_098181_(_004462_, _004592_, _004720_);
  and g_098182_(_004717_, _004720_, _004721_);
  or g_098183_(_004716_, _004719_, _004722_);
  and g_098184_(_004715_, _004721_, _004723_);
  or g_098185_(_004714_, _004722_, _004724_);
  xor g_098186_(out[101], _003246_, _004725_);
  xor g_098187_(_003123_, _003246_, _004726_);
  and g_098188_(_004474_, _004591_, _004727_);
  or g_098189_(_004473_, _004592_, _004728_);
  and g_098190_(_004481_, _004592_, _004730_);
  or g_098191_(_004480_, _004591_, _004731_);
  and g_098192_(_004728_, _004731_, _004732_);
  or g_098193_(_004727_, _004730_, _004733_);
  and g_098194_(_004726_, _004732_, _004734_);
  or g_098195_(_004725_, _004733_, _004735_);
  and g_098196_(_004724_, _004735_, _004736_);
  or g_098197_(_004723_, _004734_, _004737_);
  and g_098198_(_004725_, _004733_, _004738_);
  or g_098199_(_004726_, _004732_, _004739_);
  and g_098200_(_004714_, _004722_, _004741_);
  or g_098201_(_004715_, _004721_, _004742_);
  and g_098202_(_004739_, _004742_, _004743_);
  or g_098203_(_004738_, _004741_, _004744_);
  and g_098204_(_004736_, _004743_, _004745_);
  or g_098205_(_004737_, _004744_, _004746_);
  and g_098206_(_004710_, _004745_, _004747_);
  or g_098207_(_004711_, _004746_, _004748_);
  and g_098208_(_004689_, _004747_, _004749_);
  or g_098209_(_004690_, _004748_, _004750_);
  and g_098210_(_004599_, _004605_, _004752_);
  or g_098211_(_004598_, _004604_, _004753_);
  and g_098212_(_004749_, _004753_, _004754_);
  or g_098213_(_004750_, _004752_, _004755_);
  or g_098214_(_004628_, _004752_, _004756_);
  and g_098215_(_004631_, _004754_, _004757_);
  or g_098216_(_004632_, _004755_, _004758_);
  and g_098217_(_004710_, _004737_, _004759_);
  or g_098218_(_004711_, _004736_, _004760_);
  and g_098219_(_004739_, _004759_, _004761_);
  or g_098220_(_004738_, _004760_, _004763_);
  and g_098221_(_004698_, _004706_, _004764_);
  or g_098222_(_004697_, _004764_, _004765_);
  not g_098223_(_004765_, _004766_);
  and g_098224_(_004763_, _004766_, _004767_);
  or g_098225_(_004761_, _004765_, _004768_);
  and g_098226_(_004689_, _004768_, _004769_);
  or g_098227_(_004690_, _004767_, _004770_);
  and g_098228_(_004661_, _004678_, _004771_);
  or g_098229_(_004660_, _004679_, _004772_);
  and g_098230_(_004675_, _004772_, _004774_);
  or g_098231_(_004673_, _004771_, _004775_);
  and g_098232_(_004682_, _004775_, _004776_);
  or g_098233_(_004683_, _004774_, _004777_);
  and g_098234_(_004770_, _004777_, _004778_);
  or g_098235_(_004769_, _004776_, _004779_);
  and g_098236_(_004645_, _004649_, _004780_);
  or g_098237_(_004644_, _004648_, _004781_);
  and g_098238_(_004758_, _004781_, _004782_);
  or g_098239_(_004757_, _004780_, _004783_);
  and g_098240_(_004778_, _004782_, _004785_);
  or g_098241_(_004779_, _004783_, _004786_);
  and g_098242_(_003156_, _004618_, _004787_);
  or g_098243_(_004606_, _004787_, _004788_);
  or g_098244_(_004756_, _004788_, _004789_);
  or g_098245_(_004625_, _004789_, _004790_);
  or g_098246_(_004750_, _004790_, _004791_);
  not g_098247_(_004791_, _004792_);
  and g_098248_(_004786_, _004791_, _004793_);
  or g_098249_(_004785_, _004792_, _004794_);
  and g_098250_(_003565_, _004793_, _004796_);
  or g_098251_(_003566_, _004794_, _004797_);
  and g_098252_(_004638_, _004794_, _004798_);
  or g_098253_(_004637_, _004793_, _004799_);
  and g_098254_(_004797_, _004799_, _004800_);
  or g_098255_(_004796_, _004798_, _004801_);
  xor g_098256_(out[122], _003269_, _004802_);
  xor g_098257_(_003343_, _003269_, _004803_);
  and g_098258_(_004800_, _004802_, _004804_);
  or g_098259_(_004801_, _004803_, _004805_);
  and g_098260_(_003258_, _003273_, _004807_);
  or g_098261_(_003259_, _003272_, _004808_);
  and g_098262_(_004805_, _004808_, _004809_);
  or g_098263_(_004804_, _004807_, _004810_);
  and g_098264_(_004801_, _004803_, _004811_);
  or g_098265_(_004800_, _004802_, _004812_);
  and g_098266_(_003259_, _003272_, _004813_);
  or g_098267_(_003258_, _003273_, _004814_);
  and g_098268_(out[121], _003268_, _004815_);
  xor g_098269_(out[121], _003268_, _004816_);
  or g_098270_(_003270_, _004815_, _004818_);
  and g_098271_(_004659_, _004794_, _004819_);
  or g_098272_(_004658_, _004793_, _004820_);
  and g_098273_(_004653_, _004793_, _004821_);
  or g_098274_(_004651_, _004794_, _004822_);
  and g_098275_(_004820_, _004822_, _004823_);
  or g_098276_(_004819_, _004821_, _004824_);
  and g_098277_(_004818_, _004823_, _004825_);
  or g_098278_(_004816_, _004824_, _004826_);
  xor g_098279_(out[120], _003267_, _004827_);
  xor g_098280_(_003321_, _003267_, _004829_);
  and g_098281_(_004670_, _004794_, _004830_);
  or g_098282_(_004669_, _004793_, _004831_);
  and g_098283_(_004664_, _004793_, _004832_);
  or g_098284_(_004662_, _004794_, _004833_);
  and g_098285_(_004831_, _004833_, _004834_);
  or g_098286_(_004830_, _004832_, _004835_);
  and g_098287_(_004827_, _004835_, _004836_);
  or g_098288_(_004829_, _004834_, _004837_);
  and g_098289_(_004816_, _004824_, _004838_);
  or g_098290_(_004818_, _004823_, _004840_);
  and g_098291_(_004829_, _004834_, _004841_);
  or g_098292_(_004827_, _004835_, _004842_);
  and g_098293_(_004812_, _004814_, _004843_);
  or g_098294_(_004811_, _004813_, _004844_);
  and g_098295_(_004809_, _004843_, _004845_);
  or g_098296_(_004810_, _004844_, _004846_);
  and g_098297_(_004837_, _004840_, _004847_);
  or g_098298_(_004836_, _004838_, _004848_);
  and g_098299_(_004826_, _004842_, _004849_);
  or g_098300_(_004825_, _004841_, _004851_);
  and g_098301_(_004847_, _004849_, _004852_);
  or g_098302_(_004848_, _004851_, _004853_);
  and g_098303_(_004845_, _004852_, _004854_);
  or g_098304_(_004846_, _004853_, _004855_);
  xor g_098305_(out[118], _003264_, _004856_);
  not g_098306_(_004856_, _004857_);
  or g_098307_(_004705_, _004793_, _004858_);
  or g_098308_(_004701_, _004794_, _004859_);
  and g_098309_(_004858_, _004859_, _004860_);
  not g_098310_(_004860_, _004862_);
  xor g_098311_(out[119], _003265_, _004863_);
  xor g_098312_(_003233_, _003265_, _004864_);
  or g_098313_(_004695_, _004793_, _004865_);
  or g_098314_(_004692_, _004794_, _004866_);
  and g_098315_(_004865_, _004866_, _004867_);
  not g_098316_(_004867_, _004868_);
  and g_098317_(_004864_, _004868_, _004869_);
  or g_098318_(_004863_, _004867_, _004870_);
  and g_098319_(_004857_, _004860_, _004871_);
  or g_098320_(_004856_, _004862_, _004873_);
  and g_098321_(_004863_, _004867_, _004874_);
  not g_098322_(_004874_, _004875_);
  xor g_098323_(_004857_, _004860_, _004876_);
  xor g_098324_(_004856_, _004860_, _004877_);
  and g_098325_(_004875_, _004876_, _004878_);
  or g_098326_(_004874_, _004877_, _004879_);
  and g_098327_(_004870_, _004878_, _004880_);
  or g_098328_(_004869_, _004879_, _004881_);
  or g_098329_(_012044_, _034110_, _004882_);
  not g_098330_(_004882_, _004884_);
  and g_098331_(_003263_, _004882_, _004885_);
  or g_098332_(_003262_, _004884_, _004886_);
  and g_098333_(_004722_, _004794_, _004887_);
  or g_098334_(_004721_, _004793_, _004888_);
  and g_098335_(_004715_, _004793_, _004889_);
  or g_098336_(_004714_, _004794_, _004890_);
  and g_098337_(_004888_, _004890_, _004891_);
  or g_098338_(_004887_, _004889_, _004892_);
  and g_098339_(_004886_, _004891_, _004893_);
  or g_098340_(_004885_, _004892_, _004895_);
  xor g_098341_(out[117], _003262_, _004896_);
  xor g_098342_(_003255_, _003262_, _004897_);
  and g_098343_(_004733_, _004794_, _004898_);
  or g_098344_(_004732_, _004793_, _004899_);
  and g_098345_(_004726_, _004793_, _004900_);
  or g_098346_(_004725_, _004794_, _004901_);
  and g_098347_(_004899_, _004901_, _004902_);
  or g_098348_(_004898_, _004900_, _004903_);
  and g_098349_(_004897_, _004902_, _004904_);
  or g_098350_(_004896_, _004903_, _004906_);
  and g_098351_(_004895_, _004906_, _004907_);
  or g_098352_(_004893_, _004904_, _004908_);
  and g_098353_(_004896_, _004903_, _004909_);
  or g_098354_(_004897_, _004902_, _004910_);
  and g_098355_(_004885_, _004892_, _004911_);
  or g_098356_(_004886_, _004891_, _004912_);
  and g_098357_(_004910_, _004912_, _004913_);
  or g_098358_(_004909_, _004911_, _004914_);
  and g_098359_(_004907_, _004913_, _004915_);
  or g_098360_(_004908_, _004914_, _004917_);
  or g_098361_(_004881_, _004917_, _004918_);
  and g_098362_(_004854_, _004915_, _004919_);
  and g_098363_(_004880_, _004919_, _004920_);
  or g_098364_(_004855_, _004918_, _004921_);
  or g_098365_(_003145_, _004794_, _004922_);
  or g_098366_(_004611_, _004793_, _004923_);
  and g_098367_(_004922_, _004923_, _004924_);
  and g_098368_(out[96], _004793_, _004925_);
  not g_098369_(_004925_, _004926_);
  or g_098370_(_004617_, _004793_, _004928_);
  not g_098371_(_004928_, _004929_);
  and g_098372_(_004926_, _004928_, _004930_);
  or g_098373_(_004925_, _004929_, _004931_);
  and g_098374_(out[112], _004930_, _004932_);
  or g_098375_(_003288_, _004931_, _004933_);
  and g_098376_(out[113], _004924_, _004934_);
  not g_098377_(_004934_, _004935_);
  xor g_098378_(out[113], _004924_, _004936_);
  xor g_098379_(_003277_, _004924_, _004937_);
  and g_098380_(_004933_, _004936_, _004939_);
  or g_098381_(_004932_, _004937_, _004940_);
  and g_098382_(_031206_, _004793_, _004941_);
  not g_098383_(_004941_, _004942_);
  or g_098384_(_004595_, _004793_, _004943_);
  not g_098385_(_004943_, _004944_);
  and g_098386_(_004942_, _004943_, _004945_);
  or g_098387_(_004941_, _004944_, _004946_);
  and g_098388_(_034121_, _004945_, _004947_);
  or g_098389_(_034132_, _004946_, _004948_);
  xor g_098390_(_034121_, _004945_, _004950_);
  xor g_098391_(_034132_, _004945_, _004951_);
  xor g_098392_(out[115], _034110_, _004952_);
  xor g_098393_(_003310_, _034110_, _004953_);
  and g_098394_(_004598_, _004793_, _004954_);
  not g_098395_(_004954_, _004955_);
  or g_098396_(_004604_, _004793_, _004956_);
  not g_098397_(_004956_, _004957_);
  and g_098398_(_004955_, _004956_, _004958_);
  or g_098399_(_004954_, _004957_, _004959_);
  and g_098400_(_004953_, _004959_, _004961_);
  or g_098401_(_004952_, _004958_, _004962_);
  and g_098402_(_004952_, _004958_, _004963_);
  or g_098403_(_004953_, _004959_, _004964_);
  and g_098404_(_003288_, _004931_, _004965_);
  or g_098405_(out[112], _004930_, _004966_);
  and g_098406_(_004950_, _004962_, _004967_);
  or g_098407_(_004951_, _004961_, _004968_);
  and g_098408_(_004964_, _004966_, _004969_);
  or g_098409_(_004963_, _004965_, _004970_);
  and g_098410_(_004967_, _004969_, _004972_);
  or g_098411_(_004968_, _004970_, _004973_);
  and g_098412_(_004939_, _004972_, _004974_);
  or g_098413_(_004940_, _004973_, _004975_);
  and g_098414_(_004920_, _004974_, _004976_);
  or g_098415_(_004921_, _004975_, _004977_);
  and g_098416_(_004948_, _004964_, _004978_);
  and g_098417_(_004935_, _004940_, _004979_);
  or g_098418_(_004934_, _004939_, _004980_);
  or g_098419_(_004951_, _004979_, _004981_);
  and g_098420_(_004978_, _004981_, _004983_);
  or g_098421_(_004921_, _004961_, _004984_);
  and g_098422_(_004947_, _004962_, _004985_);
  and g_098423_(_004967_, _004980_, _004986_);
  or g_098424_(_004985_, _004986_, _004987_);
  or g_098425_(_004963_, _004987_, _004988_);
  and g_098426_(_004920_, _004988_, _004989_);
  or g_098427_(_004983_, _004984_, _004990_);
  and g_098428_(_004908_, _004910_, _004991_);
  or g_098429_(_004907_, _004909_, _004992_);
  and g_098430_(_004880_, _004991_, _004994_);
  or g_098431_(_004881_, _004992_, _004995_);
  and g_098432_(_004870_, _004871_, _004996_);
  or g_098433_(_004869_, _004873_, _004997_);
  and g_098434_(_004875_, _004997_, _004998_);
  or g_098435_(_004874_, _004996_, _004999_);
  and g_098436_(_004995_, _004998_, _005000_);
  or g_098437_(_004994_, _004999_, _005001_);
  and g_098438_(_004854_, _005001_, _005002_);
  or g_098439_(_004855_, _005000_, _005003_);
  and g_098440_(_004826_, _004841_, _005005_);
  or g_098441_(_004825_, _004842_, _005006_);
  and g_098442_(_004840_, _005006_, _005007_);
  or g_098443_(_004838_, _005005_, _005008_);
  and g_098444_(_004845_, _005008_, _005009_);
  or g_098445_(_004846_, _005007_, _005010_);
  and g_098446_(_004810_, _004814_, _005011_);
  or g_098447_(_004809_, _004813_, _005012_);
  and g_098448_(_005010_, _005012_, _005013_);
  or g_098449_(_005009_, _005011_, _005014_);
  and g_098450_(_005003_, _005013_, _005016_);
  or g_098451_(_005002_, _005014_, _005017_);
  and g_098452_(_004990_, _005016_, _005018_);
  or g_098453_(_004989_, _005017_, _005019_);
  and g_098454_(_004977_, _005019_, _005020_);
  or g_098455_(_004976_, _005018_, _005021_);
  and g_098456_(_004801_, _005021_, _005022_);
  or g_098457_(_004800_, _005020_, _005023_);
  and g_098458_(_004802_, _005020_, _005024_);
  or g_098459_(_004803_, _005021_, _005025_);
  and g_098460_(_005023_, _005025_, _005027_);
  or g_098461_(_005022_, _005024_, _005028_);
  xor g_098462_(out[138], _003285_, _005029_);
  xor g_098463_(_003475_, _003285_, _005030_);
  and g_098464_(_005027_, _005029_, _005031_);
  or g_098465_(_005028_, _005030_, _005032_);
  and g_098466_(_003274_, _003290_, _005033_);
  or g_098467_(_003275_, _003289_, _005034_);
  and g_098468_(_005032_, _005034_, _005035_);
  or g_098469_(_005031_, _005033_, _005036_);
  and g_098470_(_005028_, _005030_, _005038_);
  or g_098471_(_005027_, _005029_, _005039_);
  and g_098472_(_003275_, _003289_, _005040_);
  or g_098473_(_003274_, _003290_, _005041_);
  and g_098474_(out[137], _003284_, _005042_);
  xor g_098475_(out[137], _003284_, _005043_);
  or g_098476_(_003286_, _005042_, _005044_);
  and g_098477_(_004824_, _005021_, _005045_);
  or g_098478_(_004823_, _005020_, _005046_);
  and g_098479_(_004818_, _005020_, _005047_);
  or g_098480_(_004816_, _005021_, _005049_);
  and g_098481_(_005046_, _005049_, _005050_);
  or g_098482_(_005045_, _005047_, _005051_);
  and g_098483_(_005044_, _005050_, _005052_);
  or g_098484_(_005043_, _005051_, _005053_);
  xor g_098485_(out[136], _003283_, _005054_);
  xor g_098486_(_003453_, _003283_, _005055_);
  and g_098487_(_004829_, _005020_, _005056_);
  or g_098488_(_004827_, _005021_, _005057_);
  or g_098489_(_004834_, _005020_, _005058_);
  not g_098490_(_005058_, _005060_);
  and g_098491_(_005057_, _005058_, _005061_);
  or g_098492_(_005056_, _005060_, _005062_);
  and g_098493_(_005054_, _005062_, _005063_);
  or g_098494_(_005055_, _005061_, _005064_);
  and g_098495_(_005043_, _005051_, _005065_);
  or g_098496_(_005044_, _005050_, _005066_);
  and g_098497_(_005055_, _005061_, _005067_);
  or g_098498_(_005054_, _005062_, _005068_);
  and g_098499_(_005066_, _005068_, _005069_);
  and g_098500_(_005039_, _005041_, _005071_);
  or g_098501_(_005038_, _005040_, _005072_);
  and g_098502_(_005035_, _005071_, _005073_);
  or g_098503_(_005036_, _005072_, _005074_);
  and g_098504_(_005064_, _005066_, _005075_);
  or g_098505_(_005063_, _005065_, _005076_);
  and g_098506_(_005053_, _005068_, _005077_);
  or g_098507_(_005052_, _005067_, _005078_);
  and g_098508_(_005075_, _005077_, _005079_);
  or g_098509_(_005076_, _005078_, _005080_);
  and g_098510_(_005073_, _005079_, _005082_);
  or g_098511_(_005074_, _005080_, _005083_);
  xor g_098512_(out[135], _003282_, _005084_);
  xor g_098513_(_003365_, _003282_, _005085_);
  or g_098514_(_004864_, _005021_, _005086_);
  or g_098515_(_004867_, _005020_, _005087_);
  and g_098516_(_005086_, _005087_, _005088_);
  or g_098517_(_005084_, _005088_, _005089_);
  xor g_098518_(out[134], _003281_, _005090_);
  not g_098519_(_005090_, _005091_);
  or g_098520_(_004856_, _005021_, _005093_);
  or g_098521_(_004860_, _005020_, _005094_);
  and g_098522_(_005093_, _005094_, _005095_);
  and g_098523_(_005091_, _005095_, _005096_);
  and g_098524_(_005084_, _005088_, _005097_);
  xor g_098525_(_005084_, _005088_, _005098_);
  xor g_098526_(_005085_, _005088_, _005099_);
  xor g_098527_(_005091_, _005095_, _005100_);
  xor g_098528_(_005090_, _005095_, _005101_);
  and g_098529_(_005098_, _005100_, _005102_);
  or g_098530_(_005099_, _005101_, _005104_);
  or g_098531_(_012198_, _036178_, _005105_);
  not g_098532_(_005105_, _005106_);
  and g_098533_(_003280_, _005105_, _005107_);
  or g_098534_(_003279_, _005106_, _005108_);
  and g_098535_(_004892_, _005021_, _005109_);
  or g_098536_(_004891_, _005020_, _005110_);
  and g_098537_(_004886_, _005020_, _005111_);
  or g_098538_(_004885_, _005021_, _005112_);
  and g_098539_(_005110_, _005112_, _005113_);
  or g_098540_(_005109_, _005111_, _005115_);
  and g_098541_(_005108_, _005113_, _005116_);
  or g_098542_(_005107_, _005115_, _005117_);
  xor g_098543_(out[133], _003279_, _005118_);
  xor g_098544_(_003387_, _003279_, _005119_);
  and g_098545_(_004897_, _005020_, _005120_);
  or g_098546_(_004896_, _005021_, _005121_);
  and g_098547_(_004903_, _005021_, _005122_);
  or g_098548_(_004902_, _005020_, _005123_);
  and g_098549_(_005121_, _005123_, _005124_);
  or g_098550_(_005120_, _005122_, _005126_);
  and g_098551_(_005119_, _005124_, _005127_);
  or g_098552_(_005118_, _005126_, _005128_);
  and g_098553_(_005117_, _005128_, _005129_);
  or g_098554_(_005116_, _005127_, _005130_);
  and g_098555_(_005118_, _005126_, _005131_);
  or g_098556_(_005119_, _005124_, _005132_);
  and g_098557_(_005107_, _005115_, _005133_);
  or g_098558_(_005108_, _005113_, _005134_);
  and g_098559_(_005132_, _005134_, _005135_);
  or g_098560_(_005131_, _005133_, _005137_);
  and g_098561_(_005129_, _005135_, _005138_);
  or g_098562_(_005130_, _005137_, _005139_);
  and g_098563_(_005102_, _005138_, _005140_);
  or g_098564_(_005104_, _005139_, _005141_);
  and g_098565_(_005082_, _005140_, _005142_);
  or g_098566_(_005083_, _005141_, _005143_);
  xor g_098567_(out[131], _036178_, _005144_);
  xor g_098568_(_003442_, _036178_, _005145_);
  or g_098569_(_004958_, _005020_, _005146_);
  or g_098570_(_004953_, _005021_, _005148_);
  and g_098571_(_005146_, _005148_, _005149_);
  or g_098572_(_005144_, _005149_, _005150_);
  or g_098573_(_034132_, _005021_, _005151_);
  or g_098574_(_004945_, _005020_, _005152_);
  and g_098575_(_005151_, _005152_, _005153_);
  and g_098576_(_036189_, _005153_, _005154_);
  and g_098577_(_005144_, _005149_, _005155_);
  or g_098578_(_005154_, _005155_, _005156_);
  or g_098579_(_003277_, _005021_, _005157_);
  or g_098580_(_004924_, _005020_, _005159_);
  and g_098581_(_005157_, _005159_, _005160_);
  and g_098582_(out[129], _005160_, _005161_);
  and g_098583_(out[112], _005020_, _005162_);
  or g_098584_(_003288_, _005021_, _005163_);
  and g_098585_(_004931_, _005021_, _005164_);
  or g_098586_(_004930_, _005020_, _005165_);
  and g_098587_(_005163_, _005165_, _005166_);
  or g_098588_(_005162_, _005164_, _005167_);
  or g_098589_(_003420_, _005167_, _005168_);
  xor g_098590_(out[129], _005160_, _005170_);
  and g_098591_(_005168_, _005170_, _005171_);
  not g_098592_(_005171_, _005172_);
  or g_098593_(_005161_, _005171_, _005173_);
  xor g_098594_(_036189_, _005153_, _005174_);
  xor g_098595_(_036200_, _005153_, _005175_);
  xor g_098596_(_005144_, _005149_, _005176_);
  xor g_098597_(_005145_, _005149_, _005177_);
  and g_098598_(_005174_, _005176_, _005178_);
  or g_098599_(_005175_, _005177_, _005179_);
  and g_098600_(_005173_, _005178_, _005181_);
  and g_098601_(_005150_, _005156_, _005182_);
  or g_098602_(_005181_, _005182_, _005183_);
  not g_098603_(_005183_, _005184_);
  and g_098604_(_005142_, _005183_, _005185_);
  or g_098605_(_005143_, _005184_, _005186_);
  and g_098606_(_005102_, _005130_, _005187_);
  or g_098607_(_005104_, _005129_, _005188_);
  and g_098608_(_005132_, _005187_, _005189_);
  or g_098609_(_005131_, _005188_, _005190_);
  and g_098610_(_005089_, _005096_, _005192_);
  or g_098611_(_005097_, _005192_, _005193_);
  not g_098612_(_005193_, _005194_);
  and g_098613_(_005190_, _005194_, _005195_);
  or g_098614_(_005189_, _005193_, _005196_);
  and g_098615_(_005082_, _005196_, _005197_);
  or g_098616_(_005083_, _005195_, _005198_);
  or g_098617_(_005069_, _005074_, _005199_);
  and g_098618_(_005053_, _005067_, _005200_);
  or g_098619_(_005065_, _005200_, _005201_);
  and g_098620_(_005073_, _005201_, _005203_);
  or g_098621_(_005052_, _005199_, _005204_);
  and g_098622_(_005036_, _005041_, _005205_);
  or g_098623_(_005035_, _005040_, _005206_);
  and g_098624_(_005204_, _005206_, _005207_);
  or g_098625_(_005203_, _005205_, _005208_);
  and g_098626_(_005198_, _005207_, _005209_);
  or g_098627_(_005197_, _005208_, _005210_);
  and g_098628_(_005186_, _005209_, _005211_);
  or g_098629_(_005185_, _005210_, _005212_);
  and g_098630_(_003420_, _005167_, _005214_);
  or g_098631_(out[128], _005166_, _005215_);
  and g_098632_(_005171_, _005178_, _005216_);
  or g_098633_(_005172_, _005179_, _005217_);
  and g_098634_(_005142_, _005216_, _005218_);
  or g_098635_(_005143_, _005217_, _005219_);
  and g_098636_(_005215_, _005218_, _005220_);
  or g_098637_(_005214_, _005219_, _005221_);
  and g_098638_(_005212_, _005221_, _005222_);
  or g_098639_(_005211_, _005220_, _005223_);
  and g_098640_(_005028_, _005223_, _005225_);
  or g_098641_(_005027_, _005222_, _005226_);
  and g_098642_(_005029_, _005222_, _005227_);
  or g_098643_(_005030_, _005223_, _005228_);
  and g_098644_(_005226_, _005228_, _005229_);
  or g_098645_(_005225_, _005227_, _005230_);
  xor g_098646_(out[154], _003302_, _005231_);
  xor g_098647_(_003607_, _003302_, _005232_);
  and g_098648_(_005229_, _005231_, _005233_);
  or g_098649_(_005230_, _005232_, _005234_);
  and g_098650_(_003291_, _003306_, _005236_);
  or g_098651_(_003292_, _003305_, _005237_);
  and g_098652_(_005234_, _005237_, _005238_);
  or g_098653_(_005233_, _005236_, _005239_);
  and g_098654_(_005230_, _005232_, _005240_);
  or g_098655_(_005229_, _005231_, _005241_);
  and g_098656_(_003292_, _003305_, _005242_);
  or g_098657_(_003291_, _003306_, _005243_);
  and g_098658_(out[153], _003301_, _005244_);
  xor g_098659_(out[153], _003301_, _005245_);
  or g_098660_(_003303_, _005244_, _005247_);
  and g_098661_(_005051_, _005223_, _005248_);
  or g_098662_(_005050_, _005222_, _005249_);
  and g_098663_(_005044_, _005222_, _005250_);
  or g_098664_(_005043_, _005223_, _005251_);
  and g_098665_(_005249_, _005251_, _005252_);
  or g_098666_(_005248_, _005250_, _005253_);
  and g_098667_(_005247_, _005252_, _005254_);
  or g_098668_(_005245_, _005253_, _005255_);
  xor g_098669_(out[152], _003300_, _005256_);
  xor g_098670_(_003585_, _003300_, _005258_);
  and g_098671_(_005055_, _005222_, _005259_);
  or g_098672_(_005054_, _005223_, _005260_);
  and g_098673_(_005062_, _005223_, _005261_);
  or g_098674_(_005061_, _005222_, _005262_);
  and g_098675_(_005260_, _005262_, _005263_);
  or g_098676_(_005259_, _005261_, _005264_);
  and g_098677_(_005256_, _005264_, _005265_);
  or g_098678_(_005258_, _005263_, _005266_);
  and g_098679_(_005245_, _005253_, _005267_);
  or g_098680_(_005247_, _005252_, _005269_);
  and g_098681_(_005258_, _005263_, _005270_);
  or g_098682_(_005256_, _005264_, _005271_);
  and g_098683_(_005241_, _005243_, _005272_);
  or g_098684_(_005240_, _005242_, _005273_);
  and g_098685_(_005238_, _005272_, _005274_);
  or g_098686_(_005239_, _005273_, _005275_);
  and g_098687_(_005266_, _005269_, _005276_);
  or g_098688_(_005265_, _005267_, _005277_);
  and g_098689_(_005255_, _005271_, _005278_);
  or g_098690_(_005254_, _005270_, _005280_);
  and g_098691_(_005276_, _005278_, _005281_);
  or g_098692_(_005277_, _005280_, _005282_);
  and g_098693_(_005274_, _005281_, _005283_);
  or g_098694_(_005275_, _005282_, _005284_);
  xor g_098695_(out[151], _003298_, _005285_);
  xor g_098696_(_003497_, _003298_, _005286_);
  or g_098697_(_005085_, _005223_, _005287_);
  or g_098698_(_005088_, _005222_, _005288_);
  and g_098699_(_005287_, _005288_, _005289_);
  or g_098700_(_005285_, _005289_, _005291_);
  xor g_098701_(out[150], _003297_, _005292_);
  xor g_098702_(_003508_, _003297_, _005293_);
  or g_098703_(_005090_, _005223_, _005294_);
  or g_098704_(_005095_, _005222_, _005295_);
  and g_098705_(_005294_, _005295_, _005296_);
  and g_098706_(_005293_, _005296_, _005297_);
  and g_098707_(_005285_, _005289_, _005298_);
  xor g_098708_(_005285_, _005289_, _005299_);
  xor g_098709_(_005286_, _005289_, _005300_);
  xor g_098710_(_005293_, _005296_, _005302_);
  xor g_098711_(_005292_, _005296_, _005303_);
  and g_098712_(_005299_, _005302_, _005304_);
  or g_098713_(_005300_, _005303_, _005305_);
  or g_098714_(_012352_, _038455_, _005306_);
  not g_098715_(_005306_, _005307_);
  and g_098716_(_003296_, _005306_, _005308_);
  or g_098717_(_003295_, _005307_, _005309_);
  and g_098718_(_005115_, _005223_, _005310_);
  or g_098719_(_005113_, _005222_, _005311_);
  and g_098720_(_005108_, _005222_, _005313_);
  or g_098721_(_005107_, _005223_, _005314_);
  and g_098722_(_005311_, _005314_, _005315_);
  or g_098723_(_005310_, _005313_, _005316_);
  and g_098724_(_005309_, _005315_, _005317_);
  or g_098725_(_005308_, _005316_, _005318_);
  xor g_098726_(out[149], _003295_, _005319_);
  xor g_098727_(_003519_, _003295_, _005320_);
  and g_098728_(_005119_, _005222_, _005321_);
  or g_098729_(_005118_, _005223_, _005322_);
  and g_098730_(_005126_, _005223_, _005324_);
  or g_098731_(_005124_, _005222_, _005325_);
  and g_098732_(_005322_, _005325_, _005326_);
  or g_098733_(_005321_, _005324_, _005327_);
  and g_098734_(_005320_, _005326_, _005328_);
  or g_098735_(_005319_, _005327_, _005329_);
  and g_098736_(_005318_, _005329_, _005330_);
  or g_098737_(_005317_, _005328_, _005331_);
  and g_098738_(_005308_, _005316_, _005332_);
  or g_098739_(_005309_, _005315_, _005333_);
  and g_098740_(_005319_, _005327_, _005335_);
  or g_098741_(_005320_, _005326_, _005336_);
  and g_098742_(_005333_, _005336_, _005337_);
  or g_098743_(_005332_, _005335_, _005338_);
  and g_098744_(_005330_, _005337_, _005339_);
  or g_098745_(_005331_, _005338_, _005340_);
  and g_098746_(_005304_, _005339_, _005341_);
  or g_098747_(_005305_, _005340_, _005342_);
  and g_098748_(_005283_, _005341_, _005343_);
  or g_098749_(_005284_, _005342_, _005344_);
  or g_098750_(_003409_, _005223_, _005346_);
  or g_098751_(_005160_, _005222_, _005347_);
  and g_098752_(_005346_, _005347_, _005348_);
  and g_098753_(out[128], _005222_, _005349_);
  not g_098754_(_005349_, _005350_);
  or g_098755_(_005166_, _005222_, _005351_);
  not g_098756_(_005351_, _005352_);
  and g_098757_(_005350_, _005351_, _005353_);
  or g_098758_(_005349_, _005352_, _005354_);
  and g_098759_(out[144], _005353_, _005355_);
  or g_098760_(_003552_, _005354_, _005357_);
  and g_098761_(out[145], _005348_, _005358_);
  not g_098762_(_005358_, _005359_);
  xor g_098763_(out[145], _005348_, _005360_);
  xor g_098764_(_003541_, _005348_, _005361_);
  and g_098765_(_005357_, _005360_, _005362_);
  or g_098766_(_005355_, _005361_, _005363_);
  or g_098767_(_005153_, _005222_, _005364_);
  not g_098768_(_005364_, _005365_);
  and g_098769_(_036189_, _005222_, _005366_);
  not g_098770_(_005366_, _005368_);
  and g_098771_(_005364_, _005368_, _005369_);
  or g_098772_(_005365_, _005366_, _005370_);
  and g_098773_(_038466_, _005369_, _005371_);
  or g_098774_(_038477_, _005370_, _005372_);
  xor g_098775_(_038466_, _005369_, _005373_);
  xor g_098776_(_038477_, _005369_, _005374_);
  xor g_098777_(out[147], _038455_, _005375_);
  xor g_098778_(_003574_, _038455_, _005376_);
  and g_098779_(_005144_, _005222_, _005377_);
  not g_098780_(_005377_, _005379_);
  or g_098781_(_005149_, _005222_, _005380_);
  not g_098782_(_005380_, _005381_);
  and g_098783_(_005379_, _005380_, _005382_);
  or g_098784_(_005377_, _005381_, _005383_);
  and g_098785_(_005375_, _005382_, _005384_);
  or g_098786_(_005376_, _005383_, _005385_);
  and g_098787_(_005376_, _005383_, _005386_);
  or g_098788_(_005375_, _005382_, _005387_);
  and g_098789_(_003552_, _005354_, _005388_);
  or g_098790_(out[144], _005353_, _005390_);
  and g_098791_(_005373_, _005387_, _005391_);
  or g_098792_(_005374_, _005386_, _005392_);
  and g_098793_(_005385_, _005390_, _005393_);
  or g_098794_(_005384_, _005388_, _005394_);
  and g_098795_(_005391_, _005393_, _005395_);
  or g_098796_(_005392_, _005394_, _005396_);
  and g_098797_(_005362_, _005395_, _005397_);
  or g_098798_(_005363_, _005396_, _005398_);
  and g_098799_(_005343_, _005397_, _005399_);
  or g_098800_(_005344_, _005398_, _005401_);
  and g_098801_(_005372_, _005385_, _005402_);
  or g_098802_(_005371_, _005384_, _005403_);
  and g_098803_(_005359_, _005363_, _005404_);
  or g_098804_(_005358_, _005362_, _005405_);
  and g_098805_(_005373_, _005405_, _005406_);
  or g_098806_(_005374_, _005404_, _005407_);
  and g_098807_(_005402_, _005407_, _005408_);
  or g_098808_(_005403_, _005406_, _005409_);
  and g_098809_(_005343_, _005387_, _005410_);
  or g_098810_(_005344_, _005386_, _005412_);
  and g_098811_(_005409_, _005410_, _005413_);
  or g_098812_(_005408_, _005412_, _005414_);
  and g_098813_(_005304_, _005331_, _005415_);
  or g_098814_(_005305_, _005330_, _005416_);
  and g_098815_(_005336_, _005415_, _005417_);
  or g_098816_(_005335_, _005416_, _005418_);
  and g_098817_(_005291_, _005297_, _005419_);
  or g_098818_(_005298_, _005419_, _005420_);
  not g_098819_(_005420_, _005421_);
  and g_098820_(_005418_, _005421_, _005423_);
  or g_098821_(_005417_, _005420_, _005424_);
  and g_098822_(_005283_, _005424_, _005425_);
  or g_098823_(_005284_, _005423_, _005426_);
  and g_098824_(_005255_, _005270_, _005427_);
  or g_098825_(_005254_, _005271_, _005428_);
  and g_098826_(_005269_, _005428_, _005429_);
  or g_098827_(_005267_, _005427_, _005430_);
  and g_098828_(_005274_, _005430_, _005431_);
  or g_098829_(_005275_, _005429_, _005432_);
  and g_098830_(_005239_, _005243_, _005434_);
  or g_098831_(_005238_, _005242_, _005435_);
  and g_098832_(_005432_, _005435_, _005436_);
  or g_098833_(_005431_, _005434_, _005437_);
  and g_098834_(_005426_, _005436_, _005438_);
  or g_098835_(_005425_, _005437_, _005439_);
  and g_098836_(_005414_, _005438_, _005440_);
  or g_098837_(_005413_, _005439_, _005441_);
  and g_098838_(_005401_, _005441_, _005442_);
  or g_098839_(_005399_, _005440_, _005443_);
  and g_098840_(_005230_, _005443_, _005445_);
  or g_098841_(_005229_, _005442_, _005446_);
  and g_098842_(_005231_, _005442_, _005447_);
  or g_098843_(_005232_, _005443_, _005448_);
  and g_098844_(_005446_, _005448_, _005449_);
  or g_098845_(_005445_, _005447_, _005450_);
  xor g_098846_(out[170], _003318_, _005451_);
  not g_098847_(_005451_, _005452_);
  and g_098848_(_005449_, _005451_, _005453_);
  or g_098849_(_005450_, _005452_, _005454_);
  and g_098850_(_003307_, _003322_, _005456_);
  or g_098851_(_003308_, _003320_, _005457_);
  and g_098852_(_005454_, _005457_, _005458_);
  or g_098853_(_005453_, _005456_, _005459_);
  and g_098854_(_003308_, _003320_, _005460_);
  or g_098855_(_003307_, _003322_, _005461_);
  and g_098856_(_005459_, _005461_, _005462_);
  or g_098857_(_005458_, _005460_, _005463_);
  and g_098858_(out[169], _003317_, _005464_);
  xor g_098859_(out[169], _003317_, _005465_);
  xor g_098860_(_003728_, _003317_, _005467_);
  and g_098861_(_005253_, _005443_, _005468_);
  or g_098862_(_005252_, _005442_, _005469_);
  and g_098863_(_005247_, _005442_, _005470_);
  or g_098864_(_005245_, _005443_, _005471_);
  and g_098865_(_005469_, _005471_, _005472_);
  or g_098866_(_005468_, _005470_, _005473_);
  and g_098867_(_005467_, _005472_, _005474_);
  or g_098868_(_005465_, _005473_, _005475_);
  and g_098869_(_005450_, _005452_, _005476_);
  or g_098870_(_005449_, _005451_, _005478_);
  and g_098871_(_005465_, _005473_, _005479_);
  or g_098872_(_005467_, _005472_, _005480_);
  xor g_098873_(out[168], _003316_, _005481_);
  xor g_098874_(_003717_, _003316_, _005482_);
  or g_098875_(_005263_, _005442_, _005483_);
  not g_098876_(_005483_, _005484_);
  and g_098877_(_005258_, _005442_, _005485_);
  not g_098878_(_005485_, _005486_);
  and g_098879_(_005483_, _005486_, _005487_);
  or g_098880_(_005484_, _005485_, _005489_);
  and g_098881_(_005482_, _005487_, _005490_);
  or g_098882_(_005481_, _005489_, _005491_);
  and g_098883_(_005481_, _005489_, _005492_);
  or g_098884_(_005482_, _005487_, _005493_);
  xor g_098885_(out[167], _003315_, _005494_);
  xor g_098886_(_003629_, _003315_, _005495_);
  or g_098887_(_005286_, _005443_, _005496_);
  or g_098888_(_005289_, _005442_, _005497_);
  and g_098889_(_005496_, _005497_, _005498_);
  not g_098890_(_005498_, _005500_);
  and g_098891_(_005494_, _005498_, _005501_);
  or g_098892_(_005494_, _005498_, _005502_);
  xor g_098893_(_005494_, _005498_, _005503_);
  xor g_098894_(_005495_, _005498_, _005504_);
  xor g_098895_(out[166], _003314_, _005505_);
  xor g_098896_(_003640_, _003314_, _005506_);
  or g_098897_(_005292_, _005443_, _005507_);
  or g_098898_(_005296_, _005442_, _005508_);
  and g_098899_(_005507_, _005508_, _005509_);
  and g_098900_(_005506_, _005509_, _005511_);
  xor g_098901_(_005506_, _005509_, _005512_);
  xor g_098902_(_005505_, _005509_, _005513_);
  and g_098903_(_005503_, _005512_, _005514_);
  or g_098904_(_005504_, _005513_, _005515_);
  xor g_098905_(out[165], _003312_, _005516_);
  xor g_098906_(_003651_, _003312_, _005517_);
  and g_098907_(_005320_, _005442_, _005518_);
  or g_098908_(_005319_, _005443_, _005519_);
  and g_098909_(_005327_, _005443_, _005520_);
  or g_098910_(_005326_, _005442_, _005522_);
  and g_098911_(_005519_, _005522_, _005523_);
  or g_098912_(_005518_, _005520_, _005524_);
  and g_098913_(_005516_, _005524_, _005525_);
  or g_098914_(_005517_, _005523_, _005526_);
  or g_098915_(_012506_, _040556_, _005527_);
  not g_098916_(_005527_, _005528_);
  and g_098917_(_003313_, _005527_, _005529_);
  or g_098918_(_003312_, _005528_, _005530_);
  and g_098919_(_005316_, _005443_, _005531_);
  or g_098920_(_005315_, _005442_, _005533_);
  and g_098921_(_005309_, _005442_, _005534_);
  or g_098922_(_005308_, _005443_, _005535_);
  and g_098923_(_005533_, _005535_, _005536_);
  or g_098924_(_005531_, _005534_, _005537_);
  and g_098925_(_005530_, _005536_, _005538_);
  or g_098926_(_005529_, _005537_, _005539_);
  and g_098927_(_005517_, _005523_, _005540_);
  or g_098928_(_005516_, _005524_, _005541_);
  and g_098929_(_005539_, _005541_, _005542_);
  or g_098930_(_005538_, _005540_, _005544_);
  and g_098931_(_005514_, _005544_, _005545_);
  or g_098932_(_005515_, _005542_, _005546_);
  and g_098933_(_005526_, _005545_, _005547_);
  or g_098934_(_005525_, _005546_, _005548_);
  and g_098935_(_005502_, _005511_, _005549_);
  or g_098936_(_005501_, _005549_, _005550_);
  not g_098937_(_005550_, _005551_);
  and g_098938_(_005548_, _005551_, _005552_);
  or g_098939_(_005547_, _005550_, _005553_);
  or g_098940_(_038477_, _005443_, _005555_);
  or g_098941_(_005369_, _005442_, _005556_);
  and g_098942_(_005555_, _005556_, _005557_);
  and g_098943_(_040567_, _005557_, _005558_);
  xor g_098944_(out[163], _040556_, _005559_);
  xor g_098945_(_003706_, _040556_, _005560_);
  or g_098946_(_005382_, _005442_, _005561_);
  not g_098947_(_005561_, _005562_);
  and g_098948_(_005375_, _005442_, _005563_);
  not g_098949_(_005563_, _005564_);
  and g_098950_(_005561_, _005564_, _005566_);
  or g_098951_(_005562_, _005563_, _005567_);
  and g_098952_(_005559_, _005566_, _005568_);
  or g_098953_(_005560_, _005567_, _005569_);
  or g_098954_(_005558_, _005568_, _005570_);
  or g_098955_(_003541_, _005443_, _005571_);
  or g_098956_(_005348_, _005442_, _005572_);
  and g_098957_(_005571_, _005572_, _005573_);
  and g_098958_(out[161], _005573_, _005574_);
  and g_098959_(out[144], _005442_, _005575_);
  not g_098960_(_005575_, _005577_);
  and g_098961_(_005354_, _005443_, _005578_);
  or g_098962_(_005353_, _005442_, _005579_);
  and g_098963_(_005577_, _005579_, _005580_);
  or g_098964_(_005575_, _005578_, _005581_);
  or g_098965_(_003684_, _005581_, _005582_);
  xor g_098966_(out[161], _005573_, _005583_);
  and g_098967_(_005582_, _005583_, _005584_);
  or g_098968_(_005574_, _005584_, _005585_);
  xor g_098969_(_040567_, _005557_, _005586_);
  and g_098970_(_005569_, _005586_, _005588_);
  and g_098971_(_005585_, _005588_, _005589_);
  or g_098972_(_005570_, _005589_, _005590_);
  or g_098973_(_005530_, _005536_, _005591_);
  or g_098974_(_005559_, _005566_, _005592_);
  and g_098975_(_005458_, _005461_, _005593_);
  or g_098976_(_005459_, _005460_, _005594_);
  and g_098977_(_005478_, _005593_, _005595_);
  or g_098978_(_005476_, _005594_, _005596_);
  and g_098979_(_005480_, _005493_, _005597_);
  or g_098980_(_005479_, _005492_, _005599_);
  and g_098981_(_005475_, _005491_, _005600_);
  or g_098982_(_005474_, _005490_, _005601_);
  and g_098983_(_005597_, _005600_, _005602_);
  or g_098984_(_005599_, _005601_, _005603_);
  and g_098985_(_005595_, _005602_, _005604_);
  or g_098986_(_005596_, _005603_, _005605_);
  and g_098987_(_005526_, _005591_, _005606_);
  and g_098988_(_005542_, _005606_, _005607_);
  and g_098989_(_005514_, _005607_, _005608_);
  and g_098990_(_005604_, _005608_, _005610_);
  and g_098991_(_005590_, _005610_, _005611_);
  and g_098992_(_005592_, _005611_, _005612_);
  not g_098993_(_005612_, _005613_);
  and g_098994_(_005553_, _005604_, _005614_);
  or g_098995_(_005552_, _005605_, _005615_);
  and g_098996_(_005475_, _005490_, _005616_);
  or g_098997_(_005474_, _005491_, _005617_);
  and g_098998_(_005480_, _005617_, _005618_);
  or g_098999_(_005479_, _005616_, _005619_);
  and g_099000_(_005595_, _005619_, _005621_);
  or g_099001_(_005596_, _005618_, _005622_);
  and g_099002_(_005615_, _005622_, _005623_);
  or g_099003_(_005614_, _005621_, _005624_);
  or g_099004_(_005612_, _005624_, _005625_);
  and g_099005_(_005613_, _005623_, _005626_);
  and g_099006_(_005463_, _005626_, _005627_);
  or g_099007_(_005462_, _005625_, _005628_);
  or g_099008_(out[160], _005580_, _005629_);
  and g_099009_(_005592_, _005629_, _005630_);
  and g_099010_(_005588_, _005630_, _005632_);
  and g_099011_(_005610_, _005632_, _005633_);
  and g_099012_(_005584_, _005633_, _005634_);
  not g_099013_(_005634_, _005635_);
  and g_099014_(_005628_, _005635_, _005636_);
  or g_099015_(_005627_, _005634_, _005637_);
  and g_099016_(_005450_, _005637_, _005638_);
  or g_099017_(_005449_, _005636_, _005639_);
  and g_099018_(_005451_, _005636_, _005640_);
  or g_099019_(_005452_, _005637_, _005641_);
  and g_099020_(_005639_, _005641_, _005643_);
  or g_099021_(_005638_, _005640_, _005644_);
  xor g_099022_(out[186], _003334_, _005645_);
  not g_099023_(_005645_, _005646_);
  and g_099024_(_005644_, _005646_, _005647_);
  or g_099025_(_005643_, _005645_, _005648_);
  and g_099026_(_005643_, _005645_, _005649_);
  or g_099027_(_005644_, _005646_, _005650_);
  and g_099028_(_003323_, _003338_, _005651_);
  or g_099029_(_003324_, _003337_, _005652_);
  and g_099030_(_003324_, _003337_, _005654_);
  or g_099031_(_003323_, _003338_, _005655_);
  and g_099032_(_005648_, _005652_, _005656_);
  or g_099033_(_005647_, _005651_, _005657_);
  and g_099034_(_005650_, _005655_, _005658_);
  or g_099035_(_005649_, _005654_, _005659_);
  and g_099036_(_005656_, _005658_, _005660_);
  or g_099037_(_005657_, _005659_, _005661_);
  xor g_099038_(out[184], _003331_, _005662_);
  xor g_099039_(_003849_, _003331_, _005663_);
  and g_099040_(_005482_, _005636_, _005665_);
  or g_099041_(_005481_, _005637_, _005666_);
  and g_099042_(_005489_, _005637_, _005667_);
  or g_099043_(_005487_, _005636_, _005668_);
  and g_099044_(_005666_, _005668_, _005669_);
  or g_099045_(_005665_, _005667_, _005670_);
  and g_099046_(_005663_, _005669_, _005671_);
  or g_099047_(_005662_, _005670_, _005672_);
  and g_099048_(out[185], _003333_, _005673_);
  xor g_099049_(out[185], _003333_, _005674_);
  or g_099050_(_003335_, _005673_, _005676_);
  and g_099051_(_005473_, _005637_, _005677_);
  or g_099052_(_005472_, _005636_, _005678_);
  and g_099053_(_005467_, _005636_, _005679_);
  or g_099054_(_005465_, _005637_, _005680_);
  and g_099055_(_005678_, _005680_, _005681_);
  or g_099056_(_005677_, _005679_, _005682_);
  and g_099057_(_005674_, _005682_, _005683_);
  or g_099058_(_005676_, _005681_, _005684_);
  and g_099059_(_005672_, _005684_, _005685_);
  or g_099060_(_005671_, _005683_, _005687_);
  and g_099061_(_005676_, _005681_, _005688_);
  or g_099062_(_005674_, _005682_, _005689_);
  and g_099063_(_005662_, _005670_, _005690_);
  or g_099064_(_005663_, _005669_, _005691_);
  and g_099065_(_005689_, _005691_, _005692_);
  or g_099066_(_005688_, _005690_, _005693_);
  and g_099067_(_005685_, _005692_, _005694_);
  or g_099068_(_005687_, _005693_, _005695_);
  and g_099069_(_005660_, _005694_, _005696_);
  or g_099070_(_005661_, _005695_, _005698_);
  xor g_099071_(out[183], _003330_, _005699_);
  xor g_099072_(_003761_, _003330_, _005700_);
  and g_099073_(_005494_, _005636_, _005701_);
  or g_099074_(_005495_, _005637_, _005702_);
  and g_099075_(_005500_, _005637_, _005703_);
  or g_099076_(_005498_, _005636_, _005704_);
  and g_099077_(_005702_, _005704_, _005705_);
  or g_099078_(_005701_, _005703_, _005706_);
  and g_099079_(_005700_, _005706_, _005707_);
  or g_099080_(_005699_, _005705_, _005709_);
  and g_099081_(_005699_, _005705_, _005710_);
  or g_099082_(_005700_, _005706_, _005711_);
  and g_099083_(_005709_, _005711_, _005712_);
  or g_099084_(_005707_, _005710_, _005713_);
  xor g_099085_(out[182], _003329_, _005714_);
  not g_099086_(_005714_, _005715_);
  and g_099087_(_005506_, _005636_, _005716_);
  not g_099088_(_005716_, _005717_);
  or g_099089_(_005509_, _005636_, _005718_);
  not g_099090_(_005718_, _005720_);
  and g_099091_(_005717_, _005718_, _005721_);
  or g_099092_(_005716_, _005720_, _005722_);
  and g_099093_(_005715_, _005721_, _005723_);
  or g_099094_(_005714_, _005722_, _005724_);
  xor g_099095_(out[181], _003327_, _005725_);
  xor g_099096_(_003783_, _003327_, _005726_);
  and g_099097_(_005517_, _005636_, _005727_);
  not g_099098_(_005727_, _005728_);
  or g_099099_(_005523_, _005636_, _005729_);
  not g_099100_(_005729_, _005731_);
  and g_099101_(_005728_, _005729_, _005732_);
  or g_099102_(_005727_, _005731_, _005733_);
  and g_099103_(_005725_, _005733_, _005734_);
  or g_099104_(_005726_, _005732_, _005735_);
  xor g_099105_(_005715_, _005721_, _005736_);
  xor g_099106_(_005714_, _005721_, _005737_);
  and g_099107_(_005712_, _005736_, _005738_);
  or g_099108_(_005713_, _005737_, _005739_);
  and g_099109_(_005735_, _005738_, _005740_);
  or g_099110_(_005734_, _005739_, _005742_);
  and g_099111_(_005696_, _005740_, _005743_);
  or g_099112_(_005698_, _005742_, _005744_);
  or g_099113_(_012660_, _042679_, _005745_);
  not g_099114_(_005745_, _005746_);
  and g_099115_(_003328_, _005745_, _005747_);
  or g_099116_(_003327_, _005746_, _005748_);
  or g_099117_(_005536_, _005636_, _005749_);
  not g_099118_(_005749_, _005750_);
  and g_099119_(_005530_, _005636_, _005751_);
  not g_099120_(_005751_, _005753_);
  and g_099121_(_005749_, _005753_, _005754_);
  or g_099122_(_005750_, _005751_, _005755_);
  and g_099123_(_005748_, _005754_, _005756_);
  or g_099124_(_005747_, _005755_, _005757_);
  and g_099125_(_005726_, _005732_, _005758_);
  or g_099126_(_005725_, _005733_, _005759_);
  and g_099127_(_005757_, _005759_, _005760_);
  or g_099128_(_005756_, _005758_, _005761_);
  and g_099129_(_005747_, _005755_, _005762_);
  or g_099130_(_005748_, _005754_, _005764_);
  and g_099131_(_005760_, _005764_, _005765_);
  or g_099132_(_005761_, _005762_, _005766_);
  and g_099133_(_005743_, _005765_, _005767_);
  or g_099134_(_005744_, _005766_, _005768_);
  xor g_099135_(out[179], _042679_, _005769_);
  xor g_099136_(_003838_, _042679_, _005770_);
  and g_099137_(_005567_, _005637_, _005771_);
  or g_099138_(_005566_, _005636_, _005772_);
  and g_099139_(_005559_, _005636_, _005773_);
  or g_099140_(_005560_, _005637_, _005775_);
  and g_099141_(_005772_, _005775_, _005776_);
  or g_099142_(_005771_, _005773_, _005777_);
  and g_099143_(_005769_, _005776_, _005778_);
  or g_099144_(_005770_, _005777_, _005779_);
  and g_099145_(_040567_, _005636_, _005780_);
  not g_099146_(_005780_, _005781_);
  or g_099147_(_005557_, _005636_, _005782_);
  not g_099148_(_005782_, _005783_);
  and g_099149_(_005781_, _005782_, _005784_);
  or g_099150_(_005780_, _005783_, _005786_);
  and g_099151_(_005770_, _005777_, _005787_);
  or g_099152_(_005769_, _005776_, _005788_);
  and g_099153_(_042690_, _005784_, _005789_);
  or g_099154_(_042701_, _005786_, _005790_);
  xor g_099155_(_042690_, _005784_, _005791_);
  xor g_099156_(_042701_, _005784_, _005792_);
  and g_099157_(_005779_, _005788_, _005793_);
  or g_099158_(_005778_, _005787_, _005794_);
  and g_099159_(_005791_, _005793_, _005795_);
  or g_099160_(_005792_, _005794_, _005797_);
  and g_099161_(out[161], _005636_, _005798_);
  not g_099162_(_005798_, _005799_);
  or g_099163_(_005573_, _005636_, _005800_);
  not g_099164_(_005800_, _005801_);
  and g_099165_(_005799_, _005800_, _005802_);
  or g_099166_(_005798_, _005801_, _005803_);
  and g_099167_(out[177], _005802_, _005804_);
  or g_099168_(_003805_, _005803_, _005805_);
  and g_099169_(_005788_, _005789_, _005806_);
  or g_099170_(_005787_, _005790_, _005808_);
  and g_099171_(_005779_, _005808_, _005809_);
  or g_099172_(_005778_, _005806_, _005810_);
  and g_099173_(out[160], _005636_, _005811_);
  not g_099174_(_005811_, _005812_);
  or g_099175_(_005580_, _005636_, _005813_);
  not g_099176_(_005813_, _005814_);
  and g_099177_(_005812_, _005813_, _005815_);
  or g_099178_(_005811_, _005814_, _005816_);
  and g_099179_(out[176], _005815_, _005817_);
  or g_099180_(_003816_, _005816_, _005819_);
  xor g_099181_(out[177], _005802_, _005820_);
  xor g_099182_(_003805_, _005802_, _005821_);
  and g_099183_(_005819_, _005820_, _005822_);
  or g_099184_(_005817_, _005821_, _005823_);
  and g_099185_(_005795_, _005822_, _005824_);
  or g_099186_(_005797_, _005823_, _005825_);
  and g_099187_(_005805_, _005823_, _005826_);
  or g_099188_(_005804_, _005822_, _005827_);
  and g_099189_(_005795_, _005827_, _005828_);
  or g_099190_(_005797_, _005826_, _005830_);
  and g_099191_(_005809_, _005830_, _005831_);
  or g_099192_(_005810_, _005828_, _005832_);
  and g_099193_(_005767_, _005832_, _005833_);
  or g_099194_(_005768_, _005831_, _005834_);
  and g_099195_(_005743_, _005761_, _005835_);
  or g_099196_(_005744_, _005760_, _005836_);
  and g_099197_(_005711_, _005724_, _005837_);
  or g_099198_(_005710_, _005723_, _005838_);
  and g_099199_(_005709_, _005838_, _005839_);
  or g_099200_(_005707_, _005837_, _005841_);
  and g_099201_(_005696_, _005839_, _005842_);
  or g_099202_(_005698_, _005841_, _005843_);
  and g_099203_(_005687_, _005689_, _005844_);
  or g_099204_(_005685_, _005688_, _005845_);
  and g_099205_(_005660_, _005844_, _005846_);
  or g_099206_(_005661_, _005845_, _005847_);
  and g_099207_(_005650_, _005652_, _005848_);
  or g_099208_(_005649_, _005651_, _005849_);
  and g_099209_(_005655_, _005849_, _005850_);
  or g_099210_(_005654_, _005848_, _005852_);
  and g_099211_(_005847_, _005852_, _005853_);
  or g_099212_(_005846_, _005850_, _005854_);
  and g_099213_(_005843_, _005853_, _005855_);
  or g_099214_(_005842_, _005854_, _005856_);
  and g_099215_(_005836_, _005855_, _005857_);
  or g_099216_(_005835_, _005856_, _005858_);
  and g_099217_(_005834_, _005857_, _005859_);
  or g_099218_(_005833_, _005858_, _005860_);
  and g_099219_(_003816_, _005816_, _005861_);
  or g_099220_(out[176], _005815_, _005863_);
  and g_099221_(_005824_, _005863_, _005864_);
  or g_099222_(_005825_, _005861_, _005865_);
  and g_099223_(_005767_, _005864_, _005866_);
  or g_099224_(_005768_, _005865_, _005867_);
  and g_099225_(_005860_, _005867_, _005868_);
  or g_099226_(_005859_, _005866_, _005869_);
  and g_099227_(_005644_, _005869_, _005870_);
  and g_099228_(_005645_, _005868_, _005871_);
  or g_099229_(_005870_, _005871_, _005872_);
  xor g_099230_(out[202], _003350_, _005874_);
  xor g_099231_(out[202], _003351_, _005875_);
  or g_099232_(_005872_, _005875_, _005876_);
  or g_099233_(_003340_, _003353_, _005877_);
  and g_099234_(_005876_, _005877_, _005878_);
  and g_099235_(_003340_, _003353_, _005879_);
  xor g_099236_(_005872_, _005875_, _005880_);
  xor g_099237_(_005872_, _005874_, _005881_);
  xor g_099238_(_003340_, _003353_, _005882_);
  xor g_099239_(_003339_, _003353_, _005883_);
  and g_099240_(_005880_, _005882_, _005885_);
  or g_099241_(_005881_, _005883_, _005886_);
  xor g_099242_(out[200], _003348_, _005887_);
  xor g_099243_(_003981_, _003348_, _005888_);
  and g_099244_(_005663_, _005868_, _005889_);
  or g_099245_(_005662_, _005869_, _005890_);
  and g_099246_(_005670_, _005869_, _005891_);
  or g_099247_(_005669_, _005868_, _005892_);
  and g_099248_(_005890_, _005892_, _005893_);
  or g_099249_(_005889_, _005891_, _005894_);
  and g_099250_(_005888_, _005893_, _005896_);
  or g_099251_(_005887_, _005894_, _005897_);
  and g_099252_(out[201], _003349_, _005898_);
  xor g_099253_(out[201], _003349_, _005899_);
  or g_099254_(_003351_, _005898_, _005900_);
  and g_099255_(_005682_, _005869_, _005901_);
  or g_099256_(_005681_, _005868_, _005902_);
  and g_099257_(_005676_, _005868_, _005903_);
  or g_099258_(_005674_, _005869_, _005904_);
  and g_099259_(_005902_, _005904_, _005905_);
  or g_099260_(_005901_, _005903_, _005907_);
  and g_099261_(_005899_, _005907_, _005908_);
  or g_099262_(_005900_, _005905_, _005909_);
  and g_099263_(_005897_, _005909_, _005910_);
  or g_099264_(_005896_, _005908_, _005911_);
  and g_099265_(_005887_, _005894_, _005912_);
  or g_099266_(_005888_, _005893_, _005913_);
  and g_099267_(_005900_, _005905_, _005914_);
  or g_099268_(_005899_, _005907_, _005915_);
  and g_099269_(_005913_, _005915_, _005916_);
  or g_099270_(_005912_, _005914_, _005918_);
  and g_099271_(_005910_, _005916_, _005919_);
  or g_099272_(_005911_, _005918_, _005920_);
  and g_099273_(_005885_, _005919_, _005921_);
  or g_099274_(_005886_, _005920_, _005922_);
  xor g_099275_(out[199], _003347_, _005923_);
  xor g_099276_(_003893_, _003347_, _005924_);
  and g_099277_(_005699_, _005868_, _005925_);
  or g_099278_(_005700_, _005869_, _005926_);
  and g_099279_(_005706_, _005869_, _005927_);
  or g_099280_(_005705_, _005868_, _005929_);
  and g_099281_(_005926_, _005929_, _005930_);
  or g_099282_(_005925_, _005927_, _005931_);
  and g_099283_(_005924_, _005931_, _005932_);
  or g_099284_(_005923_, _005930_, _005933_);
  xor g_099285_(out[198], _003346_, _005934_);
  not g_099286_(_005934_, _005935_);
  or g_099287_(_005714_, _005869_, _005936_);
  or g_099288_(_005721_, _005868_, _005937_);
  and g_099289_(_005936_, _005937_, _005938_);
  not g_099290_(_005938_, _005940_);
  and g_099291_(_005935_, _005938_, _005941_);
  or g_099292_(_005934_, _005940_, _005942_);
  and g_099293_(_005923_, _005930_, _005943_);
  or g_099294_(_005924_, _005931_, _005944_);
  and g_099295_(_005933_, _005944_, _005945_);
  or g_099296_(_005932_, _005943_, _005946_);
  xor g_099297_(_005935_, _005938_, _005947_);
  xor g_099298_(_005934_, _005938_, _005948_);
  and g_099299_(_005945_, _005947_, _005949_);
  or g_099300_(_005946_, _005948_, _005951_);
  or g_099301_(_012814_, _044516_, _005952_);
  not g_099302_(_005952_, _005953_);
  and g_099303_(_003345_, _005952_, _005954_);
  or g_099304_(_003344_, _005953_, _005955_);
  and g_099305_(_005755_, _005869_, _005956_);
  or g_099306_(_005754_, _005868_, _005957_);
  and g_099307_(_005748_, _005868_, _005958_);
  or g_099308_(_005747_, _005869_, _005959_);
  and g_099309_(_005957_, _005959_, _005960_);
  or g_099310_(_005956_, _005958_, _005962_);
  and g_099311_(_005955_, _005960_, _005963_);
  or g_099312_(_005954_, _005962_, _005964_);
  xor g_099313_(out[197], _003344_, _005965_);
  xor g_099314_(_003915_, _003344_, _005966_);
  and g_099315_(_005726_, _005868_, _005967_);
  or g_099316_(_005725_, _005869_, _005968_);
  and g_099317_(_005733_, _005869_, _005969_);
  or g_099318_(_005732_, _005868_, _005970_);
  and g_099319_(_005968_, _005970_, _005971_);
  or g_099320_(_005967_, _005969_, _005973_);
  and g_099321_(_005966_, _005971_, _005974_);
  or g_099322_(_005965_, _005973_, _005975_);
  and g_099323_(_005964_, _005975_, _005976_);
  or g_099324_(_005963_, _005974_, _005977_);
  and g_099325_(_005965_, _005973_, _005978_);
  or g_099326_(_005966_, _005971_, _005979_);
  and g_099327_(_005954_, _005962_, _005980_);
  or g_099328_(_005955_, _005960_, _005981_);
  and g_099329_(_005979_, _005981_, _005982_);
  or g_099330_(_005978_, _005980_, _005984_);
  xor g_099331_(out[195], _044516_, _005985_);
  xor g_099332_(_003970_, _044516_, _005986_);
  and g_099333_(_005769_, _005868_, _005987_);
  or g_099334_(_005770_, _005869_, _005988_);
  and g_099335_(_005777_, _005869_, _005989_);
  or g_099336_(_005776_, _005868_, _005990_);
  and g_099337_(_005988_, _005990_, _005991_);
  or g_099338_(_005987_, _005989_, _005992_);
  and g_099339_(_005986_, _005992_, _005993_);
  or g_099340_(_005985_, _005991_, _005995_);
  and g_099341_(_005982_, _005995_, _005996_);
  or g_099342_(_005984_, _005993_, _005997_);
  and g_099343_(_005976_, _005996_, _005998_);
  or g_099344_(_005977_, _005997_, _005999_);
  and g_099345_(_005949_, _005998_, _006000_);
  or g_099346_(_005951_, _005999_, _006001_);
  and g_099347_(_005921_, _006000_, _006002_);
  or g_099348_(_005922_, _006001_, _006003_);
  and g_099349_(_005786_, _005869_, _006004_);
  or g_099350_(_005784_, _005868_, _006006_);
  and g_099351_(_042690_, _005868_, _006007_);
  or g_099352_(_042701_, _005869_, _006008_);
  and g_099353_(_006006_, _006008_, _006009_);
  or g_099354_(_006004_, _006007_, _006010_);
  and g_099355_(_044527_, _006009_, _006011_);
  or g_099356_(_044538_, _006010_, _006012_);
  and g_099357_(_005985_, _005991_, _006013_);
  or g_099358_(_005986_, _005992_, _006014_);
  and g_099359_(_006012_, _006014_, _006015_);
  or g_099360_(_006011_, _006013_, _006017_);
  and g_099361_(out[177], _005868_, _006018_);
  or g_099362_(_003805_, _005869_, _006019_);
  and g_099363_(_005803_, _005869_, _006020_);
  or g_099364_(_005802_, _005868_, _006021_);
  and g_099365_(_006019_, _006021_, _006022_);
  or g_099366_(_006018_, _006020_, _006023_);
  and g_099367_(out[193], _006022_, _006024_);
  or g_099368_(_003937_, _006023_, _006025_);
  and g_099369_(out[176], _005868_, _006026_);
  or g_099370_(_003816_, _005869_, _006028_);
  and g_099371_(_005816_, _005869_, _006029_);
  or g_099372_(_005815_, _005868_, _006030_);
  and g_099373_(_006028_, _006030_, _006031_);
  or g_099374_(_006026_, _006029_, _006032_);
  and g_099375_(out[192], _006031_, _006033_);
  or g_099376_(_003948_, _006032_, _006034_);
  xor g_099377_(out[193], _006022_, _006035_);
  xor g_099378_(_003937_, _006022_, _006036_);
  and g_099379_(_006034_, _006035_, _006037_);
  or g_099380_(_006033_, _006036_, _006039_);
  and g_099381_(_006025_, _006039_, _006040_);
  or g_099382_(_006024_, _006037_, _006041_);
  xor g_099383_(_044527_, _006009_, _006042_);
  xor g_099384_(_044538_, _006009_, _006043_);
  and g_099385_(_006041_, _006042_, _006044_);
  or g_099386_(_006040_, _006043_, _006045_);
  and g_099387_(_006015_, _006045_, _006046_);
  or g_099388_(_006017_, _006044_, _006047_);
  and g_099389_(_006002_, _006047_, _006048_);
  or g_099390_(_006003_, _006046_, _006050_);
  and g_099391_(_005977_, _005979_, _006051_);
  or g_099392_(_005976_, _005978_, _006052_);
  and g_099393_(_005949_, _006051_, _006053_);
  or g_099394_(_005951_, _006052_, _006054_);
  and g_099395_(_005933_, _005941_, _006055_);
  or g_099396_(_005932_, _005942_, _006056_);
  and g_099397_(_005944_, _006056_, _006057_);
  or g_099398_(_005943_, _006055_, _006058_);
  and g_099399_(_006054_, _006057_, _006059_);
  or g_099400_(_006053_, _006058_, _006061_);
  and g_099401_(_005921_, _006061_, _006062_);
  or g_099402_(_005922_, _006059_, _006063_);
  or g_099403_(_005878_, _005879_, _006064_);
  not g_099404_(_006064_, _006065_);
  and g_099405_(_005885_, _005911_, _006066_);
  or g_099406_(_005886_, _005910_, _006067_);
  and g_099407_(_005915_, _006066_, _006068_);
  or g_099408_(_005914_, _006067_, _006069_);
  and g_099409_(_006064_, _006069_, _006070_);
  or g_099410_(_006065_, _006068_, _006072_);
  and g_099411_(_006063_, _006070_, _006073_);
  or g_099412_(_006062_, _006072_, _006074_);
  and g_099413_(_006050_, _006073_, _006075_);
  or g_099414_(_006048_, _006074_, _006076_);
  and g_099415_(_003948_, _006032_, _006077_);
  or g_099416_(out[192], _006031_, _006078_);
  and g_099417_(_006014_, _006078_, _006079_);
  or g_099418_(_006013_, _006077_, _006080_);
  and g_099419_(_006042_, _006079_, _006081_);
  or g_099420_(_006043_, _006080_, _006083_);
  and g_099421_(_006037_, _006081_, _006084_);
  or g_099422_(_006039_, _006083_, _006085_);
  and g_099423_(_006002_, _006084_, _006086_);
  or g_099424_(_006003_, _006085_, _006087_);
  and g_099425_(_006076_, _006087_, _006088_);
  or g_099426_(_006075_, _006086_, _006089_);
  and g_099427_(_005872_, _006089_, _006090_);
  not g_099428_(_006090_, _006091_);
  and g_099429_(_005874_, _006088_, _006092_);
  or g_099430_(_005875_, _006089_, _006094_);
  and g_099431_(_006091_, _006094_, _006095_);
  or g_099432_(_006090_, _006092_, _006096_);
  xor g_099433_(out[218], _003364_, _006097_);
  xor g_099434_(_004113_, _003364_, _006098_);
  and g_099435_(_006095_, _006097_, _006099_);
  or g_099436_(_006096_, _006098_, _006100_);
  and g_099437_(_003356_, _003369_, _006101_);
  or g_099438_(_003357_, _003368_, _006102_);
  and g_099439_(_006100_, _006102_, _006103_);
  or g_099440_(_006099_, _006101_, _006105_);
  and g_099441_(_006096_, _006098_, _006106_);
  or g_099442_(_006095_, _006097_, _006107_);
  and g_099443_(_003357_, _003368_, _006108_);
  or g_099444_(_003356_, _003369_, _006109_);
  and g_099445_(out[217], _003363_, _006110_);
  xor g_099446_(out[217], _003363_, _006111_);
  or g_099447_(_003366_, _006110_, _006112_);
  and g_099448_(_005907_, _006089_, _006113_);
  or g_099449_(_005905_, _006088_, _006114_);
  and g_099450_(_005900_, _006088_, _006116_);
  or g_099451_(_005899_, _006089_, _006117_);
  and g_099452_(_006114_, _006117_, _006118_);
  or g_099453_(_006113_, _006116_, _006119_);
  and g_099454_(_006112_, _006118_, _006120_);
  or g_099455_(_006111_, _006119_, _006121_);
  and g_099456_(_006109_, _006121_, _006122_);
  or g_099457_(_006108_, _006120_, _006123_);
  and g_099458_(_006107_, _006122_, _006124_);
  or g_099459_(_006106_, _006123_, _006125_);
  and g_099460_(_006103_, _006124_, _006127_);
  or g_099461_(_006105_, _006125_, _006128_);
  xor g_099462_(_004091_, _003362_, _006129_);
  or g_099463_(_005887_, _006089_, _006130_);
  or g_099464_(_005893_, _006088_, _006131_);
  and g_099465_(_006130_, _006131_, _006132_);
  or g_099466_(_006129_, _006132_, _006133_);
  not g_099467_(_006133_, _006134_);
  or g_099468_(_006112_, _006118_, _006135_);
  not g_099469_(_006135_, _006136_);
  and g_099470_(_006129_, _006132_, _006138_);
  not g_099471_(_006138_, _006139_);
  and g_099472_(_006135_, _006139_, _006140_);
  or g_099473_(_006136_, _006138_, _006141_);
  and g_099474_(_006133_, _006140_, _006142_);
  or g_099475_(_006134_, _006141_, _006143_);
  and g_099476_(_006127_, _006142_, _006144_);
  or g_099477_(_006128_, _006143_, _006145_);
  xor g_099478_(out[215], _003361_, _006146_);
  xor g_099479_(_004003_, _003361_, _006147_);
  and g_099480_(_005923_, _006088_, _006149_);
  or g_099481_(_005924_, _006089_, _006150_);
  and g_099482_(_005931_, _006089_, _006151_);
  or g_099483_(_005930_, _006088_, _006152_);
  and g_099484_(_006150_, _006152_, _006153_);
  or g_099485_(_006149_, _006151_, _006154_);
  or g_099486_(_006146_, _006153_, _006155_);
  xor g_099487_(out[214], _003360_, _006156_);
  xor g_099488_(_004014_, _003360_, _006157_);
  or g_099489_(_005934_, _006089_, _006158_);
  or g_099490_(_005938_, _006088_, _006160_);
  and g_099491_(_006158_, _006160_, _006161_);
  and g_099492_(_006157_, _006161_, _006162_);
  and g_099493_(_006146_, _006153_, _006163_);
  xor g_099494_(_006146_, _006153_, _006164_);
  xor g_099495_(_006147_, _006153_, _006165_);
  xor g_099496_(_006157_, _006161_, _006166_);
  xor g_099497_(_006156_, _006161_, _006167_);
  and g_099498_(_006164_, _006166_, _006168_);
  or g_099499_(_006165_, _006167_, _006169_);
  or g_099500_(_012979_, _046870_, _006171_);
  not g_099501_(_006171_, _006172_);
  or g_099502_(_003359_, _006172_, _006173_);
  or g_099503_(_005960_, _006088_, _006174_);
  or g_099504_(_005954_, _006089_, _006175_);
  and g_099505_(_006174_, _006175_, _006176_);
  and g_099506_(_006173_, _006176_, _006177_);
  not g_099507_(_006177_, _006178_);
  xor g_099508_(out[213], _003359_, _006179_);
  xor g_099509_(_004025_, _003359_, _006180_);
  and g_099510_(_005966_, _006088_, _006182_);
  or g_099511_(_005965_, _006089_, _006183_);
  and g_099512_(_005973_, _006089_, _006184_);
  or g_099513_(_005971_, _006088_, _006185_);
  and g_099514_(_006183_, _006185_, _006186_);
  or g_099515_(_006182_, _006184_, _006187_);
  and g_099516_(_006180_, _006186_, _006188_);
  or g_099517_(_006179_, _006187_, _006189_);
  and g_099518_(_006178_, _006189_, _006190_);
  or g_099519_(_006177_, _006188_, _006191_);
  or g_099520_(_006173_, _006176_, _006193_);
  and g_099521_(_006179_, _006187_, _006194_);
  or g_099522_(_006180_, _006186_, _006195_);
  and g_099523_(_006193_, _006195_, _006196_);
  not g_099524_(_006196_, _006197_);
  and g_099525_(_006190_, _006196_, _006198_);
  or g_099526_(_006191_, _006197_, _006199_);
  and g_099527_(_006168_, _006198_, _006200_);
  or g_099528_(_006169_, _006199_, _006201_);
  and g_099529_(_006144_, _006200_, _006202_);
  or g_099530_(_006145_, _006201_, _006204_);
  or g_099531_(_003937_, _006089_, _006205_);
  or g_099532_(_006022_, _006088_, _006206_);
  and g_099533_(_006205_, _006206_, _006207_);
  or g_099534_(_003948_, _006089_, _006208_);
  or g_099535_(_006031_, _006088_, _006209_);
  and g_099536_(_006208_, _006209_, _006210_);
  and g_099537_(out[208], _006210_, _006211_);
  not g_099538_(_006211_, _006212_);
  and g_099539_(out[209], _006207_, _006213_);
  xor g_099540_(out[209], _006207_, _006215_);
  xor g_099541_(_004047_, _006207_, _006216_);
  and g_099542_(_006212_, _006215_, _006217_);
  or g_099543_(_006211_, _006216_, _006218_);
  or g_099544_(_044538_, _006089_, _006219_);
  or g_099545_(_006009_, _006088_, _006220_);
  and g_099546_(_006219_, _006220_, _006221_);
  and g_099547_(_046881_, _006221_, _006222_);
  xor g_099548_(_046881_, _006221_, _006223_);
  xor g_099549_(out[211], _046870_, _006224_);
  xor g_099550_(_004080_, _046870_, _006226_);
  and g_099551_(_005985_, _006088_, _006227_);
  or g_099552_(_005986_, _006089_, _006228_);
  and g_099553_(_005992_, _006089_, _006229_);
  or g_099554_(_005991_, _006088_, _006230_);
  and g_099555_(_006228_, _006230_, _006231_);
  or g_099556_(_006227_, _006229_, _006232_);
  and g_099557_(_006224_, _006231_, _006233_);
  and g_099558_(_006226_, _006232_, _006234_);
  or g_099559_(_006224_, _006231_, _006235_);
  xor g_099560_(_006224_, _006231_, _006237_);
  or g_099561_(out[208], _006210_, _006238_);
  and g_099562_(_006237_, _006238_, _006239_);
  and g_099563_(_006223_, _006239_, _006240_);
  not g_099564_(_006240_, _006241_);
  and g_099565_(_006217_, _006240_, _006242_);
  or g_099566_(_006218_, _006241_, _006243_);
  and g_099567_(_006202_, _006242_, _006244_);
  or g_099568_(_006204_, _006243_, _006245_);
  or g_099569_(_006222_, _006233_, _006246_);
  or g_099570_(_006213_, _006217_, _006248_);
  and g_099571_(_006223_, _006248_, _006249_);
  or g_099572_(_006246_, _006249_, _006250_);
  not g_099573_(_006250_, _006251_);
  and g_099574_(_006202_, _006235_, _006252_);
  or g_099575_(_006204_, _006234_, _006253_);
  and g_099576_(_006250_, _006252_, _006254_);
  or g_099577_(_006251_, _006253_, _006255_);
  or g_099578_(_006169_, _006190_, _006256_);
  or g_099579_(_006194_, _006256_, _006257_);
  and g_099580_(_006155_, _006162_, _006259_);
  or g_099581_(_006163_, _006259_, _006260_);
  not g_099582_(_006260_, _006261_);
  and g_099583_(_006257_, _006261_, _006262_);
  or g_099584_(_006145_, _006262_, _006263_);
  not g_099585_(_006263_, _006264_);
  and g_099586_(_006127_, _006141_, _006265_);
  or g_099587_(_006128_, _006140_, _006266_);
  and g_099588_(_006105_, _006109_, _006267_);
  or g_099589_(_006103_, _006108_, _006268_);
  and g_099590_(_006266_, _006268_, _006270_);
  or g_099591_(_006265_, _006267_, _006271_);
  and g_099592_(_006263_, _006270_, _006272_);
  or g_099593_(_006264_, _006271_, _006273_);
  and g_099594_(_006255_, _006272_, _006274_);
  or g_099595_(_006254_, _006273_, _006275_);
  and g_099596_(_006245_, _006275_, _006276_);
  or g_099597_(_006244_, _006274_, _006277_);
  and g_099598_(_006096_, _006277_, _006278_);
  or g_099599_(_006095_, _006276_, _006279_);
  and g_099600_(_006097_, _006276_, _006281_);
  or g_099601_(_006098_, _006277_, _006282_);
  and g_099602_(_006279_, _006282_, _006283_);
  or g_099603_(_006278_, _006281_, _006284_);
  and g_099604_(_046881_, _006276_, _006285_);
  or g_099605_(_006221_, _006276_, _006286_);
  not g_099606_(_006286_, _006287_);
  or g_099607_(_006285_, _006287_, _006288_);
  or g_099608_(_047827_, _006288_, _006289_);
  not g_099609_(_006289_, _006290_);
  xor g_099610_(out[227], _047805_, _006292_);
  xor g_099611_(_004212_, _047805_, _006293_);
  and g_099612_(_006224_, _006276_, _006294_);
  or g_099613_(_006226_, _006277_, _006295_);
  and g_099614_(_006232_, _006277_, _006296_);
  or g_099615_(_006231_, _006276_, _006297_);
  and g_099616_(_006295_, _006297_, _006298_);
  or g_099617_(_006294_, _006296_, _006299_);
  and g_099618_(_006292_, _006298_, _006300_);
  or g_099619_(_006293_, _006299_, _006301_);
  and g_099620_(_006289_, _006301_, _006303_);
  or g_099621_(_006290_, _006300_, _006304_);
  and g_099622_(out[209], _006276_, _006305_);
  not g_099623_(_006305_, _006306_);
  or g_099624_(_006207_, _006276_, _006307_);
  not g_099625_(_006307_, _006308_);
  and g_099626_(_006306_, _006307_, _006309_);
  or g_099627_(_006305_, _006308_, _006310_);
  and g_099628_(out[225], _006309_, _006311_);
  or g_099629_(_004179_, _006310_, _006312_);
  and g_099630_(out[208], _006276_, _006314_);
  not g_099631_(_006314_, _006315_);
  or g_099632_(_006210_, _006276_, _006316_);
  not g_099633_(_006316_, _006317_);
  and g_099634_(_006315_, _006316_, _006318_);
  or g_099635_(_006314_, _006317_, _006319_);
  and g_099636_(out[224], _006318_, _006320_);
  or g_099637_(_004190_, _006319_, _006321_);
  xor g_099638_(out[225], _006309_, _006322_);
  xor g_099639_(_004179_, _006309_, _006323_);
  and g_099640_(_006321_, _006322_, _006325_);
  or g_099641_(_006320_, _006323_, _006326_);
  and g_099642_(_006312_, _006326_, _006327_);
  or g_099643_(_006311_, _006325_, _006328_);
  xor g_099644_(_047827_, _006288_, _006329_);
  xor g_099645_(_047816_, _006288_, _006330_);
  and g_099646_(_006328_, _006329_, _006331_);
  or g_099647_(_006327_, _006330_, _006332_);
  and g_099648_(_006303_, _006332_, _006333_);
  or g_099649_(_006304_, _006331_, _006334_);
  xor g_099650_(out[234], _003381_, _006336_);
  xor g_099651_(_004234_, _003381_, _006337_);
  and g_099652_(_006283_, _006336_, _006338_);
  or g_099653_(_006284_, _006337_, _006339_);
  and g_099654_(_003370_, _003385_, _006340_);
  or g_099655_(_003371_, _003384_, _006341_);
  and g_099656_(_006339_, _006341_, _006342_);
  or g_099657_(_006338_, _006340_, _006343_);
  and g_099658_(out[233], _003380_, _006344_);
  xor g_099659_(out[233], _003380_, _006345_);
  or g_099660_(_003382_, _006344_, _006347_);
  or g_099661_(_006118_, _006276_, _006348_);
  not g_099662_(_006348_, _006349_);
  and g_099663_(_006112_, _006276_, _006350_);
  not g_099664_(_006350_, _006351_);
  and g_099665_(_006348_, _006351_, _006352_);
  or g_099666_(_006349_, _006350_, _006353_);
  and g_099667_(_006347_, _006352_, _006354_);
  or g_099668_(_006345_, _006353_, _006355_);
  and g_099669_(_003371_, _003384_, _006356_);
  or g_099670_(_003370_, _003385_, _006358_);
  and g_099671_(_006284_, _006337_, _006359_);
  or g_099672_(_006283_, _006336_, _006360_);
  and g_099673_(_006358_, _006360_, _006361_);
  or g_099674_(_006356_, _006359_, _006362_);
  and g_099675_(_006355_, _006361_, _006363_);
  or g_099676_(_006354_, _006362_, _006364_);
  and g_099677_(_006342_, _006363_, _006365_);
  or g_099678_(_006343_, _006364_, _006366_);
  xor g_099679_(out[232], _003379_, _006367_);
  xor g_099680_(_004223_, _003379_, _006369_);
  and g_099681_(_006129_, _006276_, _006370_);
  not g_099682_(_006370_, _006371_);
  or g_099683_(_006132_, _006276_, _006372_);
  not g_099684_(_006372_, _006373_);
  and g_099685_(_006371_, _006372_, _006374_);
  or g_099686_(_006370_, _006373_, _006375_);
  and g_099687_(_006367_, _006375_, _006376_);
  or g_099688_(_006369_, _006374_, _006377_);
  and g_099689_(_006345_, _006353_, _006378_);
  or g_099690_(_006347_, _006352_, _006380_);
  and g_099691_(_006369_, _006374_, _006381_);
  or g_099692_(_006367_, _006375_, _006382_);
  and g_099693_(_006380_, _006382_, _006383_);
  or g_099694_(_006378_, _006381_, _006384_);
  and g_099695_(_006377_, _006383_, _006385_);
  or g_099696_(_006376_, _006384_, _006386_);
  and g_099697_(_006365_, _006385_, _006387_);
  or g_099698_(_006366_, _006386_, _006388_);
  xor g_099699_(out[231], _003378_, _006389_);
  xor g_099700_(_004135_, _003378_, _006391_);
  and g_099701_(_006154_, _006277_, _006392_);
  or g_099702_(_006153_, _006276_, _006393_);
  and g_099703_(_006146_, _006276_, _006394_);
  or g_099704_(_006147_, _006277_, _006395_);
  and g_099705_(_006393_, _006395_, _006396_);
  or g_099706_(_006392_, _006394_, _006397_);
  and g_099707_(_006389_, _006396_, _006398_);
  or g_099708_(_006391_, _006397_, _006399_);
  and g_099709_(_006391_, _006397_, _006400_);
  or g_099710_(_006389_, _006396_, _006402_);
  and g_099711_(_006399_, _006402_, _006403_);
  or g_099712_(_006398_, _006400_, _006404_);
  xor g_099713_(out[230], _003377_, _006405_);
  not g_099714_(_006405_, _006406_);
  or g_099715_(_006161_, _006276_, _006407_);
  not g_099716_(_006407_, _006408_);
  and g_099717_(_006157_, _006276_, _006409_);
  not g_099718_(_006409_, _006410_);
  and g_099719_(_006407_, _006410_, _006411_);
  or g_099720_(_006408_, _006409_, _006413_);
  and g_099721_(_006406_, _006411_, _006414_);
  or g_099722_(_006405_, _006413_, _006415_);
  xor g_099723_(_006406_, _006411_, _006416_);
  xor g_099724_(_006405_, _006411_, _006417_);
  and g_099725_(_006403_, _006416_, _006418_);
  or g_099726_(_006404_, _006417_, _006419_);
  or g_099727_(_013133_, _047805_, _006420_);
  not g_099728_(_006420_, _006421_);
  and g_099729_(_003375_, _006420_, _006422_);
  or g_099730_(_003374_, _006421_, _006424_);
  or g_099731_(_006176_, _006276_, _006425_);
  not g_099732_(_006425_, _006426_);
  and g_099733_(_006173_, _006276_, _006427_);
  not g_099734_(_006427_, _006428_);
  and g_099735_(_006425_, _006428_, _006429_);
  or g_099736_(_006426_, _006427_, _006430_);
  and g_099737_(_006424_, _006429_, _006431_);
  or g_099738_(_006422_, _006430_, _006432_);
  xor g_099739_(out[229], _003374_, _006433_);
  xor g_099740_(_004157_, _003374_, _006435_);
  and g_099741_(_006180_, _006276_, _006436_);
  or g_099742_(_006179_, _006277_, _006437_);
  and g_099743_(_006187_, _006277_, _006438_);
  or g_099744_(_006186_, _006276_, _006439_);
  and g_099745_(_006437_, _006439_, _006440_);
  or g_099746_(_006436_, _006438_, _006441_);
  and g_099747_(_006435_, _006440_, _006442_);
  or g_099748_(_006433_, _006441_, _006443_);
  and g_099749_(_006432_, _006443_, _006444_);
  or g_099750_(_006431_, _006442_, _006446_);
  and g_099751_(_006422_, _006430_, _006447_);
  or g_099752_(_006424_, _006429_, _006448_);
  and g_099753_(_006433_, _006441_, _006449_);
  or g_099754_(_006435_, _006440_, _006450_);
  and g_099755_(_006293_, _006299_, _006451_);
  or g_099756_(_006292_, _006298_, _006452_);
  and g_099757_(_006450_, _006452_, _006453_);
  or g_099758_(_006449_, _006451_, _006454_);
  and g_099759_(_006448_, _006453_, _006455_);
  or g_099760_(_006447_, _006454_, _006457_);
  and g_099761_(_006444_, _006455_, _006458_);
  or g_099762_(_006446_, _006457_, _006459_);
  and g_099763_(_006418_, _006458_, _006460_);
  or g_099764_(_006419_, _006459_, _006461_);
  and g_099765_(_006387_, _006460_, _006462_);
  or g_099766_(_006388_, _006461_, _006463_);
  and g_099767_(_006334_, _006462_, _006464_);
  or g_099768_(_006333_, _006463_, _006465_);
  and g_099769_(_006418_, _006446_, _006466_);
  or g_099770_(_006419_, _006444_, _006468_);
  and g_099771_(_006450_, _006466_, _006469_);
  or g_099772_(_006449_, _006468_, _006470_);
  and g_099773_(_006402_, _006414_, _006471_);
  or g_099774_(_006400_, _006415_, _006472_);
  and g_099775_(_006399_, _006472_, _006473_);
  or g_099776_(_006398_, _006471_, _006474_);
  and g_099777_(_006470_, _006473_, _006475_);
  or g_099778_(_006469_, _006474_, _006476_);
  and g_099779_(_006387_, _006476_, _006477_);
  or g_099780_(_006388_, _006475_, _006479_);
  and g_099781_(_006343_, _006358_, _006480_);
  or g_099782_(_006342_, _006356_, _006481_);
  and g_099783_(_006365_, _006384_, _006482_);
  or g_099784_(_006366_, _006383_, _006483_);
  and g_099785_(_006481_, _006483_, _006484_);
  or g_099786_(_006480_, _006482_, _006485_);
  and g_099787_(_006479_, _006484_, _006486_);
  or g_099788_(_006477_, _006485_, _006487_);
  and g_099789_(_006465_, _006486_, _006488_);
  or g_099790_(_006464_, _006487_, _006490_);
  and g_099791_(_004190_, _006319_, _006491_);
  or g_099792_(out[224], _006318_, _006492_);
  and g_099793_(_006301_, _006492_, _006493_);
  or g_099794_(_006300_, _006491_, _006494_);
  and g_099795_(_006329_, _006493_, _006495_);
  or g_099796_(_006330_, _006494_, _006496_);
  and g_099797_(_006325_, _006495_, _006497_);
  or g_099798_(_006326_, _006496_, _006498_);
  and g_099799_(_006462_, _006497_, _006499_);
  or g_099800_(_006463_, _006498_, _006501_);
  and g_099801_(_006490_, _006501_, _006502_);
  or g_099802_(_006488_, _006499_, _006503_);
  and g_099803_(_006284_, _006503_, _006504_);
  not g_099804_(_006504_, _006505_);
  or g_099805_(_006337_, _006503_, _006506_);
  not g_099806_(_006506_, _006507_);
  and g_099807_(_006505_, _006506_, _006508_);
  or g_099808_(_006504_, _006507_, _006509_);
  and g_099809_(_003562_, _006508_, _006510_);
  or g_099810_(_003564_, _006509_, _006512_);
  and g_099811_(_003386_, _003400_, _006513_);
  or g_099812_(_003388_, _003399_, _006514_);
  and g_099813_(_006512_, _006514_, _006515_);
  or g_099814_(_006510_, _006513_, _006516_);
  and g_099815_(_003564_, _006509_, _006517_);
  or g_099816_(_003562_, _006508_, _006518_);
  and g_099817_(out[249], _003394_, _006519_);
  xor g_099818_(out[249], _003394_, _006520_);
  or g_099819_(_003396_, _006519_, _006521_);
  and g_099820_(_006353_, _006503_, _006523_);
  and g_099821_(_006347_, _006502_, _006524_);
  or g_099822_(_006523_, _006524_, _006525_);
  not g_099823_(_006525_, _006526_);
  and g_099824_(_006521_, _006526_, _006527_);
  or g_099825_(_006520_, _006525_, _006528_);
  xor g_099826_(out[248], _003393_, _006529_);
  xor g_099827_(_004333_, _003393_, _006530_);
  and g_099828_(_006369_, _006502_, _006531_);
  and g_099829_(_006375_, _006503_, _006532_);
  or g_099830_(_006531_, _006532_, _006534_);
  or g_099831_(_006529_, _006534_, _006535_);
  not g_099832_(_006535_, _006536_);
  and g_099833_(_006520_, _006525_, _006537_);
  or g_099834_(_006521_, _006526_, _006538_);
  and g_099835_(_006528_, _006538_, _006539_);
  or g_099836_(_006527_, _006537_, _006540_);
  xor g_099837_(_006529_, _006534_, _006541_);
  xor g_099838_(_006530_, _006534_, _006542_);
  and g_099839_(_006539_, _006541_, _006543_);
  or g_099840_(_006540_, _006542_, _006545_);
  xor g_099841_(out[247], _003392_, _006546_);
  xor g_099842_(_004256_, _003392_, _006547_);
  and g_099843_(_006389_, _006502_, _006548_);
  and g_099844_(_006397_, _006503_, _006549_);
  or g_099845_(_006548_, _006549_, _006550_);
  not g_099846_(_006550_, _006551_);
  and g_099847_(_006547_, _006550_, _006552_);
  xor g_099848_(out[246], _003391_, _006553_);
  xor g_099849_(_004267_, _003391_, _006554_);
  and g_099850_(_006406_, _006502_, _006556_);
  and g_099851_(_006413_, _006503_, _006557_);
  or g_099852_(_006556_, _006557_, _006558_);
  not g_099853_(_006558_, _006559_);
  and g_099854_(_006554_, _006559_, _006560_);
  or g_099855_(_006553_, _006558_, _006561_);
  and g_099856_(_006546_, _006551_, _006562_);
  or g_099857_(_006547_, _006550_, _006563_);
  and g_099858_(_006561_, _006563_, _006564_);
  or g_099859_(_006560_, _006562_, _006565_);
  or g_099860_(_006552_, _006564_, _006567_);
  not g_099861_(_006567_, _006568_);
  xor g_099862_(out[245], _003390_, _006569_);
  xor g_099863_(_004278_, _003390_, _006570_);
  and g_099864_(_006435_, _006502_, _006571_);
  and g_099865_(_006441_, _006503_, _006572_);
  or g_099866_(_006571_, _006572_, _006573_);
  and g_099867_(_006569_, _006573_, _006574_);
  and g_099868_(_006553_, _006558_, _006575_);
  or g_099869_(_006552_, _006575_, _006576_);
  or g_099870_(_006574_, _006576_, _006578_);
  not g_099871_(_006578_, _006579_);
  and g_099872_(_006564_, _006579_, _006580_);
  or g_099873_(_006565_, _006578_, _006581_);
  or g_099874_(_006569_, _006573_, _006582_);
  xor g_099875_(out[244], _003389_, _006583_);
  xor g_099876_(_004289_, _003389_, _006584_);
  and g_099877_(_006430_, _006503_, _006585_);
  and g_099878_(_006424_, _006502_, _006586_);
  or g_099879_(_006585_, _006586_, _006587_);
  not g_099880_(_006587_, _006589_);
  or g_099881_(_006583_, _006587_, _006590_);
  and g_099882_(_006582_, _006590_, _006591_);
  not g_099883_(_006591_, _006592_);
  and g_099884_(_006288_, _006503_, _006593_);
  and g_099885_(_047816_, _006502_, _006594_);
  or g_099886_(_006593_, _006594_, _006595_);
  not g_099887_(_006595_, _006596_);
  and g_099888_(_050478_, _006596_, _006597_);
  or g_099889_(_050489_, _006595_, _006598_);
  xor g_099890_(out[243], _050467_, _006600_);
  xor g_099891_(_004322_, _050467_, _006601_);
  and g_099892_(_006292_, _006502_, _006602_);
  and g_099893_(_006299_, _006503_, _006603_);
  or g_099894_(_006602_, _006603_, _006604_);
  not g_099895_(_006604_, _006605_);
  and g_099896_(_006600_, _006605_, _006606_);
  or g_099897_(_006601_, _006604_, _006607_);
  and g_099898_(_006598_, _006607_, _006608_);
  not g_099899_(_006608_, _006609_);
  and g_099900_(_050489_, _006595_, _006611_);
  or g_099901_(_050478_, _006596_, _006612_);
  and g_099902_(out[225], _006502_, _006613_);
  or g_099903_(_004179_, _006503_, _006614_);
  and g_099904_(_006310_, _006503_, _006615_);
  or g_099905_(_006309_, _006502_, _006616_);
  and g_099906_(_006614_, _006616_, _006617_);
  or g_099907_(_006613_, _006615_, _006618_);
  and g_099908_(out[241], _006617_, _006619_);
  or g_099909_(_053038_, _006618_, _006620_);
  and g_099910_(out[224], _006502_, _006622_);
  or g_099911_(_004190_, _006503_, _006623_);
  and g_099912_(_006319_, _006503_, _006624_);
  or g_099913_(_006318_, _006502_, _006625_);
  and g_099914_(_006623_, _006625_, _006626_);
  or g_099915_(_006622_, _006624_, _006627_);
  and g_099916_(out[240], _006626_, _006628_);
  or g_099917_(_004300_, _006627_, _006629_);
  xor g_099918_(out[241], _006617_, _006630_);
  xor g_099919_(_053038_, _006617_, _006631_);
  and g_099920_(_006629_, _006630_, _006633_);
  or g_099921_(_006628_, _006631_, _006634_);
  and g_099922_(_006620_, _006634_, _006635_);
  or g_099923_(_006619_, _006633_, _006636_);
  and g_099924_(_006612_, _006636_, _006637_);
  or g_099925_(_006611_, _006635_, _006638_);
  and g_099926_(_006608_, _006638_, _006639_);
  or g_099927_(_006609_, _006637_, _006640_);
  and g_099928_(_006583_, _006587_, _006641_);
  or g_099929_(_006584_, _006589_, _006642_);
  and g_099930_(_006601_, _006604_, _006644_);
  or g_099931_(_006600_, _006605_, _006645_);
  or g_099932_(_006641_, _006644_, _006646_);
  not g_099933_(_006646_, _006647_);
  and g_099934_(_006640_, _006647_, _006648_);
  or g_099935_(_006639_, _006646_, _006649_);
  and g_099936_(_006591_, _006649_, _006650_);
  or g_099937_(_006592_, _006648_, _006651_);
  and g_099938_(_006580_, _006651_, _006652_);
  or g_099939_(_006581_, _006650_, _006653_);
  and g_099940_(_006567_, _006653_, _006655_);
  or g_099941_(_006568_, _006652_, _006656_);
  and g_099942_(_006543_, _006656_, _006657_);
  or g_099943_(_006545_, _006655_, _006658_);
  and g_099944_(_006528_, _006536_, _006659_);
  or g_099945_(_006527_, _006535_, _006660_);
  and g_099946_(_006538_, _006660_, _006661_);
  or g_099947_(_006537_, _006659_, _006662_);
  and g_099948_(_006658_, _006661_, _006663_);
  or g_099949_(_006657_, _006662_, _006664_);
  and g_099950_(_006518_, _006664_, _006666_);
  or g_099951_(_006517_, _006663_, _006667_);
  and g_099952_(_006515_, _006667_, _006668_);
  or g_099953_(_006516_, _006666_, _006669_);
  and g_099954_(_003388_, _003399_, _006670_);
  or g_099955_(_003386_, _003400_, _006671_);
  and g_099956_(_006598_, _006645_, _006672_);
  or g_099957_(_006597_, _006644_, _006673_);
  and g_099958_(_004300_, _006627_, _006674_);
  or g_099959_(out[240], _006626_, _006675_);
  and g_099960_(_006642_, _006675_, _006677_);
  or g_099961_(_006641_, _006674_, _006678_);
  and g_099962_(_006672_, _006677_, _006679_);
  or g_099963_(_006673_, _006678_, _006680_);
  and g_099964_(_006543_, _006679_, _006681_);
  or g_099965_(_006545_, _006680_, _006682_);
  and g_099966_(_006633_, _006681_, _006683_);
  or g_099967_(_006634_, _006682_, _006684_);
  and g_099968_(_006518_, _006671_, _006685_);
  or g_099969_(_006517_, _006670_, _006686_);
  and g_099970_(_006607_, _006612_, _006688_);
  or g_099971_(_006606_, _006611_, _006689_);
  and g_099972_(_006685_, _006688_, _006690_);
  or g_099973_(_006686_, _006689_, _006691_);
  and g_099974_(_006515_, _006591_, _006692_);
  or g_099975_(_006516_, _006592_, _006693_);
  and g_099976_(_006690_, _006692_, _006694_);
  or g_099977_(_006691_, _006693_, _006695_);
  and g_099978_(_006580_, _006694_, _006696_);
  or g_099979_(_006581_, _006695_, _006697_);
  and g_099980_(_006683_, _006696_, _006699_);
  or g_099981_(_006684_, _006697_, _006700_);
  and g_099982_(_006671_, _006700_, _006701_);
  or g_099983_(_006670_, _006699_, _006702_);
  and g_099984_(_006669_, _006701_, _006703_);
  or g_099985_(_006668_, _006702_, _006704_);
  and g_099986_(_003562_, _006703_, _006705_);
  or g_099987_(_003564_, _006704_, _006706_);
  and g_099988_(_006509_, _006704_, _006707_);
  or g_099989_(_006508_, _006703_, _006708_);
  and g_099990_(_006706_, _006708_, _006710_);
  or g_099991_(_006705_, _006707_, _006711_);
  and g_099992_(_006595_, _006704_, _006712_);
  and g_099993_(_050478_, _006703_, _006713_);
  or g_099994_(_006712_, _006713_, _006714_);
  or g_099995_(_051427_, _006714_, _006715_);
  xor g_099996_(out[259], _051425_, _006716_);
  xor g_099997_(_053005_, _051425_, _006717_);
  and g_099998_(_006604_, _006704_, _006718_);
  and g_099999_(_006600_, _006703_, _006719_);
  or g_100000_(_006718_, _006719_, _006721_);
  or g_100001_(_006717_, _006721_, _006722_);
  and g_100002_(_006715_, _006722_, _006723_);
  and g_100003_(_051427_, _006714_, _006724_);
  and g_100004_(_006717_, _006721_, _006725_);
  or g_100005_(_006724_, _006725_, _006726_);
  not g_100006_(_006726_, _006727_);
  and g_100007_(_006723_, _006727_, _006728_);
  or g_100008_(_053038_, _006704_, _006729_);
  or g_100009_(_006617_, _006703_, _006730_);
  and g_100010_(_006729_, _006730_, _006732_);
  and g_100011_(out[257], _006732_, _006733_);
  and g_100012_(_006626_, _006704_, _006734_);
  or g_100013_(_006627_, _006703_, _006735_);
  or g_100014_(out[240], _006704_, _006736_);
  not g_100015_(_006736_, _006737_);
  or g_100016_(_006734_, _006737_, _006738_);
  and g_100017_(_006735_, _006736_, _006739_);
  and g_100018_(out[256], _006738_, _006740_);
  not g_100019_(_006740_, _006741_);
  xor g_100020_(out[257], _006732_, _006743_);
  xor g_100021_(_053027_, _006732_, _006744_);
  and g_100022_(_006741_, _006743_, _006745_);
  or g_100023_(_006740_, _006744_, _006746_);
  or g_100024_(_006733_, _006745_, _006747_);
  and g_100025_(_006728_, _006747_, _006748_);
  or g_100026_(_006723_, _006725_, _006749_);
  not g_100027_(_006749_, _006750_);
  or g_100028_(_006748_, _006750_, _006751_);
  xor g_100029_(out[266], _003410_, _006752_);
  xor g_100030_(_004421_, _003410_, _006754_);
  and g_100031_(_006710_, _006752_, _006755_);
  or g_100032_(_006711_, _006754_, _006756_);
  and g_100033_(_003401_, _003414_, _006757_);
  or g_100034_(_003402_, _003413_, _006758_);
  and g_100035_(_006756_, _006758_, _006759_);
  or g_100036_(_006755_, _006757_, _006760_);
  and g_100037_(_003402_, _003413_, _006761_);
  or g_100038_(_003401_, _003414_, _006762_);
  and g_100039_(_006711_, _006754_, _006763_);
  or g_100040_(_006710_, _006752_, _006765_);
  and g_100041_(_006762_, _006765_, _006766_);
  or g_100042_(_006761_, _006763_, _006767_);
  and g_100043_(_006759_, _006766_, _006768_);
  or g_100044_(_006760_, _006767_, _006769_);
  xor g_100045_(out[264], _003407_, _006770_);
  xor g_100046_(_004399_, _003407_, _006771_);
  or g_100047_(_006529_, _006704_, _006772_);
  not g_100048_(_006772_, _006773_);
  and g_100049_(_006534_, _006704_, _006774_);
  not g_100050_(_006774_, _006776_);
  and g_100051_(_006772_, _006776_, _006777_);
  or g_100052_(_006773_, _006774_, _006778_);
  and g_100053_(_006770_, _006778_, _006779_);
  and g_100054_(out[265], _003408_, _006780_);
  xor g_100055_(out[265], _003408_, _006781_);
  or g_100056_(_003411_, _006780_, _006782_);
  and g_100057_(_006525_, _006704_, _006783_);
  not g_100058_(_006783_, _006784_);
  or g_100059_(_006520_, _006704_, _006785_);
  not g_100060_(_006785_, _006787_);
  and g_100061_(_006784_, _006785_, _006788_);
  or g_100062_(_006783_, _006787_, _006789_);
  and g_100063_(_006782_, _006788_, _006790_);
  or g_100064_(_006781_, _006789_, _006791_);
  or g_100065_(_006779_, _006790_, _006792_);
  and g_100066_(_006771_, _006777_, _006793_);
  and g_100067_(_006781_, _006789_, _006794_);
  or g_100068_(_006793_, _006794_, _006795_);
  or g_100069_(_006792_, _006795_, _006796_);
  xor g_100070_(_006771_, _006777_, _006798_);
  xor g_100071_(_006782_, _006788_, _006799_);
  and g_100072_(_006768_, _006799_, _006800_);
  and g_100073_(_006798_, _006800_, _006801_);
  or g_100074_(_006769_, _006796_, _006802_);
  xor g_100075_(out[262], _003405_, _006803_);
  not g_100076_(_006803_, _006804_);
  and g_100077_(_006554_, _006703_, _006805_);
  and g_100078_(_006558_, _006704_, _006806_);
  or g_100079_(_006805_, _006806_, _006807_);
  or g_100080_(_006803_, _006807_, _006809_);
  xor g_100081_(_006803_, _006807_, _006810_);
  xor g_100082_(_006804_, _006807_, _006811_);
  xor g_100083_(out[263], _003406_, _006812_);
  xor g_100084_(_004377_, _003406_, _006813_);
  and g_100085_(_006546_, _006703_, _006814_);
  and g_100086_(_006550_, _006704_, _006815_);
  or g_100087_(_006814_, _006815_, _006816_);
  or g_100088_(_006813_, _006816_, _006817_);
  and g_100089_(_006813_, _006816_, _006818_);
  xor g_100090_(_006813_, _006816_, _006820_);
  xor g_100091_(_006812_, _006816_, _006821_);
  and g_100092_(_006810_, _006820_, _006822_);
  or g_100093_(_006811_, _006821_, _006823_);
  xor g_100094_(out[260], _003403_, _006824_);
  xor g_100095_(_052994_, _003403_, _006825_);
  and g_100096_(_006587_, _006704_, _006826_);
  and g_100097_(_006584_, _006703_, _006827_);
  or g_100098_(_006826_, _006827_, _006828_);
  or g_100099_(_006824_, _006828_, _006829_);
  not g_100100_(_006829_, _006831_);
  xor g_100101_(out[261], _003404_, _006832_);
  xor g_100102_(_052972_, _003404_, _006833_);
  and g_100103_(_006573_, _006704_, _006834_);
  and g_100104_(_006570_, _006703_, _006835_);
  or g_100105_(_006834_, _006835_, _006836_);
  or g_100106_(_006832_, _006836_, _006837_);
  not g_100107_(_006837_, _006838_);
  and g_100108_(_006829_, _006837_, _006839_);
  or g_100109_(_006831_, _006838_, _006840_);
  and g_100110_(_006832_, _006836_, _006842_);
  and g_100111_(_006824_, _006828_, _006843_);
  or g_100112_(_006842_, _006843_, _006844_);
  not g_100113_(_006844_, _006845_);
  and g_100114_(_006839_, _006845_, _006846_);
  or g_100115_(_006840_, _006844_, _006847_);
  and g_100116_(_006822_, _006846_, _006848_);
  or g_100117_(_006823_, _006847_, _006849_);
  and g_100118_(_006801_, _006848_, _006850_);
  or g_100119_(_006802_, _006849_, _006851_);
  and g_100120_(_006751_, _006850_, _006853_);
  or g_100121_(_006823_, _006839_, _006854_);
  or g_100122_(_006842_, _006854_, _006855_);
  or g_100123_(_006809_, _006818_, _006856_);
  and g_100124_(_006817_, _006856_, _006857_);
  and g_100125_(_006855_, _006857_, _006858_);
  or g_100126_(_006802_, _006858_, _006859_);
  not g_100127_(_006859_, _006860_);
  and g_100128_(_006760_, _006762_, _006861_);
  and g_100129_(_006768_, _006795_, _006862_);
  and g_100130_(_006791_, _006862_, _006864_);
  not g_100131_(_006864_, _006865_);
  and g_100132_(_006859_, _006865_, _006866_);
  or g_100133_(_006860_, _006864_, _006867_);
  or g_100134_(_006853_, _006861_, _006868_);
  not g_100135_(_006868_, _006869_);
  and g_100136_(_006866_, _006869_, _006870_);
  or g_100137_(_006867_, _006868_, _006871_);
  or g_100138_(out[256], _006738_, _006872_);
  and g_100139_(_006728_, _006872_, _006873_);
  not g_100140_(_006873_, _006875_);
  and g_100141_(_006745_, _006873_, _006876_);
  or g_100142_(_006746_, _006875_, _006877_);
  and g_100143_(_006850_, _006876_, _006878_);
  or g_100144_(_006851_, _006877_, _006879_);
  and g_100145_(_006871_, _006879_, _006880_);
  or g_100146_(_006870_, _006878_, _006881_);
  and g_100147_(_006711_, _006881_, _006882_);
  or g_100148_(_006710_, _006880_, _006883_);
  and g_100149_(_006752_, _006880_, _006884_);
  or g_100150_(_006754_, _006881_, _006886_);
  and g_100151_(_006883_, _006886_, _006887_);
  or g_100152_(_006882_, _006884_, _006888_);
  and g_100153_(_003415_, _003430_, _006889_);
  or g_100154_(_003416_, _003429_, _006890_);
  xor g_100155_(out[282], _003426_, _006891_);
  xor g_100156_(_004454_, _003426_, _006892_);
  and g_100157_(_006887_, _006891_, _006893_);
  or g_100158_(_006888_, _006892_, _006894_);
  and g_100159_(_006890_, _006894_, _006895_);
  or g_100160_(_006889_, _006893_, _006897_);
  and g_100161_(_003416_, _003429_, _006898_);
  or g_100162_(_003415_, _003430_, _006899_);
  and g_100163_(_006888_, _006892_, _006900_);
  or g_100164_(_006887_, _006891_, _006901_);
  and g_100165_(_006899_, _006901_, _006902_);
  or g_100166_(_006898_, _006900_, _006903_);
  and g_100167_(out[281], _003425_, _006904_);
  xor g_100168_(out[281], _003425_, _006905_);
  or g_100169_(_003427_, _006904_, _006906_);
  and g_100170_(_006789_, _006881_, _006908_);
  not g_100171_(_006908_, _006909_);
  or g_100172_(_006781_, _006881_, _006910_);
  not g_100173_(_006910_, _006911_);
  and g_100174_(_006909_, _006910_, _006912_);
  or g_100175_(_006908_, _006911_, _006913_);
  and g_100176_(_006906_, _006912_, _006914_);
  or g_100177_(_006905_, _006913_, _006915_);
  and g_100178_(_006902_, _006915_, _006916_);
  or g_100179_(_006903_, _006914_, _006917_);
  and g_100180_(_006895_, _006916_, _006919_);
  or g_100181_(_006897_, _006917_, _006920_);
  xor g_100182_(out[280], _003424_, _006921_);
  xor g_100183_(_053060_, _003424_, _006922_);
  or g_100184_(_006770_, _006881_, _006923_);
  not g_100185_(_006923_, _006924_);
  and g_100186_(_006778_, _006881_, _006925_);
  not g_100187_(_006925_, _006926_);
  and g_100188_(_006923_, _006926_, _006927_);
  or g_100189_(_006924_, _006925_, _006928_);
  and g_100190_(_006921_, _006928_, _006930_);
  not g_100191_(_006930_, _006931_);
  and g_100192_(_006905_, _006913_, _006932_);
  or g_100193_(_006906_, _006912_, _006933_);
  and g_100194_(_006922_, _006927_, _006934_);
  or g_100195_(_006921_, _006928_, _006935_);
  and g_100196_(_006933_, _006935_, _006936_);
  or g_100197_(_006932_, _006934_, _006937_);
  and g_100198_(_006931_, _006936_, _006938_);
  or g_100199_(_006930_, _006937_, _006939_);
  and g_100200_(_006919_, _006938_, _006941_);
  or g_100201_(_006920_, _006939_, _006942_);
  xor g_100202_(out[279], _003423_, _006943_);
  xor g_100203_(_053049_, _003423_, _006944_);
  and g_100204_(_006816_, _006881_, _006945_);
  and g_100205_(_006812_, _006880_, _006946_);
  or g_100206_(_006945_, _006946_, _006947_);
  or g_100207_(_006944_, _006947_, _006948_);
  xor g_100208_(out[278], _003422_, _006949_);
  not g_100209_(_006949_, _006950_);
  and g_100210_(_006807_, _006881_, _006952_);
  and g_100211_(_006804_, _006880_, _006953_);
  or g_100212_(_006952_, _006953_, _006954_);
  not g_100213_(_006954_, _006955_);
  or g_100214_(_006949_, _006954_, _006956_);
  and g_100215_(_006944_, _006947_, _006957_);
  xor g_100216_(_006944_, _006947_, _006958_);
  xor g_100217_(_006943_, _006947_, _006959_);
  xor g_100218_(_006949_, _006954_, _006960_);
  xor g_100219_(_006950_, _006954_, _006961_);
  and g_100220_(_006958_, _006960_, _006963_);
  or g_100221_(_006959_, _006961_, _006964_);
  or g_100222_(_013584_, _051640_, _006965_);
  not g_100223_(_006965_, _006966_);
  and g_100224_(_003421_, _006965_, _006967_);
  or g_100225_(_003419_, _006966_, _006968_);
  or g_100226_(_006824_, _006881_, _006969_);
  not g_100227_(_006969_, _006970_);
  and g_100228_(_006828_, _006881_, _006971_);
  not g_100229_(_006971_, _006972_);
  and g_100230_(_006969_, _006972_, _006974_);
  or g_100231_(_006970_, _006971_, _006975_);
  and g_100232_(_006968_, _006974_, _006976_);
  xor g_100233_(out[277], _003419_, _006977_);
  xor g_100234_(_053071_, _003419_, _006978_);
  or g_100235_(_006832_, _006881_, _006979_);
  not g_100236_(_006979_, _006980_);
  and g_100237_(_006836_, _006881_, _006981_);
  not g_100238_(_006981_, _006982_);
  and g_100239_(_006979_, _006982_, _006983_);
  or g_100240_(_006980_, _006981_, _006985_);
  and g_100241_(_006978_, _006983_, _006986_);
  or g_100242_(_006976_, _006986_, _006987_);
  and g_100243_(_006977_, _006985_, _006988_);
  or g_100244_(_006978_, _006983_, _006989_);
  and g_100245_(_006967_, _006975_, _006990_);
  or g_100246_(_006988_, _006990_, _006991_);
  or g_100247_(_006987_, _006991_, _006992_);
  or g_100248_(_006964_, _006992_, _006993_);
  or g_100249_(_006942_, _006993_, _006994_);
  xor g_100250_(out[275], _051640_, _006996_);
  xor g_100251_(_053093_, _051640_, _006997_);
  and g_100252_(_006716_, _006880_, _006998_);
  and g_100253_(_006721_, _006881_, _006999_);
  or g_100254_(_006998_, _006999_, _007000_);
  or g_100255_(_006997_, _007000_, _007001_);
  and g_100256_(_006714_, _006881_, _007002_);
  and g_100257_(_051426_, _006880_, _007003_);
  or g_100258_(_007002_, _007003_, _007004_);
  or g_100259_(_051642_, _007004_, _007005_);
  and g_100260_(_007001_, _007005_, _007007_);
  and g_100261_(_006997_, _007000_, _007008_);
  xor g_100262_(_006996_, _007000_, _007009_);
  xor g_100263_(_051641_, _007004_, _007010_);
  or g_100264_(_007009_, _007010_, _007011_);
  or g_100265_(_053027_, _006881_, _007012_);
  or g_100266_(_006732_, _006880_, _007013_);
  and g_100267_(_007012_, _007013_, _007014_);
  and g_100268_(out[273], _007014_, _007015_);
  not g_100269_(_007015_, _007016_);
  and g_100270_(out[256], _006880_, _007018_);
  or g_100271_(_004388_, _006881_, _007019_);
  and g_100272_(_006739_, _006881_, _007020_);
  or g_100273_(_006738_, _006880_, _007021_);
  and g_100274_(_007019_, _007021_, _007022_);
  or g_100275_(_007018_, _007020_, _007023_);
  and g_100276_(out[272], _007022_, _007024_);
  xor g_100277_(_053126_, _007014_, _007025_);
  or g_100278_(_007024_, _007025_, _007026_);
  and g_100279_(_007016_, _007026_, _007027_);
  or g_100280_(_007011_, _007027_, _007029_);
  or g_100281_(_007007_, _007008_, _007030_);
  and g_100282_(_007029_, _007030_, _007031_);
  or g_100283_(_006994_, _007031_, _007032_);
  and g_100284_(_006963_, _006987_, _007033_);
  and g_100285_(_006989_, _007033_, _007034_);
  or g_100286_(_006956_, _006957_, _007035_);
  and g_100287_(_006948_, _007035_, _007036_);
  not g_100288_(_007036_, _007037_);
  or g_100289_(_007034_, _007037_, _007038_);
  and g_100290_(_006941_, _007038_, _007040_);
  and g_100291_(_006919_, _006937_, _007041_);
  not g_100292_(_007041_, _007042_);
  and g_100293_(_006897_, _006899_, _007043_);
  or g_100294_(_007040_, _007043_, _007044_);
  not g_100295_(_007044_, _007045_);
  and g_100296_(_007032_, _007042_, _007046_);
  not g_100297_(_007046_, _007047_);
  and g_100298_(_007045_, _007046_, _007048_);
  or g_100299_(_007044_, _007047_, _007049_);
  and g_100300_(_004443_, _007023_, _007051_);
  or g_100301_(out[272], _007022_, _007052_);
  or g_100302_(_007011_, _007026_, _007053_);
  or g_100303_(_006994_, _007053_, _007054_);
  not g_100304_(_007054_, _007055_);
  and g_100305_(_007052_, _007055_, _007056_);
  or g_100306_(_007051_, _007054_, _007057_);
  and g_100307_(_007049_, _007057_, _007058_);
  or g_100308_(_007048_, _007056_, _007059_);
  and g_100309_(_006888_, _007059_, _007060_);
  or g_100310_(_006887_, _007058_, _007062_);
  or g_100311_(_006892_, _007059_, _007063_);
  not g_100312_(_007063_, _007064_);
  and g_100313_(_007062_, _007063_, _007065_);
  or g_100314_(_007060_, _007064_, _007066_);
  xor g_100315_(out[298], _003443_, _007067_);
  not g_100316_(_007067_, _007068_);
  or g_100317_(_007066_, _007068_, _007069_);
  not g_100318_(_007069_, _007070_);
  and g_100319_(_003432_, _003446_, _007071_);
  or g_100320_(_003433_, _003445_, _007073_);
  and g_100321_(_007069_, _007073_, _007074_);
  or g_100322_(_007070_, _007071_, _007075_);
  and g_100323_(_003433_, _003445_, _007076_);
  or g_100324_(_003432_, _003446_, _007077_);
  and g_100325_(_007066_, _007068_, _007078_);
  or g_100326_(_007065_, _007067_, _007079_);
  and g_100327_(_007077_, _007079_, _007080_);
  or g_100328_(_007076_, _007078_, _007081_);
  and g_100329_(out[297], _003441_, _007082_);
  xor g_100330_(out[297], _003441_, _007084_);
  xor g_100331_(_053236_, _003441_, _007085_);
  and g_100332_(_006913_, _007059_, _007086_);
  not g_100333_(_007086_, _007087_);
  or g_100334_(_006905_, _007059_, _007088_);
  not g_100335_(_007088_, _007089_);
  and g_100336_(_007087_, _007088_, _007090_);
  or g_100337_(_007086_, _007089_, _007091_);
  and g_100338_(_007085_, _007090_, _007092_);
  or g_100339_(_007084_, _007091_, _007093_);
  and g_100340_(_007080_, _007093_, _007095_);
  or g_100341_(_007081_, _007092_, _007096_);
  and g_100342_(_007074_, _007095_, _007097_);
  or g_100343_(_007075_, _007096_, _007098_);
  xor g_100344_(out[296], _003440_, _007099_);
  xor g_100345_(_053159_, _003440_, _007100_);
  and g_100346_(_006928_, _007059_, _007101_);
  not g_100347_(_007101_, _007102_);
  or g_100348_(_006921_, _007059_, _007103_);
  not g_100349_(_007103_, _007104_);
  and g_100350_(_007102_, _007103_, _007106_);
  or g_100351_(_007101_, _007104_, _007107_);
  or g_100352_(_007100_, _007106_, _007108_);
  not g_100353_(_007108_, _007109_);
  or g_100354_(_007085_, _007090_, _007110_);
  not g_100355_(_007110_, _007111_);
  and g_100356_(_007100_, _007106_, _007112_);
  or g_100357_(_007099_, _007107_, _007113_);
  and g_100358_(_007110_, _007113_, _007114_);
  or g_100359_(_007111_, _007112_, _007115_);
  and g_100360_(_007108_, _007114_, _007117_);
  or g_100361_(_007109_, _007115_, _007118_);
  and g_100362_(_007097_, _007117_, _007119_);
  or g_100363_(_007098_, _007118_, _007120_);
  xor g_100364_(out[295], _003439_, _007121_);
  xor g_100365_(_053148_, _003439_, _007122_);
  or g_100366_(_006944_, _007059_, _007123_);
  and g_100367_(_006947_, _007059_, _007124_);
  not g_100368_(_007124_, _007125_);
  and g_100369_(_007123_, _007125_, _007126_);
  or g_100370_(_007121_, _007126_, _007128_);
  xor g_100371_(out[294], _003438_, _007129_);
  not g_100372_(_007129_, _007130_);
  or g_100373_(_006949_, _007059_, _007131_);
  or g_100374_(_006955_, _007058_, _007132_);
  and g_100375_(_007131_, _007132_, _007133_);
  and g_100376_(_007130_, _007133_, _007134_);
  and g_100377_(_007121_, _007126_, _007135_);
  xor g_100378_(_007121_, _007126_, _007136_);
  xor g_100379_(_007122_, _007126_, _007137_);
  xor g_100380_(_007130_, _007133_, _007139_);
  xor g_100381_(_007129_, _007133_, _007140_);
  and g_100382_(_007136_, _007139_, _007141_);
  or g_100383_(_007137_, _007140_, _007142_);
  or g_100384_(_013738_, _051815_, _007143_);
  not g_100385_(_007143_, _007144_);
  and g_100386_(_003437_, _007143_, _007145_);
  or g_100387_(_003436_, _007144_, _007146_);
  or g_100388_(_006974_, _007058_, _007147_);
  or g_100389_(_006967_, _007059_, _007148_);
  and g_100390_(_007147_, _007148_, _007150_);
  and g_100391_(_007146_, _007150_, _007151_);
  not g_100392_(_007151_, _007152_);
  xor g_100393_(out[293], _003436_, _007153_);
  xor g_100394_(_053170_, _003436_, _007154_);
  or g_100395_(_006977_, _007059_, _007155_);
  or g_100396_(_006983_, _007058_, _007156_);
  and g_100397_(_007155_, _007156_, _007157_);
  and g_100398_(_007154_, _007157_, _007158_);
  not g_100399_(_007158_, _007159_);
  and g_100400_(_007152_, _007159_, _007161_);
  or g_100401_(_007151_, _007158_, _007162_);
  or g_100402_(_007154_, _007157_, _007163_);
  or g_100403_(_007146_, _007150_, _007164_);
  and g_100404_(_007163_, _007164_, _007165_);
  not g_100405_(_007165_, _007166_);
  and g_100406_(_007161_, _007165_, _007167_);
  or g_100407_(_007162_, _007166_, _007168_);
  and g_100408_(_007141_, _007167_, _007169_);
  or g_100409_(_007142_, _007168_, _007170_);
  and g_100410_(_007119_, _007169_, _007172_);
  or g_100411_(_007120_, _007170_, _007173_);
  xor g_100412_(out[291], _051815_, _007174_);
  xor g_100413_(_053192_, _051815_, _007175_);
  or g_100414_(_006997_, _007059_, _007176_);
  not g_100415_(_007176_, _007177_);
  and g_100416_(_007000_, _007059_, _007178_);
  not g_100417_(_007178_, _007179_);
  and g_100418_(_007176_, _007179_, _007180_);
  or g_100419_(_007177_, _007178_, _007181_);
  or g_100420_(_007174_, _007180_, _007183_);
  and g_100421_(_007004_, _007059_, _007184_);
  not g_100422_(_007184_, _007185_);
  or g_100423_(_051642_, _007059_, _007186_);
  and g_100424_(_007185_, _007186_, _007187_);
  and g_100425_(_051816_, _007187_, _007188_);
  and g_100426_(_007174_, _007180_, _007189_);
  or g_100427_(_007175_, _007181_, _007190_);
  or g_100428_(_007188_, _007189_, _007191_);
  or g_100429_(_053126_, _007059_, _007192_);
  or g_100430_(_007014_, _007058_, _007194_);
  and g_100431_(_007192_, _007194_, _007195_);
  and g_100432_(out[289], _007195_, _007196_);
  or g_100433_(_004443_, _007059_, _007197_);
  or g_100434_(_007022_, _007058_, _007198_);
  and g_100435_(_007197_, _007198_, _007199_);
  and g_100436_(out[288], _007199_, _007200_);
  not g_100437_(_007200_, _007201_);
  xor g_100438_(out[289], _007195_, _007202_);
  xor g_100439_(_053225_, _007195_, _007203_);
  and g_100440_(_007201_, _007202_, _007205_);
  or g_100441_(_007200_, _007203_, _007206_);
  or g_100442_(_007196_, _007205_, _007207_);
  xor g_100443_(_051816_, _007187_, _007208_);
  and g_100444_(_007183_, _007191_, _007209_);
  and g_100445_(_007183_, _007208_, _007210_);
  and g_100446_(_007207_, _007210_, _007211_);
  or g_100447_(_007209_, _007211_, _007212_);
  and g_100448_(_007172_, _007212_, _007213_);
  and g_100449_(_007162_, _007163_, _007214_);
  and g_100450_(_007141_, _007214_, _007216_);
  and g_100451_(_007128_, _007134_, _007217_);
  or g_100452_(_007135_, _007217_, _007218_);
  or g_100453_(_007216_, _007218_, _007219_);
  and g_100454_(_007119_, _007219_, _007220_);
  and g_100455_(_007075_, _007077_, _007221_);
  and g_100456_(_007097_, _007115_, _007222_);
  or g_100457_(_007221_, _007222_, _007223_);
  or g_100458_(_007220_, _007223_, _007224_);
  or g_100459_(_007213_, _007224_, _007225_);
  or g_100460_(out[288], _007199_, _007227_);
  and g_100461_(_007190_, _007227_, _007228_);
  and g_100462_(_007210_, _007228_, _007229_);
  not g_100463_(_007229_, _007230_);
  or g_100464_(_007206_, _007230_, _007231_);
  or g_100465_(_007173_, _007231_, _007232_);
  and g_100466_(_007225_, _007232_, _007233_);
  not g_100467_(_007233_, _007234_);
  or g_100468_(_007065_, _007233_, _007235_);
  not g_100469_(_007235_, _007236_);
  and g_100470_(_007067_, _007233_, _007238_);
  not g_100471_(_007238_, _007239_);
  and g_100472_(_007235_, _007239_, _007240_);
  or g_100473_(_007236_, _007238_, _007241_);
  or g_100474_(_003448_, _003458_, _007242_);
  xor g_100475_(out[314], _003456_, _007243_);
  not g_100476_(_007243_, _007244_);
  or g_100477_(_007241_, _007244_, _007245_);
  and g_100478_(_007242_, _007245_, _007246_);
  not g_100479_(_007246_, _007247_);
  and g_100480_(_003448_, _003458_, _007249_);
  and g_100481_(_007241_, _007244_, _007250_);
  or g_100482_(_007249_, _007250_, _007251_);
  and g_100483_(out[313], _003455_, _007252_);
  xor g_100484_(out[313], _003455_, _007253_);
  xor g_100485_(_053335_, _003455_, _007254_);
  or g_100486_(_007090_, _007233_, _007255_);
  or g_100487_(_007084_, _007234_, _007256_);
  and g_100488_(_007255_, _007256_, _007257_);
  and g_100489_(_007254_, _007257_, _007258_);
  or g_100490_(_007251_, _007258_, _007260_);
  or g_100491_(_007247_, _007260_, _007261_);
  not g_100492_(_007261_, _007262_);
  xor g_100493_(out[312], _003454_, _007263_);
  xor g_100494_(_053258_, _003454_, _007264_);
  or g_100495_(_007106_, _007233_, _007265_);
  not g_100496_(_007265_, _007266_);
  and g_100497_(_007100_, _007233_, _007267_);
  not g_100498_(_007267_, _007268_);
  and g_100499_(_007265_, _007268_, _007269_);
  or g_100500_(_007266_, _007267_, _007271_);
  and g_100501_(_007263_, _007271_, _007272_);
  or g_100502_(_007264_, _007269_, _007273_);
  or g_100503_(_007254_, _007257_, _007274_);
  or g_100504_(_007263_, _007271_, _007275_);
  and g_100505_(_007274_, _007275_, _007276_);
  not g_100506_(_007276_, _007277_);
  and g_100507_(_007273_, _007276_, _007278_);
  or g_100508_(_007272_, _007277_, _007279_);
  and g_100509_(_007262_, _007278_, _007280_);
  or g_100510_(_007261_, _007279_, _007282_);
  xor g_100511_(out[311], _003452_, _007283_);
  xor g_100512_(_053247_, _003452_, _007284_);
  and g_100513_(_007121_, _007233_, _007285_);
  not g_100514_(_007285_, _007286_);
  or g_100515_(_007126_, _007233_, _007287_);
  not g_100516_(_007287_, _007288_);
  and g_100517_(_007286_, _007287_, _007289_);
  or g_100518_(_007285_, _007288_, _007290_);
  or g_100519_(_007284_, _007290_, _007291_);
  xor g_100520_(out[310], _003451_, _007293_);
  not g_100521_(_007293_, _007294_);
  and g_100522_(_007130_, _007233_, _007295_);
  or g_100523_(_007133_, _007233_, _007296_);
  not g_100524_(_007296_, _007297_);
  or g_100525_(_007295_, _007297_, _007298_);
  not g_100526_(_007298_, _007299_);
  or g_100527_(_007293_, _007298_, _007300_);
  and g_100528_(_007284_, _007290_, _007301_);
  xor g_100529_(out[309], _003450_, _007302_);
  and g_100530_(_007154_, _007233_, _007304_);
  not g_100531_(_007304_, _007305_);
  or g_100532_(_007157_, _007233_, _007306_);
  not g_100533_(_007306_, _007307_);
  and g_100534_(_007305_, _007306_, _007308_);
  or g_100535_(_007304_, _007307_, _007309_);
  and g_100536_(_007302_, _007309_, _007310_);
  xor g_100537_(_007284_, _007289_, _007311_);
  xor g_100538_(_007294_, _007298_, _007312_);
  or g_100539_(_007311_, _007312_, _007313_);
  or g_100540_(_007310_, _007313_, _007315_);
  not g_100541_(_007315_, _007316_);
  xor g_100542_(out[308], _003449_, _007317_);
  xor g_100543_(_053291_, _003449_, _007318_);
  or g_100544_(_007150_, _007233_, _007319_);
  not g_100545_(_007319_, _007320_);
  and g_100546_(_007146_, _007233_, _007321_);
  not g_100547_(_007321_, _007322_);
  and g_100548_(_007319_, _007322_, _007323_);
  or g_100549_(_007320_, _007321_, _007324_);
  or g_100550_(_007317_, _007324_, _007326_);
  or g_100551_(_007302_, _007309_, _007327_);
  and g_100552_(_007326_, _007327_, _007328_);
  not g_100553_(_007328_, _007329_);
  and g_100554_(_007317_, _007324_, _007330_);
  or g_100555_(_007318_, _007323_, _007331_);
  and g_100556_(_007328_, _007331_, _007332_);
  or g_100557_(_007329_, _007330_, _007333_);
  and g_100558_(_007316_, _007332_, _007334_);
  or g_100559_(_007315_, _007333_, _007335_);
  or g_100560_(_007187_, _007233_, _007337_);
  not g_100561_(_007337_, _007338_);
  and g_100562_(_051816_, _007233_, _007339_);
  or g_100563_(_007338_, _007339_, _007340_);
  or g_100564_(_051958_, _007340_, _007341_);
  xor g_100565_(out[307], _051956_, _007342_);
  xor g_100566_(_053302_, _051956_, _007343_);
  and g_100567_(_007174_, _007233_, _007344_);
  not g_100568_(_007344_, _007345_);
  and g_100569_(_007181_, _007234_, _007346_);
  or g_100570_(_007180_, _007233_, _007348_);
  and g_100571_(_007345_, _007348_, _007349_);
  or g_100572_(_007344_, _007346_, _007350_);
  or g_100573_(_007343_, _007350_, _007351_);
  and g_100574_(_007343_, _007350_, _007352_);
  xor g_100575_(_007342_, _007349_, _007353_);
  xor g_100576_(_007343_, _007349_, _007354_);
  xor g_100577_(_051958_, _007340_, _007355_);
  xor g_100578_(_051957_, _007340_, _007356_);
  and g_100579_(_007353_, _007355_, _007357_);
  or g_100580_(_007354_, _007356_, _007359_);
  and g_100581_(out[289], _007233_, _007360_);
  or g_100582_(_007195_, _007233_, _007361_);
  not g_100583_(_007361_, _007362_);
  or g_100584_(_007360_, _007362_, _007363_);
  or g_100585_(_053324_, _007363_, _007364_);
  or g_100586_(_004476_, _007234_, _007365_);
  or g_100587_(_007199_, _007233_, _007366_);
  and g_100588_(_007365_, _007366_, _007367_);
  and g_100589_(out[304], _007367_, _007368_);
  xor g_100590_(out[305], _007363_, _007370_);
  or g_100591_(_007368_, _007370_, _007371_);
  not g_100592_(_007371_, _007372_);
  and g_100593_(_007364_, _007371_, _007373_);
  or g_100594_(_007359_, _007373_, _007374_);
  or g_100595_(_007341_, _007352_, _007375_);
  and g_100596_(_007351_, _007375_, _007376_);
  and g_100597_(_007374_, _007376_, _007377_);
  or g_100598_(_007335_, _007377_, _007378_);
  or g_100599_(_007315_, _007328_, _007379_);
  or g_100600_(_007300_, _007301_, _007381_);
  and g_100601_(_007291_, _007381_, _007382_);
  and g_100602_(_007379_, _007382_, _007383_);
  and g_100603_(_007378_, _007383_, _007384_);
  or g_100604_(_007282_, _007384_, _007385_);
  or g_100605_(_007246_, _007249_, _007386_);
  or g_100606_(_007261_, _007276_, _007387_);
  and g_100607_(_007386_, _007387_, _007388_);
  and g_100608_(_007385_, _007388_, _007389_);
  or g_100609_(out[304], _007367_, _007390_);
  and g_100610_(_007357_, _007390_, _007392_);
  and g_100611_(_007372_, _007392_, _007393_);
  and g_100612_(_007334_, _007393_, _007394_);
  and g_100613_(_007280_, _007394_, _007395_);
  or g_100614_(_007389_, _007395_, _007396_);
  not g_100615_(_007396_, _007397_);
  and g_100616_(_007241_, _007396_, _007398_);
  or g_100617_(_007240_, _007397_, _007399_);
  and g_100618_(_007243_, _007397_, _007400_);
  or g_100619_(_007244_, _007396_, _007401_);
  and g_100620_(_007399_, _007401_, _007403_);
  or g_100621_(_007398_, _007400_, _007404_);
  and g_100622_(_003460_, _003476_, _007405_);
  or g_100623_(_003461_, _003474_, _007406_);
  xor g_100624_(out[330], _003471_, _007407_);
  xor g_100625_(_004553_, _003471_, _007408_);
  and g_100626_(_007403_, _007407_, _007409_);
  or g_100627_(_007404_, _007408_, _007410_);
  and g_100628_(_007406_, _007410_, _007411_);
  or g_100629_(_007405_, _007409_, _007412_);
  and g_100630_(_007404_, _007408_, _007414_);
  or g_100631_(_007403_, _007407_, _007415_);
  and g_100632_(_003461_, _003474_, _007416_);
  or g_100633_(_003460_, _003476_, _007417_);
  and g_100634_(out[329], _003470_, _007418_);
  xor g_100635_(out[329], _003470_, _007419_);
  or g_100636_(_003472_, _007418_, _007420_);
  or g_100637_(_007257_, _007397_, _007421_);
  or g_100638_(_007253_, _007396_, _007422_);
  and g_100639_(_007421_, _007422_, _007423_);
  not g_100640_(_007423_, _007425_);
  and g_100641_(_007420_, _007423_, _007426_);
  or g_100642_(_007419_, _007425_, _007427_);
  xor g_100643_(out[328], _003469_, _007428_);
  xor g_100644_(_053357_, _003469_, _007429_);
  or g_100645_(_007263_, _007396_, _007430_);
  or g_100646_(_007269_, _007397_, _007431_);
  and g_100647_(_007430_, _007431_, _007432_);
  not g_100648_(_007432_, _007433_);
  and g_100649_(_007428_, _007433_, _007434_);
  or g_100650_(_007429_, _007432_, _007436_);
  and g_100651_(_007419_, _007425_, _007437_);
  or g_100652_(_007420_, _007423_, _007438_);
  and g_100653_(_007436_, _007438_, _007439_);
  or g_100654_(_007434_, _007437_, _007440_);
  and g_100655_(_007429_, _007432_, _007441_);
  or g_100656_(_007428_, _007433_, _007442_);
  and g_100657_(_007415_, _007417_, _007443_);
  or g_100658_(_007414_, _007416_, _007444_);
  and g_100659_(_007411_, _007443_, _007445_);
  or g_100660_(_007412_, _007444_, _007447_);
  and g_100661_(_007427_, _007442_, _007448_);
  or g_100662_(_007426_, _007441_, _007449_);
  and g_100663_(_007439_, _007448_, _007450_);
  or g_100664_(_007440_, _007449_, _007451_);
  and g_100665_(_007445_, _007450_, _007452_);
  or g_100666_(_007447_, _007451_, _007453_);
  or g_100667_(_051958_, _007396_, _007454_);
  and g_100668_(_007340_, _007396_, _007455_);
  not g_100669_(_007455_, _007456_);
  and g_100670_(_007454_, _007456_, _007458_);
  not g_100671_(_007458_, _007459_);
  and g_100672_(_052167_, _007458_, _007460_);
  or g_100673_(_052168_, _007459_, _007461_);
  xor g_100674_(out[323], _052166_, _007462_);
  xor g_100675_(_053390_, _052166_, _007463_);
  or g_100676_(_007343_, _007396_, _007464_);
  or g_100677_(_007349_, _007397_, _007465_);
  and g_100678_(_007464_, _007465_, _007466_);
  not g_100679_(_007466_, _007467_);
  and g_100680_(_007462_, _007466_, _007469_);
  not g_100681_(_007469_, _007470_);
  and g_100682_(_007461_, _007470_, _007471_);
  or g_100683_(_007460_, _007469_, _007472_);
  or g_100684_(_053324_, _007396_, _007473_);
  and g_100685_(_007363_, _007396_, _007474_);
  not g_100686_(_007474_, _007475_);
  and g_100687_(_007473_, _007475_, _007476_);
  and g_100688_(out[321], _007476_, _007477_);
  not g_100689_(_007477_, _007478_);
  or g_100690_(_004509_, _007396_, _007480_);
  or g_100691_(_007367_, _007397_, _007481_);
  and g_100692_(_007480_, _007481_, _007482_);
  and g_100693_(out[320], _007482_, _007483_);
  not g_100694_(_007483_, _007484_);
  xor g_100695_(out[321], _007476_, _007485_);
  xor g_100696_(_053423_, _007476_, _007486_);
  and g_100697_(_007484_, _007485_, _007487_);
  or g_100698_(_007483_, _007486_, _007488_);
  and g_100699_(_007478_, _007488_, _007489_);
  or g_100700_(_007477_, _007487_, _007491_);
  and g_100701_(_052168_, _007459_, _007492_);
  or g_100702_(_052167_, _007458_, _007493_);
  and g_100703_(_007491_, _007493_, _007494_);
  or g_100704_(_007489_, _007492_, _007495_);
  and g_100705_(_007471_, _007493_, _007496_);
  or g_100706_(_007472_, _007492_, _007497_);
  and g_100707_(_007471_, _007495_, _007498_);
  or g_100708_(_007472_, _007494_, _007499_);
  and g_100709_(_007463_, _007467_, _007500_);
  or g_100710_(_007462_, _007466_, _007502_);
  xor g_100711_(out[327], _003468_, _007503_);
  xor g_100712_(_053346_, _003468_, _007504_);
  and g_100713_(_007283_, _007397_, _007505_);
  or g_100714_(_007284_, _007396_, _007506_);
  and g_100715_(_007290_, _007396_, _007507_);
  or g_100716_(_007289_, _007397_, _007508_);
  and g_100717_(_007506_, _007508_, _007509_);
  or g_100718_(_007505_, _007507_, _007510_);
  and g_100719_(_007503_, _007509_, _007511_);
  or g_100720_(_007504_, _007510_, _007513_);
  xor g_100721_(out[326], _003467_, _007514_);
  not g_100722_(_007514_, _007515_);
  or g_100723_(_007293_, _007396_, _007516_);
  or g_100724_(_007299_, _007397_, _007517_);
  and g_100725_(_007516_, _007517_, _007518_);
  not g_100726_(_007518_, _007519_);
  and g_100727_(_007515_, _007518_, _007520_);
  or g_100728_(_007514_, _007519_, _007521_);
  and g_100729_(_007504_, _007510_, _007522_);
  or g_100730_(_007503_, _007509_, _007524_);
  xor g_100731_(out[325], _003465_, _007525_);
  xor g_100732_(_053368_, _003465_, _007526_);
  or g_100733_(_007302_, _007396_, _007527_);
  or g_100734_(_007308_, _007397_, _007528_);
  and g_100735_(_007527_, _007528_, _007529_);
  not g_100736_(_007529_, _007530_);
  and g_100737_(_007525_, _007530_, _007531_);
  or g_100738_(_007526_, _007529_, _007532_);
  and g_100739_(_007513_, _007524_, _007533_);
  or g_100740_(_007511_, _007522_, _007535_);
  xor g_100741_(_007515_, _007518_, _007536_);
  xor g_100742_(_007514_, _007518_, _007537_);
  and g_100743_(_007533_, _007536_, _007538_);
  or g_100744_(_007535_, _007537_, _007539_);
  and g_100745_(_007532_, _007538_, _007540_);
  or g_100746_(_007531_, _007539_, _007541_);
  or g_100747_(_014046_, _052166_, _007542_);
  not g_100748_(_007542_, _007543_);
  and g_100749_(_003466_, _007542_, _007544_);
  or g_100750_(_003465_, _007543_, _007546_);
  or g_100751_(_007317_, _007396_, _007547_);
  or g_100752_(_007323_, _007397_, _007548_);
  and g_100753_(_007547_, _007548_, _007549_);
  not g_100754_(_007549_, _007550_);
  and g_100755_(_007546_, _007549_, _007551_);
  or g_100756_(_007544_, _007550_, _007552_);
  and g_100757_(_007526_, _007529_, _007553_);
  or g_100758_(_007525_, _007530_, _007554_);
  and g_100759_(_007552_, _007554_, _007555_);
  or g_100760_(_007551_, _007553_, _007557_);
  and g_100761_(_007544_, _007550_, _007558_);
  or g_100762_(_007546_, _007549_, _007559_);
  and g_100763_(_007555_, _007559_, _007560_);
  or g_100764_(_007557_, _007558_, _007561_);
  and g_100765_(_007540_, _007560_, _007562_);
  or g_100766_(_007541_, _007561_, _007563_);
  and g_100767_(_007502_, _007562_, _007564_);
  or g_100768_(_007498_, _007563_, _007565_);
  and g_100769_(_007499_, _007564_, _007566_);
  or g_100770_(_007500_, _007565_, _007568_);
  and g_100771_(_007540_, _007557_, _007569_);
  or g_100772_(_007541_, _007555_, _007570_);
  and g_100773_(_007520_, _007524_, _007571_);
  or g_100774_(_007521_, _007522_, _007572_);
  and g_100775_(_007513_, _007572_, _007573_);
  or g_100776_(_007511_, _007571_, _007574_);
  and g_100777_(_007570_, _007573_, _007575_);
  or g_100778_(_007569_, _007574_, _007576_);
  and g_100779_(_007568_, _007575_, _007577_);
  or g_100780_(_007566_, _007576_, _007579_);
  and g_100781_(_007452_, _007579_, _007580_);
  or g_100782_(_007453_, _007577_, _007581_);
  and g_100783_(_007427_, _007441_, _007582_);
  or g_100784_(_007426_, _007442_, _007583_);
  and g_100785_(_007438_, _007583_, _007584_);
  or g_100786_(_007437_, _007582_, _007585_);
  and g_100787_(_007412_, _007417_, _007586_);
  or g_100788_(_007411_, _007416_, _007587_);
  and g_100789_(_007445_, _007585_, _007588_);
  or g_100790_(_007447_, _007584_, _007590_);
  or g_100791_(_007586_, _007588_, _007591_);
  and g_100792_(_007587_, _007590_, _007592_);
  and g_100793_(_007581_, _007592_, _007593_);
  or g_100794_(_007580_, _007591_, _007594_);
  or g_100795_(out[320], _007482_, _007595_);
  and g_100796_(_007502_, _007595_, _007596_);
  not g_100797_(_007596_, _007597_);
  and g_100798_(_007496_, _007596_, _007598_);
  or g_100799_(_007497_, _007597_, _007599_);
  and g_100800_(_007487_, _007598_, _007601_);
  or g_100801_(_007488_, _007599_, _007602_);
  and g_100802_(_007452_, _007601_, _007603_);
  or g_100803_(_007453_, _007602_, _007604_);
  and g_100804_(_007562_, _007603_, _007605_);
  or g_100805_(_007563_, _007604_, _007606_);
  and g_100806_(_007594_, _007606_, _007607_);
  or g_100807_(_007593_, _007605_, _007608_);
  and g_100808_(_007404_, _007608_, _007609_);
  or g_100809_(_007403_, _007607_, _007610_);
  and g_100810_(_007407_, _007607_, _007612_);
  or g_100811_(_007408_, _007608_, _007613_);
  and g_100812_(_007610_, _007613_, _007614_);
  or g_100813_(_007609_, _007612_, _007615_);
  xor g_100814_(out[339], _052353_, _007616_);
  xor g_100815_(_053489_, _052353_, _007617_);
  and g_100816_(_007467_, _007608_, _007618_);
  and g_100817_(_007462_, _007607_, _007619_);
  or g_100818_(_007618_, _007619_, _007620_);
  or g_100819_(_007617_, _007620_, _007621_);
  and g_100820_(_007459_, _007608_, _007623_);
  and g_100821_(_052167_, _007607_, _007624_);
  or g_100822_(_007623_, _007624_, _007625_);
  or g_100823_(_052355_, _007625_, _007626_);
  and g_100824_(_007621_, _007626_, _007627_);
  and g_100825_(_007617_, _007620_, _007628_);
  xor g_100826_(_007617_, _007620_, _007629_);
  xor g_100827_(_007616_, _007620_, _007630_);
  xor g_100828_(_052355_, _007625_, _007631_);
  xor g_100829_(_052354_, _007625_, _007632_);
  and g_100830_(_007629_, _007631_, _007634_);
  or g_100831_(_007630_, _007632_, _007635_);
  and g_100832_(out[321], _007607_, _007636_);
  not g_100833_(_007636_, _007637_);
  or g_100834_(_007476_, _007607_, _007638_);
  not g_100835_(_007638_, _007639_);
  and g_100836_(_007637_, _007638_, _007640_);
  or g_100837_(_007636_, _007639_, _007641_);
  or g_100838_(_053522_, _007641_, _007642_);
  or g_100839_(_004542_, _007608_, _007643_);
  or g_100840_(_007482_, _007607_, _007645_);
  and g_100841_(_007643_, _007645_, _007646_);
  and g_100842_(out[336], _007646_, _007647_);
  not g_100843_(_007647_, _007648_);
  xor g_100844_(out[337], _007640_, _007649_);
  xor g_100845_(_053522_, _007640_, _007650_);
  and g_100846_(_007648_, _007649_, _007651_);
  or g_100847_(_007647_, _007650_, _007652_);
  and g_100848_(_007642_, _007652_, _007653_);
  or g_100849_(_007635_, _007653_, _007654_);
  or g_100850_(_007627_, _007628_, _007656_);
  and g_100851_(_007654_, _007656_, _007657_);
  xor g_100852_(out[346], _003488_, _007658_);
  xor g_100853_(out[346], _003489_, _007659_);
  and g_100854_(_007614_, _007658_, _007660_);
  or g_100855_(_007615_, _007659_, _007661_);
  and g_100856_(_003477_, _003492_, _007662_);
  or g_100857_(_003478_, _003491_, _007663_);
  and g_100858_(_007661_, _007663_, _007664_);
  or g_100859_(_007660_, _007662_, _007665_);
  and g_100860_(_003478_, _003491_, _007667_);
  or g_100861_(_003477_, _003492_, _007668_);
  and g_100862_(_007615_, _007659_, _007669_);
  or g_100863_(_007614_, _007658_, _007670_);
  and g_100864_(_007668_, _007670_, _007671_);
  or g_100865_(_007667_, _007669_, _007672_);
  and g_100866_(out[345], _003487_, _007673_);
  xor g_100867_(out[345], _003487_, _007674_);
  or g_100868_(_003489_, _007673_, _007675_);
  and g_100869_(_007425_, _007608_, _007676_);
  and g_100870_(_007420_, _007607_, _007678_);
  or g_100871_(_007676_, _007678_, _007679_);
  or g_100872_(_007674_, _007679_, _007680_);
  xor g_100873_(out[344], _003485_, _007681_);
  xor g_100874_(_053456_, _003485_, _007682_);
  and g_100875_(_007429_, _007607_, _007683_);
  and g_100876_(_007433_, _007608_, _007684_);
  or g_100877_(_007683_, _007684_, _007685_);
  and g_100878_(_007674_, _007679_, _007686_);
  or g_100879_(_007681_, _007685_, _007687_);
  not g_100880_(_007687_, _007689_);
  or g_100881_(_007686_, _007689_, _007690_);
  xor g_100882_(_007681_, _007685_, _007691_);
  xor g_100883_(_007682_, _007685_, _007692_);
  and g_100884_(_007664_, _007671_, _007693_);
  or g_100885_(_007665_, _007672_, _007694_);
  xor g_100886_(_007674_, _007679_, _007695_);
  xor g_100887_(_007675_, _007679_, _007696_);
  and g_100888_(_007693_, _007695_, _007697_);
  or g_100889_(_007694_, _007696_, _007698_);
  and g_100890_(_007691_, _007697_, _007700_);
  or g_100891_(_007692_, _007698_, _007701_);
  xor g_100892_(out[343], _003484_, _007702_);
  xor g_100893_(_053445_, _003484_, _007703_);
  and g_100894_(_007503_, _007607_, _007704_);
  and g_100895_(_007510_, _007608_, _007705_);
  or g_100896_(_007704_, _007705_, _007706_);
  or g_100897_(_007703_, _007706_, _007707_);
  and g_100898_(_007703_, _007706_, _007708_);
  xor g_100899_(_007703_, _007706_, _007709_);
  xor g_100900_(_007702_, _007706_, _007711_);
  xor g_100901_(out[342], _003483_, _007712_);
  not g_100902_(_007712_, _007713_);
  and g_100903_(_007519_, _007608_, _007714_);
  and g_100904_(_007515_, _007607_, _007715_);
  or g_100905_(_007714_, _007715_, _007716_);
  or g_100906_(_007712_, _007716_, _007717_);
  xor g_100907_(_007712_, _007716_, _007718_);
  xor g_100908_(_007713_, _007716_, _007719_);
  and g_100909_(_007709_, _007718_, _007720_);
  or g_100910_(_007711_, _007719_, _007722_);
  or g_100911_(_014200_, _052353_, _007723_);
  not g_100912_(_007723_, _007724_);
  and g_100913_(_003482_, _007723_, _007725_);
  or g_100914_(_003481_, _007724_, _007726_);
  or g_100915_(_007549_, _007607_, _007727_);
  not g_100916_(_007727_, _007728_);
  and g_100917_(_007546_, _007607_, _007729_);
  not g_100918_(_007729_, _007730_);
  and g_100919_(_007727_, _007730_, _007731_);
  or g_100920_(_007728_, _007729_, _007733_);
  and g_100921_(_007726_, _007731_, _007734_);
  or g_100922_(_007725_, _007733_, _007735_);
  xor g_100923_(out[341], _003481_, _007736_);
  xor g_100924_(_053467_, _003481_, _007737_);
  or g_100925_(_007529_, _007607_, _007738_);
  not g_100926_(_007738_, _007739_);
  and g_100927_(_007526_, _007607_, _007740_);
  not g_100928_(_007740_, _007741_);
  and g_100929_(_007738_, _007741_, _007742_);
  or g_100930_(_007739_, _007740_, _007744_);
  and g_100931_(_007737_, _007742_, _007745_);
  or g_100932_(_007736_, _007744_, _007746_);
  and g_100933_(_007735_, _007746_, _007747_);
  or g_100934_(_007734_, _007745_, _007748_);
  and g_100935_(_007736_, _007744_, _007749_);
  and g_100936_(_007725_, _007733_, _007750_);
  or g_100937_(_007749_, _007750_, _007751_);
  not g_100938_(_007751_, _007752_);
  and g_100939_(_007747_, _007752_, _007753_);
  or g_100940_(_007748_, _007751_, _007755_);
  and g_100941_(_007720_, _007753_, _007756_);
  or g_100942_(_007722_, _007755_, _007757_);
  and g_100943_(_007700_, _007756_, _007758_);
  or g_100944_(_007701_, _007757_, _007759_);
  or g_100945_(_007657_, _007759_, _007760_);
  or g_100946_(_007722_, _007747_, _007761_);
  or g_100947_(_007749_, _007761_, _007762_);
  or g_100948_(_007708_, _007717_, _007763_);
  and g_100949_(_007707_, _007763_, _007764_);
  and g_100950_(_007762_, _007764_, _007766_);
  or g_100951_(_007701_, _007766_, _007767_);
  or g_100952_(_007664_, _007667_, _007768_);
  and g_100953_(_007690_, _007693_, _007769_);
  and g_100954_(_007680_, _007769_, _007770_);
  not g_100955_(_007770_, _007771_);
  and g_100956_(_007768_, _007771_, _007772_);
  and g_100957_(_007767_, _007772_, _007773_);
  and g_100958_(_007760_, _007773_, _007774_);
  or g_100959_(out[336], _007646_, _007775_);
  and g_100960_(_007634_, _007775_, _007777_);
  and g_100961_(_007651_, _007777_, _007778_);
  and g_100962_(_007758_, _007778_, _007779_);
  or g_100963_(_007774_, _007779_, _007780_);
  or g_100964_(_007658_, _007780_, _007781_);
  not g_100965_(_007781_, _007782_);
  and g_100966_(_007614_, _007780_, _007783_);
  or g_100967_(_007782_, _007783_, _007784_);
  xor g_100968_(out[358], _003500_, _007785_);
  xor g_100969_(_053577_, _003500_, _007786_);
  or g_100970_(_007712_, _007780_, _007788_);
  and g_100971_(_007716_, _007780_, _007789_);
  not g_100972_(_007789_, _007790_);
  and g_100973_(_007788_, _007790_, _007791_);
  not g_100974_(_007791_, _007792_);
  and g_100975_(_007786_, _007791_, _007793_);
  xor g_100976_(_007786_, _007791_, _007794_);
  xor g_100977_(_007785_, _007791_, _007795_);
  and g_100978_(_003494_, _003506_, _007796_);
  or g_100979_(_003493_, _003507_, _007797_);
  and g_100980_(out[361], _003503_, _007799_);
  xor g_100981_(out[361], _003503_, _007800_);
  xor g_100982_(_053632_, _003503_, _007801_);
  and g_100983_(_007679_, _007780_, _007802_);
  not g_100984_(_007802_, _007803_);
  or g_100985_(_007674_, _007780_, _007804_);
  not g_100986_(_007804_, _007805_);
  and g_100987_(_007803_, _007804_, _007806_);
  or g_100988_(_007802_, _007805_, _007807_);
  and g_100989_(_007801_, _007806_, _007808_);
  not g_100990_(_007808_, _007810_);
  and g_100991_(_007800_, _007807_, _007811_);
  or g_100992_(_007801_, _007806_, _007812_);
  xor g_100993_(out[360], _003502_, _007813_);
  xor g_100994_(_053555_, _003502_, _007814_);
  or g_100995_(_007681_, _007780_, _007815_);
  not g_100996_(_007815_, _007816_);
  and g_100997_(_007685_, _007780_, _007817_);
  not g_100998_(_007817_, _007818_);
  and g_100999_(_007815_, _007818_, _007819_);
  or g_101000_(_007816_, _007817_, _007821_);
  and g_101001_(_007814_, _007819_, _007822_);
  or g_101002_(_007813_, _007821_, _007823_);
  and g_101003_(_007812_, _007823_, _007824_);
  or g_101004_(_007811_, _007822_, _007825_);
  xor g_101005_(out[362], _003504_, _007826_);
  not g_101006_(_007826_, _007827_);
  and g_101007_(_007784_, _007826_, _007828_);
  not g_101008_(_007828_, _007829_);
  and g_101009_(_003493_, _003507_, _007830_);
  or g_101010_(_003494_, _003506_, _007832_);
  and g_101011_(_007829_, _007832_, _007833_);
  or g_101012_(_007828_, _007830_, _007834_);
  or g_101013_(_014354_, _052547_, _007835_);
  and g_101014_(_003499_, _007835_, _007836_);
  not g_101015_(_007836_, _007837_);
  and g_101016_(_007733_, _007780_, _007838_);
  not g_101017_(_007838_, _007839_);
  or g_101018_(_007725_, _007780_, _007840_);
  not g_101019_(_007840_, _007841_);
  and g_101020_(_007839_, _007840_, _007843_);
  or g_101021_(_007838_, _007841_, _007844_);
  and g_101022_(_007837_, _007843_, _007845_);
  or g_101023_(_007836_, _007844_, _007846_);
  xor g_101024_(_007836_, _007843_, _007847_);
  or g_101025_(_007814_, _007819_, _007848_);
  not g_101026_(_007848_, _007849_);
  xor g_101027_(out[359], _003501_, _007850_);
  xor g_101028_(_053544_, _003501_, _007851_);
  and g_101029_(_007706_, _007780_, _007852_);
  not g_101030_(_007852_, _007854_);
  or g_101031_(_007703_, _007780_, _007855_);
  not g_101032_(_007855_, _007856_);
  and g_101033_(_007854_, _007855_, _007857_);
  or g_101034_(_007852_, _007856_, _007858_);
  or g_101035_(_007850_, _007857_, _007859_);
  and g_101036_(_007850_, _007857_, _007860_);
  xor g_101037_(_007850_, _007857_, _007861_);
  xor g_101038_(_007851_, _007857_, _007862_);
  xor g_101039_(out[357], _003498_, _007863_);
  not g_101040_(_007863_, _007865_);
  or g_101041_(_007736_, _007780_, _007866_);
  not g_101042_(_007866_, _007867_);
  and g_101043_(_007744_, _007780_, _007868_);
  not g_101044_(_007868_, _007869_);
  and g_101045_(_007866_, _007869_, _007870_);
  or g_101046_(_007867_, _007868_, _007871_);
  or g_101047_(_007865_, _007870_, _007872_);
  not g_101048_(_007872_, _007873_);
  and g_101049_(_007865_, _007870_, _007874_);
  or g_101050_(_007863_, _007871_, _007876_);
  or g_101051_(_007873_, _007874_, _007877_);
  and g_101052_(_007810_, _007824_, _007878_);
  or g_101053_(_007808_, _007825_, _007879_);
  xor g_101054_(_007784_, _007826_, _007880_);
  xor g_101055_(_007784_, _007827_, _007881_);
  and g_101056_(_007797_, _007832_, _007882_);
  or g_101057_(_007796_, _007830_, _007883_);
  and g_101058_(_007880_, _007882_, _007884_);
  or g_101059_(_007881_, _007883_, _007885_);
  and g_101060_(_007848_, _007884_, _007887_);
  or g_101061_(_007849_, _007885_, _007888_);
  and g_101062_(_007878_, _007887_, _007889_);
  or g_101063_(_007879_, _007888_, _007890_);
  and g_101064_(_007794_, _007861_, _007891_);
  or g_101065_(_007795_, _007862_, _007892_);
  or g_101066_(_007847_, _007877_, _007893_);
  not g_101067_(_007893_, _007894_);
  and g_101068_(_007889_, _007894_, _007895_);
  or g_101069_(_007890_, _007893_, _007896_);
  and g_101070_(_007891_, _007895_, _007898_);
  or g_101071_(_007892_, _007896_, _007899_);
  and g_101072_(_007640_, _007780_, _007900_);
  or g_101073_(out[337], _007780_, _007901_);
  not g_101074_(_007901_, _007902_);
  or g_101075_(_007900_, _007902_, _007903_);
  and g_101076_(_007646_, _007780_, _007904_);
  or g_101077_(out[336], _007780_, _007905_);
  not g_101078_(_007905_, _007906_);
  or g_101079_(_007904_, _007906_, _007907_);
  and g_101080_(out[352], _007907_, _007909_);
  not g_101081_(_007909_, _007910_);
  and g_101082_(out[353], _007903_, _007911_);
  xor g_101083_(out[353], _007903_, _007912_);
  xor g_101084_(_053621_, _007903_, _007913_);
  and g_101085_(_007910_, _007912_, _007914_);
  or g_101086_(_007909_, _007913_, _007915_);
  or g_101087_(_052355_, _007780_, _007916_);
  and g_101088_(_007625_, _007780_, _007917_);
  not g_101089_(_007917_, _007918_);
  and g_101090_(_007916_, _007918_, _007920_);
  and g_101091_(_052548_, _007920_, _007921_);
  xor g_101092_(_052548_, _007920_, _007922_);
  xor g_101093_(out[355], _052547_, _007923_);
  xor g_101094_(_053588_, _052547_, _007924_);
  or g_101095_(_007617_, _007780_, _007925_);
  and g_101096_(_007620_, _007780_, _007926_);
  not g_101097_(_007926_, _007927_);
  and g_101098_(_007925_, _007927_, _007928_);
  not g_101099_(_007928_, _007929_);
  and g_101100_(_007924_, _007929_, _007931_);
  or g_101101_(_007923_, _007928_, _007932_);
  and g_101102_(_007923_, _007928_, _007933_);
  or g_101103_(_007924_, _007929_, _007934_);
  or g_101104_(out[352], _007907_, _007935_);
  and g_101105_(_007934_, _007935_, _007936_);
  and g_101106_(_007922_, _007932_, _007937_);
  and g_101107_(_007936_, _007937_, _007938_);
  not g_101108_(_007938_, _007939_);
  and g_101109_(_007914_, _007938_, _007940_);
  or g_101110_(_007915_, _007939_, _007942_);
  and g_101111_(_007898_, _007940_, _007943_);
  or g_101112_(_007899_, _007942_, _007944_);
  or g_101113_(_007921_, _007933_, _007945_);
  or g_101114_(_007911_, _007914_, _007946_);
  and g_101115_(_007922_, _007946_, _007947_);
  or g_101116_(_007945_, _007947_, _007948_);
  not g_101117_(_007948_, _007949_);
  and g_101118_(_007898_, _007932_, _007950_);
  or g_101119_(_007899_, _007931_, _007951_);
  and g_101120_(_007948_, _007950_, _007953_);
  or g_101121_(_007949_, _007951_, _007954_);
  and g_101122_(_007846_, _007876_, _007955_);
  or g_101123_(_007845_, _007874_, _007956_);
  and g_101124_(_007872_, _007956_, _007957_);
  or g_101125_(_007873_, _007955_, _007958_);
  and g_101126_(_007891_, _007957_, _007959_);
  or g_101127_(_007892_, _007958_, _007960_);
  and g_101128_(_007793_, _007859_, _007961_);
  or g_101129_(_007860_, _007961_, _007962_);
  not g_101130_(_007962_, _007964_);
  and g_101131_(_007960_, _007964_, _007965_);
  or g_101132_(_007959_, _007962_, _007966_);
  and g_101133_(_007889_, _007966_, _007967_);
  or g_101134_(_007890_, _007965_, _007968_);
  and g_101135_(_007825_, _007884_, _007969_);
  or g_101136_(_007824_, _007885_, _007970_);
  and g_101137_(_007810_, _007969_, _007971_);
  or g_101138_(_007808_, _007970_, _007972_);
  and g_101139_(_007797_, _007834_, _007973_);
  or g_101140_(_007796_, _007833_, _007975_);
  and g_101141_(_007972_, _007975_, _007976_);
  or g_101142_(_007971_, _007973_, _007977_);
  or g_101143_(_007967_, _007977_, _007978_);
  and g_101144_(_007968_, _007976_, _007979_);
  and g_101145_(_007954_, _007979_, _007980_);
  or g_101146_(_007953_, _007978_, _007981_);
  and g_101147_(_007944_, _007981_, _007982_);
  or g_101148_(_007943_, _007980_, _007983_);
  or g_101149_(_007784_, _007982_, _007984_);
  not g_101150_(_007984_, _007986_);
  and g_101151_(_007826_, _007982_, _007987_);
  not g_101152_(_007987_, _007988_);
  and g_101153_(_007984_, _007988_, _007989_);
  or g_101154_(_007986_, _007987_, _007990_);
  xor g_101155_(out[378], _003520_, _007991_);
  xor g_101156_(_004652_, _003520_, _007992_);
  and g_101157_(_007989_, _007991_, _007993_);
  or g_101158_(_007990_, _007992_, _007994_);
  and g_101159_(_003509_, _003524_, _007995_);
  or g_101160_(_003510_, _003523_, _007997_);
  and g_101161_(_007994_, _007997_, _007998_);
  or g_101162_(_007993_, _007995_, _007999_);
  and g_101163_(_007990_, _007992_, _008000_);
  or g_101164_(_007989_, _007991_, _008001_);
  and g_101165_(_003510_, _003523_, _008002_);
  or g_101166_(_003509_, _003524_, _008003_);
  and g_101167_(out[377], _003518_, _008004_);
  xor g_101168_(out[377], _003518_, _008005_);
  or g_101169_(_003521_, _008004_, _008006_);
  or g_101170_(_007806_, _007982_, _008008_);
  not g_101171_(_008008_, _008009_);
  and g_101172_(_007801_, _007982_, _008010_);
  not g_101173_(_008010_, _008011_);
  and g_101174_(_008008_, _008011_, _008012_);
  or g_101175_(_008009_, _008010_, _008013_);
  and g_101176_(_008006_, _008012_, _008014_);
  or g_101177_(_008005_, _008013_, _008015_);
  and g_101178_(_008003_, _008015_, _008016_);
  or g_101179_(_008002_, _008014_, _008017_);
  and g_101180_(_008001_, _008016_, _008019_);
  or g_101181_(_008000_, _008017_, _008020_);
  and g_101182_(_007998_, _008019_, _008021_);
  or g_101183_(_007999_, _008020_, _008022_);
  xor g_101184_(out[376], _003517_, _008023_);
  xor g_101185_(_053654_, _003517_, _008024_);
  and g_101186_(_007814_, _007982_, _008025_);
  not g_101187_(_008025_, _008026_);
  or g_101188_(_007819_, _007982_, _008027_);
  not g_101189_(_008027_, _008028_);
  and g_101190_(_008026_, _008027_, _008030_);
  or g_101191_(_008025_, _008028_, _008031_);
  and g_101192_(_008023_, _008031_, _008032_);
  or g_101193_(_008024_, _008030_, _008033_);
  and g_101194_(_008005_, _008013_, _008034_);
  or g_101195_(_008006_, _008012_, _008035_);
  and g_101196_(_008024_, _008030_, _008036_);
  or g_101197_(_008023_, _008031_, _008037_);
  and g_101198_(_008035_, _008037_, _008038_);
  or g_101199_(_008034_, _008036_, _008039_);
  and g_101200_(_008033_, _008038_, _008041_);
  or g_101201_(_008032_, _008039_, _008042_);
  and g_101202_(_008021_, _008041_, _008043_);
  or g_101203_(_008022_, _008042_, _008044_);
  xor g_101204_(out[374], _003515_, _008045_);
  not g_101205_(_008045_, _008046_);
  and g_101206_(_007786_, _007982_, _008047_);
  and g_101207_(_007792_, _007983_, _008048_);
  or g_101208_(_008047_, _008048_, _008049_);
  or g_101209_(_008045_, _008049_, _008050_);
  not g_101210_(_008050_, _008052_);
  xor g_101211_(out[375], _003516_, _008053_);
  xor g_101212_(_053643_, _003516_, _008054_);
  and g_101213_(_007850_, _007982_, _008055_);
  or g_101214_(_007851_, _007983_, _008056_);
  and g_101215_(_007858_, _007983_, _008057_);
  or g_101216_(_007857_, _007982_, _008058_);
  and g_101217_(_008056_, _008058_, _008059_);
  or g_101218_(_008055_, _008057_, _008060_);
  and g_101219_(_008053_, _008059_, _008061_);
  or g_101220_(_008054_, _008060_, _008063_);
  and g_101221_(_008050_, _008063_, _008064_);
  or g_101222_(_008052_, _008061_, _008065_);
  and g_101223_(_008045_, _008049_, _008066_);
  and g_101224_(_008054_, _008060_, _008067_);
  or g_101225_(_008053_, _008059_, _008068_);
  or g_101226_(_008066_, _008067_, _008069_);
  xor g_101227_(_008045_, _008049_, _008070_);
  and g_101228_(_008063_, _008070_, _008071_);
  and g_101229_(_008068_, _008071_, _008072_);
  or g_101230_(_008065_, _008069_, _008074_);
  or g_101231_(_014508_, _052741_, _008075_);
  not g_101232_(_008075_, _008076_);
  and g_101233_(_003514_, _008075_, _008077_);
  or g_101234_(_003513_, _008076_, _008078_);
  or g_101235_(_007843_, _007982_, _008079_);
  not g_101236_(_008079_, _008080_);
  and g_101237_(_007837_, _007982_, _008081_);
  not g_101238_(_008081_, _008082_);
  and g_101239_(_008079_, _008082_, _008083_);
  or g_101240_(_008080_, _008081_, _008085_);
  and g_101241_(_008078_, _008083_, _008086_);
  or g_101242_(_008077_, _008085_, _008087_);
  xor g_101243_(out[373], _003513_, _008088_);
  xor g_101244_(_053665_, _003513_, _008089_);
  and g_101245_(_007865_, _007982_, _008090_);
  not g_101246_(_008090_, _008091_);
  or g_101247_(_007870_, _007982_, _008092_);
  not g_101248_(_008092_, _008093_);
  and g_101249_(_008091_, _008092_, _008094_);
  or g_101250_(_008090_, _008093_, _008096_);
  and g_101251_(_008089_, _008094_, _008097_);
  or g_101252_(_008088_, _008096_, _008098_);
  and g_101253_(_008087_, _008098_, _008099_);
  or g_101254_(_008086_, _008097_, _008100_);
  and g_101255_(_008088_, _008096_, _008101_);
  not g_101256_(_008101_, _008102_);
  or g_101257_(_008078_, _008083_, _008103_);
  and g_101258_(_008099_, _008103_, _008104_);
  and g_101259_(_008102_, _008104_, _008105_);
  and g_101260_(_008072_, _008105_, _008107_);
  not g_101261_(_008107_, _008108_);
  and g_101262_(_008043_, _008107_, _008109_);
  or g_101263_(_008044_, _008108_, _008110_);
  xor g_101264_(out[371], _052741_, _008111_);
  xor g_101265_(_053687_, _052741_, _008112_);
  and g_101266_(_007923_, _007982_, _008113_);
  not g_101267_(_008113_, _008114_);
  or g_101268_(_007928_, _007982_, _008115_);
  not g_101269_(_008115_, _008116_);
  and g_101270_(_008114_, _008115_, _008118_);
  or g_101271_(_008113_, _008116_, _008119_);
  and g_101272_(_008111_, _008118_, _008120_);
  or g_101273_(_008112_, _008119_, _008121_);
  or g_101274_(_007920_, _007982_, _008122_);
  not g_101275_(_008122_, _008123_);
  and g_101276_(_052548_, _007982_, _008124_);
  or g_101277_(_008123_, _008124_, _008125_);
  or g_101278_(_052743_, _008125_, _008126_);
  not g_101279_(_008126_, _008127_);
  and g_101280_(_008121_, _008126_, _008129_);
  or g_101281_(_008120_, _008127_, _008130_);
  and g_101282_(_008112_, _008119_, _008131_);
  or g_101283_(_008111_, _008118_, _008132_);
  and g_101284_(_052743_, _008125_, _008133_);
  or g_101285_(_008131_, _008133_, _008134_);
  and g_101286_(_008121_, _008132_, _008135_);
  xor g_101287_(_052743_, _008125_, _008136_);
  and g_101288_(_008135_, _008136_, _008137_);
  or g_101289_(_008130_, _008134_, _008138_);
  and g_101290_(out[353], _007982_, _008140_);
  not g_101291_(_008140_, _008141_);
  or g_101292_(_007903_, _007982_, _008142_);
  not g_101293_(_008142_, _008143_);
  and g_101294_(_008141_, _008142_, _008144_);
  or g_101295_(_008140_, _008143_, _008145_);
  and g_101296_(out[369], _008144_, _008146_);
  or g_101297_(_053720_, _008145_, _008147_);
  and g_101298_(out[352], _007982_, _008148_);
  not g_101299_(_008148_, _008149_);
  or g_101300_(_007907_, _007982_, _008151_);
  not g_101301_(_008151_, _008152_);
  and g_101302_(_008149_, _008151_, _008153_);
  or g_101303_(_008148_, _008152_, _008154_);
  and g_101304_(out[368], _008153_, _008155_);
  or g_101305_(_004641_, _008154_, _008156_);
  xor g_101306_(out[369], _008144_, _008157_);
  xor g_101307_(_053720_, _008144_, _008158_);
  and g_101308_(_008156_, _008157_, _008159_);
  or g_101309_(_008155_, _008158_, _008160_);
  and g_101310_(_008147_, _008160_, _008162_);
  or g_101311_(_008146_, _008159_, _008163_);
  and g_101312_(_008137_, _008163_, _008164_);
  or g_101313_(_008138_, _008162_, _008165_);
  and g_101314_(_008130_, _008132_, _008166_);
  or g_101315_(_008129_, _008131_, _008167_);
  and g_101316_(_008165_, _008167_, _008168_);
  or g_101317_(_008164_, _008166_, _008169_);
  and g_101318_(_008109_, _008169_, _008170_);
  or g_101319_(_008110_, _008168_, _008171_);
  or g_101320_(_008099_, _008101_, _008173_);
  and g_101321_(_008072_, _008100_, _008174_);
  and g_101322_(_008102_, _008174_, _008175_);
  or g_101323_(_008074_, _008173_, _008176_);
  and g_101324_(_008065_, _008068_, _008177_);
  or g_101325_(_008064_, _008067_, _008178_);
  and g_101326_(_008176_, _008178_, _008179_);
  or g_101327_(_008175_, _008177_, _008180_);
  and g_101328_(_008043_, _008180_, _008181_);
  or g_101329_(_008044_, _008179_, _008182_);
  and g_101330_(_007999_, _008003_, _008184_);
  or g_101331_(_007998_, _008002_, _008185_);
  and g_101332_(_008021_, _008039_, _008186_);
  or g_101333_(_008022_, _008038_, _008187_);
  and g_101334_(_008185_, _008187_, _008188_);
  or g_101335_(_008184_, _008186_, _008189_);
  and g_101336_(_008182_, _008188_, _008190_);
  or g_101337_(_008181_, _008189_, _008191_);
  and g_101338_(_008171_, _008190_, _008192_);
  or g_101339_(_008170_, _008191_, _008193_);
  or g_101340_(out[368], _008153_, _008195_);
  and g_101341_(_008137_, _008195_, _008196_);
  not g_101342_(_008196_, _008197_);
  and g_101343_(_008159_, _008196_, _008198_);
  or g_101344_(_008160_, _008197_, _008199_);
  and g_101345_(_008109_, _008198_, _008200_);
  or g_101346_(_008110_, _008199_, _008201_);
  and g_101347_(_008193_, _008201_, _008202_);
  or g_101348_(_008192_, _008200_, _008203_);
  and g_101349_(_007990_, _008203_, _008204_);
  and g_101350_(_007991_, _008202_, _008206_);
  or g_101351_(_008204_, _008206_, _008207_);
  or g_101352_(_003526_, _003538_, _008208_);
  xor g_101353_(out[394], _003536_, _008209_);
  not g_101354_(_008209_, _008210_);
  or g_101355_(_008207_, _008210_, _008211_);
  and g_101356_(_008208_, _008211_, _008212_);
  and g_101357_(_003526_, _003538_, _008213_);
  xor g_101358_(_003526_, _003538_, _008214_);
  xor g_101359_(_003525_, _003538_, _008215_);
  xor g_101360_(_008207_, _008210_, _008217_);
  xor g_101361_(_008207_, _008209_, _008218_);
  and g_101362_(_008214_, _008217_, _008219_);
  or g_101363_(_008215_, _008218_, _008220_);
  xor g_101364_(out[392], _003534_, _008221_);
  xor g_101365_(_053753_, _003534_, _008222_);
  and g_101366_(_008024_, _008202_, _008223_);
  and g_101367_(_008031_, _008203_, _008224_);
  or g_101368_(_008223_, _008224_, _008225_);
  and g_101369_(_008221_, _008225_, _008226_);
  and g_101370_(out[393], _003535_, _008228_);
  xor g_101371_(out[393], _003535_, _008229_);
  xor g_101372_(_053830_, _003535_, _008230_);
  and g_101373_(_008013_, _008203_, _008231_);
  and g_101374_(_008006_, _008202_, _008232_);
  or g_101375_(_008231_, _008232_, _008233_);
  or g_101376_(_008229_, _008233_, _008234_);
  not g_101377_(_008234_, _008235_);
  or g_101378_(_008226_, _008235_, _008236_);
  or g_101379_(_008221_, _008225_, _008237_);
  not g_101380_(_008237_, _008239_);
  and g_101381_(_008229_, _008233_, _008240_);
  not g_101382_(_008240_, _008241_);
  and g_101383_(_008237_, _008241_, _008242_);
  or g_101384_(_008239_, _008240_, _008243_);
  or g_101385_(_008236_, _008243_, _008244_);
  xor g_101386_(_008221_, _008225_, _008245_);
  and g_101387_(_008234_, _008241_, _008246_);
  and g_101388_(_008219_, _008246_, _008247_);
  and g_101389_(_008245_, _008247_, _008248_);
  or g_101390_(_008220_, _008244_, _008250_);
  xor g_101391_(out[391], _003533_, _008251_);
  xor g_101392_(_053742_, _003533_, _008252_);
  and g_101393_(_008053_, _008202_, _008253_);
  or g_101394_(_008054_, _008203_, _008254_);
  and g_101395_(_008060_, _008203_, _008255_);
  or g_101396_(_008059_, _008202_, _008256_);
  and g_101397_(_008254_, _008256_, _008257_);
  or g_101398_(_008253_, _008255_, _008258_);
  and g_101399_(_008251_, _008257_, _008259_);
  or g_101400_(_008252_, _008258_, _008261_);
  xor g_101401_(out[390], _003532_, _008262_);
  xor g_101402_(_053775_, _003532_, _008263_);
  or g_101403_(_008045_, _008203_, _008264_);
  not g_101404_(_008264_, _008265_);
  and g_101405_(_008049_, _008203_, _008266_);
  not g_101406_(_008266_, _008267_);
  and g_101407_(_008264_, _008267_, _008268_);
  or g_101408_(_008265_, _008266_, _008269_);
  and g_101409_(_008263_, _008268_, _008270_);
  or g_101410_(_008262_, _008269_, _008272_);
  and g_101411_(_008252_, _008258_, _008273_);
  or g_101412_(_008251_, _008257_, _008274_);
  and g_101413_(_008261_, _008274_, _008275_);
  or g_101414_(_008259_, _008273_, _008276_);
  xor g_101415_(_008263_, _008268_, _008277_);
  xor g_101416_(_008262_, _008268_, _008278_);
  and g_101417_(_008275_, _008277_, _008279_);
  or g_101418_(_008276_, _008278_, _008280_);
  or g_101419_(_014662_, _052921_, _008281_);
  not g_101420_(_008281_, _008283_);
  and g_101421_(_003531_, _008281_, _008284_);
  or g_101422_(_003529_, _008283_, _008285_);
  and g_101423_(_008085_, _008203_, _008286_);
  not g_101424_(_008286_, _008287_);
  or g_101425_(_008077_, _008203_, _008288_);
  not g_101426_(_008288_, _008289_);
  and g_101427_(_008287_, _008288_, _008290_);
  or g_101428_(_008286_, _008289_, _008291_);
  and g_101429_(_008285_, _008290_, _008292_);
  or g_101430_(_008284_, _008291_, _008294_);
  xor g_101431_(out[389], _003529_, _008295_);
  xor g_101432_(_053764_, _003529_, _008296_);
  or g_101433_(_008088_, _008203_, _008297_);
  not g_101434_(_008297_, _008298_);
  and g_101435_(_008096_, _008203_, _008299_);
  not g_101436_(_008299_, _008300_);
  and g_101437_(_008297_, _008300_, _008301_);
  or g_101438_(_008298_, _008299_, _008302_);
  and g_101439_(_008296_, _008301_, _008303_);
  or g_101440_(_008295_, _008302_, _008305_);
  and g_101441_(_008294_, _008305_, _008306_);
  or g_101442_(_008292_, _008303_, _008307_);
  and g_101443_(_008295_, _008302_, _008308_);
  or g_101444_(_008296_, _008301_, _008309_);
  and g_101445_(_008284_, _008291_, _008310_);
  or g_101446_(_008285_, _008290_, _008311_);
  and g_101447_(_008309_, _008311_, _008312_);
  or g_101448_(_008308_, _008310_, _008313_);
  and g_101449_(_008306_, _008312_, _008314_);
  or g_101450_(_008307_, _008313_, _008316_);
  and g_101451_(_008279_, _008314_, _008317_);
  or g_101452_(_008280_, _008316_, _008318_);
  and g_101453_(_008248_, _008317_, _008319_);
  or g_101454_(_008250_, _008318_, _008320_);
  xor g_101455_(out[387], _052921_, _008321_);
  xor g_101456_(_053786_, _052921_, _008322_);
  and g_101457_(_008111_, _008202_, _008323_);
  and g_101458_(_008119_, _008203_, _008324_);
  or g_101459_(_008323_, _008324_, _008325_);
  or g_101460_(_008322_, _008325_, _008327_);
  and g_101461_(_008125_, _008203_, _008328_);
  and g_101462_(_052742_, _008202_, _008329_);
  or g_101463_(_008328_, _008329_, _008330_);
  and g_101464_(_008322_, _008325_, _008331_);
  or g_101465_(_052923_, _008330_, _008332_);
  xor g_101466_(_008322_, _008325_, _008333_);
  xor g_101467_(_008321_, _008325_, _008334_);
  xor g_101468_(_052923_, _008330_, _008335_);
  xor g_101469_(_052922_, _008330_, _008336_);
  and g_101470_(_008333_, _008335_, _008338_);
  or g_101471_(_008334_, _008336_, _008339_);
  or g_101472_(_053720_, _008203_, _008340_);
  or g_101473_(_008144_, _008202_, _008341_);
  and g_101474_(_008340_, _008341_, _008342_);
  and g_101475_(out[385], _008342_, _008343_);
  not g_101476_(_008343_, _008344_);
  or g_101477_(_004641_, _008203_, _008345_);
  not g_101478_(_008345_, _008346_);
  and g_101479_(_008154_, _008203_, _008347_);
  or g_101480_(_008153_, _008202_, _008349_);
  and g_101481_(_008345_, _008349_, _008350_);
  or g_101482_(_008346_, _008347_, _008351_);
  and g_101483_(out[384], _008350_, _008352_);
  or g_101484_(_004674_, _008351_, _008353_);
  xor g_101485_(out[385], _008342_, _008354_);
  xor g_101486_(_053819_, _008342_, _008355_);
  and g_101487_(_008353_, _008354_, _008356_);
  or g_101488_(_008352_, _008355_, _008357_);
  and g_101489_(_008344_, _008357_, _008358_);
  or g_101490_(_008343_, _008356_, _008360_);
  and g_101491_(_008338_, _008360_, _008361_);
  or g_101492_(_008339_, _008358_, _008362_);
  or g_101493_(_008331_, _008332_, _008363_);
  and g_101494_(_008327_, _008363_, _008364_);
  not g_101495_(_008364_, _008365_);
  and g_101496_(_008362_, _008364_, _008366_);
  or g_101497_(_008361_, _008365_, _008367_);
  and g_101498_(_008319_, _008367_, _008368_);
  or g_101499_(_008320_, _008366_, _008369_);
  and g_101500_(_008279_, _008307_, _008371_);
  or g_101501_(_008280_, _008306_, _008372_);
  and g_101502_(_008309_, _008371_, _008373_);
  or g_101503_(_008308_, _008372_, _008374_);
  and g_101504_(_008270_, _008274_, _008375_);
  or g_101505_(_008272_, _008273_, _008376_);
  and g_101506_(_008261_, _008376_, _008377_);
  or g_101507_(_008259_, _008375_, _008378_);
  and g_101508_(_008374_, _008377_, _008379_);
  or g_101509_(_008373_, _008378_, _008380_);
  and g_101510_(_008248_, _008380_, _008382_);
  or g_101511_(_008250_, _008379_, _008383_);
  and g_101512_(_008219_, _008243_, _008384_);
  or g_101513_(_008220_, _008242_, _008385_);
  and g_101514_(_008234_, _008384_, _008386_);
  or g_101515_(_008235_, _008385_, _008387_);
  or g_101516_(_008212_, _008213_, _008388_);
  not g_101517_(_008388_, _008389_);
  and g_101518_(_008387_, _008388_, _008390_);
  or g_101519_(_008386_, _008389_, _008391_);
  and g_101520_(_008383_, _008390_, _008393_);
  or g_101521_(_008382_, _008391_, _008394_);
  and g_101522_(_008369_, _008393_, _008395_);
  or g_101523_(_008368_, _008394_, _008396_);
  and g_101524_(_004674_, _008351_, _008397_);
  or g_101525_(_008339_, _008397_, _008398_);
  or g_101526_(_008357_, _008398_, _008399_);
  or g_101527_(_008320_, _008399_, _008400_);
  not g_101528_(_008400_, _008401_);
  and g_101529_(_008396_, _008400_, _008402_);
  or g_101530_(_008395_, _008401_, _008404_);
  and g_101531_(_008207_, _008404_, _008405_);
  not g_101532_(_008405_, _008406_);
  or g_101533_(_008210_, _008404_, _008407_);
  not g_101534_(_008407_, _008408_);
  and g_101535_(_008406_, _008407_, _008409_);
  or g_101536_(_008405_, _008408_, _008410_);
  and g_101537_(_008330_, _008404_, _008411_);
  not g_101538_(_008411_, _008412_);
  or g_101539_(_052923_, _008404_, _008413_);
  not g_101540_(_008413_, _008415_);
  and g_101541_(_008412_, _008413_, _008416_);
  or g_101542_(_008411_, _008415_, _008417_);
  and g_101543_(_053010_, _008416_, _008418_);
  xor g_101544_(out[403], _053009_, _008419_);
  xor g_101545_(_053885_, _053009_, _008420_);
  and g_101546_(_008325_, _008404_, _008421_);
  not g_101547_(_008421_, _008422_);
  or g_101548_(_008322_, _008404_, _008423_);
  not g_101549_(_008423_, _008424_);
  and g_101550_(_008422_, _008423_, _008426_);
  or g_101551_(_008421_, _008424_, _008427_);
  and g_101552_(_008419_, _008426_, _008428_);
  or g_101553_(_008418_, _008428_, _008429_);
  or g_101554_(_053819_, _008404_, _008430_);
  or g_101555_(_008342_, _008402_, _008431_);
  and g_101556_(_008430_, _008431_, _008432_);
  and g_101557_(out[401], _008432_, _008433_);
  or g_101558_(_004674_, _008404_, _008434_);
  or g_101559_(_008350_, _008402_, _008435_);
  and g_101560_(_008434_, _008435_, _008437_);
  and g_101561_(out[400], _008437_, _008438_);
  not g_101562_(_008438_, _008439_);
  xor g_101563_(out[401], _008432_, _008440_);
  xor g_101564_(_053918_, _008432_, _008441_);
  and g_101565_(_008439_, _008440_, _008442_);
  or g_101566_(_008438_, _008441_, _008443_);
  or g_101567_(_008433_, _008442_, _008444_);
  xor g_101568_(_053010_, _008416_, _008445_);
  xor g_101569_(_053011_, _008416_, _008446_);
  and g_101570_(_008444_, _008445_, _008448_);
  or g_101571_(_008429_, _008448_, _008449_);
  not g_101572_(_008449_, _008450_);
  xor g_101573_(out[410], _003551_, _008451_);
  not g_101574_(_008451_, _008452_);
  and g_101575_(_008409_, _008451_, _008453_);
  or g_101576_(_008410_, _008452_, _008454_);
  and g_101577_(_003540_, _003555_, _008455_);
  or g_101578_(_003542_, _003554_, _008456_);
  and g_101579_(_008454_, _008456_, _008457_);
  or g_101580_(_008453_, _008455_, _008459_);
  and g_101581_(_008410_, _008452_, _008460_);
  or g_101582_(_008409_, _008451_, _008461_);
  and g_101583_(_003542_, _003554_, _008462_);
  or g_101584_(_003540_, _003555_, _008463_);
  and g_101585_(_008461_, _008463_, _008464_);
  or g_101586_(_008460_, _008462_, _008465_);
  and g_101587_(_008457_, _008464_, _008466_);
  or g_101588_(_008459_, _008465_, _008467_);
  xor g_101589_(out[408], _003549_, _008468_);
  xor g_101590_(_053852_, _003549_, _008470_);
  or g_101591_(_008221_, _008404_, _008471_);
  not g_101592_(_008471_, _008472_);
  and g_101593_(_008225_, _008404_, _008473_);
  not g_101594_(_008473_, _008474_);
  and g_101595_(_008471_, _008474_, _008475_);
  or g_101596_(_008472_, _008473_, _008476_);
  and g_101597_(_008470_, _008475_, _008477_);
  or g_101598_(_008468_, _008476_, _008478_);
  and g_101599_(out[409], _003550_, _008479_);
  xor g_101600_(out[409], _003550_, _008481_);
  xor g_101601_(_053929_, _003550_, _008482_);
  and g_101602_(_008233_, _008404_, _008483_);
  not g_101603_(_008483_, _008484_);
  or g_101604_(_008229_, _008404_, _008485_);
  not g_101605_(_008485_, _008486_);
  and g_101606_(_008484_, _008485_, _008487_);
  or g_101607_(_008483_, _008486_, _008488_);
  and g_101608_(_008481_, _008488_, _008489_);
  or g_101609_(_008482_, _008487_, _008490_);
  and g_101610_(_008478_, _008490_, _008492_);
  or g_101611_(_008477_, _008489_, _008493_);
  and g_101612_(_008482_, _008487_, _008494_);
  or g_101613_(_008481_, _008488_, _008495_);
  and g_101614_(_008468_, _008476_, _008496_);
  or g_101615_(_008470_, _008475_, _008497_);
  and g_101616_(_008495_, _008497_, _008498_);
  or g_101617_(_008494_, _008496_, _008499_);
  and g_101618_(_008492_, _008498_, _008500_);
  or g_101619_(_008493_, _008499_, _008501_);
  and g_101620_(_008466_, _008500_, _008503_);
  or g_101621_(_008467_, _008501_, _008504_);
  xor g_101622_(out[406], _003547_, _008505_);
  xor g_101623_(_053874_, _003547_, _008506_);
  or g_101624_(_008262_, _008404_, _008507_);
  or g_101625_(_008268_, _008402_, _008508_);
  and g_101626_(_008507_, _008508_, _008509_);
  and g_101627_(_008506_, _008509_, _008510_);
  xor g_101628_(out[407], _003548_, _008511_);
  xor g_101629_(_053841_, _003548_, _008512_);
  or g_101630_(_008252_, _008404_, _008514_);
  or g_101631_(_008257_, _008402_, _008515_);
  and g_101632_(_008514_, _008515_, _008516_);
  or g_101633_(_008511_, _008516_, _008517_);
  not g_101634_(_008517_, _008518_);
  and g_101635_(_008511_, _008516_, _008519_);
  xor g_101636_(_008506_, _008509_, _008520_);
  xor g_101637_(_008505_, _008509_, _008521_);
  or g_101638_(_008519_, _008521_, _008522_);
  xor g_101639_(_008511_, _008516_, _008523_);
  and g_101640_(_008520_, _008523_, _008525_);
  or g_101641_(_008518_, _008522_, _008526_);
  or g_101642_(_014816_, _053009_, _008527_);
  not g_101643_(_008527_, _008528_);
  and g_101644_(_003546_, _008527_, _008529_);
  or g_101645_(_003545_, _008528_, _008530_);
  and g_101646_(_008291_, _008404_, _008531_);
  not g_101647_(_008531_, _008532_);
  or g_101648_(_008284_, _008404_, _008533_);
  not g_101649_(_008533_, _008534_);
  and g_101650_(_008532_, _008533_, _008536_);
  or g_101651_(_008531_, _008534_, _008537_);
  and g_101652_(_008530_, _008536_, _008538_);
  or g_101653_(_008529_, _008537_, _008539_);
  xor g_101654_(out[405], _003545_, _008540_);
  xor g_101655_(_053863_, _003545_, _008541_);
  or g_101656_(_008295_, _008404_, _008542_);
  not g_101657_(_008542_, _008543_);
  and g_101658_(_008302_, _008404_, _008544_);
  not g_101659_(_008544_, _008545_);
  and g_101660_(_008542_, _008545_, _008547_);
  or g_101661_(_008543_, _008544_, _008548_);
  and g_101662_(_008541_, _008547_, _008549_);
  or g_101663_(_008540_, _008548_, _008550_);
  and g_101664_(_008539_, _008550_, _008551_);
  or g_101665_(_008538_, _008549_, _008552_);
  or g_101666_(_008541_, _008547_, _008553_);
  not g_101667_(_008553_, _008554_);
  or g_101668_(_008530_, _008536_, _008555_);
  and g_101669_(_008553_, _008555_, _008556_);
  not g_101670_(_008556_, _008558_);
  and g_101671_(_008551_, _008556_, _008559_);
  or g_101672_(_008552_, _008558_, _008560_);
  and g_101673_(_008525_, _008559_, _008561_);
  or g_101674_(_008504_, _008560_, _008562_);
  and g_101675_(_008503_, _008561_, _008563_);
  or g_101676_(_008526_, _008562_, _008564_);
  and g_101677_(_008420_, _008427_, _008565_);
  or g_101678_(_008419_, _008426_, _008566_);
  and g_101679_(_008563_, _008566_, _008567_);
  or g_101680_(_008564_, _008565_, _008569_);
  or g_101681_(_008446_, _008565_, _008570_);
  xor g_101682_(_008419_, _008426_, _008571_);
  and g_101683_(_008449_, _008567_, _008572_);
  or g_101684_(_008450_, _008569_, _008573_);
  and g_101685_(_008525_, _008553_, _008574_);
  or g_101686_(_008526_, _008551_, _008575_);
  and g_101687_(_008552_, _008574_, _008576_);
  or g_101688_(_008554_, _008575_, _008577_);
  and g_101689_(_008510_, _008517_, _008578_);
  or g_101690_(_008519_, _008578_, _008580_);
  not g_101691_(_008580_, _008581_);
  and g_101692_(_008577_, _008581_, _008582_);
  or g_101693_(_008576_, _008580_, _008583_);
  and g_101694_(_008503_, _008583_, _008584_);
  or g_101695_(_008504_, _008582_, _008585_);
  and g_101696_(_008466_, _008493_, _008586_);
  not g_101697_(_008586_, _008587_);
  and g_101698_(_008495_, _008586_, _008588_);
  or g_101699_(_008494_, _008587_, _008589_);
  and g_101700_(_008459_, _008463_, _008591_);
  not g_101701_(_008591_, _008592_);
  and g_101702_(_008589_, _008592_, _008593_);
  or g_101703_(_008588_, _008591_, _008594_);
  and g_101704_(_008585_, _008593_, _008595_);
  or g_101705_(_008584_, _008594_, _008596_);
  and g_101706_(_008573_, _008595_, _008597_);
  or g_101707_(_008572_, _008596_, _008598_);
  or g_101708_(out[400], _008437_, _008599_);
  not g_101709_(_008599_, _008600_);
  and g_101710_(_008571_, _008599_, _008602_);
  or g_101711_(_008428_, _008600_, _008603_);
  and g_101712_(_008445_, _008602_, _008604_);
  or g_101713_(_008570_, _008603_, _008605_);
  and g_101714_(_008442_, _008604_, _008606_);
  or g_101715_(_008443_, _008605_, _008607_);
  and g_101716_(_008563_, _008606_, _008608_);
  or g_101717_(_008564_, _008607_, _008609_);
  and g_101718_(_008598_, _008609_, _008610_);
  or g_101719_(_008597_, _008608_, _008611_);
  or g_101720_(_008409_, _008610_, _008613_);
  not g_101721_(_008613_, _008614_);
  and g_101722_(_008451_, _008610_, _008615_);
  not g_101723_(_008615_, _008616_);
  and g_101724_(_008613_, _008616_, _008617_);
  or g_101725_(_008614_, _008615_, _008618_);
  and g_101726_(_003149_, _008617_, _008619_);
  or g_101727_(_003150_, _008618_, _008620_);
  and g_101728_(_003561_, _008620_, _008621_);
  or g_101729_(_003560_, _008619_, _008622_);
  and g_101730_(_003150_, _008618_, _008624_);
  or g_101731_(_003149_, _008617_, _008625_);
  and g_101732_(out[425], _003144_, _008626_);
  xor g_101733_(out[425], _003144_, _008627_);
  or g_101734_(_003147_, _008626_, _008628_);
  and g_101735_(_008488_, _008611_, _008629_);
  and g_101736_(_008482_, _008610_, _008630_);
  or g_101737_(_008629_, _008630_, _008631_);
  not g_101738_(_008631_, _008632_);
  and g_101739_(_008627_, _008631_, _008633_);
  or g_101740_(_008628_, _008632_, _008635_);
  and g_101741_(_008628_, _008632_, _008636_);
  or g_101742_(_008627_, _008631_, _008637_);
  and g_101743_(_008635_, _008637_, _008638_);
  xor g_101744_(out[424], _003143_, _008639_);
  xor g_101745_(_053951_, _003143_, _008640_);
  and g_101746_(_008470_, _008610_, _008641_);
  and g_101747_(_008476_, _008611_, _008642_);
  or g_101748_(_008641_, _008642_, _008643_);
  and g_101749_(_008639_, _008643_, _008644_);
  or g_101750_(_008639_, _008643_, _008646_);
  not g_101751_(_008646_, _008647_);
  xor g_101752_(_008639_, _008643_, _008648_);
  or g_101753_(_008633_, _008644_, _008649_);
  or g_101754_(_008636_, _008647_, _008650_);
  and g_101755_(_008638_, _008648_, _008651_);
  or g_101756_(_008649_, _008650_, _008652_);
  xor g_101757_(out[422], _003141_, _008653_);
  not g_101758_(_008653_, _008654_);
  and g_101759_(_008506_, _008610_, _008655_);
  not g_101760_(_008655_, _008657_);
  or g_101761_(_008509_, _008610_, _008658_);
  not g_101762_(_008658_, _008659_);
  and g_101763_(_008657_, _008658_, _008660_);
  or g_101764_(_008655_, _008659_, _008661_);
  and g_101765_(_008654_, _008660_, _008662_);
  or g_101766_(_008653_, _008661_, _008663_);
  xor g_101767_(out[423], _003142_, _008664_);
  xor g_101768_(_053940_, _003142_, _008665_);
  and g_101769_(_008511_, _008610_, _008666_);
  not g_101770_(_008666_, _008668_);
  or g_101771_(_008516_, _008610_, _008669_);
  not g_101772_(_008669_, _008670_);
  and g_101773_(_008668_, _008669_, _008671_);
  or g_101774_(_008666_, _008670_, _008672_);
  and g_101775_(_008664_, _008671_, _008673_);
  or g_101776_(_008665_, _008672_, _008674_);
  and g_101777_(_008663_, _008674_, _008675_);
  or g_101778_(_008662_, _008673_, _008676_);
  and g_101779_(_008653_, _008661_, _008677_);
  and g_101780_(_008665_, _008672_, _008679_);
  or g_101781_(_008677_, _008679_, _008680_);
  not g_101782_(_008680_, _008681_);
  and g_101783_(_008675_, _008681_, _008682_);
  or g_101784_(_008676_, _008680_, _008683_);
  or g_101785_(_014970_, _053270_, _008684_);
  not g_101786_(_008684_, _008685_);
  and g_101787_(_003140_, _008684_, _008686_);
  or g_101788_(_003139_, _008685_, _008687_);
  and g_101789_(_008537_, _008611_, _008688_);
  and g_101790_(_008530_, _008610_, _008690_);
  or g_101791_(_008688_, _008690_, _008691_);
  or g_101792_(_008686_, _008691_, _008692_);
  not g_101793_(_008692_, _008693_);
  xor g_101794_(out[421], _003139_, _008694_);
  xor g_101795_(_053962_, _003139_, _008695_);
  and g_101796_(_008541_, _008610_, _008696_);
  and g_101797_(_008548_, _008611_, _008697_);
  or g_101798_(_008696_, _008697_, _008698_);
  or g_101799_(_008694_, _008698_, _008699_);
  not g_101800_(_008699_, _008701_);
  and g_101801_(_008692_, _008699_, _008702_);
  or g_101802_(_008693_, _008701_, _008703_);
  and g_101803_(_008694_, _008698_, _008704_);
  and g_101804_(_008686_, _008691_, _008705_);
  or g_101805_(_008704_, _008705_, _008706_);
  not g_101806_(_008706_, _008707_);
  and g_101807_(_008702_, _008707_, _008708_);
  or g_101808_(_008703_, _008706_, _008709_);
  and g_101809_(_008682_, _008708_, _008710_);
  or g_101810_(_008683_, _008709_, _008712_);
  and g_101811_(out[401], _008610_, _008713_);
  not g_101812_(_008713_, _008714_);
  or g_101813_(_008432_, _008610_, _008715_);
  not g_101814_(_008715_, _008716_);
  and g_101815_(_008714_, _008715_, _008717_);
  or g_101816_(_008713_, _008716_, _008718_);
  and g_101817_(out[417], _008717_, _008719_);
  or g_101818_(_054017_, _008718_, _008720_);
  and g_101819_(_053010_, _008610_, _008721_);
  and g_101820_(_008417_, _008611_, _008723_);
  or g_101821_(_008721_, _008723_, _008724_);
  or g_101822_(_053272_, _008724_, _008725_);
  xor g_101823_(_053272_, _008724_, _008726_);
  xor g_101824_(_053271_, _008724_, _008727_);
  xor g_101825_(out[419], _053270_, _008728_);
  xor g_101826_(_053984_, _053270_, _008729_);
  and g_101827_(_008419_, _008610_, _008730_);
  and g_101828_(_008427_, _008611_, _008731_);
  or g_101829_(_008730_, _008731_, _008732_);
  or g_101830_(_008729_, _008732_, _008734_);
  and g_101831_(_008729_, _008732_, _008735_);
  xor g_101832_(_008729_, _008732_, _008736_);
  xor g_101833_(_008728_, _008732_, _008737_);
  and g_101834_(_008726_, _008736_, _008738_);
  or g_101835_(_008727_, _008737_, _008739_);
  and g_101836_(_008719_, _008738_, _008740_);
  or g_101837_(_008720_, _008739_, _008741_);
  and g_101838_(out[400], _008610_, _008742_);
  not g_101839_(_008742_, _008743_);
  or g_101840_(_008437_, _008610_, _008745_);
  not g_101841_(_008745_, _008746_);
  and g_101842_(_008743_, _008745_, _008747_);
  or g_101843_(_008742_, _008746_, _008748_);
  and g_101844_(out[416], _008747_, _008749_);
  or g_101845_(_004740_, _008748_, _008750_);
  xor g_101846_(out[417], _008717_, _008751_);
  xor g_101847_(_054017_, _008717_, _008752_);
  and g_101848_(_008750_, _008751_, _008753_);
  or g_101849_(_008749_, _008752_, _008754_);
  and g_101850_(_008738_, _008753_, _008756_);
  or g_101851_(_008739_, _008754_, _008757_);
  and g_101852_(_008725_, _008734_, _008758_);
  or g_101853_(_008735_, _008758_, _008759_);
  not g_101854_(_008759_, _008760_);
  and g_101855_(_008741_, _008759_, _008761_);
  or g_101856_(_008740_, _008760_, _008762_);
  and g_101857_(_008757_, _008761_, _008763_);
  or g_101858_(_008756_, _008762_, _008764_);
  and g_101859_(_008710_, _008764_, _008765_);
  or g_101860_(_008712_, _008763_, _008767_);
  or g_101861_(_008702_, _008704_, _008768_);
  not g_101862_(_008768_, _008769_);
  and g_101863_(_008682_, _008769_, _008770_);
  or g_101864_(_008675_, _008679_, _008771_);
  not g_101865_(_008771_, _008772_);
  or g_101866_(_008770_, _008772_, _008773_);
  not g_101867_(_008773_, _008774_);
  and g_101868_(_008767_, _008774_, _008775_);
  or g_101869_(_008765_, _008773_, _008776_);
  and g_101870_(_008651_, _008776_, _008778_);
  or g_101871_(_008652_, _008775_, _008779_);
  and g_101872_(_008637_, _008647_, _008780_);
  or g_101873_(_008636_, _008646_, _008781_);
  or g_101874_(_008633_, _008780_, _008782_);
  and g_101875_(_008635_, _008781_, _008783_);
  and g_101876_(_008779_, _008783_, _008784_);
  or g_101877_(_008778_, _008782_, _008785_);
  and g_101878_(_008625_, _008785_, _008786_);
  or g_101879_(_008624_, _008784_, _008787_);
  and g_101880_(_008621_, _008787_, _008789_);
  or g_101881_(_008622_, _008786_, _008790_);
  and g_101882_(_003557_, _003558_, _008791_);
  or g_101883_(_003556_, _003559_, _008792_);
  or g_101884_(out[416], _008747_, _008793_);
  and g_101885_(_008625_, _008793_, _008794_);
  and g_101886_(_008621_, _008794_, _008795_);
  and g_101887_(_008651_, _008795_, _008796_);
  and g_101888_(_008710_, _008796_, _008797_);
  not g_101889_(_008797_, _008798_);
  and g_101890_(_008756_, _008797_, _008800_);
  or g_101891_(_008757_, _008798_, _008801_);
  and g_101892_(_008792_, _008801_, _008802_);
  or g_101893_(_008791_, _008800_, _008803_);
  and g_101894_(_008790_, _008802_, _008804_);
  or g_101895_(_008789_, _008803_, _008805_);
  and g_101896_(_003149_, _008804_, _008806_);
  or g_101897_(_003150_, _008805_, _008807_);
  and g_101898_(_008618_, _008805_, _008808_);
  not g_101899_(_008808_, _008809_);
  and g_101900_(_008807_, _008809_, _008811_);
  or g_101901_(_008806_, _008808_, _008812_);
  or g_101902_(out[435], _053386_, _008813_);
  not g_101903_(_008813_, _008814_);
  and g_101904_(out[436], _008813_, _008815_);
  or g_101905_(_054094_, _008814_, _008816_);
  and g_101906_(out[437], _008815_, _008817_);
  and g_101907_(out[438], _008817_, _008818_);
  or g_101908_(out[439], _008818_, _008819_);
  and g_101909_(out[440], _008819_, _008820_);
  or g_101910_(out[441], _008820_, _008822_);
  not g_101911_(_008822_, _008823_);
  or g_101912_(out[442], _008822_, _008824_);
  xor g_101913_(out[442], _008822_, _008825_);
  xor g_101914_(_004784_, _008822_, _008826_);
  and g_101915_(_008811_, _008825_, _008827_);
  or g_101916_(_008812_, _008826_, _008828_);
  and g_101917_(_003556_, _003558_, _008829_);
  or g_101918_(_003557_, _003559_, _008830_);
  xor g_101919_(out[443], _008824_, _008831_);
  xor g_101920_(_004762_, _008824_, _008833_);
  and g_101921_(_008829_, _008833_, _008834_);
  or g_101922_(_008830_, _008831_, _008835_);
  and g_101923_(_008828_, _008835_, _008836_);
  or g_101924_(_008827_, _008834_, _008837_);
  or g_101925_(_008829_, _008833_, _008838_);
  or g_101926_(_008811_, _008825_, _008839_);
  and g_101927_(_008838_, _008839_, _008840_);
  not g_101928_(_008840_, _008841_);
  and g_101929_(_008836_, _008840_, _008842_);
  or g_101930_(_008837_, _008841_, _008844_);
  xor g_101931_(out[440], _008819_, _008845_);
  xor g_101932_(_054050_, _008819_, _008846_);
  and g_101933_(_008643_, _008805_, _008847_);
  and g_101934_(_008640_, _008804_, _008848_);
  or g_101935_(_008847_, _008848_, _008849_);
  or g_101936_(_008845_, _008849_, _008850_);
  not g_101937_(_008850_, _008851_);
  xor g_101938_(_008845_, _008849_, _008852_);
  and g_101939_(out[441], _008820_, _008853_);
  xor g_101940_(out[441], _008820_, _008855_);
  or g_101941_(_008823_, _008853_, _008856_);
  and g_101942_(_008631_, _008805_, _008857_);
  and g_101943_(_008628_, _008804_, _008858_);
  or g_101944_(_008857_, _008858_, _008859_);
  and g_101945_(_008855_, _008859_, _008860_);
  or g_101946_(_008855_, _008859_, _008861_);
  xor g_101947_(_008855_, _008859_, _008862_);
  and g_101948_(_008852_, _008862_, _008863_);
  not g_101949_(_008863_, _008864_);
  and g_101950_(_008842_, _008863_, _008866_);
  or g_101951_(_008844_, _008864_, _008867_);
  xor g_101952_(out[438], _008817_, _008868_);
  not g_101953_(_008868_, _008869_);
  and g_101954_(_008654_, _008804_, _008870_);
  and g_101955_(_008661_, _008805_, _008871_);
  or g_101956_(_008870_, _008871_, _008872_);
  not g_101957_(_008872_, _008873_);
  or g_101958_(_008868_, _008872_, _008874_);
  xor g_101959_(_008868_, _008872_, _008875_);
  xor g_101960_(_008869_, _008872_, _008877_);
  xor g_101961_(out[439], _008818_, _008878_);
  xor g_101962_(_054039_, _008818_, _008879_);
  and g_101963_(_008664_, _008804_, _008880_);
  and g_101964_(_008672_, _008805_, _008881_);
  or g_101965_(_008880_, _008881_, _008882_);
  or g_101966_(_008879_, _008882_, _008883_);
  and g_101967_(_008879_, _008882_, _008884_);
  xor g_101968_(_008879_, _008882_, _008885_);
  xor g_101969_(_008878_, _008882_, _008886_);
  and g_101970_(_008875_, _008885_, _008888_);
  or g_101971_(_008877_, _008886_, _008889_);
  or g_101972_(_015124_, _053386_, _008890_);
  not g_101973_(_008890_, _008891_);
  and g_101974_(_008816_, _008890_, _008892_);
  or g_101975_(_008815_, _008891_, _008893_);
  and g_101976_(_008691_, _008805_, _008894_);
  and g_101977_(_008687_, _008804_, _008895_);
  or g_101978_(_008894_, _008895_, _008896_);
  or g_101979_(_008892_, _008896_, _008897_);
  xor g_101980_(out[437], _008815_, _008899_);
  xor g_101981_(_054061_, _008815_, _008900_);
  and g_101982_(_008695_, _008804_, _008901_);
  and g_101983_(_008698_, _008805_, _008902_);
  or g_101984_(_008901_, _008902_, _008903_);
  or g_101985_(_008899_, _008903_, _008904_);
  and g_101986_(_008897_, _008904_, _008905_);
  and g_101987_(_008899_, _008903_, _008906_);
  and g_101988_(_008892_, _008896_, _008907_);
  or g_101989_(_008906_, _008907_, _008908_);
  not g_101990_(_008908_, _008910_);
  and g_101991_(_008905_, _008910_, _008911_);
  and g_101992_(_008888_, _008911_, _008912_);
  and g_101993_(_008866_, _008912_, _008913_);
  and g_101994_(_008728_, _008804_, _008914_);
  and g_101995_(_008732_, _008805_, _008915_);
  or g_101996_(_008914_, _008915_, _008916_);
  not g_101997_(_008916_, _008917_);
  xor g_101998_(out[435], _053386_, _008918_);
  xor g_101999_(_054083_, _053386_, _008919_);
  and g_102000_(_008917_, _008918_, _008921_);
  not g_102001_(_008921_, _008922_);
  or g_102002_(_008917_, _008918_, _008923_);
  and g_102003_(_053271_, _008804_, _008924_);
  and g_102004_(_008724_, _008805_, _008925_);
  or g_102005_(_008924_, _008925_, _008926_);
  not g_102006_(_008926_, _008927_);
  and g_102007_(_053387_, _008927_, _008928_);
  and g_102008_(_008923_, _008928_, _008929_);
  or g_102009_(_008921_, _008929_, _008930_);
  or g_102010_(_054017_, _008805_, _008932_);
  or g_102011_(_008717_, _008804_, _008933_);
  and g_102012_(_008932_, _008933_, _008934_);
  not g_102013_(_008934_, _008935_);
  and g_102014_(out[433], _008934_, _008936_);
  or g_102015_(_004740_, _008805_, _008937_);
  or g_102016_(_008747_, _008804_, _008938_);
  and g_102017_(_008937_, _008938_, _008939_);
  and g_102018_(out[432], _008939_, _008940_);
  not g_102019_(_008940_, _008941_);
  xor g_102020_(out[433], _008934_, _008943_);
  and g_102021_(_008941_, _008943_, _008944_);
  or g_102022_(_008936_, _008944_, _008945_);
  xor g_102023_(_053388_, _008926_, _008946_);
  and g_102024_(_008923_, _008946_, _008947_);
  and g_102025_(_008945_, _008947_, _008948_);
  or g_102026_(_008930_, _008948_, _008949_);
  and g_102027_(_008913_, _008949_, _008950_);
  or g_102028_(_008905_, _008906_, _008951_);
  not g_102029_(_008951_, _008952_);
  and g_102030_(_008888_, _008952_, _008954_);
  or g_102031_(_008889_, _008951_, _008955_);
  or g_102032_(_008874_, _008884_, _008956_);
  and g_102033_(_008883_, _008956_, _008957_);
  not g_102034_(_008957_, _008958_);
  and g_102035_(_008955_, _008957_, _008959_);
  or g_102036_(_008954_, _008958_, _008960_);
  and g_102037_(_008866_, _008960_, _008961_);
  or g_102038_(_008867_, _008959_, _008962_);
  and g_102039_(_008837_, _008838_, _008963_);
  or g_102040_(_008851_, _008860_, _008965_);
  and g_102041_(_008861_, _008965_, _008966_);
  not g_102042_(_008966_, _008967_);
  and g_102043_(_008842_, _008966_, _008968_);
  or g_102044_(_008844_, _008967_, _008969_);
  and g_102045_(_008962_, _008969_, _008970_);
  or g_102046_(_008961_, _008968_, _008971_);
  or g_102047_(_008950_, _008963_, _008972_);
  not g_102048_(_008972_, _008973_);
  and g_102049_(_008970_, _008973_, _008974_);
  or g_102050_(_008971_, _008972_, _008976_);
  or g_102051_(out[432], _008939_, _008977_);
  and g_102052_(_008922_, _008977_, _008978_);
  and g_102053_(_008944_, _008978_, _008979_);
  and g_102054_(_008947_, _008979_, _008980_);
  and g_102055_(_008913_, _008980_, _008981_);
  not g_102056_(_008981_, _008982_);
  and g_102057_(_008976_, _008982_, _008983_);
  or g_102058_(_008974_, _008981_, _008984_);
  and g_102059_(_008812_, _008984_, _008985_);
  or g_102060_(_008811_, _008983_, _008987_);
  or g_102061_(_008826_, _008984_, _008988_);
  not g_102062_(_008988_, _008989_);
  and g_102063_(_008987_, _008988_, _008990_);
  or g_102064_(_008985_, _008989_, _008991_);
  and g_102065_(_053387_, _008983_, _008992_);
  and g_102066_(_008926_, _008984_, _008993_);
  or g_102067_(_008992_, _008993_, _008994_);
  or g_102068_(out[451], _053560_, _008995_);
  not g_102069_(_008995_, _008996_);
  xor g_102070_(out[451], _053560_, _008998_);
  xor g_102071_(_054182_, _053560_, _008999_);
  and g_102072_(_008916_, _008984_, _009000_);
  and g_102073_(_008918_, _008983_, _009001_);
  or g_102074_(_009000_, _009001_, _009002_);
  or g_102075_(_008999_, _009002_, _009003_);
  or g_102076_(_053562_, _008994_, _009004_);
  and g_102077_(_008999_, _009002_, _009005_);
  xor g_102078_(_053562_, _008994_, _009006_);
  xor g_102079_(_053561_, _008994_, _009007_);
  xor g_102080_(_008999_, _009002_, _009009_);
  xor g_102081_(_008998_, _009002_, _009010_);
  and g_102082_(_009006_, _009009_, _009011_);
  or g_102083_(_009007_, _009010_, _009012_);
  or g_102084_(_054116_, _008984_, _009013_);
  not g_102085_(_009013_, _009014_);
  and g_102086_(_008935_, _008984_, _009015_);
  or g_102087_(_008934_, _008983_, _009016_);
  and g_102088_(_009013_, _009016_, _009017_);
  or g_102089_(_009014_, _009015_, _009018_);
  and g_102090_(out[449], _009017_, _009020_);
  not g_102091_(_009020_, _009021_);
  or g_102092_(_004773_, _008984_, _009022_);
  or g_102093_(_008939_, _008983_, _009023_);
  and g_102094_(_009022_, _009023_, _009024_);
  and g_102095_(out[448], _009024_, _009025_);
  not g_102096_(_009025_, _009026_);
  xor g_102097_(out[449], _009017_, _009027_);
  xor g_102098_(_054215_, _009017_, _009028_);
  and g_102099_(_009026_, _009027_, _009029_);
  or g_102100_(_009025_, _009028_, _009031_);
  and g_102101_(_009021_, _009031_, _009032_);
  or g_102102_(_009012_, _009032_, _009033_);
  or g_102103_(_009004_, _009005_, _009034_);
  and g_102104_(_009003_, _009034_, _009035_);
  and g_102105_(_009033_, _009035_, _009036_);
  and g_102106_(out[452], _008995_, _009037_);
  or g_102107_(_054193_, _008996_, _009038_);
  and g_102108_(out[453], _009037_, _009039_);
  and g_102109_(out[454], _009039_, _009040_);
  or g_102110_(out[455], _009040_, _009042_);
  and g_102111_(out[456], _009042_, _009043_);
  or g_102112_(out[457], _009043_, _009044_);
  or g_102113_(out[458], _009044_, _009045_);
  xor g_102114_(out[458], _009044_, _009046_);
  not g_102115_(_009046_, _009047_);
  and g_102116_(_008990_, _009046_, _009048_);
  or g_102117_(_008991_, _009047_, _009049_);
  and g_102118_(_008829_, _008831_, _009050_);
  or g_102119_(_008830_, _008833_, _009051_);
  xor g_102120_(out[459], _009045_, _009053_);
  not g_102121_(_009053_, _009054_);
  and g_102122_(_009050_, _009054_, _009055_);
  or g_102123_(_009051_, _009053_, _009056_);
  and g_102124_(_009049_, _009056_, _009057_);
  or g_102125_(_009048_, _009055_, _009058_);
  and g_102126_(_009051_, _009053_, _009059_);
  and g_102127_(_008991_, _009047_, _009060_);
  or g_102128_(_009059_, _009060_, _009061_);
  not g_102129_(_009061_, _009062_);
  and g_102130_(_009057_, _009062_, _009064_);
  or g_102131_(_009058_, _009061_, _009065_);
  xor g_102132_(out[456], _009042_, _009066_);
  xor g_102133_(_054149_, _009042_, _009067_);
  or g_102134_(_008845_, _008984_, _009068_);
  not g_102135_(_009068_, _009069_);
  and g_102136_(_008849_, _008984_, _009070_);
  not g_102137_(_009070_, _009071_);
  and g_102138_(_009068_, _009071_, _009072_);
  or g_102139_(_009069_, _009070_, _009073_);
  and g_102140_(_009066_, _009073_, _009075_);
  or g_102141_(_009067_, _009072_, _009076_);
  and g_102142_(out[457], _009043_, _009077_);
  xor g_102143_(out[457], _009043_, _009078_);
  xor g_102144_(_054226_, _009043_, _009079_);
  and g_102145_(_008859_, _008984_, _009080_);
  not g_102146_(_009080_, _009081_);
  or g_102147_(_008855_, _008984_, _009082_);
  not g_102148_(_009082_, _009083_);
  and g_102149_(_009081_, _009082_, _009084_);
  or g_102150_(_009080_, _009083_, _009086_);
  and g_102151_(_009079_, _009084_, _009087_);
  or g_102152_(_009078_, _009086_, _009088_);
  and g_102153_(_009076_, _009088_, _009089_);
  or g_102154_(_009075_, _009087_, _009090_);
  and g_102155_(_009078_, _009086_, _009091_);
  and g_102156_(_009067_, _009072_, _009092_);
  or g_102157_(_009091_, _009092_, _009093_);
  not g_102158_(_009093_, _009094_);
  and g_102159_(_009089_, _009094_, _009095_);
  or g_102160_(_009090_, _009093_, _009097_);
  and g_102161_(_009064_, _009095_, _009098_);
  or g_102162_(_009065_, _009097_, _009099_);
  xor g_102163_(out[455], _009040_, _009100_);
  xor g_102164_(_054138_, _009040_, _009101_);
  and g_102165_(_008878_, _008983_, _009102_);
  and g_102166_(_008882_, _008984_, _009103_);
  or g_102167_(_009102_, _009103_, _009104_);
  or g_102168_(_009101_, _009104_, _009105_);
  and g_102169_(_009101_, _009104_, _009106_);
  xor g_102170_(_009101_, _009104_, _009108_);
  xor g_102171_(_009100_, _009104_, _009109_);
  xor g_102172_(out[454], _009039_, _009110_);
  xor g_102173_(_054171_, _009039_, _009111_);
  or g_102174_(_008868_, _008984_, _009112_);
  or g_102175_(_008873_, _008983_, _009113_);
  and g_102176_(_009112_, _009113_, _009114_);
  not g_102177_(_009114_, _009115_);
  or g_102178_(_009110_, _009115_, _009116_);
  xor g_102179_(_009111_, _009114_, _009117_);
  xor g_102180_(_009110_, _009114_, _009119_);
  and g_102181_(_009108_, _009117_, _009120_);
  or g_102182_(_009109_, _009119_, _009121_);
  or g_102183_(_015278_, _053560_, _009122_);
  not g_102184_(_009122_, _009123_);
  and g_102185_(_009038_, _009122_, _009124_);
  or g_102186_(_009037_, _009123_, _009125_);
  and g_102187_(_008896_, _008984_, _009126_);
  and g_102188_(_008893_, _008983_, _009127_);
  or g_102189_(_009126_, _009127_, _009128_);
  or g_102190_(_009124_, _009128_, _009130_);
  not g_102191_(_009130_, _009131_);
  xor g_102192_(out[453], _009037_, _009132_);
  xor g_102193_(_054160_, _009037_, _009133_);
  and g_102194_(_008900_, _008983_, _009134_);
  and g_102195_(_008903_, _008984_, _009135_);
  or g_102196_(_009134_, _009135_, _009136_);
  or g_102197_(_009132_, _009136_, _009137_);
  not g_102198_(_009137_, _009138_);
  and g_102199_(_009130_, _009137_, _009139_);
  or g_102200_(_009131_, _009138_, _009141_);
  and g_102201_(_009132_, _009136_, _009142_);
  and g_102202_(_009124_, _009128_, _009143_);
  or g_102203_(_009142_, _009143_, _009144_);
  not g_102204_(_009144_, _009145_);
  and g_102205_(_009139_, _009145_, _009146_);
  or g_102206_(_009141_, _009144_, _009147_);
  and g_102207_(_009120_, _009146_, _009148_);
  or g_102208_(_009121_, _009147_, _009149_);
  and g_102209_(_009098_, _009148_, _009150_);
  or g_102210_(_009099_, _009149_, _009152_);
  or g_102211_(_009036_, _009152_, _009153_);
  or g_102212_(_009121_, _009139_, _009154_);
  or g_102213_(_009142_, _009154_, _009155_);
  or g_102214_(_009106_, _009116_, _009156_);
  and g_102215_(_009105_, _009156_, _009157_);
  and g_102216_(_009155_, _009157_, _009158_);
  or g_102217_(_009099_, _009158_, _009159_);
  or g_102218_(_009057_, _009059_, _009160_);
  and g_102219_(_009088_, _009093_, _009161_);
  and g_102220_(_009064_, _009161_, _009163_);
  not g_102221_(_009163_, _009164_);
  and g_102222_(_009160_, _009164_, _009165_);
  and g_102223_(_009159_, _009165_, _009166_);
  and g_102224_(_009153_, _009166_, _009167_);
  or g_102225_(out[448], _009024_, _009168_);
  and g_102226_(_009011_, _009168_, _009169_);
  and g_102227_(_009029_, _009169_, _009170_);
  and g_102228_(_009150_, _009170_, _009171_);
  or g_102229_(_009167_, _009171_, _009172_);
  not g_102230_(_009172_, _009174_);
  and g_102231_(_008991_, _009172_, _009175_);
  and g_102232_(_009046_, _009174_, _009176_);
  or g_102233_(_009175_, _009176_, _009177_);
  not g_102234_(_009177_, _009178_);
  and g_102235_(_003135_, _009178_, _009179_);
  or g_102236_(_003136_, _009177_, _009180_);
  and g_102237_(_009050_, _009053_, _009181_);
  not g_102238_(_009181_, _009182_);
  xor g_102239_(out[475], _003133_, _009183_);
  not g_102240_(_009183_, _009185_);
  and g_102241_(_009181_, _009185_, _009186_);
  or g_102242_(_009182_, _009183_, _009187_);
  and g_102243_(_009180_, _009187_, _009188_);
  or g_102244_(_009179_, _009186_, _009189_);
  and g_102245_(out[473], _003131_, _009190_);
  xor g_102246_(out[473], _003131_, _009191_);
  xor g_102247_(_054325_, _003131_, _009192_);
  and g_102248_(_009086_, _009172_, _009193_);
  not g_102249_(_009193_, _009194_);
  or g_102250_(_009078_, _009172_, _009196_);
  not g_102251_(_009196_, _009197_);
  and g_102252_(_009194_, _009196_, _009198_);
  or g_102253_(_009193_, _009197_, _009199_);
  and g_102254_(_009192_, _009198_, _009200_);
  or g_102255_(_009191_, _009199_, _009201_);
  and g_102256_(_009182_, _009183_, _009202_);
  or g_102257_(_009181_, _009185_, _009203_);
  xor g_102258_(out[472], _003128_, _009204_);
  xor g_102259_(_054248_, _003128_, _009205_);
  or g_102260_(_009066_, _009172_, _009207_);
  or g_102261_(_009072_, _009174_, _009208_);
  and g_102262_(_009207_, _009208_, _009209_);
  not g_102263_(_009209_, _009210_);
  and g_102264_(_009204_, _009210_, _009211_);
  or g_102265_(_009205_, _009209_, _009212_);
  and g_102266_(_009191_, _009199_, _009213_);
  or g_102267_(_009192_, _009198_, _009214_);
  and g_102268_(_009205_, _009209_, _009215_);
  or g_102269_(_009204_, _009210_, _009216_);
  xor g_102270_(_003136_, _009177_, _009218_);
  xor g_102271_(_003135_, _009177_, _009219_);
  and g_102272_(_009187_, _009203_, _009220_);
  or g_102273_(_009186_, _009202_, _009221_);
  and g_102274_(_009218_, _009220_, _009222_);
  or g_102275_(_009219_, _009221_, _009223_);
  and g_102276_(_009212_, _009214_, _009224_);
  or g_102277_(_009211_, _009213_, _009225_);
  and g_102278_(_009201_, _009216_, _009226_);
  or g_102279_(_009200_, _009215_, _009227_);
  and g_102280_(_009224_, _009226_, _009229_);
  or g_102281_(_009225_, _009227_, _009230_);
  and g_102282_(_009222_, _009229_, _009231_);
  or g_102283_(_009223_, _009230_, _009232_);
  xor g_102284_(out[470], _003126_, _009233_);
  or g_102285_(_009110_, _009172_, _009234_);
  or g_102286_(_009114_, _009174_, _009235_);
  and g_102287_(_009234_, _009235_, _009236_);
  not g_102288_(_009236_, _009237_);
  or g_102289_(_009233_, _009237_, _009238_);
  xor g_102290_(_009233_, _009237_, _009240_);
  xor g_102291_(_009233_, _009236_, _009241_);
  and g_102292_(_009100_, _009174_, _009242_);
  and g_102293_(_009104_, _009172_, _009243_);
  or g_102294_(_009242_, _009243_, _009244_);
  and g_102295_(_003130_, _009244_, _009245_);
  or g_102296_(_003130_, _009244_, _009246_);
  xor g_102297_(_003130_, _009244_, _009247_);
  xor g_102298_(_003129_, _009244_, _009248_);
  and g_102299_(_009240_, _009247_, _009249_);
  or g_102300_(_009241_, _009248_, _009251_);
  or g_102301_(_015432_, _053880_, _009252_);
  not g_102302_(_009252_, _009253_);
  and g_102303_(_003125_, _009252_, _009254_);
  or g_102304_(_003124_, _009253_, _009255_);
  and g_102305_(_009128_, _009172_, _009256_);
  not g_102306_(_009256_, _009257_);
  or g_102307_(_009124_, _009172_, _009258_);
  and g_102308_(_009257_, _009258_, _009259_);
  not g_102309_(_009259_, _009260_);
  and g_102310_(_009255_, _009259_, _009262_);
  or g_102311_(_009254_, _009260_, _009263_);
  xor g_102312_(out[469], _003124_, _009264_);
  xor g_102313_(_054259_, _003124_, _009265_);
  or g_102314_(_009132_, _009172_, _009266_);
  not g_102315_(_009266_, _009267_);
  and g_102316_(_009136_, _009172_, _009268_);
  not g_102317_(_009268_, _009269_);
  and g_102318_(_009266_, _009269_, _009270_);
  or g_102319_(_009267_, _009268_, _009271_);
  and g_102320_(_009265_, _009270_, _009273_);
  or g_102321_(_009264_, _009271_, _009274_);
  and g_102322_(_009263_, _009274_, _009275_);
  or g_102323_(_009262_, _009273_, _009276_);
  and g_102324_(_009264_, _009271_, _009277_);
  or g_102325_(_009265_, _009270_, _009278_);
  and g_102326_(_009254_, _009260_, _009279_);
  or g_102327_(_009255_, _009259_, _009280_);
  and g_102328_(_009278_, _009280_, _009281_);
  or g_102329_(_009276_, _009279_, _009282_);
  and g_102330_(_009275_, _009281_, _009284_);
  or g_102331_(_009277_, _009282_, _009285_);
  and g_102332_(_009249_, _009284_, _009286_);
  or g_102333_(_009251_, _009285_, _009287_);
  and g_102334_(_009231_, _009286_, _009288_);
  or g_102335_(_009232_, _009287_, _009289_);
  xor g_102336_(out[467], _053880_, _009290_);
  xor g_102337_(_054281_, _053880_, _009291_);
  or g_102338_(_008999_, _009172_, _009292_);
  and g_102339_(_009002_, _009172_, _009293_);
  not g_102340_(_009293_, _009295_);
  and g_102341_(_009292_, _009295_, _009296_);
  not g_102342_(_009296_, _009297_);
  and g_102343_(_009290_, _009296_, _009298_);
  or g_102344_(_009291_, _009297_, _009299_);
  and g_102345_(_008994_, _009172_, _009300_);
  and g_102346_(_053561_, _009174_, _009301_);
  or g_102347_(_009300_, _009301_, _009302_);
  not g_102348_(_009302_, _009303_);
  and g_102349_(_053882_, _009302_, _009304_);
  or g_102350_(_053881_, _009303_, _009306_);
  and g_102351_(_009299_, _009306_, _009307_);
  or g_102352_(_009298_, _009304_, _009308_);
  and g_102353_(_053881_, _009303_, _009309_);
  or g_102354_(_053882_, _009302_, _009310_);
  and g_102355_(_009291_, _009297_, _009311_);
  or g_102356_(_009290_, _009296_, _009312_);
  and g_102357_(_009310_, _009312_, _009313_);
  or g_102358_(_009309_, _009311_, _009314_);
  and g_102359_(_009307_, _009313_, _009315_);
  or g_102360_(_009308_, _009314_, _009317_);
  and g_102361_(out[449], _009174_, _009318_);
  and g_102362_(_009018_, _009172_, _009319_);
  or g_102363_(_009318_, _009319_, _009320_);
  not g_102364_(_009320_, _009321_);
  and g_102365_(out[465], _009321_, _009322_);
  or g_102366_(_054314_, _009320_, _009323_);
  and g_102367_(_009024_, _009172_, _009324_);
  not g_102368_(_009324_, _009325_);
  or g_102369_(out[448], _009172_, _009326_);
  and g_102370_(_009325_, _009326_, _009328_);
  not g_102371_(_009328_, _009329_);
  and g_102372_(out[464], _009329_, _009330_);
  or g_102373_(_004839_, _009328_, _009331_);
  xor g_102374_(_054314_, _009320_, _009332_);
  xor g_102375_(out[465], _009320_, _009333_);
  and g_102376_(_009331_, _009332_, _009334_);
  or g_102377_(_009330_, _009333_, _009335_);
  and g_102378_(_009323_, _009335_, _009336_);
  or g_102379_(_009322_, _009334_, _009337_);
  and g_102380_(_009315_, _009337_, _009339_);
  or g_102381_(_009317_, _009336_, _009340_);
  and g_102382_(_009309_, _009312_, _009341_);
  or g_102383_(_009310_, _009311_, _009342_);
  and g_102384_(_009299_, _009342_, _009343_);
  or g_102385_(_009298_, _009341_, _009344_);
  and g_102386_(_009340_, _009343_, _009345_);
  or g_102387_(_009339_, _009344_, _009346_);
  and g_102388_(_009288_, _009346_, _009347_);
  or g_102389_(_009289_, _009345_, _009348_);
  or g_102390_(_009251_, _009277_, _009350_);
  or g_102391_(_009275_, _009350_, _009351_);
  or g_102392_(_009238_, _009245_, _009352_);
  and g_102393_(_009246_, _009352_, _009353_);
  and g_102394_(_009351_, _009353_, _009354_);
  or g_102395_(_009232_, _009354_, _009355_);
  not g_102396_(_009355_, _009356_);
  and g_102397_(_009189_, _009203_, _009357_);
  or g_102398_(_009188_, _009202_, _009358_);
  and g_102399_(_009348_, _009358_, _009359_);
  or g_102400_(_009347_, _009357_, _009361_);
  and g_102401_(_009201_, _009215_, _009362_);
  or g_102402_(_009200_, _009216_, _009363_);
  and g_102403_(_009214_, _009363_, _009364_);
  or g_102404_(_009213_, _009362_, _009365_);
  and g_102405_(_009222_, _009365_, _009366_);
  or g_102406_(_009223_, _009364_, _009367_);
  and g_102407_(_009355_, _009367_, _009368_);
  or g_102408_(_009356_, _009366_, _009369_);
  and g_102409_(_009359_, _009368_, _009370_);
  or g_102410_(_009361_, _009369_, _009372_);
  and g_102411_(_004839_, _009328_, _009373_);
  or g_102412_(_009317_, _009373_, _009374_);
  or g_102413_(_009335_, _009374_, _009375_);
  or g_102414_(_009289_, _009375_, _009376_);
  not g_102415_(_009376_, _009377_);
  and g_102416_(_009372_, _009376_, _009378_);
  or g_102417_(_009370_, _009377_, _009379_);
  and g_102418_(_003129_, _009378_, _009380_);
  and g_102419_(_009244_, _009379_, _009381_);
  or g_102420_(_009380_, _009381_, _009383_);
  or g_102421_(out[947], _002904_, _009384_);
  and g_102422_(out[948], _009384_, _009385_);
  and g_102423_(out[949], _009385_, _009386_);
  and g_102424_(out[950], _009386_, _009387_);
  or g_102425_(out[951], _009387_, _009388_);
  xor g_102426_(out[951], _009387_, _009389_);
  xor g_102427_(_002188_, _009387_, _009390_);
  and g_102428_(out[952], _009388_, _009391_);
  or g_102429_(out[953], _009391_, _009392_);
  not g_102430_(_009392_, _009394_);
  or g_102431_(out[954], _009392_, _009395_);
  xor g_102432_(out[955], _009395_, _009396_);
  not g_102433_(_009396_, _009397_);
  or g_102434_(out[931], _002719_, _009398_);
  not g_102435_(_009398_, _009399_);
  and g_102436_(out[932], _009398_, _009400_);
  or g_102437_(_002100_, _009399_, _009401_);
  and g_102438_(out[933], _009400_, _009402_);
  and g_102439_(out[934], _009402_, _009403_);
  or g_102440_(out[935], _009403_, _009405_);
  and g_102441_(out[936], _009405_, _009406_);
  or g_102442_(out[937], _009406_, _009407_);
  or g_102443_(out[938], _009407_, _009408_);
  xor g_102444_(out[939], _009408_, _009409_);
  not g_102445_(_009409_, _009410_);
  or g_102446_(out[483], _016389_, _009411_);
  and g_102447_(out[484], _009411_, _009412_);
  not g_102448_(_009412_, _009413_);
  and g_102449_(out[485], _009412_, _009414_);
  and g_102450_(out[486], _009414_, _009416_);
  or g_102451_(out[487], _009416_, _009417_);
  and g_102452_(out[488], _009417_, _009418_);
  or g_102453_(out[489], _009418_, _009419_);
  or g_102454_(out[490], _009419_, _009420_);
  xor g_102455_(out[491], _009420_, _009421_);
  xor g_102456_(_054358_, _009420_, _009422_);
  or g_102457_(out[499], _016356_, _009423_);
  and g_102458_(out[500], _009423_, _009424_);
  not g_102459_(_009424_, _009425_);
  and g_102460_(out[501], _009424_, _009427_);
  and g_102461_(out[502], _009427_, _009428_);
  or g_102462_(out[503], _009428_, _009429_);
  and g_102463_(out[504], _009429_, _009430_);
  or g_102464_(out[505], _009430_, _009431_);
  or g_102465_(out[506], _009431_, _009432_);
  xor g_102466_(out[507], _009432_, _009433_);
  xor g_102467_(_054479_, _009432_, _009434_);
  and g_102468_(_009421_, _009433_, _009435_);
  or g_102469_(_009422_, _009434_, _009436_);
  or g_102470_(out[515], _019073_, _009438_);
  not g_102471_(_009438_, _009439_);
  and g_102472_(out[516], _009438_, _009440_);
  or g_102473_(_054655_, _009439_, _009441_);
  and g_102474_(out[517], _009440_, _009442_);
  and g_102475_(out[518], _009442_, _009443_);
  or g_102476_(out[519], _009443_, _009444_);
  and g_102477_(out[520], _009444_, _009445_);
  or g_102478_(out[521], _009445_, _009446_);
  not g_102479_(_009446_, _009447_);
  or g_102480_(out[522], _009446_, _009449_);
  xor g_102481_(out[523], _009449_, _009450_);
  xor g_102482_(_054611_, _009449_, _009451_);
  and g_102483_(_009435_, _009450_, _009452_);
  or g_102484_(_009436_, _009451_, _009453_);
  or g_102485_(out[531], _020976_, _009454_);
  not g_102486_(_009454_, _009455_);
  and g_102487_(out[532], _009454_, _009456_);
  or g_102488_(_054787_, _009455_, _009457_);
  and g_102489_(out[533], _009456_, _009458_);
  and g_102490_(out[534], _009458_, _009460_);
  or g_102491_(out[535], _009460_, _009461_);
  and g_102492_(out[536], _009461_, _009462_);
  or g_102493_(out[537], _009462_, _009463_);
  not g_102494_(_009463_, _009464_);
  or g_102495_(out[538], _009463_, _009465_);
  xor g_102496_(out[539], _009465_, _009466_);
  xor g_102497_(_054743_, _009465_, _009467_);
  and g_102498_(_009452_, _009466_, _009468_);
  or g_102499_(_009453_, _009467_, _009469_);
  or g_102500_(out[547], _054003_, _009471_);
  not g_102501_(_009471_, _009472_);
  and g_102502_(out[548], _009471_, _009473_);
  or g_102503_(_054919_, _009472_, _009474_);
  and g_102504_(out[549], _009473_, _009475_);
  and g_102505_(out[550], _009475_, _009476_);
  or g_102506_(out[551], _009476_, _009477_);
  and g_102507_(out[552], _009477_, _009478_);
  or g_102508_(out[553], _009478_, _009479_);
  not g_102509_(_009479_, _009480_);
  or g_102510_(out[554], _009479_, _009482_);
  xor g_102511_(out[555], _009482_, _009483_);
  xor g_102512_(_054875_, _009482_, _009484_);
  and g_102513_(_009468_, _009483_, _009485_);
  or g_102514_(_009469_, _009484_, _009486_);
  or g_102515_(out[563], _054260_, _009487_);
  not g_102516_(_009487_, _009488_);
  and g_102517_(out[564], _009487_, _009489_);
  or g_102518_(_055051_, _009488_, _009490_);
  and g_102519_(out[565], _009489_, _009491_);
  and g_102520_(out[566], _009491_, _009493_);
  or g_102521_(out[567], _009493_, _009494_);
  and g_102522_(out[568], _009494_, _009495_);
  or g_102523_(out[569], _009495_, _009496_);
  not g_102524_(_009496_, _009497_);
  or g_102525_(out[570], _009496_, _009498_);
  xor g_102526_(out[571], _009498_, _009499_);
  xor g_102527_(_055007_, _009498_, _009500_);
  and g_102528_(_009485_, _009499_, _009501_);
  or g_102529_(_009486_, _009500_, _009502_);
  or g_102530_(out[579], _054570_, _009504_);
  not g_102531_(_009504_, _009505_);
  and g_102532_(out[580], _009504_, _009506_);
  or g_102533_(_055183_, _009505_, _009507_);
  and g_102534_(out[581], _009506_, _009508_);
  and g_102535_(out[582], _009508_, _009509_);
  or g_102536_(out[583], _009509_, _009510_);
  and g_102537_(out[584], _009510_, _009511_);
  or g_102538_(out[585], _009511_, _009512_);
  or g_102539_(out[586], _009512_, _009513_);
  xor g_102540_(out[587], _009513_, _009515_);
  not g_102541_(_009515_, _009516_);
  and g_102542_(_009501_, _009515_, _009517_);
  or g_102543_(_009502_, _009516_, _009518_);
  or g_102544_(out[595], _054791_, _009519_);
  not g_102545_(_009519_, _009520_);
  and g_102546_(out[596], _009519_, _009521_);
  or g_102547_(_055315_, _009520_, _009522_);
  and g_102548_(out[597], _009521_, _009523_);
  and g_102549_(out[598], _009523_, _009524_);
  or g_102550_(out[599], _009524_, _009526_);
  and g_102551_(out[600], _009526_, _009527_);
  or g_102552_(out[601], _009527_, _009528_);
  or g_102553_(out[602], _009528_, _009529_);
  xor g_102554_(out[603], _009529_, _009530_);
  xor g_102555_(_055271_, _009529_, _009531_);
  and g_102556_(_009517_, _009530_, _009532_);
  or g_102557_(_009518_, _009531_, _009533_);
  or g_102558_(out[611], _054977_, _009534_);
  not g_102559_(_009534_, _009535_);
  and g_102560_(out[612], _009534_, _009537_);
  or g_102561_(_055447_, _009535_, _009538_);
  and g_102562_(out[613], _009537_, _009539_);
  and g_102563_(out[614], _009539_, _009540_);
  or g_102564_(out[615], _009540_, _009541_);
  and g_102565_(out[616], _009541_, _009542_);
  or g_102566_(out[617], _009542_, _009543_);
  or g_102567_(out[618], _009543_, _009544_);
  xor g_102568_(out[619], _009544_, _009545_);
  xor g_102569_(_055403_, _009544_, _009546_);
  and g_102570_(_009532_, _009545_, _009548_);
  or g_102571_(_009533_, _009546_, _009549_);
  or g_102572_(out[627], _055090_, _009550_);
  not g_102573_(_009550_, _009551_);
  and g_102574_(out[628], _009550_, _009552_);
  or g_102575_(_055579_, _009551_, _009553_);
  and g_102576_(out[629], _009552_, _009554_);
  and g_102577_(out[630], _009554_, _009555_);
  or g_102578_(out[631], _009555_, _009556_);
  and g_102579_(out[632], _009556_, _009557_);
  or g_102580_(out[633], _009557_, _009559_);
  not g_102581_(_009559_, _009560_);
  or g_102582_(out[634], _009559_, _009561_);
  xor g_102583_(out[635], _009561_, _009562_);
  xor g_102584_(_055535_, _009561_, _009563_);
  and g_102585_(_009548_, _009562_, _009564_);
  or g_102586_(_009549_, _009563_, _009565_);
  or g_102587_(out[643], _055356_, _009566_);
  not g_102588_(_009566_, _009567_);
  and g_102589_(out[644], _009566_, _009568_);
  or g_102590_(_055711_, _009567_, _009570_);
  and g_102591_(out[645], _009568_, _009571_);
  and g_102592_(out[646], _009571_, _009572_);
  or g_102593_(out[647], _009572_, _009573_);
  and g_102594_(out[648], _009573_, _009574_);
  or g_102595_(out[649], _009574_, _009575_);
  or g_102596_(out[650], _009575_, _009576_);
  xor g_102597_(out[651], _009576_, _009577_);
  not g_102598_(_009577_, _009578_);
  and g_102599_(_009564_, _009577_, _009579_);
  or g_102600_(_009565_, _009578_, _009581_);
  or g_102601_(out[659], _055437_, _009582_);
  not g_102602_(_009582_, _009583_);
  and g_102603_(out[660], _009582_, _009584_);
  or g_102604_(_055843_, _009583_, _009585_);
  and g_102605_(out[661], _009584_, _009586_);
  and g_102606_(out[662], _009586_, _009587_);
  or g_102607_(out[663], _009587_, _009588_);
  and g_102608_(out[664], _009588_, _009589_);
  or g_102609_(out[665], _009589_, _009590_);
  or g_102610_(out[666], _009590_, _009592_);
  xor g_102611_(out[667], _009592_, _009593_);
  xor g_102612_(_055799_, _009592_, _009594_);
  and g_102613_(_009579_, _009593_, _009595_);
  or g_102614_(_009581_, _009594_, _009596_);
  or g_102615_(out[675], _055741_, _009597_);
  not g_102616_(_009597_, _009598_);
  and g_102617_(out[676], _009597_, _009599_);
  or g_102618_(_000010_, _009598_, _009600_);
  and g_102619_(out[677], _009599_, _009601_);
  and g_102620_(out[678], _009601_, _009603_);
  or g_102621_(out[679], _009603_, _009604_);
  and g_102622_(out[680], _009604_, _009605_);
  or g_102623_(out[681], _009605_, _009606_);
  or g_102624_(out[682], _009606_, _009607_);
  xor g_102625_(out[683], _009607_, _009608_);
  xor g_102626_(_055931_, _009607_, _009609_);
  and g_102627_(_009595_, _009608_, _009610_);
  or g_102628_(_009596_, _009609_, _009611_);
  or g_102629_(out[691], _055929_, _009612_);
  not g_102630_(_009612_, _009614_);
  and g_102631_(out[692], _009612_, _009615_);
  or g_102632_(_000142_, _009614_, _009616_);
  and g_102633_(out[693], _009615_, _009617_);
  and g_102634_(out[694], _009617_, _009618_);
  or g_102635_(out[695], _009618_, _009619_);
  and g_102636_(out[696], _009619_, _009620_);
  or g_102637_(out[697], _009620_, _009621_);
  not g_102638_(_009621_, _009622_);
  or g_102639_(out[698], _009621_, _009623_);
  xor g_102640_(out[699], _009623_, _009625_);
  xor g_102641_(_000098_, _009623_, _009626_);
  and g_102642_(_009610_, _009625_, _009627_);
  or g_102643_(_009611_, _009626_, _009628_);
  or g_102644_(out[707], _000140_, _009629_);
  not g_102645_(_009629_, _009630_);
  and g_102646_(out[708], _009629_, _009631_);
  or g_102647_(_000274_, _009630_, _009632_);
  and g_102648_(out[709], _009631_, _009633_);
  and g_102649_(out[710], _009633_, _009634_);
  or g_102650_(out[711], _009634_, _009636_);
  and g_102651_(out[712], _009636_, _009637_);
  or g_102652_(out[713], _009637_, _009638_);
  or g_102653_(out[714], _009638_, _009639_);
  xor g_102654_(out[715], _009639_, _009640_);
  not g_102655_(_009640_, _009641_);
  and g_102656_(_009627_, _009640_, _009642_);
  or g_102657_(_009628_, _009641_, _009643_);
  or g_102658_(out[723], _000239_, _009644_);
  not g_102659_(_009644_, _009645_);
  and g_102660_(out[724], _009644_, _009647_);
  or g_102661_(_000406_, _009645_, _009648_);
  and g_102662_(out[725], _009647_, _009649_);
  and g_102663_(out[726], _009649_, _009650_);
  or g_102664_(out[727], _009650_, _009651_);
  and g_102665_(out[728], _009651_, _009652_);
  or g_102666_(out[729], _009652_, _009653_);
  not g_102667_(_009653_, _009654_);
  or g_102668_(out[730], _009653_, _009655_);
  xor g_102669_(out[731], _009655_, _009656_);
  xor g_102670_(_000362_, _009655_, _009658_);
  and g_102671_(_009642_, _009656_, _009659_);
  or g_102672_(_009643_, _009658_, _009660_);
  or g_102673_(out[739], _000361_, _009661_);
  not g_102674_(_009661_, _009662_);
  and g_102675_(out[740], _009661_, _009663_);
  or g_102676_(_000538_, _009662_, _009664_);
  and g_102677_(out[741], _009663_, _009665_);
  and g_102678_(out[742], _009665_, _009666_);
  or g_102679_(out[743], _009666_, _009667_);
  and g_102680_(out[744], _009667_, _009669_);
  or g_102681_(out[745], _009669_, _009670_);
  or g_102682_(out[746], _009670_, _009671_);
  xor g_102683_(out[747], _009671_, _009672_);
  xor g_102684_(_000494_, _009671_, _009673_);
  and g_102685_(_009659_, _009672_, _009674_);
  or g_102686_(_009660_, _009673_, _009675_);
  or g_102687_(out[755], _000650_, _009676_);
  not g_102688_(_009676_, _009677_);
  and g_102689_(out[756], _009676_, _009678_);
  or g_102690_(_000670_, _009677_, _009680_);
  and g_102691_(out[757], _009678_, _009681_);
  and g_102692_(out[758], _009681_, _009682_);
  or g_102693_(out[759], _009682_, _009683_);
  and g_102694_(out[760], _009683_, _009684_);
  or g_102695_(out[761], _009684_, _009685_);
  not g_102696_(_009685_, _009686_);
  or g_102697_(out[762], _009685_, _009687_);
  xor g_102698_(out[763], _009687_, _009688_);
  xor g_102699_(_000626_, _009687_, _009689_);
  and g_102700_(_009674_, _009688_, _009691_);
  or g_102701_(_009675_, _009689_, _009692_);
  or g_102702_(out[771], _000827_, _009693_);
  not g_102703_(_009693_, _009694_);
  and g_102704_(out[772], _009693_, _009695_);
  or g_102705_(_000802_, _009694_, _009696_);
  and g_102706_(out[773], _009695_, _009697_);
  and g_102707_(out[774], _009697_, _009698_);
  or g_102708_(out[775], _009698_, _009699_);
  and g_102709_(out[776], _009699_, _009700_);
  or g_102710_(out[777], _009700_, _009702_);
  or g_102711_(out[778], _009702_, _009703_);
  xor g_102712_(out[779], _009703_, _009704_);
  xor g_102713_(_000758_, _009703_, _009705_);
  and g_102714_(_009691_, _009704_, _009706_);
  or g_102715_(_009692_, _009705_, _009707_);
  or g_102716_(out[787], _001009_, _009708_);
  not g_102717_(_009708_, _009709_);
  and g_102718_(out[788], _009708_, _009710_);
  or g_102719_(_000934_, _009709_, _009711_);
  and g_102720_(out[789], _009710_, _009713_);
  and g_102721_(out[790], _009713_, _009714_);
  or g_102722_(out[791], _009714_, _009715_);
  and g_102723_(out[792], _009715_, _009716_);
  or g_102724_(out[793], _009716_, _009717_);
  or g_102725_(out[794], _009717_, _009718_);
  xor g_102726_(out[795], _009718_, _009719_);
  not g_102727_(_009719_, _009720_);
  and g_102728_(_009706_, _009719_, _009721_);
  or g_102729_(_009707_, _009720_, _009722_);
  or g_102730_(out[803], _001210_, _009724_);
  not g_102731_(_009724_, _009725_);
  and g_102732_(out[804], _009724_, _009726_);
  or g_102733_(_001066_, _009725_, _009727_);
  and g_102734_(out[805], _009726_, _009728_);
  and g_102735_(out[806], _009728_, _009729_);
  or g_102736_(out[807], _009729_, _009730_);
  and g_102737_(out[808], _009730_, _009731_);
  or g_102738_(out[809], _009731_, _009732_);
  not g_102739_(_009732_, _009733_);
  or g_102740_(out[810], _009732_, _009735_);
  xor g_102741_(out[811], _009735_, _009736_);
  xor g_102742_(_001022_, _009735_, _009737_);
  and g_102743_(_009721_, _009736_, _009738_);
  or g_102744_(_009722_, _009737_, _009739_);
  or g_102745_(out[819], _001338_, _009740_);
  not g_102746_(_009740_, _009741_);
  and g_102747_(out[820], _009740_, _009742_);
  or g_102748_(_001198_, _009741_, _009743_);
  and g_102749_(out[821], _009742_, _009744_);
  and g_102750_(out[822], _009744_, _009746_);
  or g_102751_(out[823], _009746_, _009747_);
  and g_102752_(out[824], _009747_, _009748_);
  or g_102753_(out[825], _009748_, _009749_);
  not g_102754_(_009749_, _009750_);
  or g_102755_(out[826], _009749_, _009751_);
  xor g_102756_(out[827], _009751_, _009752_);
  xor g_102757_(_001154_, _009751_, _009753_);
  and g_102758_(_009738_, _009752_, _009754_);
  or g_102759_(_009739_, _009753_, _009755_);
  or g_102760_(out[835], _001514_, _009757_);
  not g_102761_(_009757_, _009758_);
  and g_102762_(out[836], _009757_, _009759_);
  or g_102763_(_001330_, _009758_, _009760_);
  and g_102764_(out[837], _009759_, _009761_);
  and g_102765_(out[838], _009761_, _009762_);
  or g_102766_(out[839], _009762_, _009763_);
  and g_102767_(out[840], _009763_, _009764_);
  or g_102768_(out[841], _009764_, _009765_);
  or g_102769_(out[842], _009765_, _009766_);
  xor g_102770_(out[843], _009766_, _009768_);
  not g_102771_(_009768_, _009769_);
  and g_102772_(_009754_, _009768_, _009770_);
  or g_102773_(_009755_, _009769_, _009771_);
  or g_102774_(out[851], _001844_, _009772_);
  not g_102775_(_009772_, _009773_);
  and g_102776_(out[852], _009772_, _009774_);
  or g_102777_(_001462_, _009773_, _009775_);
  and g_102778_(out[853], _009774_, _009776_);
  and g_102779_(out[854], _009776_, _009777_);
  or g_102780_(out[855], _009777_, _009779_);
  and g_102781_(out[856], _009779_, _009780_);
  or g_102782_(out[857], _009780_, _009781_);
  not g_102783_(_009781_, _009782_);
  or g_102784_(out[858], _009781_, _009783_);
  xor g_102785_(out[859], _009783_, _009784_);
  xor g_102786_(_001418_, _009783_, _009785_);
  and g_102787_(_009770_, _009784_, _009786_);
  or g_102788_(_009771_, _009785_, _009787_);
  or g_102789_(out[867], _002016_, _009788_);
  not g_102790_(_009788_, _009790_);
  and g_102791_(out[868], _009788_, _009791_);
  or g_102792_(_001594_, _009790_, _009792_);
  and g_102793_(out[869], _009791_, _009793_);
  and g_102794_(out[870], _009793_, _009794_);
  or g_102795_(out[871], _009794_, _009795_);
  and g_102796_(out[872], _009795_, _009796_);
  or g_102797_(out[873], _009796_, _009797_);
  not g_102798_(_009797_, _009798_);
  or g_102799_(out[874], _009797_, _009799_);
  xor g_102800_(out[875], _009799_, _009801_);
  xor g_102801_(_001550_, _009799_, _009802_);
  and g_102802_(_009786_, _009801_, _009803_);
  or g_102803_(_009787_, _009802_, _009804_);
  or g_102804_(out[883], _002075_, _009805_);
  not g_102805_(_009805_, _009806_);
  and g_102806_(out[884], _009805_, _009807_);
  or g_102807_(_001726_, _009806_, _009808_);
  and g_102808_(out[885], _009807_, _009809_);
  and g_102809_(out[886], _009809_, _009810_);
  or g_102810_(out[887], _009810_, _009812_);
  and g_102811_(out[888], _009812_, _009813_);
  or g_102812_(out[889], _009813_, _009814_);
  not g_102813_(_009814_, _009815_);
  or g_102814_(out[890], _009814_, _009816_);
  xor g_102815_(out[891], _009816_, _009817_);
  xor g_102816_(_001682_, _009816_, _009818_);
  and g_102817_(_009803_, _009817_, _009819_);
  or g_102818_(_009804_, _009818_, _009820_);
  or g_102819_(out[899], _002332_, _009821_);
  not g_102820_(_009821_, _009823_);
  and g_102821_(out[900], _009821_, _009824_);
  or g_102822_(_001858_, _009823_, _009825_);
  and g_102823_(out[901], _009824_, _009826_);
  and g_102824_(out[902], _009826_, _009827_);
  or g_102825_(out[903], _009827_, _009828_);
  and g_102826_(out[904], _009828_, _009829_);
  or g_102827_(out[905], _009829_, _009830_);
  not g_102828_(_009830_, _009831_);
  or g_102829_(out[906], _009830_, _009832_);
  xor g_102830_(out[907], _009832_, _009834_);
  xor g_102831_(_001814_, _009832_, _009835_);
  and g_102832_(_009819_, _009834_, _009836_);
  or g_102833_(_009820_, _009835_, _009837_);
  or g_102834_(out[915], _002528_, _009838_);
  not g_102835_(_009838_, _009839_);
  and g_102836_(out[916], _009838_, _009840_);
  or g_102837_(_001990_, _009839_, _009841_);
  and g_102838_(out[917], _009840_, _009842_);
  and g_102839_(out[918], _009842_, _009843_);
  or g_102840_(out[919], _009843_, _009845_);
  and g_102841_(out[920], _009845_, _009846_);
  or g_102842_(out[921], _009846_, _009847_);
  not g_102843_(_009847_, _009848_);
  or g_102844_(out[922], _009847_, _009849_);
  xor g_102845_(out[923], _009849_, _009850_);
  xor g_102846_(_001946_, _009849_, _009851_);
  and g_102847_(_009836_, _009850_, _009852_);
  or g_102848_(_009837_, _009851_, _009853_);
  or g_102849_(_009409_, _009853_, _009854_);
  not g_102850_(_009854_, _009856_);
  xor g_102851_(out[938], _009407_, _009857_);
  not g_102852_(_009857_, _009858_);
  xor g_102853_(out[522], _009446_, _009859_);
  xor g_102854_(_054732_, _009446_, _009860_);
  xor g_102855_(out[506], _009431_, _009861_);
  xor g_102856_(_054600_, _009431_, _009862_);
  and g_102857_(_009421_, _009434_, _009863_);
  or g_102858_(_009422_, _009433_, _009864_);
  xor g_102859_(out[490], _009419_, _009865_);
  xor g_102860_(_054468_, _009419_, _009867_);
  or g_102861_(_009862_, _009865_, _009868_);
  not g_102862_(_009868_, _009869_);
  and g_102863_(_009864_, _009868_, _009870_);
  or g_102864_(_009863_, _009869_, _009871_);
  and g_102865_(out[489], _009418_, _009872_);
  xor g_102866_(out[489], _009418_, _009873_);
  xor g_102867_(_054457_, _009418_, _009874_);
  and g_102868_(out[505], _009430_, _009875_);
  xor g_102869_(out[505], _009430_, _009876_);
  xor g_102870_(_054589_, _009430_, _009878_);
  and g_102871_(_009873_, _009878_, _009879_);
  or g_102872_(_009874_, _009876_, _009880_);
  and g_102873_(_009874_, _009876_, _009881_);
  or g_102874_(_009873_, _009878_, _009882_);
  xor g_102875_(_009874_, _009876_, _009883_);
  xor g_102876_(_009873_, _009876_, _009884_);
  xor g_102877_(out[488], _009417_, _009885_);
  xor g_102878_(_054446_, _009417_, _009886_);
  xor g_102879_(out[504], _009429_, _009887_);
  xor g_102880_(_054578_, _009429_, _009889_);
  and g_102881_(_009885_, _009889_, _009890_);
  or g_102882_(_009886_, _009887_, _009891_);
  xor g_102883_(_009886_, _009887_, _009892_);
  xor g_102884_(_009885_, _009887_, _009893_);
  and g_102885_(_009883_, _009892_, _009894_);
  or g_102886_(_009884_, _009893_, _009895_);
  and g_102887_(_009422_, _009433_, _009896_);
  or g_102888_(_009421_, _009434_, _009897_);
  and g_102889_(_009864_, _009897_, _009898_);
  or g_102890_(_009863_, _009896_, _009900_);
  xor g_102891_(_009862_, _009865_, _009901_);
  xor g_102892_(_009861_, _009865_, _009902_);
  and g_102893_(_009898_, _009901_, _009903_);
  or g_102894_(_009900_, _009902_, _009904_);
  and g_102895_(_009894_, _009903_, _009905_);
  or g_102896_(_009895_, _009904_, _009906_);
  xor g_102897_(out[487], _009416_, _009907_);
  xor g_102898_(_054369_, _009416_, _009908_);
  xor g_102899_(out[503], _009428_, _009909_);
  xor g_102900_(_054490_, _009428_, _009911_);
  and g_102901_(_009908_, _009909_, _009912_);
  or g_102902_(_009907_, _009911_, _009913_);
  xor g_102903_(out[486], _009414_, _009914_);
  xor g_102904_(_054380_, _009414_, _009915_);
  xor g_102905_(out[502], _009427_, _009916_);
  xor g_102906_(_054501_, _009427_, _009917_);
  and g_102907_(_009914_, _009917_, _009918_);
  or g_102908_(_009915_, _009916_, _009919_);
  and g_102909_(_009913_, _009919_, _009920_);
  or g_102910_(_009912_, _009918_, _009922_);
  and g_102911_(_009915_, _009916_, _009923_);
  or g_102912_(_009914_, _009917_, _009924_);
  and g_102913_(_009907_, _009911_, _009925_);
  or g_102914_(_009908_, _009909_, _009926_);
  and g_102915_(_009924_, _009926_, _009927_);
  or g_102916_(_009923_, _009925_, _009928_);
  and g_102917_(_009920_, _009927_, _009929_);
  or g_102918_(_009922_, _009928_, _009930_);
  or g_102919_(_016103_, _016389_, _009931_);
  not g_102920_(_009931_, _009933_);
  and g_102921_(_009413_, _009931_, _009934_);
  or g_102922_(_009412_, _009933_, _009935_);
  or g_102923_(_015971_, _016356_, _009936_);
  not g_102924_(_009936_, _009937_);
  and g_102925_(_009425_, _009936_, _009938_);
  or g_102926_(_009424_, _009937_, _009939_);
  and g_102927_(_009934_, _009939_, _009940_);
  or g_102928_(_009935_, _009938_, _009941_);
  xor g_102929_(out[501], _009424_, _009942_);
  xor g_102930_(_054512_, _009424_, _009944_);
  xor g_102931_(out[485], _009412_, _009945_);
  xor g_102932_(_054391_, _009412_, _009946_);
  and g_102933_(_009944_, _009945_, _009947_);
  or g_102934_(_009942_, _009946_, _009948_);
  and g_102935_(_009941_, _009948_, _009949_);
  or g_102936_(_009940_, _009947_, _009950_);
  and g_102937_(_009942_, _009946_, _009951_);
  or g_102938_(_009944_, _009945_, _009952_);
  and g_102939_(_009935_, _009938_, _009953_);
  or g_102940_(_009934_, _009939_, _009955_);
  and g_102941_(_009952_, _009955_, _009956_);
  or g_102942_(_009951_, _009953_, _009957_);
  and g_102943_(_009949_, _009956_, _009958_);
  or g_102944_(_009950_, _009957_, _009959_);
  and g_102945_(_009929_, _009958_, _009960_);
  or g_102946_(_009930_, _009959_, _009961_);
  and g_102947_(_016884_, _009960_, _009962_);
  or g_102948_(_016895_, _009961_, _009963_);
  and g_102949_(_009905_, _009962_, _009964_);
  or g_102950_(_009906_, _009963_, _009966_);
  xor g_102951_(out[499], _016356_, _009967_);
  xor g_102952_(_054567_, _016356_, _009968_);
  xor g_102953_(out[483], _016389_, _009969_);
  xor g_102954_(_054435_, _016389_, _009970_);
  and g_102955_(_009968_, _009969_, _009971_);
  or g_102956_(_009967_, _009970_, _009972_);
  and g_102957_(_009967_, _009970_, _009973_);
  or g_102958_(_009968_, _009969_, _009974_);
  and g_102959_(_016455_, _009974_, _009975_);
  or g_102960_(_016444_, _009973_, _009977_);
  and g_102961_(_009972_, _009977_, _009978_);
  or g_102962_(_009971_, _009975_, _009979_);
  and g_102963_(_016697_, _009979_, _009980_);
  or g_102964_(_016686_, _009978_, _009981_);
  and g_102965_(_009960_, _009981_, _009982_);
  or g_102966_(_009961_, _009980_, _009983_);
  and g_102967_(_009950_, _009952_, _009984_);
  or g_102968_(_009949_, _009951_, _009985_);
  and g_102969_(_009929_, _009984_, _009986_);
  or g_102970_(_009930_, _009985_, _009988_);
  and g_102971_(_009922_, _009926_, _009989_);
  or g_102972_(_009920_, _009925_, _009990_);
  and g_102973_(_009988_, _009990_, _009991_);
  or g_102974_(_009986_, _009989_, _009992_);
  and g_102975_(_009983_, _009991_, _009993_);
  or g_102976_(_009982_, _009992_, _009994_);
  and g_102977_(_009905_, _009994_, _009995_);
  or g_102978_(_009906_, _009993_, _009996_);
  and g_102979_(_009871_, _009897_, _009997_);
  or g_102980_(_009870_, _009896_, _009999_);
  and g_102981_(_009883_, _009890_, _010000_);
  or g_102982_(_009884_, _009891_, _010001_);
  and g_102983_(_009882_, _010001_, _010002_);
  or g_102984_(_009881_, _010000_, _010003_);
  and g_102985_(_009903_, _010003_, _010004_);
  or g_102986_(_009904_, _010002_, _010005_);
  and g_102987_(_009999_, _010005_, _010006_);
  or g_102988_(_009997_, _010004_, _010007_);
  and g_102989_(_009996_, _010006_, _010008_);
  or g_102990_(_009995_, _010007_, _010010_);
  and g_102991_(_009966_, _010010_, _010011_);
  or g_102992_(_009964_, _010008_, _010012_);
  and g_102993_(_009861_, _010011_, _010013_);
  or g_102994_(_009862_, _010012_, _010014_);
  and g_102995_(_009865_, _010012_, _010015_);
  or g_102996_(_009867_, _010011_, _010016_);
  and g_102997_(_010014_, _010016_, _010017_);
  or g_102998_(_010013_, _010015_, _010018_);
  and g_102999_(_009859_, _010017_, _010019_);
  or g_103000_(_009860_, _010018_, _010021_);
  and g_103001_(_009435_, _009451_, _010022_);
  or g_103002_(_009436_, _009450_, _010023_);
  and g_103003_(_010021_, _010023_, _010024_);
  or g_103004_(_010019_, _010022_, _010025_);
  and g_103005_(_009436_, _009450_, _010026_);
  or g_103006_(_009435_, _009451_, _010027_);
  and g_103007_(_009860_, _010018_, _010028_);
  or g_103008_(_009859_, _010017_, _010029_);
  and g_103009_(_010027_, _010029_, _010030_);
  or g_103010_(_010026_, _010028_, _010032_);
  and g_103011_(_010024_, _010030_, _010033_);
  or g_103012_(_010025_, _010032_, _010034_);
  and g_103013_(out[521], _009445_, _010035_);
  xor g_103014_(out[521], _009445_, _010036_);
  or g_103015_(_009447_, _010035_, _010037_);
  and g_103016_(_009876_, _010011_, _010038_);
  or g_103017_(_009878_, _010012_, _010039_);
  and g_103018_(_009873_, _010012_, _010040_);
  or g_103019_(_009874_, _010011_, _010041_);
  and g_103020_(_010039_, _010041_, _010043_);
  or g_103021_(_010038_, _010040_, _010044_);
  and g_103022_(_010036_, _010043_, _010045_);
  or g_103023_(_010037_, _010044_, _010046_);
  and g_103024_(_009889_, _010011_, _010047_);
  or g_103025_(_009887_, _010012_, _010048_);
  and g_103026_(_009886_, _010012_, _010049_);
  or g_103027_(_009885_, _010011_, _010050_);
  and g_103028_(_010048_, _010050_, _010051_);
  or g_103029_(_010047_, _010049_, _010052_);
  xor g_103030_(out[520], _009444_, _010054_);
  xor g_103031_(_054710_, _009444_, _010055_);
  and g_103032_(_010051_, _010055_, _010056_);
  or g_103033_(_010052_, _010054_, _010057_);
  and g_103034_(_010046_, _010057_, _010058_);
  or g_103035_(_010045_, _010056_, _010059_);
  and g_103036_(_010037_, _010044_, _010060_);
  or g_103037_(_010036_, _010043_, _010061_);
  and g_103038_(_010052_, _010054_, _010062_);
  or g_103039_(_010051_, _010055_, _010063_);
  and g_103040_(_010061_, _010063_, _010065_);
  or g_103041_(_010060_, _010062_, _010066_);
  and g_103042_(_010058_, _010065_, _010067_);
  or g_103043_(_010059_, _010066_, _010068_);
  and g_103044_(_010033_, _010067_, _010069_);
  or g_103045_(_010034_, _010068_, _010070_);
  xor g_103046_(out[518], _009442_, _010071_);
  not g_103047_(_010071_, _010072_);
  or g_103048_(_009916_, _010012_, _010073_);
  or g_103049_(_009914_, _010011_, _010074_);
  and g_103050_(_010073_, _010074_, _010076_);
  and g_103051_(_010072_, _010076_, _010077_);
  xor g_103052_(_010072_, _010076_, _010078_);
  xor g_103053_(_010071_, _010076_, _010079_);
  xor g_103054_(out[519], _009443_, _010080_);
  xor g_103055_(_054622_, _009443_, _010081_);
  or g_103056_(_009911_, _010012_, _010082_);
  or g_103057_(_009908_, _010011_, _010083_);
  and g_103058_(_010082_, _010083_, _010084_);
  and g_103059_(_010080_, _010084_, _010085_);
  or g_103060_(_010080_, _010084_, _010087_);
  xor g_103061_(_010080_, _010084_, _010088_);
  xor g_103062_(_010081_, _010084_, _010089_);
  and g_103063_(_010078_, _010088_, _010090_);
  or g_103064_(_010079_, _010089_, _010091_);
  or g_103065_(_015839_, _019073_, _010092_);
  not g_103066_(_010092_, _010093_);
  and g_103067_(_009441_, _010092_, _010094_);
  or g_103068_(_009440_, _010093_, _010095_);
  and g_103069_(_009935_, _010012_, _010096_);
  or g_103070_(_009934_, _010011_, _010098_);
  and g_103071_(_009939_, _010011_, _010099_);
  or g_103072_(_009938_, _010012_, _010100_);
  and g_103073_(_010098_, _010100_, _010101_);
  or g_103074_(_010096_, _010099_, _010102_);
  and g_103075_(_010095_, _010101_, _010103_);
  or g_103076_(_010094_, _010102_, _010104_);
  xor g_103077_(out[517], _009440_, _010105_);
  xor g_103078_(_054644_, _009440_, _010106_);
  and g_103079_(_009944_, _010011_, _010107_);
  or g_103080_(_009942_, _010012_, _010109_);
  and g_103081_(_009946_, _010012_, _010110_);
  or g_103082_(_009945_, _010011_, _010111_);
  and g_103083_(_010109_, _010111_, _010112_);
  or g_103084_(_010107_, _010110_, _010113_);
  and g_103085_(_010106_, _010112_, _010114_);
  or g_103086_(_010105_, _010113_, _010115_);
  and g_103087_(_010104_, _010115_, _010116_);
  or g_103088_(_010103_, _010114_, _010117_);
  and g_103089_(_010105_, _010113_, _010118_);
  or g_103090_(_010106_, _010112_, _010120_);
  and g_103091_(_010094_, _010102_, _010121_);
  or g_103092_(_010095_, _010101_, _010122_);
  and g_103093_(_010120_, _010122_, _010123_);
  or g_103094_(_010118_, _010121_, _010124_);
  and g_103095_(_010116_, _010123_, _010125_);
  or g_103096_(_010117_, _010124_, _010126_);
  and g_103097_(_010090_, _010125_, _010127_);
  or g_103098_(_010091_, _010126_, _010128_);
  and g_103099_(_010069_, _010127_, _010129_);
  or g_103100_(_010070_, _010128_, _010131_);
  xor g_103101_(out[515], _019073_, _010132_);
  xor g_103102_(_054699_, _019073_, _010133_);
  and g_103103_(_009967_, _010011_, _010134_);
  or g_103104_(_009968_, _010012_, _010135_);
  and g_103105_(_009969_, _010012_, _010136_);
  not g_103106_(_010136_, _010137_);
  and g_103107_(_010135_, _010137_, _010138_);
  or g_103108_(_010134_, _010136_, _010139_);
  and g_103109_(_010132_, _010138_, _010140_);
  or g_103110_(_010133_, _010139_, _010142_);
  and g_103111_(_016400_, _010012_, _010143_);
  and g_103112_(_016367_, _010011_, _010144_);
  or g_103113_(_010143_, _010144_, _010145_);
  not g_103114_(_010145_, _010146_);
  and g_103115_(_019084_, _010146_, _010147_);
  or g_103116_(_019095_, _010145_, _010148_);
  and g_103117_(_010142_, _010148_, _010149_);
  or g_103118_(_010140_, _010147_, _010150_);
  and g_103119_(_010133_, _010139_, _010151_);
  or g_103120_(_010132_, _010138_, _010153_);
  and g_103121_(_019095_, _010145_, _010154_);
  or g_103122_(_019084_, _010146_, _010155_);
  and g_103123_(_010153_, _010155_, _010156_);
  or g_103124_(_010151_, _010154_, _010157_);
  and g_103125_(_010149_, _010156_, _010158_);
  or g_103126_(_010150_, _010157_, _010159_);
  or g_103127_(_054534_, _010012_, _010160_);
  or g_103128_(_054413_, _010011_, _010161_);
  and g_103129_(_010160_, _010161_, _010162_);
  and g_103130_(out[513], _010162_, _010164_);
  not g_103131_(_010164_, _010165_);
  and g_103132_(_054347_, _010012_, _010166_);
  or g_103133_(out[480], _010011_, _010167_);
  or g_103134_(out[496], _010012_, _010168_);
  not g_103135_(_010168_, _010169_);
  and g_103136_(_010167_, _010168_, _010170_);
  or g_103137_(_010166_, _010169_, _010171_);
  and g_103138_(out[512], _010171_, _010172_);
  or g_103139_(_054677_, _010170_, _010173_);
  xor g_103140_(out[513], _010162_, _010175_);
  xor g_103141_(_054666_, _010162_, _010176_);
  and g_103142_(_010173_, _010175_, _010177_);
  or g_103143_(_010172_, _010176_, _010178_);
  and g_103144_(_010165_, _010178_, _010179_);
  or g_103145_(_010164_, _010177_, _010180_);
  and g_103146_(_010158_, _010180_, _010181_);
  or g_103147_(_010159_, _010179_, _010182_);
  and g_103148_(_010150_, _010153_, _010183_);
  or g_103149_(_010149_, _010151_, _010184_);
  and g_103150_(_010182_, _010184_, _010186_);
  or g_103151_(_010181_, _010183_, _010187_);
  and g_103152_(_010129_, _010187_, _010188_);
  or g_103153_(_010131_, _010186_, _010189_);
  and g_103154_(_010090_, _010117_, _010190_);
  or g_103155_(_010091_, _010116_, _010191_);
  and g_103156_(_010120_, _010190_, _010192_);
  or g_103157_(_010118_, _010191_, _010193_);
  and g_103158_(_010077_, _010087_, _010194_);
  or g_103159_(_010085_, _010194_, _010195_);
  not g_103160_(_010195_, _010197_);
  and g_103161_(_010193_, _010197_, _010198_);
  or g_103162_(_010192_, _010195_, _010199_);
  and g_103163_(_010069_, _010199_, _010200_);
  or g_103164_(_010070_, _010198_, _010201_);
  and g_103165_(_010025_, _010027_, _010202_);
  or g_103166_(_010024_, _010026_, _010203_);
  and g_103167_(_010059_, _010061_, _010204_);
  or g_103168_(_010058_, _010060_, _010205_);
  and g_103169_(_010033_, _010204_, _010206_);
  or g_103170_(_010034_, _010205_, _010208_);
  and g_103171_(_010203_, _010208_, _010209_);
  or g_103172_(_010202_, _010206_, _010210_);
  and g_103173_(_010201_, _010209_, _010211_);
  or g_103174_(_010200_, _010210_, _010212_);
  and g_103175_(_010189_, _010211_, _010213_);
  or g_103176_(_010188_, _010212_, _010214_);
  and g_103177_(_054677_, _010170_, _010215_);
  or g_103178_(out[512], _010171_, _010216_);
  and g_103179_(_010158_, _010177_, _010217_);
  or g_103180_(_010159_, _010178_, _010219_);
  and g_103181_(_010129_, _010217_, _010220_);
  or g_103182_(_010131_, _010219_, _010221_);
  and g_103183_(_010216_, _010220_, _010222_);
  or g_103184_(_010215_, _010221_, _010223_);
  and g_103185_(_010214_, _010223_, _010224_);
  or g_103186_(_010213_, _010222_, _010225_);
  and g_103187_(_009859_, _010224_, _010226_);
  or g_103188_(_009860_, _010225_, _010227_);
  and g_103189_(_010018_, _010225_, _010228_);
  or g_103190_(_010017_, _010224_, _010230_);
  and g_103191_(_010227_, _010230_, _010231_);
  or g_103192_(_010226_, _010228_, _010232_);
  xor g_103193_(out[538], _009463_, _010233_);
  xor g_103194_(_054864_, _009463_, _010234_);
  and g_103195_(_010231_, _010233_, _010235_);
  or g_103196_(_010232_, _010234_, _010236_);
  and g_103197_(_009452_, _009467_, _010237_);
  or g_103198_(_009453_, _009466_, _010238_);
  and g_103199_(_010236_, _010238_, _010239_);
  or g_103200_(_010235_, _010237_, _010241_);
  and g_103201_(_010232_, _010234_, _010242_);
  or g_103202_(_010231_, _010233_, _010243_);
  and g_103203_(_010055_, _010224_, _010244_);
  or g_103204_(_010054_, _010225_, _010245_);
  and g_103205_(_010052_, _010225_, _010246_);
  or g_103206_(_010051_, _010224_, _010247_);
  and g_103207_(_010245_, _010247_, _010248_);
  or g_103208_(_010244_, _010246_, _010249_);
  xor g_103209_(out[536], _009461_, _010250_);
  xor g_103210_(_054842_, _009461_, _010252_);
  and g_103211_(_010248_, _010252_, _010253_);
  or g_103212_(_010249_, _010250_, _010254_);
  and g_103213_(out[537], _009462_, _010255_);
  xor g_103214_(out[537], _009462_, _010256_);
  or g_103215_(_009464_, _010255_, _010257_);
  and g_103216_(_010037_, _010224_, _010258_);
  or g_103217_(_010036_, _010225_, _010259_);
  and g_103218_(_010043_, _010225_, _010260_);
  or g_103219_(_010044_, _010224_, _010261_);
  and g_103220_(_010259_, _010261_, _010263_);
  or g_103221_(_010258_, _010260_, _010264_);
  and g_103222_(_010257_, _010263_, _010265_);
  or g_103223_(_010256_, _010264_, _010266_);
  and g_103224_(_010254_, _010266_, _010267_);
  or g_103225_(_010253_, _010265_, _010268_);
  and g_103226_(_010249_, _010250_, _010269_);
  or g_103227_(_010248_, _010252_, _010270_);
  and g_103228_(_009453_, _009466_, _010271_);
  or g_103229_(_009452_, _009467_, _010272_);
  and g_103230_(_010256_, _010264_, _010274_);
  or g_103231_(_010257_, _010263_, _010275_);
  and g_103232_(_010243_, _010272_, _010276_);
  or g_103233_(_010242_, _010271_, _010277_);
  and g_103234_(_010239_, _010276_, _010278_);
  or g_103235_(_010241_, _010277_, _010279_);
  and g_103236_(_010270_, _010275_, _010280_);
  or g_103237_(_010269_, _010274_, _010281_);
  and g_103238_(_010267_, _010280_, _010282_);
  or g_103239_(_010268_, _010281_, _010283_);
  and g_103240_(_010278_, _010282_, _010285_);
  or g_103241_(_010279_, _010283_, _010286_);
  xor g_103242_(out[534], _009458_, _010287_);
  xor g_103243_(_054765_, _009458_, _010288_);
  or g_103244_(_010071_, _010225_, _010289_);
  or g_103245_(_010076_, _010224_, _010290_);
  and g_103246_(_010289_, _010290_, _010291_);
  and g_103247_(_010288_, _010291_, _010292_);
  xor g_103248_(_010288_, _010291_, _010293_);
  xor g_103249_(_010287_, _010291_, _010294_);
  xor g_103250_(out[535], _009460_, _010296_);
  xor g_103251_(_054754_, _009460_, _010297_);
  or g_103252_(_010081_, _010225_, _010298_);
  or g_103253_(_010084_, _010224_, _010299_);
  and g_103254_(_010298_, _010299_, _010300_);
  not g_103255_(_010300_, _010301_);
  and g_103256_(_010297_, _010301_, _010302_);
  not g_103257_(_010302_, _010303_);
  and g_103258_(_010296_, _010300_, _010304_);
  xor g_103259_(_010296_, _010300_, _010305_);
  or g_103260_(_010294_, _010304_, _010307_);
  and g_103261_(_010293_, _010305_, _010308_);
  or g_103262_(_010302_, _010307_, _010309_);
  or g_103263_(_015707_, _020976_, _010310_);
  not g_103264_(_010310_, _010311_);
  and g_103265_(_009457_, _010310_, _010312_);
  or g_103266_(_009456_, _010311_, _010313_);
  and g_103267_(_010102_, _010225_, _010314_);
  or g_103268_(_010101_, _010224_, _010315_);
  and g_103269_(_010095_, _010224_, _010316_);
  or g_103270_(_010094_, _010225_, _010318_);
  and g_103271_(_010315_, _010318_, _010319_);
  or g_103272_(_010314_, _010316_, _010320_);
  and g_103273_(_010313_, _010319_, _010321_);
  or g_103274_(_010312_, _010320_, _010322_);
  xor g_103275_(out[533], _009456_, _010323_);
  xor g_103276_(_054776_, _009456_, _010324_);
  and g_103277_(_010106_, _010224_, _010325_);
  or g_103278_(_010105_, _010225_, _010326_);
  and g_103279_(_010113_, _010225_, _010327_);
  or g_103280_(_010112_, _010224_, _010329_);
  and g_103281_(_010326_, _010329_, _010330_);
  or g_103282_(_010325_, _010327_, _010331_);
  and g_103283_(_010324_, _010330_, _010332_);
  or g_103284_(_010323_, _010331_, _010333_);
  and g_103285_(_010322_, _010333_, _010334_);
  or g_103286_(_010321_, _010332_, _010335_);
  and g_103287_(_010323_, _010331_, _010336_);
  or g_103288_(_010324_, _010330_, _010337_);
  and g_103289_(_010312_, _010320_, _010338_);
  or g_103290_(_010313_, _010319_, _010340_);
  and g_103291_(_010337_, _010340_, _010341_);
  or g_103292_(_010336_, _010338_, _010342_);
  and g_103293_(_010334_, _010341_, _010343_);
  or g_103294_(_010335_, _010342_, _010344_);
  and g_103295_(_010308_, _010343_, _010345_);
  or g_103296_(_010309_, _010344_, _010346_);
  and g_103297_(_010285_, _010345_, _010347_);
  or g_103298_(_010286_, _010346_, _010348_);
  xor g_103299_(out[531], _020976_, _010349_);
  xor g_103300_(_054831_, _020976_, _010351_);
  and g_103301_(_010132_, _010224_, _010352_);
  or g_103302_(_010133_, _010225_, _010353_);
  and g_103303_(_010139_, _010225_, _010354_);
  or g_103304_(_010138_, _010224_, _010355_);
  and g_103305_(_010353_, _010355_, _010356_);
  or g_103306_(_010352_, _010354_, _010357_);
  and g_103307_(_010351_, _010357_, _010358_);
  or g_103308_(_010349_, _010356_, _010359_);
  and g_103309_(_019084_, _010224_, _010360_);
  and g_103310_(_010145_, _010225_, _010362_);
  or g_103311_(_010360_, _010362_, _010363_);
  not g_103312_(_010363_, _010364_);
  or g_103313_(_020998_, _010363_, _010365_);
  not g_103314_(_010365_, _010366_);
  and g_103315_(_010349_, _010356_, _010367_);
  or g_103316_(_010351_, _010357_, _010368_);
  and g_103317_(_010365_, _010368_, _010369_);
  or g_103318_(_010366_, _010367_, _010370_);
  or g_103319_(_054666_, _010225_, _010371_);
  or g_103320_(_010162_, _010224_, _010373_);
  and g_103321_(_010371_, _010373_, _010374_);
  and g_103322_(out[529], _010374_, _010375_);
  not g_103323_(_010375_, _010376_);
  and g_103324_(out[512], _010224_, _010377_);
  or g_103325_(_054677_, _010225_, _010378_);
  and g_103326_(_010170_, _010225_, _010379_);
  or g_103327_(_010171_, _010224_, _010380_);
  and g_103328_(_010378_, _010380_, _010381_);
  or g_103329_(_010377_, _010379_, _010382_);
  and g_103330_(out[528], _010381_, _010384_);
  or g_103331_(_054809_, _010382_, _010385_);
  xor g_103332_(out[529], _010374_, _010386_);
  xor g_103333_(_054798_, _010374_, _010387_);
  and g_103334_(_010385_, _010386_, _010388_);
  or g_103335_(_010384_, _010387_, _010389_);
  and g_103336_(_010376_, _010389_, _010390_);
  or g_103337_(_010375_, _010388_, _010391_);
  xor g_103338_(_020998_, _010363_, _010392_);
  not g_103339_(_010392_, _010393_);
  and g_103340_(_010391_, _010392_, _010395_);
  or g_103341_(_010370_, _010395_, _010396_);
  and g_103342_(_010359_, _010392_, _010397_);
  or g_103343_(_010358_, _010367_, _010398_);
  or g_103344_(_010393_, _010398_, _010399_);
  or g_103345_(_010390_, _010399_, _010400_);
  or g_103346_(_010358_, _010369_, _010401_);
  and g_103347_(_010359_, _010396_, _010402_);
  and g_103348_(_010400_, _010401_, _010403_);
  and g_103349_(_010347_, _010402_, _010404_);
  or g_103350_(_010348_, _010403_, _010406_);
  or g_103351_(_010334_, _010336_, _010407_);
  and g_103352_(_010308_, _010335_, _010408_);
  and g_103353_(_010337_, _010408_, _010409_);
  or g_103354_(_010309_, _010407_, _010410_);
  or g_103355_(_010292_, _010304_, _010411_);
  not g_103356_(_010411_, _010412_);
  and g_103357_(_010303_, _010411_, _010413_);
  or g_103358_(_010302_, _010412_, _010414_);
  and g_103359_(_010410_, _010414_, _010415_);
  or g_103360_(_010409_, _010413_, _010417_);
  and g_103361_(_010285_, _010417_, _010418_);
  or g_103362_(_010286_, _010415_, _010419_);
  and g_103363_(_010254_, _010275_, _010420_);
  or g_103364_(_010253_, _010274_, _010421_);
  and g_103365_(_010266_, _010421_, _010422_);
  or g_103366_(_010265_, _010420_, _010423_);
  and g_103367_(_010278_, _010422_, _010424_);
  or g_103368_(_010279_, _010423_, _010425_);
  and g_103369_(_010241_, _010272_, _010426_);
  or g_103370_(_010239_, _010271_, _010428_);
  and g_103371_(_010406_, _010425_, _010429_);
  or g_103372_(_010404_, _010424_, _010430_);
  and g_103373_(_010419_, _010428_, _010431_);
  or g_103374_(_010418_, _010426_, _010432_);
  and g_103375_(_010429_, _010431_, _010433_);
  or g_103376_(_010430_, _010432_, _010434_);
  and g_103377_(_054809_, _010382_, _010435_);
  or g_103378_(out[528], _010381_, _010436_);
  and g_103379_(_010368_, _010436_, _010437_);
  and g_103380_(_010397_, _010437_, _010439_);
  and g_103381_(_010388_, _010439_, _010440_);
  or g_103382_(_010348_, _010435_, _010441_);
  or g_103383_(_010389_, _010441_, _010442_);
  and g_103384_(_010347_, _010440_, _010443_);
  or g_103385_(_010399_, _010442_, _010444_);
  and g_103386_(_010434_, _010444_, _010445_);
  or g_103387_(_010433_, _010443_, _010446_);
  and g_103388_(_010232_, _010446_, _010447_);
  or g_103389_(_010231_, _010445_, _010448_);
  and g_103390_(_010233_, _010445_, _010450_);
  or g_103391_(_010234_, _010446_, _010451_);
  and g_103392_(_010448_, _010451_, _010452_);
  or g_103393_(_010447_, _010450_, _010453_);
  xor g_103394_(out[550], _009475_, _010454_);
  xor g_103395_(_054897_, _009475_, _010455_);
  or g_103396_(_010287_, _010446_, _010456_);
  or g_103397_(_010291_, _010445_, _010457_);
  and g_103398_(_010456_, _010457_, _010458_);
  xor g_103399_(out[549], _009473_, _010459_);
  xor g_103400_(_054908_, _009473_, _010461_);
  and g_103401_(_010324_, _010445_, _010462_);
  or g_103402_(_010323_, _010446_, _010463_);
  and g_103403_(_010331_, _010446_, _010464_);
  or g_103404_(_010330_, _010445_, _010465_);
  and g_103405_(_010463_, _010465_, _010466_);
  or g_103406_(_010462_, _010464_, _010467_);
  and g_103407_(_010459_, _010467_, _010468_);
  or g_103408_(_010461_, _010466_, _010469_);
  xor g_103409_(out[551], _009476_, _010470_);
  xor g_103410_(_054886_, _009476_, _010472_);
  or g_103411_(_010297_, _010446_, _010473_);
  or g_103412_(_010300_, _010445_, _010474_);
  and g_103413_(_010473_, _010474_, _010475_);
  and g_103414_(_010470_, _010475_, _010476_);
  and g_103415_(_010455_, _010458_, _010477_);
  or g_103416_(_010470_, _010475_, _010478_);
  xor g_103417_(_010455_, _010458_, _010479_);
  xor g_103418_(_010454_, _010458_, _010480_);
  xor g_103419_(_010470_, _010475_, _010481_);
  xor g_103420_(_010472_, _010475_, _010483_);
  and g_103421_(_010479_, _010481_, _010484_);
  or g_103422_(_010480_, _010483_, _010485_);
  and g_103423_(_010469_, _010484_, _010486_);
  or g_103424_(_010468_, _010485_, _010487_);
  or g_103425_(_015575_, _054003_, _010488_);
  not g_103426_(_010488_, _010489_);
  and g_103427_(_009474_, _010488_, _010490_);
  or g_103428_(_009473_, _010489_, _010491_);
  and g_103429_(_010320_, _010446_, _010492_);
  or g_103430_(_010319_, _010445_, _010494_);
  and g_103431_(_010313_, _010445_, _010495_);
  or g_103432_(_010312_, _010446_, _010496_);
  and g_103433_(_010494_, _010496_, _010497_);
  or g_103434_(_010492_, _010495_, _010498_);
  and g_103435_(_010491_, _010497_, _010499_);
  or g_103436_(_010490_, _010498_, _010500_);
  and g_103437_(_010461_, _010466_, _010501_);
  or g_103438_(_010459_, _010467_, _010502_);
  and g_103439_(_010500_, _010502_, _010503_);
  or g_103440_(_010499_, _010501_, _010505_);
  and g_103441_(_010490_, _010498_, _010506_);
  or g_103442_(_010491_, _010497_, _010507_);
  and g_103443_(_010503_, _010507_, _010508_);
  or g_103444_(_010505_, _010506_, _010509_);
  and g_103445_(_010486_, _010508_, _010510_);
  or g_103446_(_010487_, _010509_, _010511_);
  xor g_103447_(out[554], _009479_, _010512_);
  xor g_103448_(_054996_, _009479_, _010513_);
  and g_103449_(_010452_, _010512_, _010514_);
  or g_103450_(_010453_, _010513_, _010516_);
  and g_103451_(_009468_, _009484_, _010517_);
  or g_103452_(_009469_, _009483_, _010518_);
  and g_103453_(_010516_, _010518_, _010519_);
  or g_103454_(_010514_, _010517_, _010520_);
  and g_103455_(_010453_, _010513_, _010521_);
  or g_103456_(_010452_, _010512_, _010522_);
  and g_103457_(_009469_, _009483_, _010523_);
  or g_103458_(_009468_, _009484_, _010524_);
  and g_103459_(out[553], _009478_, _010525_);
  xor g_103460_(out[553], _009478_, _010527_);
  or g_103461_(_009480_, _010525_, _010528_);
  and g_103462_(_010264_, _010446_, _010529_);
  or g_103463_(_010263_, _010445_, _010530_);
  and g_103464_(_010257_, _010445_, _010531_);
  or g_103465_(_010256_, _010446_, _010532_);
  and g_103466_(_010530_, _010532_, _010533_);
  or g_103467_(_010529_, _010531_, _010534_);
  and g_103468_(_010528_, _010533_, _010535_);
  or g_103469_(_010527_, _010534_, _010536_);
  and g_103470_(_010252_, _010445_, _010538_);
  or g_103471_(_010250_, _010446_, _010539_);
  and g_103472_(_010249_, _010446_, _010540_);
  or g_103473_(_010248_, _010445_, _010541_);
  and g_103474_(_010539_, _010541_, _010542_);
  or g_103475_(_010538_, _010540_, _010543_);
  xor g_103476_(out[552], _009477_, _010544_);
  xor g_103477_(_054974_, _009477_, _010545_);
  and g_103478_(_010543_, _010544_, _010546_);
  or g_103479_(_010542_, _010545_, _010547_);
  and g_103480_(_010527_, _010534_, _010549_);
  or g_103481_(_010528_, _010533_, _010550_);
  and g_103482_(_010542_, _010545_, _010551_);
  or g_103483_(_010543_, _010544_, _010552_);
  and g_103484_(_010522_, _010524_, _010553_);
  or g_103485_(_010521_, _010523_, _010554_);
  and g_103486_(_010519_, _010553_, _010555_);
  or g_103487_(_010520_, _010554_, _010556_);
  and g_103488_(_010547_, _010550_, _010557_);
  or g_103489_(_010546_, _010549_, _010558_);
  and g_103490_(_010536_, _010552_, _010560_);
  or g_103491_(_010535_, _010551_, _010561_);
  and g_103492_(_010557_, _010560_, _010562_);
  or g_103493_(_010558_, _010561_, _010563_);
  and g_103494_(_010555_, _010562_, _010564_);
  or g_103495_(_010556_, _010563_, _010565_);
  xor g_103496_(out[547], _054003_, _010566_);
  xor g_103497_(_054963_, _054003_, _010567_);
  or g_103498_(_010356_, _010445_, _010568_);
  or g_103499_(_010351_, _010446_, _010569_);
  and g_103500_(_010568_, _010569_, _010571_);
  and g_103501_(_010566_, _010571_, _010572_);
  and g_103502_(_010363_, _010446_, _010573_);
  or g_103503_(_010364_, _010445_, _010574_);
  and g_103504_(_020987_, _010445_, _010575_);
  or g_103505_(_020998_, _010446_, _010576_);
  and g_103506_(_010574_, _010576_, _010577_);
  or g_103507_(_010573_, _010575_, _010578_);
  or g_103508_(_010566_, _010571_, _010579_);
  and g_103509_(_054004_, _010577_, _010580_);
  xor g_103510_(_010566_, _010571_, _010582_);
  xor g_103511_(_010567_, _010571_, _010583_);
  xor g_103512_(_054004_, _010577_, _010584_);
  xor g_103513_(_054005_, _010577_, _010585_);
  and g_103514_(_010582_, _010584_, _010586_);
  or g_103515_(_010583_, _010585_, _010587_);
  or g_103516_(_054798_, _010446_, _010588_);
  or g_103517_(_010374_, _010445_, _010589_);
  and g_103518_(_010588_, _010589_, _010590_);
  and g_103519_(out[528], _010445_, _010591_);
  or g_103520_(_054809_, _010446_, _010593_);
  and g_103521_(_010382_, _010446_, _010594_);
  or g_103522_(_010381_, _010445_, _010595_);
  and g_103523_(_010593_, _010595_, _010596_);
  or g_103524_(_010591_, _010594_, _010597_);
  and g_103525_(out[544], _010596_, _010598_);
  or g_103526_(_054941_, _010597_, _010599_);
  and g_103527_(out[545], _010590_, _010600_);
  not g_103528_(_010600_, _010601_);
  xor g_103529_(out[545], _010590_, _010602_);
  xor g_103530_(_054930_, _010590_, _010604_);
  and g_103531_(_010599_, _010602_, _010605_);
  or g_103532_(_010598_, _010604_, _010606_);
  and g_103533_(_054941_, _010597_, _010607_);
  or g_103534_(out[544], _010596_, _010608_);
  and g_103535_(_010605_, _010608_, _010609_);
  or g_103536_(_010606_, _010607_, _010610_);
  and g_103537_(_010586_, _010609_, _010611_);
  or g_103538_(_010587_, _010610_, _010612_);
  and g_103539_(_010564_, _010611_, _010613_);
  or g_103540_(_010565_, _010612_, _010615_);
  and g_103541_(_010510_, _010613_, _010616_);
  or g_103542_(_010511_, _010615_, _010617_);
  and g_103543_(_010601_, _010606_, _010618_);
  or g_103544_(_010600_, _010605_, _010619_);
  and g_103545_(_010586_, _010619_, _010620_);
  or g_103546_(_010587_, _010618_, _010621_);
  and g_103547_(_010579_, _010580_, _010622_);
  or g_103548_(_010572_, _010622_, _010623_);
  not g_103549_(_010623_, _010624_);
  and g_103550_(_010621_, _010624_, _010626_);
  or g_103551_(_010620_, _010623_, _010627_);
  and g_103552_(_010510_, _010627_, _010628_);
  or g_103553_(_010511_, _010626_, _010629_);
  and g_103554_(_010486_, _010505_, _010630_);
  and g_103555_(_010477_, _010478_, _010631_);
  or g_103556_(_010476_, _010631_, _010632_);
  or g_103557_(_010630_, _010632_, _010633_);
  not g_103558_(_010633_, _010634_);
  and g_103559_(_010629_, _010634_, _010635_);
  or g_103560_(_010628_, _010633_, _010637_);
  and g_103561_(_010564_, _010637_, _010638_);
  or g_103562_(_010565_, _010635_, _010639_);
  and g_103563_(_010536_, _010551_, _010640_);
  or g_103564_(_010535_, _010552_, _010641_);
  and g_103565_(_010550_, _010641_, _010642_);
  or g_103566_(_010549_, _010640_, _010643_);
  and g_103567_(_010555_, _010643_, _010644_);
  or g_103568_(_010556_, _010642_, _010645_);
  and g_103569_(_010520_, _010524_, _010646_);
  or g_103570_(_010519_, _010523_, _010648_);
  and g_103571_(_010645_, _010648_, _010649_);
  or g_103572_(_010644_, _010646_, _010650_);
  and g_103573_(_010639_, _010649_, _010651_);
  or g_103574_(_010638_, _010650_, _010652_);
  and g_103575_(_010617_, _010652_, _010653_);
  or g_103576_(_010616_, _010651_, _010654_);
  and g_103577_(_010453_, _010654_, _010655_);
  or g_103578_(_010452_, _010653_, _010656_);
  and g_103579_(_010512_, _010653_, _010657_);
  or g_103580_(_010513_, _010654_, _010659_);
  and g_103581_(_010656_, _010659_, _010660_);
  or g_103582_(_010655_, _010657_, _010661_);
  xor g_103583_(out[570], _009496_, _010662_);
  xor g_103584_(_055128_, _009496_, _010663_);
  and g_103585_(_010660_, _010662_, _010664_);
  or g_103586_(_010661_, _010663_, _010665_);
  and g_103587_(_009485_, _009500_, _010666_);
  or g_103588_(_009486_, _009499_, _010667_);
  and g_103589_(_010665_, _010667_, _010668_);
  or g_103590_(_010664_, _010666_, _010670_);
  and g_103591_(_009486_, _009499_, _010671_);
  or g_103592_(_009485_, _009500_, _010672_);
  and g_103593_(_010661_, _010663_, _010673_);
  or g_103594_(_010660_, _010662_, _010674_);
  and g_103595_(_010672_, _010674_, _010675_);
  or g_103596_(_010671_, _010673_, _010676_);
  and g_103597_(out[569], _009495_, _010677_);
  xor g_103598_(out[569], _009495_, _010678_);
  or g_103599_(_009497_, _010677_, _010679_);
  or g_103600_(_010533_, _010653_, _010681_);
  not g_103601_(_010681_, _010682_);
  and g_103602_(_010528_, _010653_, _010683_);
  not g_103603_(_010683_, _010684_);
  and g_103604_(_010681_, _010684_, _010685_);
  or g_103605_(_010682_, _010683_, _010686_);
  and g_103606_(_010679_, _010685_, _010687_);
  or g_103607_(_010678_, _010686_, _010688_);
  and g_103608_(_010675_, _010688_, _010689_);
  or g_103609_(_010676_, _010687_, _010690_);
  and g_103610_(_010668_, _010689_, _010692_);
  or g_103611_(_010670_, _010690_, _010693_);
  and g_103612_(_010545_, _010653_, _010694_);
  not g_103613_(_010694_, _010695_);
  or g_103614_(_010542_, _010653_, _010696_);
  not g_103615_(_010696_, _010697_);
  and g_103616_(_010695_, _010696_, _010698_);
  or g_103617_(_010694_, _010697_, _010699_);
  xor g_103618_(out[568], _009494_, _010700_);
  xor g_103619_(_055106_, _009494_, _010701_);
  and g_103620_(_010699_, _010700_, _010703_);
  or g_103621_(_010698_, _010701_, _010704_);
  and g_103622_(_010678_, _010686_, _010705_);
  or g_103623_(_010679_, _010685_, _010706_);
  and g_103624_(_010698_, _010701_, _010707_);
  or g_103625_(_010699_, _010700_, _010708_);
  and g_103626_(_010706_, _010708_, _010709_);
  or g_103627_(_010705_, _010707_, _010710_);
  and g_103628_(_010704_, _010709_, _010711_);
  or g_103629_(_010703_, _010710_, _010712_);
  and g_103630_(_010692_, _010711_, _010714_);
  or g_103631_(_010693_, _010712_, _010715_);
  xor g_103632_(out[567], _009493_, _010716_);
  xor g_103633_(_055018_, _009493_, _010717_);
  or g_103634_(_010472_, _010654_, _010718_);
  or g_103635_(_010475_, _010653_, _010719_);
  and g_103636_(_010718_, _010719_, _010720_);
  and g_103637_(_010716_, _010720_, _010721_);
  or g_103638_(_010716_, _010720_, _010722_);
  xor g_103639_(_010716_, _010720_, _010723_);
  xor g_103640_(_010717_, _010720_, _010725_);
  xor g_103641_(out[566], _009491_, _010726_);
  xor g_103642_(_055029_, _009491_, _010727_);
  or g_103643_(_010454_, _010654_, _010728_);
  or g_103644_(_010458_, _010653_, _010729_);
  and g_103645_(_010728_, _010729_, _010730_);
  and g_103646_(_010727_, _010730_, _010731_);
  xor g_103647_(_010727_, _010730_, _010732_);
  xor g_103648_(_010726_, _010730_, _010733_);
  and g_103649_(_010723_, _010732_, _010734_);
  or g_103650_(_010725_, _010733_, _010736_);
  or g_103651_(_022307_, _054260_, _010737_);
  not g_103652_(_010737_, _010738_);
  and g_103653_(_009490_, _010737_, _010739_);
  or g_103654_(_009489_, _010738_, _010740_);
  and g_103655_(_010498_, _010654_, _010741_);
  or g_103656_(_010497_, _010653_, _010742_);
  and g_103657_(_010491_, _010653_, _010743_);
  or g_103658_(_010490_, _010654_, _010744_);
  and g_103659_(_010742_, _010744_, _010745_);
  or g_103660_(_010741_, _010743_, _010747_);
  and g_103661_(_010740_, _010745_, _010748_);
  or g_103662_(_010739_, _010747_, _010749_);
  xor g_103663_(out[565], _009489_, _010750_);
  xor g_103664_(_055040_, _009489_, _010751_);
  and g_103665_(_010461_, _010653_, _010752_);
  or g_103666_(_010459_, _010654_, _010753_);
  and g_103667_(_010467_, _010654_, _010754_);
  or g_103668_(_010466_, _010653_, _010755_);
  and g_103669_(_010753_, _010755_, _010756_);
  or g_103670_(_010752_, _010754_, _010758_);
  and g_103671_(_010751_, _010756_, _010759_);
  or g_103672_(_010750_, _010758_, _010760_);
  and g_103673_(_010749_, _010760_, _010761_);
  or g_103674_(_010748_, _010759_, _010762_);
  and g_103675_(_010750_, _010758_, _010763_);
  or g_103676_(_010751_, _010756_, _010764_);
  and g_103677_(_010739_, _010747_, _010765_);
  or g_103678_(_010740_, _010745_, _010766_);
  and g_103679_(_010764_, _010766_, _010767_);
  or g_103680_(_010763_, _010765_, _010769_);
  and g_103681_(_010761_, _010767_, _010770_);
  or g_103682_(_010762_, _010769_, _010771_);
  and g_103683_(_010734_, _010770_, _010772_);
  or g_103684_(_010736_, _010771_, _010773_);
  and g_103685_(_010714_, _010772_, _010774_);
  or g_103686_(_010715_, _010773_, _010775_);
  xor g_103687_(out[563], _054260_, _010776_);
  xor g_103688_(_055095_, _054260_, _010777_);
  and g_103689_(_010566_, _010653_, _010778_);
  not g_103690_(_010778_, _010780_);
  or g_103691_(_010571_, _010653_, _010781_);
  not g_103692_(_010781_, _010782_);
  and g_103693_(_010780_, _010781_, _010783_);
  or g_103694_(_010778_, _010782_, _010784_);
  and g_103695_(_010776_, _010783_, _010785_);
  or g_103696_(_010777_, _010784_, _010786_);
  and g_103697_(_010777_, _010784_, _010787_);
  or g_103698_(_010776_, _010783_, _010788_);
  and g_103699_(_054004_, _010653_, _010789_);
  and g_103700_(_010578_, _010654_, _010791_);
  or g_103701_(_010789_, _010791_, _010792_);
  not g_103702_(_010792_, _010793_);
  or g_103703_(_054262_, _010792_, _010794_);
  not g_103704_(_010794_, _010795_);
  and g_103705_(_010788_, _010795_, _010796_);
  or g_103706_(_010787_, _010794_, _010797_);
  and g_103707_(_010786_, _010797_, _010798_);
  or g_103708_(_010785_, _010796_, _010799_);
  or g_103709_(_054930_, _010654_, _010800_);
  or g_103710_(_010590_, _010653_, _010802_);
  and g_103711_(_010800_, _010802_, _010803_);
  and g_103712_(out[561], _010803_, _010804_);
  not g_103713_(_010804_, _010805_);
  and g_103714_(out[544], _010653_, _010806_);
  not g_103715_(_010806_, _010807_);
  or g_103716_(_010596_, _010653_, _010808_);
  not g_103717_(_010808_, _010809_);
  and g_103718_(_010807_, _010808_, _010810_);
  or g_103719_(_010806_, _010809_, _010811_);
  and g_103720_(out[560], _010810_, _010813_);
  or g_103721_(_055073_, _010811_, _010814_);
  xor g_103722_(out[561], _010803_, _010815_);
  xor g_103723_(_055062_, _010803_, _010816_);
  and g_103724_(_010814_, _010815_, _010817_);
  or g_103725_(_010813_, _010816_, _010818_);
  and g_103726_(_010805_, _010818_, _010819_);
  or g_103727_(_010804_, _010817_, _010820_);
  xor g_103728_(_054262_, _010792_, _010821_);
  xor g_103729_(_054261_, _010792_, _010822_);
  and g_103730_(_010788_, _010821_, _010824_);
  or g_103731_(_010787_, _010822_, _010825_);
  and g_103732_(_010820_, _010824_, _010826_);
  or g_103733_(_010819_, _010825_, _010827_);
  and g_103734_(_010798_, _010827_, _010828_);
  or g_103735_(_010799_, _010826_, _010829_);
  and g_103736_(_010774_, _010829_, _010830_);
  or g_103737_(_010775_, _010828_, _010831_);
  and g_103738_(_010734_, _010762_, _010832_);
  or g_103739_(_010736_, _010761_, _010833_);
  and g_103740_(_010764_, _010832_, _010835_);
  or g_103741_(_010763_, _010833_, _010836_);
  and g_103742_(_010722_, _010731_, _010837_);
  or g_103743_(_010721_, _010837_, _010838_);
  not g_103744_(_010838_, _010839_);
  and g_103745_(_010836_, _010839_, _010840_);
  or g_103746_(_010835_, _010838_, _010841_);
  and g_103747_(_010714_, _010841_, _010842_);
  or g_103748_(_010715_, _010840_, _010843_);
  and g_103749_(_010670_, _010672_, _010844_);
  or g_103750_(_010668_, _010671_, _010846_);
  and g_103751_(_010692_, _010710_, _010847_);
  or g_103752_(_010693_, _010709_, _010848_);
  and g_103753_(_010846_, _010848_, _010849_);
  or g_103754_(_010844_, _010847_, _010850_);
  and g_103755_(_010843_, _010849_, _010851_);
  or g_103756_(_010842_, _010850_, _010852_);
  and g_103757_(_010831_, _010851_, _010853_);
  or g_103758_(_010830_, _010852_, _010854_);
  and g_103759_(_055073_, _010811_, _010855_);
  or g_103760_(out[560], _010810_, _010857_);
  and g_103761_(_010786_, _010857_, _010858_);
  or g_103762_(_010785_, _010855_, _010859_);
  and g_103763_(_010817_, _010858_, _010860_);
  or g_103764_(_010818_, _010859_, _010861_);
  and g_103765_(_010824_, _010860_, _010862_);
  or g_103766_(_010825_, _010861_, _010863_);
  and g_103767_(_010774_, _010862_, _010864_);
  or g_103768_(_010775_, _010863_, _010865_);
  and g_103769_(_010854_, _010865_, _010866_);
  or g_103770_(_010853_, _010864_, _010868_);
  and g_103771_(_010661_, _010868_, _010869_);
  or g_103772_(_010660_, _010866_, _010870_);
  and g_103773_(_010662_, _010866_, _010871_);
  or g_103774_(_010663_, _010868_, _010872_);
  and g_103775_(_010870_, _010872_, _010873_);
  or g_103776_(_010869_, _010871_, _010874_);
  and g_103777_(_009502_, _009515_, _010875_);
  or g_103778_(_009501_, _009516_, _010876_);
  and g_103779_(_009501_, _009516_, _010877_);
  or g_103780_(_009502_, _009515_, _010879_);
  xor g_103781_(out[586], _009512_, _010880_);
  not g_103782_(_010880_, _010881_);
  and g_103783_(_010873_, _010880_, _010882_);
  or g_103784_(_010874_, _010881_, _010883_);
  and g_103785_(_010879_, _010883_, _010884_);
  or g_103786_(_010877_, _010882_, _010885_);
  and g_103787_(_010874_, _010881_, _010886_);
  or g_103788_(_010873_, _010880_, _010887_);
  and g_103789_(out[585], _009511_, _010888_);
  xor g_103790_(out[585], _009511_, _010890_);
  xor g_103791_(_055249_, _009511_, _010891_);
  and g_103792_(_010686_, _010868_, _010892_);
  or g_103793_(_010685_, _010866_, _010893_);
  and g_103794_(_010679_, _010866_, _010894_);
  or g_103795_(_010678_, _010868_, _010895_);
  and g_103796_(_010893_, _010895_, _010896_);
  or g_103797_(_010892_, _010894_, _010897_);
  and g_103798_(_010890_, _010897_, _010898_);
  or g_103799_(_010891_, _010896_, _010899_);
  and g_103800_(_010701_, _010866_, _010901_);
  or g_103801_(_010700_, _010868_, _010902_);
  and g_103802_(_010699_, _010868_, _010903_);
  or g_103803_(_010698_, _010866_, _010904_);
  and g_103804_(_010902_, _010904_, _010905_);
  or g_103805_(_010901_, _010903_, _010906_);
  xor g_103806_(out[584], _009510_, _010907_);
  xor g_103807_(_055238_, _009510_, _010908_);
  and g_103808_(_010905_, _010908_, _010909_);
  or g_103809_(_010906_, _010907_, _010910_);
  and g_103810_(_010891_, _010896_, _010912_);
  or g_103811_(_010890_, _010897_, _010913_);
  and g_103812_(_010909_, _010913_, _010914_);
  or g_103813_(_010910_, _010912_, _010915_);
  and g_103814_(_010899_, _010915_, _010916_);
  or g_103815_(_010898_, _010914_, _010917_);
  and g_103816_(_010910_, _010913_, _010918_);
  or g_103817_(_010909_, _010912_, _010919_);
  and g_103818_(_010906_, _010907_, _010920_);
  or g_103819_(_010905_, _010908_, _010921_);
  and g_103820_(_010876_, _010887_, _010923_);
  or g_103821_(_010875_, _010886_, _010924_);
  and g_103822_(_010884_, _010923_, _010925_);
  or g_103823_(_010885_, _010924_, _010926_);
  and g_103824_(_010899_, _010921_, _010927_);
  or g_103825_(_010898_, _010920_, _010928_);
  and g_103826_(_010918_, _010927_, _010929_);
  or g_103827_(_010919_, _010928_, _010930_);
  and g_103828_(_010925_, _010929_, _010931_);
  or g_103829_(_010926_, _010930_, _010932_);
  xor g_103830_(out[583], _009509_, _010934_);
  xor g_103831_(_055150_, _009509_, _010935_);
  or g_103832_(_010717_, _010868_, _010936_);
  or g_103833_(_010720_, _010866_, _010937_);
  and g_103834_(_010936_, _010937_, _010938_);
  and g_103835_(_010934_, _010938_, _010939_);
  xor g_103836_(out[582], _009508_, _010940_);
  xor g_103837_(_055161_, _009508_, _010941_);
  or g_103838_(_010730_, _010866_, _010942_);
  or g_103839_(_010726_, _010868_, _010943_);
  and g_103840_(_010942_, _010943_, _010945_);
  and g_103841_(_010941_, _010945_, _010946_);
  or g_103842_(_010934_, _010938_, _010947_);
  xor g_103843_(_010934_, _010938_, _010948_);
  xor g_103844_(_010935_, _010938_, _010949_);
  xor g_103845_(_010941_, _010945_, _010950_);
  xor g_103846_(_010940_, _010945_, _010951_);
  and g_103847_(_010948_, _010950_, _010952_);
  or g_103848_(_010949_, _010951_, _010953_);
  xor g_103849_(out[581], _009506_, _010954_);
  xor g_103850_(_055172_, _009506_, _010956_);
  and g_103851_(_010751_, _010866_, _010957_);
  or g_103852_(_010750_, _010868_, _010958_);
  and g_103853_(_010758_, _010868_, _010959_);
  or g_103854_(_010756_, _010866_, _010960_);
  and g_103855_(_010958_, _010960_, _010961_);
  or g_103856_(_010957_, _010959_, _010962_);
  and g_103857_(_010954_, _010962_, _010963_);
  or g_103858_(_010956_, _010961_, _010964_);
  or g_103859_(_022461_, _054570_, _010965_);
  not g_103860_(_010965_, _010967_);
  and g_103861_(_009507_, _010965_, _010968_);
  or g_103862_(_009506_, _010967_, _010969_);
  and g_103863_(_010747_, _010868_, _010970_);
  or g_103864_(_010745_, _010866_, _010971_);
  and g_103865_(_010740_, _010866_, _010972_);
  or g_103866_(_010739_, _010868_, _010973_);
  and g_103867_(_010971_, _010973_, _010974_);
  or g_103868_(_010970_, _010972_, _010975_);
  and g_103869_(_010969_, _010974_, _010976_);
  or g_103870_(_010968_, _010975_, _010978_);
  and g_103871_(_010956_, _010961_, _010979_);
  or g_103872_(_010954_, _010962_, _010980_);
  and g_103873_(_010978_, _010980_, _010981_);
  or g_103874_(_010976_, _010979_, _010982_);
  and g_103875_(_010952_, _010982_, _010983_);
  or g_103876_(_010953_, _010981_, _010984_);
  and g_103877_(_010964_, _010983_, _010985_);
  or g_103878_(_010963_, _010984_, _010986_);
  and g_103879_(_010946_, _010947_, _010987_);
  or g_103880_(_010939_, _010987_, _010989_);
  not g_103881_(_010989_, _010990_);
  and g_103882_(_010986_, _010990_, _010991_);
  or g_103883_(_010985_, _010989_, _010992_);
  and g_103884_(_054261_, _010866_, _010993_);
  or g_103885_(_054262_, _010868_, _010994_);
  and g_103886_(_010792_, _010868_, _010995_);
  or g_103887_(_010793_, _010866_, _010996_);
  and g_103888_(_010994_, _010996_, _010997_);
  or g_103889_(_010993_, _010995_, _010998_);
  and g_103890_(_054571_, _010997_, _011000_);
  or g_103891_(_054572_, _010998_, _011001_);
  xor g_103892_(out[579], _054570_, _011002_);
  xor g_103893_(_055227_, _054570_, _011003_);
  and g_103894_(_010776_, _010866_, _011004_);
  or g_103895_(_010777_, _010868_, _011005_);
  and g_103896_(_010784_, _010868_, _011006_);
  or g_103897_(_010783_, _010866_, _011007_);
  and g_103898_(_011005_, _011007_, _011008_);
  or g_103899_(_011004_, _011006_, _011009_);
  and g_103900_(_011002_, _011008_, _011011_);
  or g_103901_(_011003_, _011009_, _011012_);
  and g_103902_(_011001_, _011012_, _011013_);
  or g_103903_(_011000_, _011011_, _011014_);
  or g_103904_(_055062_, _010868_, _011015_);
  or g_103905_(_010803_, _010866_, _011016_);
  and g_103906_(_011015_, _011016_, _011017_);
  and g_103907_(out[577], _011017_, _011018_);
  not g_103908_(_011018_, _011019_);
  and g_103909_(out[560], _010866_, _011020_);
  or g_103910_(_055073_, _010868_, _011022_);
  and g_103911_(_010811_, _010868_, _011023_);
  or g_103912_(_010810_, _010866_, _011024_);
  and g_103913_(_011022_, _011024_, _011025_);
  or g_103914_(_011020_, _011023_, _011026_);
  and g_103915_(out[576], _011025_, _011027_);
  or g_103916_(_055205_, _011026_, _011028_);
  xor g_103917_(out[577], _011017_, _011029_);
  xor g_103918_(_055194_, _011017_, _011030_);
  and g_103919_(_011028_, _011029_, _011031_);
  or g_103920_(_011027_, _011030_, _011033_);
  and g_103921_(_011019_, _011033_, _011034_);
  or g_103922_(_011018_, _011031_, _011035_);
  xor g_103923_(_054571_, _010997_, _011036_);
  xor g_103924_(_054572_, _010997_, _011037_);
  and g_103925_(_010968_, _010975_, _011038_);
  or g_103926_(_010969_, _010974_, _011039_);
  and g_103927_(_011003_, _011009_, _011040_);
  or g_103928_(_011002_, _011008_, _011041_);
  and g_103929_(_010917_, _010925_, _011042_);
  or g_103930_(_010916_, _010926_, _011044_);
  and g_103931_(_010964_, _011039_, _011045_);
  or g_103932_(_010963_, _011038_, _011046_);
  and g_103933_(_010981_, _011045_, _011047_);
  or g_103934_(_010982_, _011046_, _011048_);
  and g_103935_(_010952_, _011047_, _011049_);
  or g_103936_(_010953_, _011048_, _011050_);
  and g_103937_(_010931_, _011049_, _011051_);
  or g_103938_(_010932_, _011050_, _011052_);
  and g_103939_(_011012_, _011041_, _011053_);
  or g_103940_(_011011_, _011040_, _011055_);
  and g_103941_(_011036_, _011053_, _011056_);
  or g_103942_(_011037_, _011055_, _011057_);
  and g_103943_(_011035_, _011056_, _011058_);
  or g_103944_(_011034_, _011057_, _011059_);
  and g_103945_(_011014_, _011041_, _011060_);
  or g_103946_(_011013_, _011040_, _011061_);
  and g_103947_(_011059_, _011061_, _011062_);
  or g_103948_(_011058_, _011060_, _011063_);
  and g_103949_(_011051_, _011063_, _011064_);
  or g_103950_(_011052_, _011062_, _011066_);
  and g_103951_(_011044_, _011066_, _011067_);
  or g_103952_(_011042_, _011064_, _011068_);
  and g_103953_(_010876_, _010885_, _011069_);
  or g_103954_(_010875_, _010884_, _011070_);
  and g_103955_(_010931_, _010992_, _011071_);
  or g_103956_(_010932_, _010991_, _011072_);
  and g_103957_(_011070_, _011072_, _011073_);
  or g_103958_(_011069_, _011071_, _011074_);
  and g_103959_(_011067_, _011073_, _011075_);
  or g_103960_(_011068_, _011074_, _011077_);
  and g_103961_(_055205_, _011026_, _011078_);
  or g_103962_(out[576], _011025_, _011079_);
  and g_103963_(_011051_, _011079_, _011080_);
  or g_103964_(_011052_, _011078_, _011081_);
  and g_103965_(_011031_, _011080_, _011082_);
  or g_103966_(_011033_, _011081_, _011083_);
  and g_103967_(_011056_, _011082_, _011084_);
  or g_103968_(_011057_, _011083_, _011085_);
  and g_103969_(_011077_, _011085_, _011086_);
  or g_103970_(_011075_, _011084_, _011088_);
  and g_103971_(_010874_, _011088_, _011089_);
  or g_103972_(_010873_, _011086_, _011090_);
  and g_103973_(_010880_, _011086_, _011091_);
  or g_103974_(_010881_, _011088_, _011092_);
  and g_103975_(_011090_, _011092_, _011093_);
  or g_103976_(_011089_, _011091_, _011094_);
  xor g_103977_(out[602], _009528_, _011095_);
  not g_103978_(_011095_, _011096_);
  and g_103979_(_011093_, _011095_, _011097_);
  or g_103980_(_011094_, _011096_, _011099_);
  and g_103981_(_009517_, _009531_, _011100_);
  or g_103982_(_009518_, _009530_, _011101_);
  and g_103983_(_011099_, _011101_, _011102_);
  or g_103984_(_011097_, _011100_, _011103_);
  and g_103985_(_009518_, _009530_, _011104_);
  or g_103986_(_009517_, _009531_, _011105_);
  and g_103987_(_011094_, _011096_, _011106_);
  or g_103988_(_011093_, _011095_, _011107_);
  and g_103989_(_011105_, _011107_, _011108_);
  or g_103990_(_011104_, _011106_, _011110_);
  and g_103991_(out[601], _009527_, _011111_);
  xor g_103992_(out[601], _009527_, _011112_);
  xor g_103993_(_055381_, _009527_, _011113_);
  or g_103994_(_010896_, _011086_, _011114_);
  not g_103995_(_011114_, _011115_);
  and g_103996_(_010891_, _011086_, _011116_);
  not g_103997_(_011116_, _011117_);
  and g_103998_(_011114_, _011117_, _011118_);
  or g_103999_(_011115_, _011116_, _011119_);
  and g_104000_(_011113_, _011118_, _011121_);
  or g_104001_(_011112_, _011119_, _011122_);
  or g_104002_(_011110_, _011121_, _011123_);
  or g_104003_(_011103_, _011123_, _011124_);
  and g_104004_(_010908_, _011086_, _011125_);
  not g_104005_(_011125_, _011126_);
  or g_104006_(_010905_, _011086_, _011127_);
  not g_104007_(_011127_, _011128_);
  and g_104008_(_011126_, _011127_, _011129_);
  or g_104009_(_011125_, _011128_, _011130_);
  xor g_104010_(out[600], _009526_, _011132_);
  xor g_104011_(_055370_, _009526_, _011133_);
  and g_104012_(_011130_, _011132_, _011134_);
  and g_104013_(_011112_, _011119_, _011135_);
  and g_104014_(_011129_, _011133_, _011136_);
  or g_104015_(_011135_, _011136_, _011137_);
  or g_104016_(_011134_, _011137_, _011138_);
  xor g_104017_(_011130_, _011132_, _011139_);
  and g_104018_(_011102_, _011108_, _011140_);
  xor g_104019_(_011113_, _011118_, _011141_);
  and g_104020_(_011140_, _011141_, _011143_);
  and g_104021_(_011139_, _011143_, _011144_);
  or g_104022_(_011124_, _011138_, _011145_);
  xor g_104023_(out[599], _009524_, _011146_);
  xor g_104024_(_055282_, _009524_, _011147_);
  or g_104025_(_010935_, _011088_, _011148_);
  or g_104026_(_010938_, _011086_, _011149_);
  and g_104027_(_011148_, _011149_, _011150_);
  or g_104028_(_011146_, _011150_, _011151_);
  xor g_104029_(out[598], _009523_, _011152_);
  xor g_104030_(_055293_, _009523_, _011154_);
  or g_104031_(_010940_, _011088_, _011155_);
  or g_104032_(_010945_, _011086_, _011156_);
  and g_104033_(_011155_, _011156_, _011157_);
  and g_104034_(_011154_, _011157_, _011158_);
  and g_104035_(_011146_, _011150_, _011159_);
  xor g_104036_(_011146_, _011150_, _011160_);
  xor g_104037_(_011147_, _011150_, _011161_);
  xor g_104038_(_011154_, _011157_, _011162_);
  xor g_104039_(_011152_, _011157_, _011163_);
  and g_104040_(_011160_, _011162_, _011165_);
  or g_104041_(_011161_, _011163_, _011166_);
  xor g_104042_(out[597], _009521_, _011167_);
  xor g_104043_(_055304_, _009521_, _011168_);
  and g_104044_(_010956_, _011086_, _011169_);
  or g_104045_(_010954_, _011088_, _011170_);
  and g_104046_(_010962_, _011088_, _011171_);
  or g_104047_(_010961_, _011086_, _011172_);
  and g_104048_(_011170_, _011172_, _011173_);
  or g_104049_(_011169_, _011171_, _011174_);
  or g_104050_(_011168_, _011173_, _011176_);
  not g_104051_(_011176_, _011177_);
  or g_104052_(_022615_, _054791_, _011178_);
  not g_104053_(_011178_, _011179_);
  and g_104054_(_009522_, _011178_, _011180_);
  or g_104055_(_009521_, _011179_, _011181_);
  and g_104056_(_010975_, _011088_, _011182_);
  or g_104057_(_010974_, _011086_, _011183_);
  and g_104058_(_010969_, _011086_, _011184_);
  or g_104059_(_010968_, _011088_, _011185_);
  and g_104060_(_011183_, _011185_, _011187_);
  or g_104061_(_011182_, _011184_, _011188_);
  or g_104062_(_011181_, _011187_, _011189_);
  and g_104063_(_011176_, _011189_, _011190_);
  not g_104064_(_011190_, _011191_);
  and g_104065_(_011181_, _011187_, _011192_);
  or g_104066_(_011180_, _011188_, _011193_);
  and g_104067_(_011168_, _011173_, _011194_);
  or g_104068_(_011167_, _011174_, _011195_);
  and g_104069_(_011193_, _011195_, _011196_);
  or g_104070_(_011192_, _011194_, _011198_);
  and g_104071_(_011190_, _011196_, _011199_);
  or g_104072_(_011191_, _011198_, _011200_);
  and g_104073_(_011165_, _011199_, _011201_);
  or g_104074_(_011166_, _011200_, _011202_);
  and g_104075_(_011144_, _011201_, _011203_);
  or g_104076_(_011145_, _011202_, _011204_);
  or g_104077_(_055194_, _011088_, _011205_);
  or g_104078_(_011017_, _011086_, _011206_);
  and g_104079_(_011205_, _011206_, _011207_);
  and g_104080_(out[576], _011086_, _011209_);
  not g_104081_(_011209_, _011210_);
  or g_104082_(_011025_, _011086_, _011211_);
  not g_104083_(_011211_, _011212_);
  and g_104084_(_011210_, _011211_, _011213_);
  or g_104085_(_011209_, _011212_, _011214_);
  and g_104086_(out[592], _011213_, _011215_);
  or g_104087_(_055337_, _011214_, _011216_);
  and g_104088_(out[593], _011207_, _011217_);
  not g_104089_(_011217_, _011218_);
  xor g_104090_(out[593], _011207_, _011220_);
  xor g_104091_(_055326_, _011207_, _011221_);
  and g_104092_(_011216_, _011220_, _011222_);
  or g_104093_(_011215_, _011221_, _011223_);
  or g_104094_(_054572_, _011088_, _011224_);
  or g_104095_(_010997_, _011086_, _011225_);
  and g_104096_(_011224_, _011225_, _011226_);
  not g_104097_(_011226_, _011227_);
  and g_104098_(_054792_, _011226_, _011228_);
  or g_104099_(_054793_, _011227_, _011229_);
  xor g_104100_(out[595], _054791_, _011231_);
  xor g_104101_(_055359_, _054791_, _011232_);
  or g_104102_(_011003_, _011088_, _011233_);
  or g_104103_(_011008_, _011086_, _011234_);
  and g_104104_(_011233_, _011234_, _011235_);
  not g_104105_(_011235_, _011236_);
  and g_104106_(_011231_, _011235_, _011237_);
  or g_104107_(_011232_, _011236_, _011238_);
  and g_104108_(_011229_, _011238_, _011239_);
  or g_104109_(_011228_, _011237_, _011240_);
  or g_104110_(out[592], _011213_, _011242_);
  or g_104111_(_054792_, _011226_, _011243_);
  and g_104112_(_011232_, _011236_, _011244_);
  or g_104113_(_011231_, _011235_, _011245_);
  xor g_104114_(_054793_, _011226_, _011246_);
  or g_104115_(_011237_, _011246_, _011247_);
  and g_104116_(_011242_, _011245_, _011248_);
  not g_104117_(_011248_, _011249_);
  or g_104118_(_011247_, _011249_, _011250_);
  or g_104119_(_011223_, _011250_, _011251_);
  or g_104120_(_011204_, _011251_, _011253_);
  not g_104121_(_011253_, _011254_);
  and g_104122_(_011218_, _011223_, _011255_);
  or g_104123_(_011217_, _011222_, _011256_);
  and g_104124_(_011243_, _011256_, _011257_);
  or g_104125_(_011247_, _011255_, _011258_);
  and g_104126_(_011239_, _011258_, _011259_);
  or g_104127_(_011240_, _011257_, _011260_);
  and g_104128_(_011203_, _011260_, _011261_);
  or g_104129_(_011204_, _011259_, _011262_);
  and g_104130_(_011245_, _011261_, _011264_);
  or g_104131_(_011244_, _011262_, _011265_);
  and g_104132_(_011165_, _011198_, _011266_);
  or g_104133_(_011166_, _011196_, _011267_);
  and g_104134_(_011176_, _011266_, _011268_);
  or g_104135_(_011177_, _011267_, _011269_);
  and g_104136_(_011151_, _011158_, _011270_);
  or g_104137_(_011159_, _011270_, _011271_);
  not g_104138_(_011271_, _011272_);
  and g_104139_(_011269_, _011272_, _011273_);
  or g_104140_(_011268_, _011271_, _011275_);
  and g_104141_(_011144_, _011275_, _011276_);
  or g_104142_(_011145_, _011273_, _011277_);
  and g_104143_(_011103_, _011105_, _011278_);
  and g_104144_(_011137_, _011140_, _011279_);
  and g_104145_(_011122_, _011279_, _011280_);
  or g_104146_(_011278_, _011280_, _011281_);
  not g_104147_(_011281_, _011282_);
  and g_104148_(_011277_, _011282_, _011283_);
  or g_104149_(_011276_, _011281_, _011284_);
  and g_104150_(_011265_, _011283_, _011286_);
  or g_104151_(_011264_, _011284_, _011287_);
  and g_104152_(_011253_, _011287_, _011288_);
  or g_104153_(_011254_, _011286_, _011289_);
  or g_104154_(_011093_, _011288_, _011290_);
  not g_104155_(_011290_, _011291_);
  and g_104156_(_011095_, _011288_, _011292_);
  not g_104157_(_011292_, _011293_);
  and g_104158_(_011290_, _011293_, _011294_);
  or g_104159_(_011291_, _011292_, _011295_);
  xor g_104160_(out[618], _009543_, _011297_);
  not g_104161_(_011297_, _011298_);
  and g_104162_(_009532_, _009546_, _011299_);
  or g_104163_(_009533_, _009545_, _011300_);
  and g_104164_(_009533_, _009545_, _011301_);
  or g_104165_(_009532_, _009546_, _011302_);
  and g_104166_(_011300_, _011302_, _011303_);
  or g_104167_(_011299_, _011301_, _011304_);
  and g_104168_(_011294_, _011297_, _011305_);
  or g_104169_(_011295_, _011298_, _011306_);
  xor g_104170_(_011294_, _011297_, _011308_);
  xor g_104171_(_011295_, _011297_, _011309_);
  and g_104172_(_011303_, _011308_, _011310_);
  or g_104173_(_011304_, _011309_, _011311_);
  and g_104174_(_011133_, _011288_, _011312_);
  or g_104175_(_011132_, _011289_, _011313_);
  and g_104176_(_011130_, _011289_, _011314_);
  or g_104177_(_011129_, _011288_, _011315_);
  and g_104178_(_011313_, _011315_, _011316_);
  or g_104179_(_011312_, _011314_, _011317_);
  xor g_104180_(out[616], _009541_, _011319_);
  xor g_104181_(_055502_, _009541_, _011320_);
  and g_104182_(out[617], _009542_, _011321_);
  xor g_104183_(out[617], _009542_, _011322_);
  xor g_104184_(_055513_, _009542_, _011323_);
  or g_104185_(_011118_, _011288_, _011324_);
  or g_104186_(_011112_, _011289_, _011325_);
  and g_104187_(_011324_, _011325_, _011326_);
  and g_104188_(_011323_, _011326_, _011327_);
  or g_104189_(_011317_, _011319_, _011328_);
  or g_104190_(_011323_, _011326_, _011330_);
  and g_104191_(_011328_, _011330_, _011331_);
  xor g_104192_(_011317_, _011319_, _011332_);
  xor g_104193_(_011316_, _011319_, _011333_);
  xor g_104194_(_011323_, _011326_, _011334_);
  xor g_104195_(_011322_, _011326_, _011335_);
  and g_104196_(_011310_, _011334_, _011336_);
  or g_104197_(_011311_, _011335_, _011337_);
  and g_104198_(_011332_, _011336_, _011338_);
  or g_104199_(_011333_, _011337_, _011339_);
  xor g_104200_(out[615], _009540_, _011341_);
  xor g_104201_(_055414_, _009540_, _011342_);
  or g_104202_(_011147_, _011289_, _011343_);
  or g_104203_(_011150_, _011288_, _011344_);
  and g_104204_(_011343_, _011344_, _011345_);
  and g_104205_(_011341_, _011345_, _011346_);
  or g_104206_(_011341_, _011345_, _011347_);
  xor g_104207_(_011341_, _011345_, _011348_);
  xor g_104208_(_011342_, _011345_, _011349_);
  xor g_104209_(out[614], _009539_, _011350_);
  xor g_104210_(_055425_, _009539_, _011352_);
  or g_104211_(_011152_, _011289_, _011353_);
  or g_104212_(_011157_, _011288_, _011354_);
  and g_104213_(_011353_, _011354_, _011355_);
  and g_104214_(_011352_, _011355_, _011356_);
  xor g_104215_(_011352_, _011355_, _011357_);
  xor g_104216_(_011350_, _011355_, _011358_);
  and g_104217_(_011348_, _011357_, _011359_);
  or g_104218_(_011349_, _011358_, _011360_);
  or g_104219_(_022769_, _054977_, _011361_);
  not g_104220_(_011361_, _011363_);
  and g_104221_(_009538_, _011361_, _011364_);
  or g_104222_(_009537_, _011363_, _011365_);
  or g_104223_(_011187_, _011288_, _011366_);
  not g_104224_(_011366_, _011367_);
  and g_104225_(_011181_, _011288_, _011368_);
  not g_104226_(_011368_, _011369_);
  and g_104227_(_011366_, _011369_, _011370_);
  or g_104228_(_011367_, _011368_, _011371_);
  and g_104229_(_011365_, _011370_, _011372_);
  or g_104230_(_011364_, _011371_, _011374_);
  xor g_104231_(out[613], _009537_, _011375_);
  xor g_104232_(_055436_, _009537_, _011376_);
  and g_104233_(_011168_, _011288_, _011377_);
  not g_104234_(_011377_, _011378_);
  or g_104235_(_011173_, _011288_, _011379_);
  not g_104236_(_011379_, _011380_);
  and g_104237_(_011378_, _011379_, _011381_);
  or g_104238_(_011377_, _011380_, _011382_);
  and g_104239_(_011376_, _011381_, _011383_);
  or g_104240_(_011375_, _011382_, _011385_);
  and g_104241_(_011374_, _011385_, _011386_);
  or g_104242_(_011372_, _011383_, _011387_);
  and g_104243_(_011375_, _011382_, _011388_);
  or g_104244_(_011376_, _011381_, _011389_);
  and g_104245_(_011364_, _011371_, _011390_);
  or g_104246_(_011365_, _011370_, _011391_);
  and g_104247_(_011389_, _011391_, _011392_);
  or g_104248_(_011388_, _011390_, _011393_);
  and g_104249_(_011386_, _011392_, _011394_);
  or g_104250_(_011387_, _011393_, _011396_);
  or g_104251_(_011360_, _011396_, _011397_);
  and g_104252_(_011338_, _011394_, _011398_);
  and g_104253_(_011359_, _011398_, _011399_);
  or g_104254_(_011339_, _011397_, _011400_);
  xor g_104255_(out[611], _054977_, _011401_);
  xor g_104256_(_055491_, _054977_, _011402_);
  or g_104257_(_011232_, _011289_, _011403_);
  or g_104258_(_011235_, _011288_, _011404_);
  and g_104259_(_011403_, _011404_, _011405_);
  and g_104260_(_011401_, _011405_, _011407_);
  or g_104261_(_011226_, _011288_, _011408_);
  or g_104262_(_054793_, _011289_, _011409_);
  and g_104263_(_011408_, _011409_, _011410_);
  and g_104264_(_054978_, _011410_, _011411_);
  or g_104265_(_011407_, _011411_, _011412_);
  or g_104266_(_011401_, _011405_, _011413_);
  xor g_104267_(_011401_, _011405_, _011414_);
  xor g_104268_(_011402_, _011405_, _011415_);
  xor g_104269_(_054978_, _011410_, _011416_);
  xor g_104270_(_054979_, _011410_, _011418_);
  and g_104271_(_011414_, _011416_, _011419_);
  or g_104272_(_011415_, _011418_, _011420_);
  or g_104273_(_055326_, _011289_, _011421_);
  or g_104274_(_011207_, _011288_, _011422_);
  and g_104275_(_011421_, _011422_, _011423_);
  and g_104276_(out[609], _011423_, _011424_);
  not g_104277_(_011424_, _011425_);
  and g_104278_(out[592], _011288_, _011426_);
  not g_104279_(_011426_, _011427_);
  or g_104280_(_011213_, _011288_, _011429_);
  not g_104281_(_011429_, _011430_);
  and g_104282_(_011427_, _011429_, _011431_);
  or g_104283_(_011426_, _011430_, _011432_);
  and g_104284_(out[608], _011431_, _011433_);
  or g_104285_(_055469_, _011432_, _011434_);
  xor g_104286_(out[609], _011423_, _011435_);
  xor g_104287_(_055458_, _011423_, _011436_);
  and g_104288_(_011434_, _011435_, _011437_);
  or g_104289_(_011433_, _011436_, _011438_);
  and g_104290_(_011425_, _011438_, _011440_);
  or g_104291_(_011424_, _011437_, _011441_);
  and g_104292_(_011419_, _011441_, _011442_);
  or g_104293_(_011420_, _011440_, _011443_);
  and g_104294_(_011412_, _011413_, _011444_);
  not g_104295_(_011444_, _011445_);
  and g_104296_(_011443_, _011445_, _011446_);
  or g_104297_(_011442_, _011444_, _011447_);
  and g_104298_(_011399_, _011447_, _011448_);
  or g_104299_(_011400_, _011446_, _011449_);
  and g_104300_(_011359_, _011387_, _011451_);
  and g_104301_(_011389_, _011451_, _011452_);
  and g_104302_(_011347_, _011356_, _011453_);
  or g_104303_(_011346_, _011453_, _011454_);
  or g_104304_(_011452_, _011454_, _011455_);
  and g_104305_(_011338_, _011455_, _011456_);
  not g_104306_(_011456_, _011457_);
  or g_104307_(_011311_, _011331_, _011458_);
  or g_104308_(_011327_, _011458_, _011459_);
  not g_104309_(_011459_, _011460_);
  and g_104310_(_011302_, _011305_, _011462_);
  or g_104311_(_011301_, _011306_, _011463_);
  and g_104312_(_011300_, _011463_, _011464_);
  or g_104313_(_011299_, _011462_, _011465_);
  and g_104314_(_011449_, _011464_, _011466_);
  or g_104315_(_011448_, _011465_, _011467_);
  and g_104316_(_011457_, _011459_, _011468_);
  or g_104317_(_011456_, _011460_, _011469_);
  and g_104318_(_011466_, _011468_, _011470_);
  or g_104319_(_011467_, _011469_, _011471_);
  or g_104320_(out[608], _011431_, _011473_);
  and g_104321_(_011399_, _011473_, _011474_);
  not g_104322_(_011474_, _011475_);
  and g_104323_(_011437_, _011474_, _011476_);
  or g_104324_(_011438_, _011475_, _011477_);
  and g_104325_(_011419_, _011476_, _011478_);
  or g_104326_(_011420_, _011477_, _011479_);
  and g_104327_(_011471_, _011479_, _011480_);
  or g_104328_(_011470_, _011478_, _011481_);
  and g_104329_(_011295_, _011481_, _011482_);
  or g_104330_(_011294_, _011480_, _011484_);
  and g_104331_(_011297_, _011480_, _011485_);
  or g_104332_(_011298_, _011481_, _011486_);
  and g_104333_(_011484_, _011486_, _011487_);
  or g_104334_(_011482_, _011485_, _011488_);
  xor g_104335_(out[634], _009559_, _011489_);
  xor g_104336_(_055656_, _009559_, _011490_);
  and g_104337_(_011487_, _011489_, _011491_);
  or g_104338_(_011488_, _011490_, _011492_);
  and g_104339_(_009548_, _009563_, _011493_);
  or g_104340_(_009549_, _009562_, _011495_);
  and g_104341_(_011492_, _011495_, _011496_);
  or g_104342_(_011491_, _011493_, _011497_);
  and g_104343_(_009549_, _009562_, _011498_);
  or g_104344_(_009548_, _009563_, _011499_);
  and g_104345_(_011488_, _011490_, _011500_);
  or g_104346_(_011487_, _011489_, _011501_);
  and g_104347_(_011499_, _011501_, _011502_);
  or g_104348_(_011498_, _011500_, _011503_);
  and g_104349_(out[633], _009557_, _011504_);
  xor g_104350_(out[633], _009557_, _011506_);
  or g_104351_(_009560_, _011504_, _011507_);
  or g_104352_(_011326_, _011480_, _011508_);
  not g_104353_(_011508_, _011509_);
  and g_104354_(_011323_, _011480_, _011510_);
  not g_104355_(_011510_, _011511_);
  and g_104356_(_011508_, _011511_, _011512_);
  or g_104357_(_011509_, _011510_, _011513_);
  and g_104358_(_011507_, _011512_, _011514_);
  or g_104359_(_011506_, _011513_, _011515_);
  and g_104360_(_011502_, _011515_, _011517_);
  or g_104361_(_011503_, _011514_, _011518_);
  and g_104362_(_011496_, _011517_, _011519_);
  or g_104363_(_011497_, _011518_, _011520_);
  and g_104364_(_011320_, _011480_, _011521_);
  not g_104365_(_011521_, _011522_);
  or g_104366_(_011316_, _011480_, _011523_);
  not g_104367_(_011523_, _011524_);
  and g_104368_(_011522_, _011523_, _011525_);
  or g_104369_(_011521_, _011524_, _011526_);
  xor g_104370_(out[632], _009556_, _011528_);
  xor g_104371_(_055634_, _009556_, _011529_);
  and g_104372_(_011526_, _011528_, _011530_);
  or g_104373_(_011525_, _011529_, _011531_);
  and g_104374_(_011506_, _011513_, _011532_);
  or g_104375_(_011507_, _011512_, _011533_);
  and g_104376_(_011525_, _011529_, _011534_);
  or g_104377_(_011526_, _011528_, _011535_);
  and g_104378_(_011533_, _011535_, _011536_);
  or g_104379_(_011532_, _011534_, _011537_);
  and g_104380_(_011531_, _011536_, _011539_);
  or g_104381_(_011530_, _011537_, _011540_);
  and g_104382_(_011519_, _011539_, _011541_);
  or g_104383_(_011520_, _011540_, _011542_);
  xor g_104384_(out[630], _009554_, _011543_);
  xor g_104385_(_055557_, _009554_, _011544_);
  and g_104386_(_011352_, _011480_, _011545_);
  not g_104387_(_011545_, _011546_);
  or g_104388_(_011355_, _011480_, _011547_);
  not g_104389_(_011547_, _011548_);
  and g_104390_(_011546_, _011547_, _011550_);
  or g_104391_(_011545_, _011548_, _011551_);
  and g_104392_(_011544_, _011550_, _011552_);
  or g_104393_(_011543_, _011551_, _011553_);
  xor g_104394_(_011544_, _011550_, _011554_);
  xor g_104395_(_011543_, _011550_, _011555_);
  xor g_104396_(out[631], _009555_, _011556_);
  xor g_104397_(_055546_, _009555_, _011557_);
  and g_104398_(_011341_, _011480_, _011558_);
  not g_104399_(_011558_, _011559_);
  or g_104400_(_011345_, _011480_, _011561_);
  not g_104401_(_011561_, _011562_);
  and g_104402_(_011559_, _011561_, _011563_);
  or g_104403_(_011558_, _011562_, _011564_);
  and g_104404_(_011556_, _011563_, _011565_);
  or g_104405_(_011557_, _011564_, _011566_);
  and g_104406_(_011557_, _011564_, _011567_);
  or g_104407_(_011556_, _011563_, _011568_);
  and g_104408_(_011554_, _011566_, _011569_);
  or g_104409_(_011555_, _011565_, _011570_);
  and g_104410_(_011568_, _011569_, _011572_);
  or g_104411_(_011567_, _011570_, _011573_);
  or g_104412_(_022923_, _055090_, _011574_);
  not g_104413_(_011574_, _011575_);
  and g_104414_(_009553_, _011574_, _011576_);
  or g_104415_(_009552_, _011575_, _011577_);
  or g_104416_(_011370_, _011480_, _011578_);
  not g_104417_(_011578_, _011579_);
  and g_104418_(_011365_, _011480_, _011580_);
  not g_104419_(_011580_, _011581_);
  and g_104420_(_011578_, _011581_, _011583_);
  or g_104421_(_011579_, _011580_, _011584_);
  and g_104422_(_011577_, _011583_, _011585_);
  or g_104423_(_011576_, _011584_, _011586_);
  xor g_104424_(out[629], _009552_, _011587_);
  xor g_104425_(_055568_, _009552_, _011588_);
  and g_104426_(_011376_, _011480_, _011589_);
  not g_104427_(_011589_, _011590_);
  or g_104428_(_011381_, _011480_, _011591_);
  not g_104429_(_011591_, _011592_);
  and g_104430_(_011590_, _011591_, _011594_);
  or g_104431_(_011589_, _011592_, _011595_);
  and g_104432_(_011588_, _011594_, _011596_);
  or g_104433_(_011587_, _011595_, _011597_);
  and g_104434_(_011586_, _011597_, _011598_);
  or g_104435_(_011585_, _011596_, _011599_);
  and g_104436_(_011587_, _011595_, _011600_);
  or g_104437_(_011588_, _011594_, _011601_);
  and g_104438_(_011576_, _011584_, _011602_);
  or g_104439_(_011577_, _011583_, _011603_);
  and g_104440_(_011601_, _011603_, _011605_);
  or g_104441_(_011600_, _011602_, _011606_);
  and g_104442_(_011598_, _011605_, _011607_);
  or g_104443_(_011599_, _011606_, _011608_);
  and g_104444_(_011572_, _011607_, _011609_);
  or g_104445_(_011573_, _011608_, _011610_);
  and g_104446_(_011541_, _011609_, _011611_);
  or g_104447_(_011542_, _011610_, _011612_);
  xor g_104448_(out[627], _055090_, _011613_);
  xor g_104449_(_055623_, _055090_, _011614_);
  and g_104450_(_011401_, _011480_, _011616_);
  not g_104451_(_011616_, _011617_);
  or g_104452_(_011405_, _011480_, _011618_);
  not g_104453_(_011618_, _011619_);
  and g_104454_(_011617_, _011618_, _011620_);
  or g_104455_(_011616_, _011619_, _011621_);
  and g_104456_(_011613_, _011620_, _011622_);
  or g_104457_(_011410_, _011480_, _011623_);
  not g_104458_(_011623_, _011624_);
  and g_104459_(_054978_, _011480_, _011625_);
  not g_104460_(_011625_, _011627_);
  and g_104461_(_011623_, _011627_, _011628_);
  or g_104462_(_011624_, _011625_, _011629_);
  and g_104463_(_055091_, _011628_, _011630_);
  or g_104464_(_011622_, _011630_, _011631_);
  and g_104465_(_011614_, _011621_, _011632_);
  or g_104466_(_011613_, _011620_, _011633_);
  and g_104467_(_055092_, _011629_, _011634_);
  or g_104468_(_011632_, _011634_, _011635_);
  xor g_104469_(_011613_, _011620_, _011636_);
  xor g_104470_(_055091_, _011628_, _011638_);
  and g_104471_(_011636_, _011638_, _011639_);
  or g_104472_(_011631_, _011635_, _011640_);
  and g_104473_(out[609], _011480_, _011641_);
  not g_104474_(_011641_, _011642_);
  or g_104475_(_011423_, _011480_, _011643_);
  not g_104476_(_011643_, _011644_);
  and g_104477_(_011642_, _011643_, _011645_);
  or g_104478_(_011641_, _011644_, _011646_);
  and g_104479_(out[625], _011645_, _011647_);
  and g_104480_(out[608], _011480_, _011649_);
  not g_104481_(_011649_, _011650_);
  or g_104482_(_011431_, _011480_, _011651_);
  not g_104483_(_011651_, _011652_);
  and g_104484_(_011650_, _011651_, _011653_);
  or g_104485_(_011649_, _011652_, _011654_);
  and g_104486_(out[624], _011653_, _011655_);
  or g_104487_(_055601_, _011654_, _011656_);
  xor g_104488_(out[625], _011645_, _011657_);
  xor g_104489_(_055590_, _011645_, _011658_);
  and g_104490_(_011656_, _011657_, _011660_);
  or g_104491_(_011655_, _011658_, _011661_);
  or g_104492_(_011647_, _011660_, _011662_);
  and g_104493_(_011639_, _011662_, _011663_);
  and g_104494_(_011631_, _011633_, _011664_);
  or g_104495_(_011663_, _011664_, _011665_);
  not g_104496_(_011665_, _011666_);
  and g_104497_(_011611_, _011665_, _011667_);
  or g_104498_(_011612_, _011666_, _011668_);
  and g_104499_(_011599_, _011601_, _011669_);
  or g_104500_(_011598_, _011600_, _011671_);
  and g_104501_(_011572_, _011669_, _011672_);
  or g_104502_(_011573_, _011671_, _011673_);
  and g_104503_(_011552_, _011568_, _011674_);
  or g_104504_(_011553_, _011567_, _011675_);
  and g_104505_(_011566_, _011675_, _011676_);
  or g_104506_(_011565_, _011674_, _011677_);
  and g_104507_(_011673_, _011676_, _011678_);
  or g_104508_(_011672_, _011677_, _011679_);
  and g_104509_(_011541_, _011679_, _011680_);
  or g_104510_(_011542_, _011678_, _011682_);
  and g_104511_(_011497_, _011499_, _011683_);
  or g_104512_(_011496_, _011498_, _011684_);
  and g_104513_(_011519_, _011537_, _011685_);
  or g_104514_(_011520_, _011536_, _011686_);
  and g_104515_(_011684_, _011686_, _011687_);
  or g_104516_(_011683_, _011685_, _011688_);
  and g_104517_(_011682_, _011687_, _011689_);
  or g_104518_(_011680_, _011688_, _011690_);
  and g_104519_(_011668_, _011689_, _011691_);
  or g_104520_(_011667_, _011690_, _011693_);
  and g_104521_(_055601_, _011654_, _011694_);
  or g_104522_(out[624], _011653_, _011695_);
  and g_104523_(_011639_, _011695_, _011696_);
  or g_104524_(_011640_, _011694_, _011697_);
  and g_104525_(_011660_, _011696_, _011698_);
  or g_104526_(_011661_, _011697_, _011699_);
  and g_104527_(_011611_, _011698_, _011700_);
  or g_104528_(_011612_, _011699_, _011701_);
  and g_104529_(_011693_, _011701_, _011702_);
  or g_104530_(_011691_, _011700_, _011704_);
  and g_104531_(_011488_, _011704_, _011705_);
  or g_104532_(_011487_, _011702_, _011706_);
  and g_104533_(_011489_, _011702_, _011707_);
  or g_104534_(_011490_, _011704_, _011708_);
  and g_104535_(_011706_, _011708_, _011709_);
  or g_104536_(_011705_, _011707_, _011710_);
  xor g_104537_(out[643], _055356_, _011711_);
  xor g_104538_(_055755_, _055356_, _011712_);
  and g_104539_(_011613_, _011702_, _011713_);
  or g_104540_(_011614_, _011704_, _011715_);
  and g_104541_(_011621_, _011704_, _011716_);
  or g_104542_(_011620_, _011702_, _011717_);
  and g_104543_(_011715_, _011717_, _011718_);
  or g_104544_(_011713_, _011716_, _011719_);
  and g_104545_(_011711_, _011718_, _011720_);
  or g_104546_(_011712_, _011719_, _011721_);
  and g_104547_(_011629_, _011704_, _011722_);
  or g_104548_(_011628_, _011702_, _011723_);
  and g_104549_(_055091_, _011702_, _011724_);
  or g_104550_(_055092_, _011704_, _011726_);
  and g_104551_(_011723_, _011726_, _011727_);
  or g_104552_(_011722_, _011724_, _011728_);
  and g_104553_(_055357_, _011727_, _011729_);
  or g_104554_(_055358_, _011728_, _011730_);
  and g_104555_(_011721_, _011730_, _011731_);
  or g_104556_(_011720_, _011729_, _011732_);
  and g_104557_(_011712_, _011719_, _011733_);
  or g_104558_(_011711_, _011718_, _011734_);
  and g_104559_(_055358_, _011728_, _011735_);
  or g_104560_(_055357_, _011727_, _011737_);
  and g_104561_(_011734_, _011737_, _011738_);
  or g_104562_(_011733_, _011735_, _011739_);
  and g_104563_(_011731_, _011738_, _011740_);
  or g_104564_(_011732_, _011739_, _011741_);
  and g_104565_(out[625], _011702_, _011742_);
  or g_104566_(_055590_, _011704_, _011743_);
  and g_104567_(_011646_, _011704_, _011744_);
  or g_104568_(_011645_, _011702_, _011745_);
  and g_104569_(_011743_, _011745_, _011746_);
  or g_104570_(_011742_, _011744_, _011748_);
  and g_104571_(out[641], _011746_, _011749_);
  or g_104572_(_055722_, _011748_, _011750_);
  and g_104573_(out[624], _011702_, _011751_);
  or g_104574_(_055601_, _011704_, _011752_);
  and g_104575_(_011654_, _011704_, _011753_);
  or g_104576_(_011653_, _011702_, _011754_);
  and g_104577_(_011752_, _011754_, _011755_);
  or g_104578_(_011751_, _011753_, _011756_);
  and g_104579_(out[640], _011755_, _011757_);
  or g_104580_(_055733_, _011756_, _011759_);
  xor g_104581_(out[641], _011746_, _011760_);
  xor g_104582_(_055722_, _011746_, _011761_);
  and g_104583_(_011759_, _011760_, _011762_);
  or g_104584_(_011757_, _011761_, _011763_);
  and g_104585_(_011750_, _011763_, _011764_);
  or g_104586_(_011749_, _011762_, _011765_);
  and g_104587_(_011740_, _011765_, _011766_);
  or g_104588_(_011741_, _011764_, _011767_);
  and g_104589_(_011732_, _011734_, _011768_);
  or g_104590_(_011731_, _011733_, _011770_);
  and g_104591_(_011767_, _011770_, _011771_);
  or g_104592_(_011766_, _011768_, _011772_);
  or g_104593_(_009565_, _009577_, _011773_);
  xor g_104594_(out[650], _009575_, _011774_);
  not g_104595_(_011774_, _011775_);
  or g_104596_(_011710_, _011775_, _011776_);
  and g_104597_(_011773_, _011776_, _011777_);
  and g_104598_(_009565_, _009577_, _011778_);
  or g_104599_(_009564_, _009578_, _011779_);
  or g_104600_(_011709_, _011774_, _011781_);
  and g_104601_(_011779_, _011781_, _011782_);
  xor g_104602_(_009564_, _009577_, _011783_);
  xor g_104603_(_011710_, _011774_, _011784_);
  and g_104604_(_011777_, _011782_, _011785_);
  or g_104605_(_011783_, _011784_, _011786_);
  xor g_104606_(out[648], _009573_, _011787_);
  xor g_104607_(_055766_, _009573_, _011788_);
  and g_104608_(_011529_, _011702_, _011789_);
  or g_104609_(_011528_, _011704_, _011790_);
  and g_104610_(_011526_, _011704_, _011792_);
  or g_104611_(_011525_, _011702_, _011793_);
  and g_104612_(_011790_, _011793_, _011794_);
  or g_104613_(_011789_, _011792_, _011795_);
  and g_104614_(_011788_, _011794_, _011796_);
  or g_104615_(_011787_, _011795_, _011797_);
  and g_104616_(out[649], _009574_, _011798_);
  xor g_104617_(out[649], _009574_, _011799_);
  xor g_104618_(_055777_, _009574_, _011800_);
  and g_104619_(_011513_, _011704_, _011801_);
  or g_104620_(_011512_, _011702_, _011803_);
  and g_104621_(_011507_, _011702_, _011804_);
  or g_104622_(_011506_, _011704_, _011805_);
  and g_104623_(_011803_, _011805_, _011806_);
  or g_104624_(_011801_, _011804_, _011807_);
  and g_104625_(_011799_, _011807_, _011808_);
  or g_104626_(_011800_, _011806_, _011809_);
  and g_104627_(_011797_, _011809_, _011810_);
  or g_104628_(_011796_, _011808_, _011811_);
  and g_104629_(_011800_, _011806_, _011812_);
  or g_104630_(_011799_, _011807_, _011814_);
  and g_104631_(_011787_, _011795_, _011815_);
  or g_104632_(_011788_, _011794_, _011816_);
  and g_104633_(_011814_, _011816_, _011817_);
  or g_104634_(_011812_, _011815_, _011818_);
  and g_104635_(_011810_, _011817_, _011819_);
  or g_104636_(_011786_, _011818_, _011820_);
  and g_104637_(_011785_, _011819_, _011821_);
  or g_104638_(_011811_, _011820_, _011822_);
  xor g_104639_(out[646], _009571_, _011823_);
  not g_104640_(_011823_, _011825_);
  or g_104641_(_011543_, _011704_, _011826_);
  or g_104642_(_011550_, _011702_, _011827_);
  and g_104643_(_011826_, _011827_, _011828_);
  and g_104644_(_011825_, _011828_, _011829_);
  xor g_104645_(_011825_, _011828_, _011830_);
  xor g_104646_(_011823_, _011828_, _011831_);
  xor g_104647_(out[647], _009572_, _011832_);
  xor g_104648_(_055678_, _009572_, _011833_);
  or g_104649_(_011557_, _011704_, _011834_);
  or g_104650_(_011563_, _011702_, _011836_);
  and g_104651_(_011834_, _011836_, _011837_);
  and g_104652_(_011832_, _011837_, _011838_);
  or g_104653_(_011832_, _011837_, _011839_);
  xor g_104654_(_011832_, _011837_, _011840_);
  xor g_104655_(_011833_, _011837_, _011841_);
  and g_104656_(_011830_, _011840_, _011842_);
  or g_104657_(_011831_, _011841_, _011843_);
  or g_104658_(_023077_, _055356_, _011844_);
  not g_104659_(_011844_, _011845_);
  and g_104660_(_009570_, _011844_, _011847_);
  or g_104661_(_009568_, _011845_, _011848_);
  and g_104662_(_011584_, _011704_, _011849_);
  or g_104663_(_011583_, _011702_, _011850_);
  and g_104664_(_011577_, _011702_, _011851_);
  or g_104665_(_011576_, _011704_, _011852_);
  and g_104666_(_011850_, _011852_, _011853_);
  or g_104667_(_011849_, _011851_, _011854_);
  or g_104668_(_011847_, _011854_, _011855_);
  xor g_104669_(out[645], _009568_, _011856_);
  xor g_104670_(_055700_, _009568_, _011858_);
  and g_104671_(_011588_, _011702_, _011859_);
  or g_104672_(_011587_, _011704_, _011860_);
  and g_104673_(_011595_, _011704_, _011861_);
  or g_104674_(_011594_, _011702_, _011862_);
  and g_104675_(_011860_, _011862_, _011863_);
  or g_104676_(_011859_, _011861_, _011864_);
  or g_104677_(_011856_, _011864_, _011865_);
  and g_104678_(_011855_, _011865_, _011866_);
  and g_104679_(_011856_, _011864_, _011867_);
  or g_104680_(_011858_, _011863_, _011869_);
  or g_104681_(_011848_, _011853_, _011870_);
  xor g_104682_(_011847_, _011853_, _011871_);
  xor g_104683_(_011856_, _011863_, _011872_);
  or g_104684_(_011871_, _011872_, _011873_);
  or g_104685_(_011843_, _011873_, _011874_);
  and g_104686_(_011866_, _011869_, _011875_);
  and g_104687_(_011842_, _011870_, _011876_);
  and g_104688_(_011821_, _011876_, _011877_);
  and g_104689_(_011875_, _011877_, _011878_);
  or g_104690_(_011822_, _011874_, _011880_);
  and g_104691_(_011772_, _011878_, _011881_);
  or g_104692_(_011771_, _011880_, _011882_);
  or g_104693_(_011843_, _011866_, _011883_);
  or g_104694_(_011867_, _011883_, _011884_);
  and g_104695_(_011829_, _011839_, _011885_);
  or g_104696_(_011838_, _011885_, _011886_);
  not g_104697_(_011886_, _011887_);
  and g_104698_(_011884_, _011887_, _011888_);
  or g_104699_(_011822_, _011888_, _011889_);
  or g_104700_(_011777_, _011778_, _011891_);
  or g_104701_(_011786_, _011810_, _011892_);
  or g_104702_(_011812_, _011892_, _011893_);
  and g_104703_(_011891_, _011893_, _011894_);
  and g_104704_(_011889_, _011894_, _011895_);
  not g_104705_(_011895_, _011896_);
  and g_104706_(_011882_, _011895_, _011897_);
  or g_104707_(_011881_, _011896_, _011898_);
  and g_104708_(_055733_, _011756_, _011899_);
  or g_104709_(out[640], _011755_, _011900_);
  and g_104710_(_011740_, _011900_, _011902_);
  or g_104711_(_011741_, _011899_, _011903_);
  and g_104712_(_011762_, _011902_, _011904_);
  or g_104713_(_011763_, _011903_, _011905_);
  and g_104714_(_011878_, _011904_, _011906_);
  or g_104715_(_011880_, _011905_, _011907_);
  and g_104716_(_011898_, _011907_, _011908_);
  or g_104717_(_011897_, _011906_, _011909_);
  and g_104718_(_011710_, _011909_, _011910_);
  or g_104719_(_011709_, _011908_, _011911_);
  and g_104720_(_011774_, _011908_, _011913_);
  or g_104721_(_011775_, _011909_, _011914_);
  and g_104722_(_011911_, _011914_, _011915_);
  or g_104723_(_011910_, _011913_, _011916_);
  xor g_104724_(out[666], _009590_, _011917_);
  not g_104725_(_011917_, _011918_);
  and g_104726_(_011915_, _011917_, _011919_);
  or g_104727_(_011916_, _011918_, _011920_);
  and g_104728_(_009579_, _009594_, _011921_);
  or g_104729_(_009581_, _009593_, _011922_);
  and g_104730_(_011920_, _011922_, _011924_);
  or g_104731_(_011919_, _011921_, _011925_);
  or g_104732_(_009579_, _009594_, _011926_);
  or g_104733_(_011915_, _011917_, _011927_);
  and g_104734_(_011926_, _011927_, _011928_);
  not g_104735_(_011928_, _011929_);
  and g_104736_(_011924_, _011928_, _011930_);
  or g_104737_(_011925_, _011929_, _011931_);
  xor g_104738_(out[664], _009588_, _011932_);
  xor g_104739_(_055898_, _009588_, _011933_);
  and g_104740_(_011788_, _011908_, _011935_);
  or g_104741_(_011787_, _011909_, _011936_);
  and g_104742_(_011795_, _011909_, _011937_);
  or g_104743_(_011794_, _011908_, _011938_);
  and g_104744_(_011936_, _011938_, _011939_);
  or g_104745_(_011935_, _011937_, _011940_);
  or g_104746_(_011932_, _011940_, _011941_);
  and g_104747_(out[665], _009589_, _011942_);
  xor g_104748_(out[665], _009589_, _011943_);
  xor g_104749_(_055909_, _009589_, _011944_);
  and g_104750_(_011807_, _011909_, _011946_);
  or g_104751_(_011806_, _011908_, _011947_);
  and g_104752_(_011800_, _011908_, _011948_);
  or g_104753_(_011799_, _011909_, _011949_);
  and g_104754_(_011947_, _011949_, _011950_);
  or g_104755_(_011946_, _011948_, _011951_);
  and g_104756_(_011943_, _011951_, _011952_);
  or g_104757_(_011944_, _011950_, _011953_);
  and g_104758_(_011941_, _011953_, _011954_);
  and g_104759_(_011944_, _011950_, _011955_);
  or g_104760_(_011943_, _011951_, _011957_);
  or g_104761_(_011933_, _011939_, _011958_);
  and g_104762_(_011957_, _011958_, _011959_);
  and g_104763_(_011954_, _011959_, _011960_);
  xor g_104764_(_011932_, _011939_, _011961_);
  or g_104765_(_011955_, _011961_, _011962_);
  or g_104766_(_011931_, _011952_, _011963_);
  and g_104767_(_011930_, _011960_, _011964_);
  or g_104768_(_011962_, _011963_, _011965_);
  xor g_104769_(out[662], _009586_, _011966_);
  xor g_104770_(_055821_, _009586_, _011968_);
  or g_104771_(_011823_, _011909_, _011969_);
  or g_104772_(_011828_, _011908_, _011970_);
  and g_104773_(_011969_, _011970_, _011971_);
  and g_104774_(_011968_, _011971_, _011972_);
  xor g_104775_(out[663], _009587_, _011973_);
  xor g_104776_(_055810_, _009587_, _011974_);
  or g_104777_(_011833_, _011909_, _011975_);
  or g_104778_(_011837_, _011908_, _011976_);
  and g_104779_(_011975_, _011976_, _011977_);
  or g_104780_(_011973_, _011977_, _011979_);
  and g_104781_(_011973_, _011977_, _011980_);
  xor g_104782_(_011968_, _011971_, _011981_);
  xor g_104783_(_011966_, _011971_, _011982_);
  xor g_104784_(_011973_, _011977_, _011983_);
  xor g_104785_(_011974_, _011977_, _011984_);
  and g_104786_(_011981_, _011983_, _011985_);
  or g_104787_(_011982_, _011984_, _011986_);
  or g_104788_(_023231_, _055437_, _011987_);
  not g_104789_(_011987_, _011988_);
  and g_104790_(_009585_, _011987_, _011990_);
  or g_104791_(_009584_, _011988_, _011991_);
  and g_104792_(_011854_, _011909_, _011992_);
  or g_104793_(_011853_, _011908_, _011993_);
  and g_104794_(_011848_, _011908_, _011994_);
  or g_104795_(_011847_, _011909_, _011995_);
  and g_104796_(_011993_, _011995_, _011996_);
  or g_104797_(_011992_, _011994_, _011997_);
  and g_104798_(_011991_, _011996_, _011998_);
  or g_104799_(_011990_, _011997_, _011999_);
  xor g_104800_(out[661], _009584_, _012001_);
  xor g_104801_(_055832_, _009584_, _012002_);
  and g_104802_(_011858_, _011908_, _012003_);
  or g_104803_(_011856_, _011909_, _012004_);
  and g_104804_(_011864_, _011909_, _012005_);
  or g_104805_(_011863_, _011908_, _012006_);
  and g_104806_(_012004_, _012006_, _012007_);
  or g_104807_(_012003_, _012005_, _012008_);
  and g_104808_(_012002_, _012007_, _012009_);
  or g_104809_(_012001_, _012008_, _012010_);
  and g_104810_(_011999_, _012010_, _012012_);
  or g_104811_(_011998_, _012009_, _012013_);
  and g_104812_(_012001_, _012008_, _012014_);
  or g_104813_(_012002_, _012007_, _012015_);
  and g_104814_(_011990_, _011997_, _012016_);
  or g_104815_(_011991_, _011996_, _012017_);
  and g_104816_(_012015_, _012017_, _012018_);
  or g_104817_(_012014_, _012016_, _012019_);
  and g_104818_(_012012_, _012018_, _012020_);
  or g_104819_(_012013_, _012019_, _012021_);
  and g_104820_(_011985_, _012020_, _012023_);
  or g_104821_(_011986_, _012021_, _012024_);
  and g_104822_(_011964_, _012023_, _012025_);
  or g_104823_(_011965_, _012024_, _012026_);
  or g_104824_(_055722_, _011909_, _012027_);
  or g_104825_(_011746_, _011908_, _012028_);
  and g_104826_(_012027_, _012028_, _012029_);
  or g_104827_(_055733_, _011909_, _012030_);
  or g_104828_(_011755_, _011908_, _012031_);
  and g_104829_(_012030_, _012031_, _012032_);
  and g_104830_(out[656], _012032_, _012034_);
  not g_104831_(_012034_, _012035_);
  and g_104832_(out[657], _012029_, _012036_);
  xor g_104833_(out[657], _012029_, _012037_);
  xor g_104834_(_055854_, _012029_, _012038_);
  and g_104835_(_012035_, _012037_, _012039_);
  or g_104836_(_012034_, _012038_, _012040_);
  or g_104837_(_055358_, _011909_, _012041_);
  or g_104838_(_011727_, _011908_, _012042_);
  and g_104839_(_012041_, _012042_, _012043_);
  and g_104840_(_055438_, _012043_, _012045_);
  xor g_104841_(_055438_, _012043_, _012046_);
  xor g_104842_(out[659], _055437_, _012047_);
  xor g_104843_(_055887_, _055437_, _012048_);
  or g_104844_(_011712_, _011909_, _012049_);
  or g_104845_(_011718_, _011908_, _012050_);
  and g_104846_(_012049_, _012050_, _012051_);
  not g_104847_(_012051_, _012052_);
  and g_104848_(_012048_, _012052_, _012053_);
  or g_104849_(_012047_, _012051_, _012054_);
  and g_104850_(_012047_, _012051_, _012056_);
  xor g_104851_(_012047_, _012051_, _012057_);
  or g_104852_(out[656], _012032_, _012058_);
  and g_104853_(_012057_, _012058_, _012059_);
  and g_104854_(_012046_, _012059_, _012060_);
  not g_104855_(_012060_, _012061_);
  and g_104856_(_012039_, _012060_, _012062_);
  or g_104857_(_012040_, _012061_, _012063_);
  and g_104858_(_012025_, _012062_, _012064_);
  or g_104859_(_012026_, _012063_, _012065_);
  or g_104860_(_012045_, _012056_, _012067_);
  or g_104861_(_012036_, _012039_, _012068_);
  and g_104862_(_012046_, _012068_, _012069_);
  or g_104863_(_012067_, _012069_, _012070_);
  not g_104864_(_012070_, _012071_);
  and g_104865_(_012025_, _012054_, _012072_);
  or g_104866_(_012026_, _012053_, _012073_);
  and g_104867_(_012070_, _012072_, _012074_);
  or g_104868_(_012071_, _012073_, _012075_);
  or g_104869_(_011986_, _012012_, _012076_);
  or g_104870_(_012014_, _012076_, _012078_);
  or g_104871_(_011972_, _011980_, _012079_);
  and g_104872_(_011979_, _012079_, _012080_);
  not g_104873_(_012080_, _012081_);
  and g_104874_(_012078_, _012081_, _012082_);
  or g_104875_(_011965_, _012082_, _012083_);
  or g_104876_(_011954_, _011955_, _012084_);
  or g_104877_(_011931_, _012084_, _012085_);
  and g_104878_(_011925_, _011926_, _012086_);
  not g_104879_(_012086_, _012087_);
  and g_104880_(_012083_, _012085_, _012089_);
  not g_104881_(_012089_, _012090_);
  and g_104882_(_012075_, _012089_, _012091_);
  or g_104883_(_012074_, _012090_, _012092_);
  and g_104884_(_012087_, _012091_, _012093_);
  or g_104885_(_012086_, _012092_, _012094_);
  and g_104886_(_012065_, _012094_, _012095_);
  or g_104887_(_012064_, _012093_, _012096_);
  or g_104888_(_011915_, _012095_, _012097_);
  not g_104889_(_012097_, _012098_);
  and g_104890_(_011917_, _012095_, _012100_);
  not g_104891_(_012100_, _012101_);
  and g_104892_(_012097_, _012101_, _012102_);
  or g_104893_(_012098_, _012100_, _012103_);
  xor g_104894_(out[682], _009606_, _012104_);
  not g_104895_(_012104_, _012105_);
  and g_104896_(_012102_, _012104_, _012106_);
  or g_104897_(_009596_, _009608_, _012107_);
  not g_104898_(_012107_, _012108_);
  or g_104899_(_009595_, _009609_, _012109_);
  and g_104900_(_012107_, _012109_, _012111_);
  xor g_104901_(_009595_, _009608_, _012112_);
  xor g_104902_(_012102_, _012104_, _012113_);
  xor g_104903_(_012103_, _012104_, _012114_);
  and g_104904_(_012111_, _012113_, _012115_);
  or g_104905_(_012112_, _012114_, _012116_);
  xor g_104906_(out[680], _009604_, _012117_);
  xor g_104907_(_000065_, _009604_, _012118_);
  and g_104908_(_011933_, _012095_, _012119_);
  or g_104909_(_011932_, _012096_, _012120_);
  and g_104910_(_011940_, _012096_, _012122_);
  or g_104911_(_011939_, _012095_, _012123_);
  and g_104912_(_012120_, _012123_, _012124_);
  or g_104913_(_012119_, _012122_, _012125_);
  and g_104914_(_012118_, _012124_, _012126_);
  and g_104915_(out[681], _009605_, _012127_);
  xor g_104916_(out[681], _009605_, _012128_);
  xor g_104917_(_000076_, _009605_, _012129_);
  and g_104918_(_011951_, _012096_, _012130_);
  or g_104919_(_011950_, _012095_, _012131_);
  and g_104920_(_011944_, _012095_, _012133_);
  or g_104921_(_011943_, _012096_, _012134_);
  and g_104922_(_012131_, _012134_, _012135_);
  or g_104923_(_012130_, _012133_, _012136_);
  and g_104924_(_012128_, _012136_, _012137_);
  or g_104925_(_012129_, _012135_, _012138_);
  or g_104926_(_012126_, _012137_, _012139_);
  and g_104927_(_012129_, _012135_, _012140_);
  or g_104928_(_012128_, _012136_, _012141_);
  and g_104929_(_012117_, _012125_, _012142_);
  or g_104930_(_012140_, _012142_, _012144_);
  or g_104931_(_012139_, _012144_, _012145_);
  xor g_104932_(_012118_, _012124_, _012146_);
  and g_104933_(_012141_, _012146_, _012147_);
  and g_104934_(_012115_, _012138_, _012148_);
  and g_104935_(_012147_, _012148_, _012149_);
  or g_104936_(_012116_, _012145_, _012150_);
  xor g_104937_(out[678], _009601_, _012151_);
  not g_104938_(_012151_, _012152_);
  and g_104939_(_011968_, _012095_, _012153_);
  or g_104940_(_011971_, _012095_, _012155_);
  not g_104941_(_012155_, _012156_);
  or g_104942_(_012153_, _012156_, _012157_);
  or g_104943_(_012151_, _012157_, _012158_);
  xor g_104944_(out[679], _009603_, _012159_);
  xor g_104945_(_055942_, _009603_, _012160_);
  and g_104946_(_011973_, _012095_, _012161_);
  not g_104947_(_012161_, _012162_);
  or g_104948_(_011977_, _012095_, _012163_);
  not g_104949_(_012163_, _012164_);
  and g_104950_(_012162_, _012163_, _012166_);
  or g_104951_(_012161_, _012164_, _012167_);
  or g_104952_(_012160_, _012167_, _012168_);
  and g_104953_(_012158_, _012168_, _012169_);
  and g_104954_(_012160_, _012167_, _012170_);
  xor g_104955_(_012151_, _012157_, _012171_);
  xor g_104956_(_012152_, _012157_, _012172_);
  xor g_104957_(_012159_, _012166_, _012173_);
  xor g_104958_(_012160_, _012166_, _012174_);
  and g_104959_(_012171_, _012173_, _012175_);
  or g_104960_(_012172_, _012174_, _012177_);
  or g_104961_(_023374_, _055741_, _012178_);
  not g_104962_(_012178_, _012179_);
  and g_104963_(_009600_, _012178_, _012180_);
  or g_104964_(_009599_, _012179_, _012181_);
  and g_104965_(_011997_, _012096_, _012182_);
  or g_104966_(_011996_, _012095_, _012183_);
  and g_104967_(_011991_, _012095_, _012184_);
  or g_104968_(_011990_, _012096_, _012185_);
  and g_104969_(_012183_, _012185_, _012186_);
  or g_104970_(_012182_, _012184_, _012188_);
  and g_104971_(_012181_, _012186_, _012189_);
  or g_104972_(_012180_, _012188_, _012190_);
  xor g_104973_(out[677], _009599_, _012191_);
  xor g_104974_(_055964_, _009599_, _012192_);
  and g_104975_(_012002_, _012095_, _012193_);
  or g_104976_(_012001_, _012096_, _012194_);
  and g_104977_(_012008_, _012096_, _012195_);
  or g_104978_(_012007_, _012095_, _012196_);
  and g_104979_(_012194_, _012196_, _012197_);
  or g_104980_(_012193_, _012195_, _012199_);
  and g_104981_(_012192_, _012197_, _012200_);
  or g_104982_(_012191_, _012199_, _012201_);
  and g_104983_(_012190_, _012201_, _012202_);
  or g_104984_(_012189_, _012200_, _012203_);
  and g_104985_(_012191_, _012199_, _012204_);
  and g_104986_(_012180_, _012188_, _012205_);
  or g_104987_(_012204_, _012205_, _012206_);
  not g_104988_(_012206_, _012207_);
  and g_104989_(_012202_, _012207_, _012208_);
  or g_104990_(_012203_, _012206_, _012210_);
  and g_104991_(_012175_, _012208_, _012211_);
  or g_104992_(_012177_, _012210_, _012212_);
  and g_104993_(_012149_, _012211_, _012213_);
  or g_104994_(_012150_, _012212_, _012214_);
  xor g_104995_(out[675], _055741_, _012215_);
  xor g_104996_(_000054_, _055741_, _012216_);
  or g_104997_(_012051_, _012095_, _012217_);
  not g_104998_(_012217_, _012218_);
  and g_104999_(_012047_, _012095_, _012219_);
  not g_105000_(_012219_, _012221_);
  and g_105001_(_012217_, _012221_, _012222_);
  or g_105002_(_012218_, _012219_, _012223_);
  and g_105003_(_012215_, _012222_, _012224_);
  or g_105004_(_012216_, _012223_, _012225_);
  or g_105005_(_012043_, _012095_, _012226_);
  not g_105006_(_012226_, _012227_);
  and g_105007_(_055438_, _012095_, _012228_);
  or g_105008_(_012227_, _012228_, _012229_);
  and g_105009_(_055742_, _012229_, _012230_);
  or g_105010_(_012224_, _012230_, _012232_);
  or g_105011_(_055742_, _012229_, _012233_);
  not g_105012_(_012233_, _012234_);
  and g_105013_(_012216_, _012223_, _012235_);
  or g_105014_(_012215_, _012222_, _012236_);
  or g_105015_(_012234_, _012235_, _012237_);
  xor g_105016_(_055742_, _012229_, _012238_);
  and g_105017_(_012225_, _012236_, _012239_);
  and g_105018_(_012238_, _012239_, _012240_);
  or g_105019_(_012232_, _012237_, _012241_);
  and g_105020_(out[657], _012095_, _012243_);
  not g_105021_(_012243_, _012244_);
  or g_105022_(_012029_, _012095_, _012245_);
  not g_105023_(_012245_, _012246_);
  and g_105024_(_012244_, _012245_, _012247_);
  or g_105025_(_012243_, _012246_, _012248_);
  and g_105026_(out[673], _012247_, _012249_);
  or g_105027_(_000021_, _012248_, _012250_);
  and g_105028_(out[656], _012095_, _012251_);
  not g_105029_(_012251_, _012252_);
  or g_105030_(_012032_, _012095_, _012254_);
  not g_105031_(_012254_, _012255_);
  and g_105032_(_012252_, _012254_, _012256_);
  or g_105033_(_012251_, _012255_, _012257_);
  and g_105034_(out[672], _012256_, _012258_);
  or g_105035_(_000032_, _012257_, _012259_);
  xor g_105036_(out[673], _012247_, _012260_);
  xor g_105037_(_000021_, _012247_, _012261_);
  and g_105038_(_012259_, _012260_, _012262_);
  or g_105039_(_012258_, _012261_, _012263_);
  and g_105040_(_012250_, _012263_, _012265_);
  or g_105041_(_012249_, _012262_, _012266_);
  and g_105042_(_012240_, _012266_, _012267_);
  or g_105043_(_012241_, _012265_, _012268_);
  and g_105044_(_012225_, _012233_, _012269_);
  or g_105045_(_012224_, _012234_, _012270_);
  and g_105046_(_012236_, _012270_, _012271_);
  or g_105047_(_012235_, _012269_, _012272_);
  and g_105048_(_012268_, _012272_, _012273_);
  or g_105049_(_012267_, _012271_, _012274_);
  and g_105050_(_012213_, _012274_, _012276_);
  or g_105051_(_012214_, _012273_, _012277_);
  or g_105052_(_012202_, _012204_, _012278_);
  not g_105053_(_012278_, _012279_);
  and g_105054_(_012175_, _012279_, _012280_);
  or g_105055_(_012177_, _012278_, _012281_);
  or g_105056_(_012169_, _012170_, _012282_);
  not g_105057_(_012282_, _012283_);
  and g_105058_(_012281_, _012282_, _012284_);
  or g_105059_(_012280_, _012283_, _012285_);
  and g_105060_(_012149_, _012285_, _012287_);
  or g_105061_(_012150_, _012284_, _012288_);
  and g_105062_(_012139_, _012141_, _012289_);
  and g_105063_(_012115_, _012289_, _012290_);
  not g_105064_(_012290_, _012291_);
  and g_105065_(_012106_, _012109_, _012292_);
  not g_105066_(_012292_, _012293_);
  and g_105067_(_012107_, _012293_, _012294_);
  or g_105068_(_012108_, _012292_, _012295_);
  and g_105069_(_012291_, _012294_, _012296_);
  or g_105070_(_012290_, _012295_, _012298_);
  and g_105071_(_012288_, _012296_, _012299_);
  or g_105072_(_012287_, _012298_, _012300_);
  and g_105073_(_012277_, _012299_, _012301_);
  or g_105074_(_012276_, _012300_, _012302_);
  or g_105075_(out[672], _012256_, _012303_);
  and g_105076_(_012240_, _012303_, _012304_);
  and g_105077_(_012262_, _012304_, _012305_);
  and g_105078_(_012213_, _012305_, _012306_);
  not g_105079_(_012306_, _012307_);
  and g_105080_(_012302_, _012307_, _012309_);
  or g_105081_(_012301_, _012306_, _012310_);
  and g_105082_(_012103_, _012310_, _012311_);
  or g_105083_(_012102_, _012309_, _012312_);
  and g_105084_(_012104_, _012309_, _012313_);
  or g_105085_(_012105_, _012310_, _012314_);
  and g_105086_(_012312_, _012314_, _012315_);
  or g_105087_(_012311_, _012313_, _012316_);
  xor g_105088_(out[698], _009621_, _012317_);
  xor g_105089_(_000219_, _009621_, _012318_);
  and g_105090_(_012315_, _012317_, _012320_);
  or g_105091_(_012316_, _012318_, _012321_);
  and g_105092_(_009610_, _009626_, _012322_);
  or g_105093_(_009611_, _009625_, _012323_);
  and g_105094_(_012321_, _012323_, _012324_);
  or g_105095_(_012320_, _012322_, _012325_);
  and g_105096_(_009611_, _009625_, _012326_);
  or g_105097_(_009610_, _009626_, _012327_);
  and g_105098_(_012316_, _012318_, _012328_);
  or g_105099_(_012315_, _012317_, _012329_);
  and g_105100_(_012327_, _012329_, _012331_);
  or g_105101_(_012326_, _012328_, _012332_);
  and g_105102_(out[697], _009620_, _012333_);
  xor g_105103_(out[697], _009620_, _012334_);
  or g_105104_(_009622_, _012333_, _012335_);
  and g_105105_(_012136_, _012310_, _012336_);
  and g_105106_(_012129_, _012309_, _012337_);
  or g_105107_(_012336_, _012337_, _012338_);
  or g_105108_(_012334_, _012338_, _012339_);
  not g_105109_(_012339_, _012340_);
  xor g_105110_(out[696], _009619_, _012342_);
  xor g_105111_(_000197_, _009619_, _012343_);
  and g_105112_(_012118_, _012309_, _012344_);
  and g_105113_(_012125_, _012310_, _012345_);
  or g_105114_(_012344_, _012345_, _012346_);
  and g_105115_(_012334_, _012338_, _012347_);
  not g_105116_(_012347_, _012348_);
  or g_105117_(_012342_, _012346_, _012349_);
  and g_105118_(_012348_, _012349_, _012350_);
  xor g_105119_(_012342_, _012346_, _012351_);
  xor g_105120_(_012343_, _012346_, _012353_);
  and g_105121_(_012324_, _012331_, _012354_);
  or g_105122_(_012325_, _012332_, _012355_);
  and g_105123_(_012339_, _012348_, _012356_);
  or g_105124_(_012340_, _012347_, _012357_);
  and g_105125_(_012354_, _012356_, _012358_);
  or g_105126_(_012355_, _012357_, _012359_);
  and g_105127_(_012351_, _012358_, _012360_);
  or g_105128_(_012353_, _012359_, _012361_);
  xor g_105129_(out[695], _009618_, _012362_);
  xor g_105130_(_000109_, _009618_, _012364_);
  and g_105131_(_012159_, _012309_, _012365_);
  or g_105132_(_012160_, _012310_, _012366_);
  and g_105133_(_012167_, _012310_, _012367_);
  or g_105134_(_012166_, _012309_, _012368_);
  and g_105135_(_012366_, _012368_, _012369_);
  or g_105136_(_012365_, _012367_, _012370_);
  and g_105137_(_012362_, _012369_, _012371_);
  or g_105138_(_012364_, _012370_, _012372_);
  xor g_105139_(out[694], _009617_, _012373_);
  not g_105140_(_012373_, _012375_);
  and g_105141_(_012152_, _012309_, _012376_);
  and g_105142_(_012157_, _012310_, _012377_);
  or g_105143_(_012376_, _012377_, _012378_);
  or g_105144_(_012373_, _012378_, _012379_);
  not g_105145_(_012379_, _012380_);
  and g_105146_(_012364_, _012370_, _012381_);
  or g_105147_(_012362_, _012369_, _012382_);
  and g_105148_(_012372_, _012382_, _012383_);
  or g_105149_(_012371_, _012381_, _012384_);
  xor g_105150_(_012373_, _012378_, _012386_);
  xor g_105151_(_012375_, _012378_, _012387_);
  and g_105152_(_012383_, _012386_, _012388_);
  or g_105153_(_012384_, _012387_, _012389_);
  or g_105154_(_023528_, _055929_, _012390_);
  not g_105155_(_012390_, _012391_);
  and g_105156_(_009616_, _012390_, _012392_);
  or g_105157_(_009615_, _012391_, _012393_);
  and g_105158_(_012188_, _012310_, _012394_);
  not g_105159_(_012394_, _012395_);
  or g_105160_(_012180_, _012310_, _012397_);
  not g_105161_(_012397_, _012398_);
  and g_105162_(_012395_, _012397_, _012399_);
  or g_105163_(_012394_, _012398_, _012400_);
  and g_105164_(_012393_, _012399_, _012401_);
  or g_105165_(_012392_, _012400_, _012402_);
  xor g_105166_(out[693], _009615_, _012403_);
  xor g_105167_(_000131_, _009615_, _012404_);
  or g_105168_(_012191_, _012310_, _012405_);
  not g_105169_(_012405_, _012406_);
  and g_105170_(_012199_, _012310_, _012408_);
  not g_105171_(_012408_, _012409_);
  and g_105172_(_012405_, _012409_, _012410_);
  or g_105173_(_012406_, _012408_, _012411_);
  and g_105174_(_012404_, _012410_, _012412_);
  or g_105175_(_012403_, _012411_, _012413_);
  and g_105176_(_012402_, _012413_, _012414_);
  or g_105177_(_012401_, _012412_, _012415_);
  and g_105178_(_012403_, _012411_, _012416_);
  or g_105179_(_012404_, _012410_, _012417_);
  and g_105180_(_012392_, _012400_, _012419_);
  or g_105181_(_012416_, _012419_, _012420_);
  or g_105182_(_012415_, _012420_, _012421_);
  or g_105183_(_012389_, _012421_, _012422_);
  or g_105184_(_012361_, _012422_, _012423_);
  xor g_105185_(out[691], _055929_, _012424_);
  xor g_105186_(_000186_, _055929_, _012425_);
  and g_105187_(_012215_, _012309_, _012426_);
  and g_105188_(_012223_, _012310_, _012427_);
  or g_105189_(_012426_, _012427_, _012428_);
  or g_105190_(_012425_, _012428_, _012430_);
  and g_105191_(_012229_, _012310_, _012431_);
  and g_105192_(_055743_, _012309_, _012432_);
  or g_105193_(_012431_, _012432_, _012433_);
  and g_105194_(_012425_, _012428_, _012434_);
  or g_105195_(_055932_, _012433_, _012435_);
  xor g_105196_(_012424_, _012428_, _012436_);
  xor g_105197_(_055930_, _012433_, _012437_);
  or g_105198_(_012436_, _012437_, _012438_);
  or g_105199_(_000021_, _012310_, _012439_);
  or g_105200_(_012247_, _012309_, _012441_);
  and g_105201_(_012439_, _012441_, _012442_);
  and g_105202_(out[689], _012442_, _012443_);
  not g_105203_(_012443_, _012444_);
  and g_105204_(_012256_, _012310_, _012445_);
  or g_105205_(_012257_, _012309_, _012446_);
  or g_105206_(out[672], _012310_, _012447_);
  not g_105207_(_012447_, _012448_);
  or g_105208_(_012445_, _012448_, _012449_);
  and g_105209_(_012446_, _012447_, _012450_);
  and g_105210_(out[688], _012449_, _012452_);
  xor g_105211_(_000153_, _012442_, _012453_);
  or g_105212_(_012452_, _012453_, _012454_);
  and g_105213_(_012444_, _012454_, _012455_);
  or g_105214_(_012438_, _012455_, _012456_);
  or g_105215_(_012434_, _012435_, _012457_);
  and g_105216_(_012430_, _012457_, _012458_);
  and g_105217_(_012456_, _012458_, _012459_);
  or g_105218_(_012423_, _012459_, _012460_);
  and g_105219_(_012388_, _012415_, _012461_);
  or g_105220_(_012389_, _012414_, _012463_);
  and g_105221_(_012417_, _012461_, _012464_);
  or g_105222_(_012416_, _012463_, _012465_);
  and g_105223_(_012380_, _012382_, _012466_);
  or g_105224_(_012379_, _012381_, _012467_);
  and g_105225_(_012372_, _012467_, _012468_);
  or g_105226_(_012371_, _012466_, _012469_);
  and g_105227_(_012465_, _012468_, _012470_);
  or g_105228_(_012464_, _012469_, _012471_);
  and g_105229_(_012360_, _012471_, _012472_);
  or g_105230_(_012361_, _012470_, _012474_);
  or g_105231_(_012324_, _012326_, _012475_);
  or g_105232_(_012350_, _012355_, _012476_);
  not g_105233_(_012476_, _012477_);
  and g_105234_(_012339_, _012477_, _012478_);
  or g_105235_(_012340_, _012476_, _012479_);
  and g_105236_(_012474_, _012479_, _012480_);
  or g_105237_(_012472_, _012478_, _012481_);
  and g_105238_(_012460_, _012475_, _012482_);
  not g_105239_(_012482_, _012483_);
  and g_105240_(_012480_, _012482_, _012485_);
  or g_105241_(_012481_, _012483_, _012486_);
  and g_105242_(_000164_, _012450_, _012487_);
  or g_105243_(out[688], _012449_, _012488_);
  or g_105244_(_012438_, _012454_, _012489_);
  or g_105245_(_012423_, _012489_, _012490_);
  not g_105246_(_012490_, _012491_);
  and g_105247_(_012488_, _012491_, _012492_);
  or g_105248_(_012487_, _012490_, _012493_);
  and g_105249_(_012486_, _012493_, _012494_);
  or g_105250_(_012485_, _012492_, _012496_);
  and g_105251_(_012316_, _012496_, _012497_);
  not g_105252_(_012497_, _012498_);
  or g_105253_(_012318_, _012496_, _012499_);
  not g_105254_(_012499_, _012500_);
  and g_105255_(_012498_, _012499_, _012501_);
  or g_105256_(_012497_, _012500_, _012502_);
  xor g_105257_(out[714], _009638_, _012503_);
  not g_105258_(_012503_, _012504_);
  and g_105259_(_012501_, _012503_, _012505_);
  or g_105260_(_012502_, _012504_, _012507_);
  and g_105261_(_009627_, _009641_, _012508_);
  or g_105262_(_009628_, _009640_, _012509_);
  and g_105263_(_012507_, _012509_, _012510_);
  or g_105264_(_012505_, _012508_, _012511_);
  and g_105265_(_009628_, _009640_, _012512_);
  or g_105266_(_009627_, _009641_, _012513_);
  and g_105267_(_012502_, _012504_, _012514_);
  or g_105268_(_012501_, _012503_, _012515_);
  and g_105269_(_012513_, _012515_, _012516_);
  or g_105270_(_012512_, _012514_, _012518_);
  and g_105271_(_012510_, _012516_, _012519_);
  or g_105272_(_012511_, _012518_, _012520_);
  xor g_105273_(out[712], _009636_, _012521_);
  xor g_105274_(_000329_, _009636_, _012522_);
  or g_105275_(_012342_, _012496_, _012523_);
  not g_105276_(_012523_, _012524_);
  and g_105277_(_012346_, _012496_, _012525_);
  not g_105278_(_012525_, _012526_);
  and g_105279_(_012523_, _012526_, _012527_);
  or g_105280_(_012524_, _012525_, _012529_);
  and g_105281_(_012521_, _012529_, _012530_);
  or g_105282_(_012522_, _012527_, _012531_);
  and g_105283_(out[713], _009637_, _012532_);
  xor g_105284_(out[713], _009637_, _012533_);
  xor g_105285_(_000340_, _009637_, _012534_);
  and g_105286_(_012338_, _012496_, _012535_);
  not g_105287_(_012535_, _012536_);
  or g_105288_(_012334_, _012496_, _012537_);
  not g_105289_(_012537_, _012538_);
  and g_105290_(_012536_, _012537_, _012540_);
  or g_105291_(_012535_, _012538_, _012541_);
  and g_105292_(_012534_, _012540_, _012542_);
  or g_105293_(_012533_, _012541_, _012543_);
  and g_105294_(_012531_, _012543_, _012544_);
  or g_105295_(_012530_, _012542_, _012545_);
  and g_105296_(_012522_, _012527_, _012546_);
  or g_105297_(_012521_, _012529_, _012547_);
  and g_105298_(_012533_, _012541_, _012548_);
  or g_105299_(_012534_, _012540_, _012549_);
  and g_105300_(_012547_, _012549_, _012551_);
  or g_105301_(_012546_, _012548_, _012552_);
  and g_105302_(_012544_, _012551_, _012553_);
  or g_105303_(_012545_, _012552_, _012554_);
  and g_105304_(_012519_, _012553_, _012555_);
  or g_105305_(_012520_, _012554_, _012556_);
  xor g_105306_(out[711], _009634_, _012557_);
  xor g_105307_(_000241_, _009634_, _012558_);
  and g_105308_(_012362_, _012494_, _012559_);
  or g_105309_(_012364_, _012496_, _012560_);
  and g_105310_(_012370_, _012496_, _012562_);
  or g_105311_(_012369_, _012494_, _012563_);
  and g_105312_(_012560_, _012563_, _012564_);
  or g_105313_(_012559_, _012562_, _012565_);
  and g_105314_(_012557_, _012564_, _012566_);
  or g_105315_(_012558_, _012565_, _012567_);
  and g_105316_(_012558_, _012565_, _012568_);
  or g_105317_(_012557_, _012564_, _012569_);
  and g_105318_(_012567_, _012569_, _012570_);
  or g_105319_(_012566_, _012568_, _012571_);
  xor g_105320_(out[710], _009633_, _012573_);
  not g_105321_(_012573_, _012574_);
  and g_105322_(_012375_, _012494_, _012575_);
  and g_105323_(_012378_, _012496_, _012576_);
  or g_105324_(_012575_, _012576_, _012577_);
  or g_105325_(_012573_, _012577_, _012578_);
  not g_105326_(_012578_, _012579_);
  xor g_105327_(_012573_, _012577_, _012580_);
  xor g_105328_(_012574_, _012577_, _012581_);
  and g_105329_(_012570_, _012580_, _012582_);
  or g_105330_(_012571_, _012581_, _012584_);
  or g_105331_(_023682_, _000140_, _012585_);
  not g_105332_(_012585_, _012586_);
  and g_105333_(_009632_, _012585_, _012587_);
  or g_105334_(_009631_, _012586_, _012588_);
  and g_105335_(_012400_, _012496_, _012589_);
  not g_105336_(_012589_, _012590_);
  or g_105337_(_012392_, _012496_, _012591_);
  not g_105338_(_012591_, _012592_);
  and g_105339_(_012590_, _012591_, _012593_);
  or g_105340_(_012589_, _012592_, _012595_);
  and g_105341_(_012588_, _012593_, _012596_);
  or g_105342_(_012587_, _012595_, _012597_);
  xor g_105343_(out[709], _009631_, _012598_);
  xor g_105344_(_000263_, _009631_, _012599_);
  or g_105345_(_012403_, _012496_, _012600_);
  not g_105346_(_012600_, _012601_);
  and g_105347_(_012411_, _012496_, _012602_);
  not g_105348_(_012602_, _012603_);
  and g_105349_(_012600_, _012603_, _012604_);
  or g_105350_(_012601_, _012602_, _012606_);
  and g_105351_(_012599_, _012604_, _012607_);
  or g_105352_(_012598_, _012606_, _012608_);
  and g_105353_(_012597_, _012608_, _012609_);
  or g_105354_(_012596_, _012607_, _012610_);
  and g_105355_(_012598_, _012606_, _012611_);
  not g_105356_(_012611_, _012612_);
  or g_105357_(_012588_, _012593_, _012613_);
  and g_105358_(_012612_, _012613_, _012614_);
  and g_105359_(_012609_, _012614_, _012615_);
  and g_105360_(_012582_, _012615_, _012617_);
  not g_105361_(_012617_, _012618_);
  and g_105362_(_012555_, _012617_, _012619_);
  or g_105363_(_012556_, _012618_, _012620_);
  xor g_105364_(out[707], _000140_, _012621_);
  xor g_105365_(_000318_, _000140_, _012622_);
  and g_105366_(_012424_, _012494_, _012623_);
  and g_105367_(_012428_, _012496_, _012624_);
  or g_105368_(_012623_, _012624_, _012625_);
  not g_105369_(_012625_, _012626_);
  or g_105370_(_012622_, _012625_, _012628_);
  and g_105371_(_012622_, _012625_, _012629_);
  or g_105372_(_012621_, _012626_, _012630_);
  and g_105373_(_012433_, _012496_, _012631_);
  and g_105374_(_055930_, _012494_, _012632_);
  or g_105375_(_012631_, _012632_, _012633_);
  or g_105376_(_000143_, _012633_, _012634_);
  or g_105377_(_012629_, _012634_, _012635_);
  and g_105378_(_012628_, _012635_, _012636_);
  not g_105379_(_012636_, _012637_);
  or g_105380_(_000153_, _012496_, _012639_);
  or g_105381_(_012442_, _012494_, _012640_);
  and g_105382_(_012639_, _012640_, _012641_);
  and g_105383_(out[705], _012641_, _012642_);
  or g_105384_(_000164_, _012496_, _012643_);
  or g_105385_(_012449_, _012494_, _012644_);
  and g_105386_(_012643_, _012644_, _012645_);
  and g_105387_(out[704], _012645_, _012646_);
  not g_105388_(_012646_, _012647_);
  xor g_105389_(out[705], _012641_, _012648_);
  xor g_105390_(_000285_, _012641_, _012650_);
  and g_105391_(_012647_, _012648_, _012651_);
  or g_105392_(_012646_, _012650_, _012652_);
  or g_105393_(_012642_, _012651_, _012653_);
  xor g_105394_(_000143_, _012633_, _012654_);
  and g_105395_(_012630_, _012654_, _012655_);
  and g_105396_(_012653_, _012655_, _012656_);
  not g_105397_(_012656_, _012657_);
  and g_105398_(_012636_, _012657_, _012658_);
  or g_105399_(_012637_, _012656_, _012659_);
  and g_105400_(_012619_, _012659_, _012661_);
  or g_105401_(_012620_, _012658_, _012662_);
  and g_105402_(_012610_, _012612_, _012663_);
  or g_105403_(_012609_, _012611_, _012664_);
  and g_105404_(_012582_, _012663_, _012665_);
  or g_105405_(_012584_, _012664_, _012666_);
  and g_105406_(_012569_, _012579_, _012667_);
  or g_105407_(_012568_, _012578_, _012668_);
  and g_105408_(_012567_, _012668_, _012669_);
  or g_105409_(_012566_, _012667_, _012670_);
  and g_105410_(_012666_, _012669_, _012672_);
  or g_105411_(_012665_, _012670_, _012673_);
  and g_105412_(_012555_, _012673_, _012674_);
  or g_105413_(_012556_, _012672_, _012675_);
  and g_105414_(_012511_, _012513_, _012676_);
  or g_105415_(_012510_, _012512_, _012677_);
  and g_105416_(_012519_, _012552_, _012678_);
  or g_105417_(_012520_, _012551_, _012679_);
  and g_105418_(_012543_, _012678_, _012680_);
  or g_105419_(_012542_, _012679_, _012681_);
  and g_105420_(_012677_, _012681_, _012683_);
  or g_105421_(_012676_, _012680_, _012684_);
  and g_105422_(_012675_, _012683_, _012685_);
  or g_105423_(_012674_, _012684_, _012686_);
  and g_105424_(_012662_, _012685_, _012687_);
  or g_105425_(_012661_, _012686_, _012688_);
  or g_105426_(out[704], _012645_, _012689_);
  and g_105427_(_012628_, _012689_, _012690_);
  and g_105428_(_012655_, _012690_, _012691_);
  and g_105429_(_012619_, _012691_, _012692_);
  not g_105430_(_012692_, _012694_);
  and g_105431_(_012651_, _012692_, _012695_);
  or g_105432_(_012652_, _012694_, _012696_);
  and g_105433_(_012688_, _012696_, _012697_);
  or g_105434_(_012687_, _012695_, _012698_);
  and g_105435_(_012502_, _012698_, _012699_);
  or g_105436_(_012501_, _012697_, _012700_);
  and g_105437_(_012503_, _012697_, _012701_);
  or g_105438_(_012504_, _012698_, _012702_);
  and g_105439_(_012700_, _012702_, _012703_);
  or g_105440_(_012699_, _012701_, _012705_);
  xor g_105441_(out[730], _009653_, _012706_);
  xor g_105442_(_000483_, _009653_, _012707_);
  and g_105443_(_012703_, _012706_, _012708_);
  or g_105444_(_012705_, _012707_, _012709_);
  and g_105445_(_009642_, _009658_, _012710_);
  or g_105446_(_009643_, _009656_, _012711_);
  and g_105447_(_012709_, _012711_, _012712_);
  or g_105448_(_012708_, _012710_, _012713_);
  and g_105449_(_009643_, _009656_, _012714_);
  or g_105450_(_009642_, _009658_, _012716_);
  xor g_105451_(out[728], _009651_, _012717_);
  xor g_105452_(_000461_, _009651_, _012718_);
  or g_105453_(_012521_, _012698_, _012719_);
  not g_105454_(_012719_, _012720_);
  and g_105455_(_012529_, _012698_, _012721_);
  not g_105456_(_012721_, _012722_);
  and g_105457_(_012719_, _012722_, _012723_);
  or g_105458_(_012720_, _012721_, _012724_);
  and g_105459_(_012717_, _012724_, _012725_);
  or g_105460_(_012718_, _012723_, _012727_);
  and g_105461_(_012716_, _012727_, _012728_);
  or g_105462_(_012714_, _012725_, _012729_);
  and g_105463_(_012712_, _012728_, _012730_);
  or g_105464_(_012713_, _012729_, _012731_);
  and g_105465_(out[729], _009652_, _012732_);
  xor g_105466_(out[729], _009652_, _012733_);
  or g_105467_(_009654_, _012732_, _012734_);
  and g_105468_(_012541_, _012698_, _012735_);
  not g_105469_(_012735_, _012736_);
  or g_105470_(_012533_, _012698_, _012738_);
  not g_105471_(_012738_, _012739_);
  and g_105472_(_012736_, _012738_, _012740_);
  or g_105473_(_012735_, _012739_, _012741_);
  and g_105474_(_012733_, _012741_, _012742_);
  or g_105475_(_012734_, _012740_, _012743_);
  and g_105476_(_012718_, _012723_, _012744_);
  or g_105477_(_012717_, _012724_, _012745_);
  and g_105478_(_012743_, _012745_, _012746_);
  or g_105479_(_012742_, _012744_, _012747_);
  and g_105480_(_012705_, _012707_, _012749_);
  or g_105481_(_012703_, _012706_, _012750_);
  and g_105482_(_012734_, _012740_, _012751_);
  or g_105483_(_012733_, _012741_, _012752_);
  and g_105484_(_012750_, _012752_, _012753_);
  or g_105485_(_012749_, _012751_, _012754_);
  and g_105486_(_012746_, _012753_, _012755_);
  or g_105487_(_012747_, _012754_, _012756_);
  and g_105488_(_012730_, _012755_, _012757_);
  or g_105489_(_012731_, _012756_, _012758_);
  xor g_105490_(out[727], _009650_, _012760_);
  xor g_105491_(_000373_, _009650_, _012761_);
  and g_105492_(_012557_, _012697_, _012762_);
  and g_105493_(_012565_, _012698_, _012763_);
  or g_105494_(_012762_, _012763_, _012764_);
  or g_105495_(_012761_, _012764_, _012765_);
  xor g_105496_(out[726], _009649_, _012766_);
  xor g_105497_(_000384_, _009649_, _012767_);
  and g_105498_(_012574_, _012697_, _012768_);
  and g_105499_(_012577_, _012698_, _012769_);
  or g_105500_(_012768_, _012769_, _012771_);
  or g_105501_(_012766_, _012771_, _012772_);
  and g_105502_(_012761_, _012764_, _012773_);
  xor g_105503_(_012761_, _012764_, _012774_);
  xor g_105504_(_012760_, _012764_, _012775_);
  xor g_105505_(_012766_, _012771_, _012776_);
  xor g_105506_(_012767_, _012771_, _012777_);
  and g_105507_(_012774_, _012776_, _012778_);
  or g_105508_(_012775_, _012777_, _012779_);
  or g_105509_(_023836_, _000239_, _012780_);
  not g_105510_(_012780_, _012782_);
  and g_105511_(_009648_, _012780_, _012783_);
  or g_105512_(_009647_, _012782_, _012784_);
  and g_105513_(_012595_, _012698_, _012785_);
  not g_105514_(_012785_, _012786_);
  or g_105515_(_012587_, _012698_, _012787_);
  not g_105516_(_012787_, _012788_);
  and g_105517_(_012786_, _012787_, _012789_);
  or g_105518_(_012785_, _012788_, _012790_);
  and g_105519_(_012784_, _012789_, _012791_);
  or g_105520_(_012783_, _012790_, _012793_);
  xor g_105521_(out[725], _009647_, _012794_);
  xor g_105522_(_000395_, _009647_, _012795_);
  or g_105523_(_012598_, _012698_, _012796_);
  not g_105524_(_012796_, _012797_);
  and g_105525_(_012606_, _012698_, _012798_);
  not g_105526_(_012798_, _012799_);
  and g_105527_(_012796_, _012799_, _012800_);
  or g_105528_(_012797_, _012798_, _012801_);
  and g_105529_(_012795_, _012800_, _012802_);
  or g_105530_(_012794_, _012801_, _012804_);
  and g_105531_(_012793_, _012804_, _012805_);
  or g_105532_(_012791_, _012802_, _012806_);
  and g_105533_(_012794_, _012801_, _012807_);
  or g_105534_(_012795_, _012800_, _012808_);
  and g_105535_(_012783_, _012790_, _012809_);
  or g_105536_(_012784_, _012789_, _012810_);
  and g_105537_(_012808_, _012810_, _012811_);
  or g_105538_(_012807_, _012809_, _012812_);
  and g_105539_(_012805_, _012811_, _012813_);
  or g_105540_(_012806_, _012812_, _012815_);
  and g_105541_(_012778_, _012813_, _012816_);
  or g_105542_(_012779_, _012815_, _012817_);
  and g_105543_(_012757_, _012816_, _012818_);
  or g_105544_(_012758_, _012817_, _012819_);
  xor g_105545_(out[723], _000239_, _012820_);
  xor g_105546_(_000450_, _000239_, _012821_);
  and g_105547_(_012621_, _012697_, _012822_);
  and g_105548_(_012625_, _012698_, _012823_);
  or g_105549_(_012822_, _012823_, _012824_);
  or g_105550_(_012821_, _012824_, _012826_);
  and g_105551_(_012633_, _012698_, _012827_);
  and g_105552_(_000141_, _012697_, _012828_);
  or g_105553_(_012827_, _012828_, _012829_);
  or g_105554_(_000242_, _012829_, _012830_);
  and g_105555_(_012821_, _012824_, _012831_);
  xor g_105556_(_000242_, _012829_, _012832_);
  xor g_105557_(_000240_, _012829_, _012833_);
  xor g_105558_(_012821_, _012824_, _012834_);
  xor g_105559_(_012820_, _012824_, _012835_);
  and g_105560_(_012832_, _012834_, _012837_);
  or g_105561_(_012833_, _012835_, _012838_);
  or g_105562_(_000285_, _012698_, _012839_);
  or g_105563_(_012641_, _012697_, _012840_);
  and g_105564_(_012839_, _012840_, _012841_);
  and g_105565_(out[721], _012841_, _012842_);
  not g_105566_(_012842_, _012843_);
  and g_105567_(_012645_, _012698_, _012844_);
  not g_105568_(_012844_, _012845_);
  or g_105569_(out[704], _012698_, _012846_);
  not g_105570_(_012846_, _012848_);
  or g_105571_(_012844_, _012848_, _012849_);
  and g_105572_(_012845_, _012846_, _012850_);
  and g_105573_(out[720], _012849_, _012851_);
  or g_105574_(_000428_, _012850_, _012852_);
  xor g_105575_(out[721], _012841_, _012853_);
  xor g_105576_(_000417_, _012841_, _012854_);
  and g_105577_(_012852_, _012853_, _012855_);
  or g_105578_(_012851_, _012854_, _012856_);
  and g_105579_(_012843_, _012856_, _012857_);
  or g_105580_(_012842_, _012855_, _012859_);
  and g_105581_(_012837_, _012859_, _012860_);
  or g_105582_(_012838_, _012857_, _012861_);
  and g_105583_(_012826_, _012830_, _012862_);
  or g_105584_(_012831_, _012862_, _012863_);
  not g_105585_(_012863_, _012864_);
  and g_105586_(_012861_, _012863_, _012865_);
  or g_105587_(_012860_, _012864_, _012866_);
  and g_105588_(_012818_, _012866_, _012867_);
  or g_105589_(_012819_, _012865_, _012868_);
  and g_105590_(_012778_, _012806_, _012870_);
  or g_105591_(_012779_, _012805_, _012871_);
  and g_105592_(_012808_, _012870_, _012872_);
  or g_105593_(_012807_, _012871_, _012873_);
  or g_105594_(_012772_, _012773_, _012874_);
  and g_105595_(_012765_, _012874_, _012875_);
  not g_105596_(_012875_, _012876_);
  and g_105597_(_012873_, _012875_, _012877_);
  or g_105598_(_012872_, _012876_, _012878_);
  and g_105599_(_012757_, _012878_, _012879_);
  or g_105600_(_012758_, _012877_, _012881_);
  and g_105601_(_012747_, _012753_, _012882_);
  or g_105602_(_012746_, _012754_, _012883_);
  and g_105603_(_012712_, _012883_, _012884_);
  or g_105604_(_012713_, _012882_, _012885_);
  and g_105605_(_012716_, _012885_, _012886_);
  or g_105606_(_012714_, _012884_, _012887_);
  and g_105607_(_012881_, _012887_, _012888_);
  or g_105608_(_012879_, _012886_, _012889_);
  and g_105609_(_012868_, _012888_, _012890_);
  or g_105610_(_012867_, _012889_, _012892_);
  or g_105611_(out[720], _012849_, _012893_);
  not g_105612_(_012893_, _012894_);
  or g_105613_(_012838_, _012894_, _012895_);
  or g_105614_(_012856_, _012895_, _012896_);
  or g_105615_(_012819_, _012896_, _012897_);
  not g_105616_(_012897_, _012898_);
  and g_105617_(_012892_, _012897_, _012899_);
  or g_105618_(_012890_, _012898_, _012900_);
  and g_105619_(_012705_, _012900_, _012901_);
  or g_105620_(_012703_, _012899_, _012903_);
  and g_105621_(_012706_, _012899_, _012904_);
  or g_105622_(_012707_, _012900_, _012905_);
  and g_105623_(_012903_, _012905_, _012906_);
  or g_105624_(_012901_, _012904_, _012907_);
  or g_105625_(_009660_, _009672_, _012908_);
  and g_105626_(_009660_, _009672_, _012909_);
  xor g_105627_(_009659_, _009672_, _012910_);
  xor g_105628_(out[746], _009670_, _012911_);
  not g_105629_(_012911_, _012912_);
  and g_105630_(_012906_, _012911_, _012914_);
  or g_105631_(_012907_, _012912_, _012915_);
  or g_105632_(_012910_, _012914_, _012916_);
  and g_105633_(_012907_, _012912_, _012917_);
  and g_105634_(out[745], _009669_, _012918_);
  xor g_105635_(out[745], _009669_, _012919_);
  xor g_105636_(_000604_, _009669_, _012920_);
  and g_105637_(_012741_, _012900_, _012921_);
  or g_105638_(_012740_, _012899_, _012922_);
  and g_105639_(_012734_, _012899_, _012923_);
  or g_105640_(_012733_, _012900_, _012925_);
  and g_105641_(_012922_, _012925_, _012926_);
  or g_105642_(_012921_, _012923_, _012927_);
  and g_105643_(_012920_, _012926_, _012928_);
  or g_105644_(_012917_, _012928_, _012929_);
  or g_105645_(_012916_, _012929_, _012930_);
  xor g_105646_(out[744], _009667_, _012931_);
  xor g_105647_(_000593_, _009667_, _012932_);
  or g_105648_(_012717_, _012900_, _012933_);
  not g_105649_(_012933_, _012934_);
  and g_105650_(_012724_, _012900_, _012936_);
  or g_105651_(_012723_, _012899_, _012937_);
  and g_105652_(_012933_, _012937_, _012938_);
  or g_105653_(_012934_, _012936_, _012939_);
  and g_105654_(_012931_, _012939_, _012940_);
  and g_105655_(_012919_, _012927_, _012941_);
  or g_105656_(_012920_, _012926_, _012942_);
  and g_105657_(_012932_, _012938_, _012943_);
  or g_105658_(_012931_, _012939_, _012944_);
  and g_105659_(_012942_, _012944_, _012945_);
  or g_105660_(_012941_, _012943_, _012947_);
  or g_105661_(_012940_, _012947_, _012948_);
  or g_105662_(_012930_, _012948_, _012949_);
  xor g_105663_(out[743], _009666_, _012950_);
  xor g_105664_(_000505_, _009666_, _012951_);
  and g_105665_(_012760_, _012899_, _012952_);
  and g_105666_(_012764_, _012900_, _012953_);
  or g_105667_(_012952_, _012953_, _012954_);
  or g_105668_(_012951_, _012954_, _012955_);
  xor g_105669_(out[742], _009665_, _012956_);
  not g_105670_(_012956_, _012958_);
  and g_105671_(_012767_, _012899_, _012959_);
  and g_105672_(_012771_, _012900_, _012960_);
  or g_105673_(_012959_, _012960_, _012961_);
  or g_105674_(_012956_, _012961_, _012962_);
  and g_105675_(_012951_, _012954_, _012963_);
  xor g_105676_(_012950_, _012954_, _012964_);
  xor g_105677_(_012958_, _012961_, _012965_);
  or g_105678_(_012964_, _012965_, _012966_);
  or g_105679_(_023990_, _000361_, _012967_);
  not g_105680_(_012967_, _012969_);
  and g_105681_(_009664_, _012967_, _012970_);
  or g_105682_(_009663_, _012969_, _012971_);
  and g_105683_(_012790_, _012900_, _012972_);
  not g_105684_(_012972_, _012973_);
  or g_105685_(_012783_, _012900_, _012974_);
  not g_105686_(_012974_, _012975_);
  and g_105687_(_012973_, _012974_, _012976_);
  or g_105688_(_012972_, _012975_, _012977_);
  and g_105689_(_012971_, _012976_, _012978_);
  or g_105690_(_012970_, _012977_, _012980_);
  xor g_105691_(out[741], _009663_, _012981_);
  xor g_105692_(_000527_, _009663_, _012982_);
  or g_105693_(_012794_, _012900_, _012983_);
  not g_105694_(_012983_, _012984_);
  and g_105695_(_012801_, _012900_, _012985_);
  not g_105696_(_012985_, _012986_);
  and g_105697_(_012983_, _012986_, _012987_);
  or g_105698_(_012984_, _012985_, _012988_);
  and g_105699_(_012982_, _012987_, _012989_);
  or g_105700_(_012981_, _012988_, _012991_);
  and g_105701_(_012980_, _012991_, _012992_);
  or g_105702_(_012978_, _012989_, _012993_);
  and g_105703_(_012981_, _012988_, _012994_);
  and g_105704_(_012970_, _012977_, _012995_);
  or g_105705_(_012994_, _012995_, _012996_);
  or g_105706_(_012993_, _012996_, _012997_);
  or g_105707_(_012949_, _012997_, _012998_);
  or g_105708_(_012966_, _012998_, _012999_);
  and g_105709_(_012829_, _012900_, _013000_);
  and g_105710_(_000240_, _012899_, _013002_);
  or g_105711_(_013000_, _013002_, _013003_);
  not g_105712_(_013003_, _013004_);
  xor g_105713_(out[739], _000361_, _013005_);
  xor g_105714_(_000582_, _000361_, _013006_);
  and g_105715_(_012820_, _012899_, _013007_);
  and g_105716_(_012824_, _012900_, _013008_);
  or g_105717_(_013007_, _013008_, _013009_);
  or g_105718_(_013006_, _013009_, _013010_);
  or g_105719_(_000363_, _013003_, _013011_);
  and g_105720_(_013006_, _013009_, _013013_);
  xor g_105721_(_000363_, _013003_, _013014_);
  xor g_105722_(_000363_, _013004_, _013015_);
  xor g_105723_(_013006_, _013009_, _013016_);
  xor g_105724_(_013005_, _013009_, _013017_);
  and g_105725_(_013014_, _013016_, _013018_);
  or g_105726_(_013015_, _013017_, _013019_);
  or g_105727_(_000417_, _012900_, _013020_);
  or g_105728_(_012841_, _012899_, _013021_);
  and g_105729_(_013020_, _013021_, _013022_);
  and g_105730_(out[737], _013022_, _013024_);
  not g_105731_(_013024_, _013025_);
  and g_105732_(out[720], _012899_, _013026_);
  or g_105733_(_000428_, _012900_, _013027_);
  and g_105734_(_012850_, _012900_, _013028_);
  or g_105735_(_012849_, _012899_, _013029_);
  and g_105736_(_013027_, _013029_, _013030_);
  or g_105737_(_013026_, _013028_, _013031_);
  and g_105738_(out[736], _013030_, _013032_);
  xor g_105739_(_000549_, _013022_, _013033_);
  or g_105740_(_013032_, _013033_, _013035_);
  and g_105741_(_013025_, _013035_, _013036_);
  or g_105742_(_013019_, _013036_, _013037_);
  or g_105743_(_013011_, _013013_, _013038_);
  and g_105744_(_013010_, _013038_, _013039_);
  and g_105745_(_013037_, _013039_, _013040_);
  or g_105746_(_012999_, _013040_, _013041_);
  or g_105747_(_012966_, _012992_, _013042_);
  or g_105748_(_012994_, _013042_, _013043_);
  or g_105749_(_012962_, _012963_, _013044_);
  and g_105750_(_012955_, _013044_, _013046_);
  and g_105751_(_013043_, _013046_, _013047_);
  or g_105752_(_012949_, _013047_, _013048_);
  or g_105753_(_012930_, _012945_, _013049_);
  and g_105754_(_012908_, _012915_, _013050_);
  or g_105755_(_012909_, _013050_, _013051_);
  and g_105756_(_013041_, _013051_, _013052_);
  and g_105757_(_013048_, _013049_, _013053_);
  and g_105758_(_013052_, _013053_, _013054_);
  and g_105759_(_000560_, _013031_, _013055_);
  or g_105760_(_012999_, _013055_, _013057_);
  or g_105761_(_013035_, _013057_, _013058_);
  not g_105762_(_013058_, _013059_);
  and g_105763_(_013018_, _013059_, _013060_);
  or g_105764_(_013054_, _013060_, _013061_);
  not g_105765_(_013061_, _013062_);
  and g_105766_(_012907_, _013061_, _013063_);
  and g_105767_(_012911_, _013062_, _013064_);
  or g_105768_(_013063_, _013064_, _013065_);
  not g_105769_(_013065_, _013066_);
  xor g_105770_(out[762], _009685_, _013068_);
  xor g_105771_(_000747_, _009685_, _013069_);
  or g_105772_(_013065_, _013069_, _013070_);
  or g_105773_(_009675_, _009688_, _013071_);
  and g_105774_(_013070_, _013071_, _013072_);
  and g_105775_(_013065_, _013069_, _013073_);
  or g_105776_(_013066_, _013068_, _013074_);
  and g_105777_(out[761], _009684_, _013075_);
  xor g_105778_(out[761], _009684_, _013076_);
  or g_105779_(_009686_, _013075_, _013077_);
  and g_105780_(_012927_, _013061_, _013079_);
  and g_105781_(_012920_, _013062_, _013080_);
  or g_105782_(_013079_, _013080_, _013081_);
  not g_105783_(_013081_, _013082_);
  or g_105784_(_013077_, _013082_, _013083_);
  and g_105785_(_013077_, _013082_, _013084_);
  xor g_105786_(_013077_, _013081_, _013085_);
  xor g_105787_(out[760], _009683_, _013086_);
  and g_105788_(_012932_, _013062_, _013087_);
  and g_105789_(_012939_, _013061_, _013088_);
  or g_105790_(_013087_, _013088_, _013090_);
  not g_105791_(_013090_, _013091_);
  or g_105792_(_013086_, _013090_, _013092_);
  xor g_105793_(_013086_, _013091_, _013093_);
  or g_105794_(_013085_, _013093_, _013094_);
  xor g_105795_(out[759], _009682_, _013095_);
  xor g_105796_(_000637_, _009682_, _013096_);
  and g_105797_(_012950_, _013062_, _013097_);
  and g_105798_(_012954_, _013061_, _013098_);
  or g_105799_(_013097_, _013098_, _013099_);
  or g_105800_(_013096_, _013099_, _013101_);
  xor g_105801_(out[758], _009681_, _013102_);
  not g_105802_(_013102_, _013103_);
  and g_105803_(_012958_, _013062_, _013104_);
  and g_105804_(_012961_, _013061_, _013105_);
  or g_105805_(_013104_, _013105_, _013106_);
  or g_105806_(_013102_, _013106_, _013107_);
  and g_105807_(_013101_, _013107_, _013108_);
  xor g_105808_(out[757], _009678_, _013109_);
  and g_105809_(_012982_, _013062_, _013110_);
  and g_105810_(_012988_, _013061_, _013112_);
  or g_105811_(_013110_, _013112_, _013113_);
  and g_105812_(_013109_, _013113_, _013114_);
  not g_105813_(_013114_, _013115_);
  and g_105814_(_013096_, _013099_, _013116_);
  xor g_105815_(_013096_, _013099_, _013117_);
  xor g_105816_(_013095_, _013099_, _013118_);
  xor g_105817_(_013102_, _013106_, _013119_);
  xor g_105818_(_013103_, _013106_, _013120_);
  and g_105819_(_013117_, _013119_, _013121_);
  or g_105820_(_013118_, _013120_, _013123_);
  and g_105821_(_013115_, _013121_, _013124_);
  or g_105822_(_013114_, _013123_, _013125_);
  or g_105823_(_024144_, _000650_, _013126_);
  and g_105824_(_009680_, _013126_, _013127_);
  and g_105825_(_012977_, _013061_, _013128_);
  and g_105826_(_012971_, _013062_, _013129_);
  or g_105827_(_013128_, _013129_, _013130_);
  and g_105828_(_013127_, _013130_, _013131_);
  or g_105829_(_013127_, _013130_, _013132_);
  not g_105830_(_013132_, _013134_);
  or g_105831_(_013109_, _013113_, _013135_);
  not g_105832_(_013135_, _013136_);
  and g_105833_(_013132_, _013135_, _013137_);
  or g_105834_(_013134_, _013136_, _013138_);
  xor g_105835_(_013127_, _013130_, _013139_);
  and g_105836_(_013135_, _013139_, _013140_);
  or g_105837_(_013131_, _013138_, _013141_);
  and g_105838_(_013124_, _013140_, _013142_);
  or g_105839_(_013125_, _013141_, _013143_);
  xor g_105840_(out[755], _000650_, _013145_);
  xor g_105841_(_000714_, _000650_, _013146_);
  and g_105842_(_013005_, _013062_, _013147_);
  and g_105843_(_013009_, _013061_, _013148_);
  or g_105844_(_013147_, _013148_, _013149_);
  or g_105845_(_013146_, _013149_, _013150_);
  and g_105846_(_013003_, _013061_, _013151_);
  or g_105847_(_000363_, _013061_, _013152_);
  not g_105848_(_013152_, _013153_);
  or g_105849_(_013151_, _013153_, _013154_);
  or g_105850_(_000652_, _013154_, _013156_);
  and g_105851_(_013150_, _013156_, _013157_);
  and g_105852_(_013146_, _013149_, _013158_);
  xor g_105853_(_013146_, _013149_, _013159_);
  xor g_105854_(_013145_, _013149_, _013160_);
  xor g_105855_(_000652_, _013154_, _013161_);
  xor g_105856_(_000651_, _013154_, _013162_);
  and g_105857_(_013159_, _013161_, _013163_);
  or g_105858_(_013160_, _013162_, _013164_);
  and g_105859_(_013022_, _013061_, _013165_);
  not g_105860_(_013165_, _013167_);
  or g_105861_(out[737], _013061_, _013168_);
  not g_105862_(_013168_, _013169_);
  or g_105863_(_013165_, _013169_, _013170_);
  and g_105864_(_013167_, _013168_, _013171_);
  or g_105865_(_000681_, _013171_, _013172_);
  or g_105866_(_000560_, _013061_, _013173_);
  or g_105867_(_013030_, _013062_, _013174_);
  and g_105868_(_013173_, _013174_, _013175_);
  and g_105869_(out[752], _013175_, _013176_);
  xor g_105870_(_000681_, _013170_, _013178_);
  or g_105871_(_013176_, _013178_, _013179_);
  and g_105872_(_013172_, _013179_, _013180_);
  or g_105873_(_013164_, _013180_, _013181_);
  or g_105874_(_013157_, _013158_, _013182_);
  and g_105875_(_013181_, _013182_, _013183_);
  or g_105876_(_013143_, _013183_, _013184_);
  or g_105877_(_013108_, _013116_, _013185_);
  or g_105878_(_013125_, _013137_, _013186_);
  and g_105879_(_013185_, _013186_, _013187_);
  and g_105880_(_013184_, _013187_, _013189_);
  or g_105881_(_013094_, _013189_, _013190_);
  or g_105882_(_013084_, _013092_, _013191_);
  and g_105883_(_013083_, _013191_, _013192_);
  and g_105884_(_013190_, _013192_, _013193_);
  or g_105885_(_013073_, _013193_, _013194_);
  and g_105886_(_013072_, _013194_, _013195_);
  and g_105887_(_009675_, _009688_, _013196_);
  or g_105888_(_009674_, _009689_, _013197_);
  or g_105889_(_013094_, _013179_, _013198_);
  not g_105890_(_013198_, _013200_);
  and g_105891_(_013163_, _013200_, _013201_);
  and g_105892_(_013074_, _013197_, _013202_);
  or g_105893_(out[752], _013175_, _013203_);
  and g_105894_(_013202_, _013203_, _013204_);
  and g_105895_(_013072_, _013204_, _013205_);
  and g_105896_(_013201_, _013205_, _013206_);
  and g_105897_(_013142_, _013206_, _013207_);
  or g_105898_(_013196_, _013207_, _013208_);
  or g_105899_(_013195_, _013208_, _013209_);
  and g_105900_(_013065_, _013209_, _013211_);
  not g_105901_(_013211_, _013212_);
  or g_105902_(_013069_, _013209_, _013213_);
  and g_105903_(_013212_, _013213_, _013214_);
  or g_105904_(_009692_, _009704_, _013215_);
  xor g_105905_(out[778], _009702_, _013216_);
  not g_105906_(_013216_, _013217_);
  and g_105907_(_013214_, _013216_, _013218_);
  not g_105908_(_013218_, _013219_);
  and g_105909_(_013215_, _013219_, _013220_);
  and g_105910_(_009692_, _009704_, _013222_);
  and g_105911_(out[777], _009700_, _013223_);
  xor g_105912_(out[777], _009700_, _013224_);
  xor g_105913_(_000868_, _009700_, _013225_);
  and g_105914_(_013081_, _013209_, _013226_);
  not g_105915_(_013226_, _013227_);
  or g_105916_(_013076_, _013209_, _013228_);
  and g_105917_(_013227_, _013228_, _013229_);
  and g_105918_(_013225_, _013229_, _013230_);
  xor g_105919_(out[776], _009699_, _013231_);
  xor g_105920_(_000857_, _009699_, _013233_);
  or g_105921_(_013086_, _013209_, _013234_);
  not g_105922_(_013234_, _013235_);
  and g_105923_(_013090_, _013209_, _013236_);
  or g_105924_(_013235_, _013236_, _013237_);
  or g_105925_(_013225_, _013229_, _013238_);
  or g_105926_(_013231_, _013237_, _013239_);
  and g_105927_(_013238_, _013239_, _013240_);
  xor g_105928_(_013233_, _013237_, _013241_);
  xor g_105929_(_009691_, _009704_, _013242_);
  xor g_105930_(_013214_, _013217_, _013244_);
  or g_105931_(_013242_, _013244_, _013245_);
  xor g_105932_(_013224_, _013229_, _013246_);
  or g_105933_(_013245_, _013246_, _013247_);
  or g_105934_(_013241_, _013247_, _013248_);
  xor g_105935_(out[774], _009697_, _013249_);
  not g_105936_(_013249_, _013250_);
  and g_105937_(_013106_, _013209_, _013251_);
  or g_105938_(_013102_, _013209_, _013252_);
  not g_105939_(_013252_, _013253_);
  or g_105940_(_013251_, _013253_, _013255_);
  not g_105941_(_013255_, _013256_);
  or g_105942_(_013249_, _013255_, _013257_);
  xor g_105943_(_013250_, _013255_, _013258_);
  xor g_105944_(out[775], _009698_, _013259_);
  xor g_105945_(_000769_, _009698_, _013260_);
  and g_105946_(_013099_, _013209_, _013261_);
  or g_105947_(_013096_, _013209_, _013262_);
  not g_105948_(_013262_, _013263_);
  or g_105949_(_013261_, _013263_, _013264_);
  and g_105950_(_013260_, _013264_, _013266_);
  or g_105951_(_013260_, _013264_, _013267_);
  xor g_105952_(_013259_, _013264_, _013268_);
  or g_105953_(_013258_, _013268_, _013269_);
  or g_105954_(_024298_, _000827_, _013270_);
  not g_105955_(_013270_, _013271_);
  and g_105956_(_009696_, _013270_, _013272_);
  or g_105957_(_009695_, _013271_, _013273_);
  and g_105958_(_013130_, _013209_, _013274_);
  or g_105959_(_013127_, _013209_, _013275_);
  not g_105960_(_013275_, _013277_);
  or g_105961_(_013274_, _013277_, _013278_);
  or g_105962_(_013272_, _013278_, _013279_);
  xor g_105963_(out[773], _009695_, _013280_);
  xor g_105964_(_000791_, _009695_, _013281_);
  and g_105965_(_013113_, _013209_, _013282_);
  or g_105966_(_013109_, _013209_, _013283_);
  not g_105967_(_013283_, _013284_);
  or g_105968_(_013282_, _013284_, _013285_);
  or g_105969_(_013280_, _013285_, _013286_);
  and g_105970_(_013279_, _013286_, _013288_);
  not g_105971_(_013288_, _013289_);
  and g_105972_(_013272_, _013278_, _013290_);
  and g_105973_(_013280_, _013285_, _013291_);
  or g_105974_(_013290_, _013291_, _013292_);
  or g_105975_(_013289_, _013292_, _013293_);
  or g_105976_(_013248_, _013293_, _013294_);
  or g_105977_(_013269_, _013294_, _013295_);
  not g_105978_(_013295_, _013296_);
  and g_105979_(_013154_, _013209_, _013297_);
  or g_105980_(_000652_, _013209_, _013299_);
  not g_105981_(_013299_, _013300_);
  or g_105982_(_013297_, _013300_, _013301_);
  or g_105983_(_000829_, _013301_, _013302_);
  xor g_105984_(out[771], _000827_, _013303_);
  xor g_105985_(_000846_, _000827_, _013304_);
  and g_105986_(_013149_, _013209_, _013305_);
  or g_105987_(_013146_, _013209_, _013306_);
  not g_105988_(_013306_, _013307_);
  or g_105989_(_013305_, _013307_, _013308_);
  and g_105990_(_013304_, _013308_, _013310_);
  not g_105991_(_013310_, _013311_);
  xor g_105992_(_000829_, _013301_, _013312_);
  xor g_105993_(_000828_, _013301_, _013313_);
  and g_105994_(_013311_, _013312_, _013314_);
  or g_105995_(_013310_, _013313_, _013315_);
  or g_105996_(out[753], _013209_, _013316_);
  not g_105997_(_013316_, _013317_);
  and g_105998_(_013170_, _013209_, _013318_);
  or g_105999_(_013317_, _013318_, _013319_);
  and g_106000_(_013175_, _013209_, _013321_);
  or g_106001_(out[752], _013209_, _013322_);
  not g_106002_(_013322_, _013323_);
  or g_106003_(_013321_, _013323_, _013324_);
  and g_106004_(out[768], _013324_, _013325_);
  not g_106005_(_013325_, _013326_);
  and g_106006_(out[769], _013319_, _013327_);
  not g_106007_(_013327_, _013328_);
  xor g_106008_(out[769], _013319_, _013329_);
  xor g_106009_(_000813_, _013319_, _013330_);
  and g_106010_(_013326_, _013329_, _013332_);
  or g_106011_(_013325_, _013330_, _013333_);
  or g_106012_(_013304_, _013308_, _013334_);
  or g_106013_(out[768], _013324_, _013335_);
  and g_106014_(_013334_, _013335_, _013336_);
  and g_106015_(_013332_, _013336_, _013337_);
  and g_106016_(_013314_, _013337_, _013338_);
  and g_106017_(_013296_, _013338_, _013339_);
  or g_106018_(_013302_, _013310_, _013340_);
  and g_106019_(_013334_, _013340_, _013341_);
  and g_106020_(_013328_, _013333_, _013343_);
  or g_106021_(_013315_, _013343_, _013344_);
  and g_106022_(_013341_, _013344_, _013345_);
  or g_106023_(_013295_, _013345_, _013346_);
  or g_106024_(_013269_, _013288_, _013347_);
  or g_106025_(_013291_, _013347_, _013348_);
  or g_106026_(_013257_, _013266_, _013349_);
  and g_106027_(_013267_, _013349_, _013350_);
  and g_106028_(_013348_, _013350_, _013351_);
  or g_106029_(_013248_, _013351_, _013352_);
  or g_106030_(_013220_, _013222_, _013354_);
  or g_106031_(_013240_, _013245_, _013355_);
  or g_106032_(_013230_, _013355_, _013356_);
  and g_106033_(_013354_, _013356_, _013357_);
  and g_106034_(_013352_, _013357_, _013358_);
  and g_106035_(_013346_, _013358_, _013359_);
  or g_106036_(_013339_, _013359_, _013360_);
  not g_106037_(_013360_, _013361_);
  or g_106038_(_013216_, _013360_, _013362_);
  and g_106039_(_013214_, _013360_, _013363_);
  not g_106040_(_013363_, _013365_);
  and g_106041_(_013362_, _013365_, _013366_);
  not g_106042_(_013366_, _013367_);
  or g_106043_(_024452_, _001009_, _013368_);
  not g_106044_(_013368_, _013369_);
  and g_106045_(_009711_, _013368_, _013370_);
  or g_106046_(_009710_, _013369_, _013371_);
  and g_106047_(_013278_, _013360_, _013372_);
  and g_106048_(_013273_, _013361_, _013373_);
  or g_106049_(_013372_, _013373_, _013374_);
  or g_106050_(_013370_, _013374_, _013376_);
  and g_106051_(_013285_, _013360_, _013377_);
  and g_106052_(_013281_, _013361_, _013378_);
  or g_106053_(_013377_, _013378_, _013379_);
  xor g_106054_(out[789], _009710_, _013380_);
  xor g_106055_(_000923_, _009710_, _013381_);
  or g_106056_(_013379_, _013380_, _013382_);
  and g_106057_(_013376_, _013382_, _013383_);
  and g_106058_(_013370_, _013374_, _013384_);
  xor g_106059_(out[787], _001009_, _013385_);
  xor g_106060_(_000978_, _001009_, _013387_);
  and g_106061_(_013308_, _013360_, _013388_);
  and g_106062_(_013303_, _013361_, _013389_);
  or g_106063_(_013388_, _013389_, _013390_);
  and g_106064_(_013387_, _013390_, _013391_);
  or g_106065_(_013384_, _013391_, _013392_);
  or g_106066_(_013387_, _013390_, _013393_);
  and g_106067_(_000828_, _013361_, _013394_);
  and g_106068_(_013301_, _013360_, _013395_);
  or g_106069_(_013394_, _013395_, _013396_);
  or g_106070_(_001012_, _013396_, _013398_);
  and g_106071_(_013393_, _013398_, _013399_);
  and g_106072_(_001012_, _013396_, _013400_);
  and g_106073_(_013319_, _013360_, _013401_);
  not g_106074_(_013401_, _013402_);
  or g_106075_(out[769], _013360_, _013403_);
  and g_106076_(_013402_, _013403_, _013404_);
  or g_106077_(_000945_, _013404_, _013405_);
  or g_106078_(_000824_, _013360_, _013406_);
  or g_106079_(_013324_, _013361_, _013407_);
  and g_106080_(_013406_, _013407_, _013409_);
  or g_106081_(out[784], _013409_, _013410_);
  and g_106082_(out[784], _013409_, _013411_);
  and g_106083_(_000945_, _013404_, _013412_);
  or g_106084_(_013411_, _013412_, _013413_);
  or g_106085_(_013410_, _013413_, _013414_);
  and g_106086_(_013405_, _013414_, _013415_);
  or g_106087_(_013400_, _013415_, _013416_);
  and g_106088_(_013399_, _013416_, _013417_);
  or g_106089_(_013392_, _013417_, _013418_);
  and g_106090_(_013383_, _013418_, _013420_);
  and g_106091_(out[793], _009716_, _013421_);
  xor g_106092_(out[793], _009716_, _013422_);
  xor g_106093_(_001000_, _009716_, _013423_);
  or g_106094_(_013229_, _013361_, _013424_);
  or g_106095_(_013224_, _013360_, _013425_);
  and g_106096_(_013424_, _013425_, _013426_);
  not g_106097_(_013426_, _013427_);
  or g_106098_(_013423_, _013426_, _013428_);
  xor g_106099_(out[792], _009715_, _013429_);
  not g_106100_(_013429_, _013431_);
  and g_106101_(_013233_, _013361_, _013432_);
  and g_106102_(_013237_, _013360_, _013433_);
  or g_106103_(_013432_, _013433_, _013434_);
  or g_106104_(_013429_, _013434_, _013435_);
  and g_106105_(_013423_, _013426_, _013436_);
  and g_106106_(_009707_, _009719_, _013437_);
  xor g_106107_(out[794], _009717_, _013438_);
  not g_106108_(_013438_, _013439_);
  and g_106109_(_013366_, _013439_, _013440_);
  or g_106110_(_013437_, _013440_, _013442_);
  or g_106111_(_009707_, _009719_, _013443_);
  not g_106112_(_013443_, _013444_);
  and g_106113_(_013367_, _013438_, _013445_);
  or g_106114_(_013366_, _013439_, _013446_);
  and g_106115_(_013443_, _013446_, _013447_);
  or g_106116_(_013444_, _013445_, _013448_);
  xor g_106117_(_013422_, _013426_, _013449_);
  or g_106118_(_013442_, _013449_, _013450_);
  xor g_106119_(_013431_, _013434_, _013451_);
  or g_106120_(_013448_, _013451_, _013453_);
  or g_106121_(_013450_, _013453_, _013454_);
  xor g_106122_(out[790], _009713_, _013455_);
  not g_106123_(_013455_, _013456_);
  or g_106124_(_013256_, _013361_, _013457_);
  or g_106125_(_013249_, _013360_, _013458_);
  and g_106126_(_013457_, _013458_, _013459_);
  not g_106127_(_013459_, _013460_);
  or g_106128_(_013455_, _013460_, _013461_);
  xor g_106129_(out[791], _009714_, _013462_);
  xor g_106130_(_000901_, _009714_, _013464_);
  and g_106131_(_013259_, _013361_, _013465_);
  and g_106132_(_013264_, _013360_, _013466_);
  or g_106133_(_013465_, _013466_, _013467_);
  or g_106134_(_013464_, _013467_, _013468_);
  and g_106135_(_013379_, _013380_, _013469_);
  and g_106136_(_013464_, _013467_, _013470_);
  xor g_106137_(_013455_, _013459_, _013471_);
  xor g_106138_(_013462_, _013467_, _013472_);
  or g_106139_(_013471_, _013472_, _013473_);
  or g_106140_(_013469_, _013473_, _013475_);
  or g_106141_(_013454_, _013475_, _013476_);
  or g_106142_(_013420_, _013476_, _013477_);
  or g_106143_(_013435_, _013436_, _013478_);
  and g_106144_(_013428_, _013478_, _013479_);
  or g_106145_(_013442_, _013479_, _013480_);
  or g_106146_(_013437_, _013447_, _013481_);
  and g_106147_(_013480_, _013481_, _013482_);
  or g_106148_(_013461_, _013470_, _013483_);
  and g_106149_(_013468_, _013483_, _013484_);
  or g_106150_(_013454_, _013484_, _013486_);
  and g_106151_(_013482_, _013486_, _013487_);
  and g_106152_(_013477_, _013487_, _013488_);
  not g_106153_(_013488_, _013489_);
  and g_106154_(_013366_, _013488_, _013490_);
  not g_106155_(_013490_, _013491_);
  and g_106156_(_013438_, _013489_, _013492_);
  or g_106157_(_013439_, _013488_, _013493_);
  and g_106158_(_013491_, _013493_, _013494_);
  or g_106159_(_013490_, _013492_, _013495_);
  xor g_106160_(out[806], _009728_, _013497_);
  xor g_106161_(_001044_, _009728_, _013498_);
  or g_106162_(_013455_, _013488_, _013499_);
  or g_106163_(_013459_, _013489_, _013500_);
  and g_106164_(_013499_, _013500_, _013501_);
  not g_106165_(_013501_, _013502_);
  and g_106166_(_013498_, _013501_, _013503_);
  or g_106167_(_013497_, _013502_, _013504_);
  xor g_106168_(out[807], _009729_, _013505_);
  xor g_106169_(_001033_, _009729_, _013506_);
  and g_106170_(_013462_, _013489_, _013508_);
  or g_106171_(_013464_, _013488_, _013509_);
  and g_106172_(_013467_, _013488_, _013510_);
  not g_106173_(_013510_, _013511_);
  and g_106174_(_013509_, _013511_, _013512_);
  or g_106175_(_013508_, _013510_, _013513_);
  and g_106176_(_013505_, _013512_, _013514_);
  or g_106177_(_013506_, _013513_, _013515_);
  xor g_106178_(out[805], _009726_, _013516_);
  and g_106179_(_013381_, _013489_, _013517_);
  and g_106180_(_013379_, _013488_, _013519_);
  or g_106181_(_013517_, _013519_, _013520_);
  and g_106182_(_013516_, _013520_, _013521_);
  not g_106183_(_013521_, _013522_);
  and g_106184_(_013506_, _013513_, _013523_);
  or g_106185_(_013505_, _013512_, _013524_);
  xor g_106186_(_013498_, _013501_, _013525_);
  xor g_106187_(_013497_, _013501_, _013526_);
  and g_106188_(_013515_, _013525_, _013527_);
  or g_106189_(_013514_, _013526_, _013528_);
  and g_106190_(_013524_, _013527_, _013530_);
  or g_106191_(_013523_, _013528_, _013531_);
  and g_106192_(_013522_, _013530_, _013532_);
  or g_106193_(_013521_, _013531_, _013533_);
  xor g_106194_(out[810], _009732_, _013534_);
  xor g_106195_(_001143_, _009732_, _013535_);
  and g_106196_(_013495_, _013535_, _013536_);
  xor g_106197_(out[808], _009730_, _013537_);
  and g_106198_(_013431_, _013489_, _013538_);
  and g_106199_(_013434_, _013488_, _013539_);
  or g_106200_(_013538_, _013539_, _013541_);
  or g_106201_(_013537_, _013541_, _013542_);
  not g_106202_(_013542_, _013543_);
  and g_106203_(_013537_, _013541_, _013544_);
  and g_106204_(out[809], _009731_, _013545_);
  xor g_106205_(out[809], _009731_, _013546_);
  or g_106206_(_009733_, _013545_, _013547_);
  and g_106207_(_013427_, _013488_, _013548_);
  and g_106208_(_013423_, _013489_, _013549_);
  or g_106209_(_013548_, _013549_, _013550_);
  not g_106210_(_013550_, _013552_);
  and g_106211_(_013547_, _013552_, _013553_);
  or g_106212_(_013546_, _013550_, _013554_);
  and g_106213_(_013494_, _013534_, _013555_);
  or g_106214_(_013495_, _013535_, _013556_);
  and g_106215_(_009721_, _009737_, _013557_);
  or g_106216_(_009722_, _009736_, _013558_);
  and g_106217_(_013556_, _013558_, _013559_);
  or g_106218_(_013555_, _013557_, _013560_);
  and g_106219_(_009722_, _009736_, _013561_);
  and g_106220_(_013546_, _013550_, _013563_);
  xor g_106221_(_013537_, _013541_, _013564_);
  or g_106222_(_013536_, _013561_, _013565_);
  not g_106223_(_013565_, _013566_);
  and g_106224_(_013559_, _013566_, _013567_);
  or g_106225_(_013560_, _013565_, _013568_);
  xor g_106226_(_013546_, _013550_, _013569_);
  and g_106227_(_013567_, _013569_, _013570_);
  or g_106228_(_013544_, _013563_, _013571_);
  or g_106229_(_013543_, _013553_, _013572_);
  or g_106230_(_013571_, _013572_, _013574_);
  and g_106231_(_013564_, _013570_, _013575_);
  or g_106232_(_013568_, _013574_, _013576_);
  or g_106233_(_024606_, _001210_, _013577_);
  and g_106234_(_009727_, _013577_, _013578_);
  and g_106235_(_013374_, _013488_, _013579_);
  and g_106236_(_013371_, _013489_, _013580_);
  or g_106237_(_013579_, _013580_, _013581_);
  and g_106238_(_013578_, _013581_, _013582_);
  not g_106239_(_013582_, _013583_);
  or g_106240_(_013578_, _013581_, _013585_);
  not g_106241_(_013585_, _013586_);
  or g_106242_(_013516_, _013520_, _013587_);
  not g_106243_(_013587_, _013588_);
  and g_106244_(_013585_, _013587_, _013589_);
  or g_106245_(_013586_, _013588_, _013590_);
  and g_106246_(_013583_, _013589_, _013591_);
  or g_106247_(_013582_, _013590_, _013592_);
  and g_106248_(_013575_, _013591_, _013593_);
  or g_106249_(_013576_, _013592_, _013594_);
  and g_106250_(_013532_, _013593_, _013596_);
  or g_106251_(_013533_, _013594_, _013597_);
  xor g_106252_(out[803], _001210_, _013598_);
  xor g_106253_(_001110_, _001210_, _013599_);
  and g_106254_(_013385_, _013489_, _013600_);
  and g_106255_(_013390_, _013488_, _013601_);
  or g_106256_(_013600_, _013601_, _013602_);
  and g_106257_(_013599_, _013602_, _013603_);
  and g_106258_(_013396_, _013488_, _013604_);
  and g_106259_(_001010_, _013489_, _013605_);
  or g_106260_(_013604_, _013605_, _013607_);
  or g_106261_(_001212_, _013607_, _013608_);
  or g_106262_(_013599_, _013602_, _013609_);
  xor g_106263_(_013599_, _013602_, _013610_);
  xor g_106264_(_013598_, _013602_, _013611_);
  xor g_106265_(_001212_, _013607_, _013612_);
  xor g_106266_(_001211_, _013607_, _013613_);
  and g_106267_(_013610_, _013612_, _013614_);
  or g_106268_(_013611_, _013613_, _013615_);
  or g_106269_(_000956_, _013488_, _013616_);
  or g_106270_(_013409_, _013489_, _013618_);
  and g_106271_(_013616_, _013618_, _013619_);
  and g_106272_(out[800], _013619_, _013620_);
  and g_106273_(out[785], _013489_, _013621_);
  or g_106274_(_000945_, _013488_, _013622_);
  and g_106275_(_013404_, _013488_, _013623_);
  not g_106276_(_013623_, _013624_);
  and g_106277_(_013622_, _013624_, _013625_);
  or g_106278_(_013621_, _013623_, _013626_);
  and g_106279_(out[801], _013625_, _013627_);
  or g_106280_(_001077_, _013626_, _013629_);
  xor g_106281_(_001077_, _013625_, _013630_);
  or g_106282_(_013620_, _013630_, _013631_);
  not g_106283_(_013631_, _013632_);
  and g_106284_(_013614_, _013632_, _013633_);
  or g_106285_(_013615_, _013631_, _013634_);
  and g_106286_(_013614_, _013627_, _013635_);
  or g_106287_(_013615_, _013629_, _013636_);
  and g_106288_(_013608_, _013609_, _013637_);
  or g_106289_(_013603_, _013637_, _013638_);
  and g_106290_(_013634_, _013638_, _013640_);
  not g_106291_(_013640_, _013641_);
  and g_106292_(_013636_, _013640_, _013642_);
  or g_106293_(_013635_, _013641_, _013643_);
  and g_106294_(_013596_, _013643_, _013644_);
  or g_106295_(_013597_, _013642_, _013645_);
  or g_106296_(_013533_, _013589_, _013646_);
  not g_106297_(_013646_, _013647_);
  and g_106298_(_013503_, _013524_, _013648_);
  or g_106299_(_013504_, _013523_, _013649_);
  and g_106300_(_013515_, _013649_, _013651_);
  or g_106301_(_013514_, _013648_, _013652_);
  and g_106302_(_013646_, _013651_, _013653_);
  or g_106303_(_013647_, _013652_, _013654_);
  and g_106304_(_013575_, _013654_, _013655_);
  or g_106305_(_013576_, _013653_, _013656_);
  and g_106306_(_013543_, _013554_, _013657_);
  or g_106307_(_013563_, _013657_, _013658_);
  and g_106308_(_013567_, _013658_, _013659_);
  not g_106309_(_013659_, _013660_);
  or g_106310_(_013559_, _013561_, _013662_);
  not g_106311_(_013662_, _013663_);
  and g_106312_(_013645_, _013660_, _013664_);
  or g_106313_(_013644_, _013659_, _013665_);
  and g_106314_(_013656_, _013662_, _013666_);
  or g_106315_(_013655_, _013663_, _013667_);
  and g_106316_(_013664_, _013666_, _013668_);
  or g_106317_(_013665_, _013667_, _013669_);
  or g_106318_(out[800], _013619_, _013670_);
  and g_106319_(_013596_, _013670_, _013671_);
  not g_106320_(_013671_, _013673_);
  and g_106321_(_013633_, _013671_, _013674_);
  or g_106322_(_013634_, _013673_, _013675_);
  and g_106323_(_013669_, _013675_, _013676_);
  or g_106324_(_013668_, _013674_, _013677_);
  and g_106325_(_013495_, _013677_, _013678_);
  not g_106326_(_013678_, _013679_);
  or g_106327_(_013535_, _013677_, _013680_);
  not g_106328_(_013680_, _013681_);
  and g_106329_(_013679_, _013680_, _013682_);
  or g_106330_(_013678_, _013681_, _013684_);
  xor g_106331_(out[826], _009749_, _013685_);
  xor g_106332_(_001275_, _009749_, _013686_);
  and g_106333_(_013682_, _013685_, _013687_);
  or g_106334_(_013684_, _013686_, _013688_);
  and g_106335_(_009738_, _009753_, _013689_);
  or g_106336_(_009739_, _009752_, _013690_);
  and g_106337_(_013688_, _013690_, _013691_);
  or g_106338_(_013687_, _013689_, _013692_);
  and g_106339_(_013684_, _013686_, _013693_);
  or g_106340_(_013682_, _013685_, _013695_);
  and g_106341_(_009739_, _009752_, _013696_);
  or g_106342_(_009738_, _009753_, _013697_);
  and g_106343_(out[825], _009748_, _013698_);
  xor g_106344_(out[825], _009748_, _013699_);
  or g_106345_(_009750_, _013698_, _013700_);
  and g_106346_(_013550_, _013677_, _013701_);
  not g_106347_(_013701_, _013702_);
  or g_106348_(_013546_, _013677_, _013703_);
  not g_106349_(_013703_, _013704_);
  and g_106350_(_013702_, _013703_, _013706_);
  or g_106351_(_013701_, _013704_, _013707_);
  and g_106352_(_013700_, _013706_, _013708_);
  or g_106353_(_013699_, _013707_, _013709_);
  and g_106354_(_013697_, _013709_, _013710_);
  or g_106355_(_013696_, _013708_, _013711_);
  and g_106356_(_013695_, _013710_, _013712_);
  or g_106357_(_013693_, _013711_, _013713_);
  and g_106358_(_013691_, _013712_, _013714_);
  or g_106359_(_013692_, _013713_, _013715_);
  xor g_106360_(out[824], _009747_, _013717_);
  xor g_106361_(_001253_, _009747_, _013718_);
  or g_106362_(_013537_, _013677_, _013719_);
  not g_106363_(_013719_, _013720_);
  and g_106364_(_013541_, _013677_, _013721_);
  not g_106365_(_013721_, _013722_);
  and g_106366_(_013719_, _013722_, _013723_);
  or g_106367_(_013720_, _013721_, _013724_);
  and g_106368_(_013717_, _013724_, _013725_);
  or g_106369_(_013718_, _013723_, _013726_);
  and g_106370_(_013699_, _013707_, _013728_);
  or g_106371_(_013700_, _013706_, _013729_);
  and g_106372_(_013718_, _013723_, _013730_);
  or g_106373_(_013717_, _013724_, _013731_);
  and g_106374_(_013729_, _013731_, _013732_);
  or g_106375_(_013728_, _013730_, _013733_);
  and g_106376_(_013726_, _013732_, _013734_);
  or g_106377_(_013725_, _013733_, _013735_);
  and g_106378_(_013714_, _013734_, _013736_);
  or g_106379_(_013715_, _013735_, _013737_);
  xor g_106380_(out[823], _009746_, _013739_);
  xor g_106381_(_001165_, _009746_, _013740_);
  and g_106382_(_013505_, _013676_, _013741_);
  or g_106383_(_013506_, _013677_, _013742_);
  and g_106384_(_013513_, _013677_, _013743_);
  or g_106385_(_013512_, _013676_, _013744_);
  and g_106386_(_013742_, _013744_, _013745_);
  or g_106387_(_013741_, _013743_, _013746_);
  and g_106388_(_013739_, _013745_, _013747_);
  or g_106389_(_013740_, _013746_, _013748_);
  xor g_106390_(out[822], _009744_, _013750_);
  not g_106391_(_013750_, _013751_);
  and g_106392_(_013498_, _013676_, _013752_);
  and g_106393_(_013502_, _013677_, _013753_);
  or g_106394_(_013752_, _013753_, _013754_);
  or g_106395_(_013750_, _013754_, _013755_);
  not g_106396_(_013755_, _013756_);
  and g_106397_(_013740_, _013746_, _013757_);
  or g_106398_(_013739_, _013745_, _013758_);
  and g_106399_(_013748_, _013758_, _013759_);
  or g_106400_(_013747_, _013757_, _013761_);
  xor g_106401_(_013750_, _013754_, _013762_);
  xor g_106402_(_013751_, _013754_, _013763_);
  and g_106403_(_013759_, _013762_, _013764_);
  or g_106404_(_013761_, _013763_, _013765_);
  or g_106405_(_024760_, _001338_, _013766_);
  not g_106406_(_013766_, _013767_);
  and g_106407_(_009743_, _013766_, _013768_);
  or g_106408_(_009742_, _013767_, _013769_);
  and g_106409_(_013581_, _013677_, _013770_);
  not g_106410_(_013770_, _013772_);
  or g_106411_(_013578_, _013677_, _013773_);
  not g_106412_(_013773_, _013774_);
  and g_106413_(_013772_, _013773_, _013775_);
  or g_106414_(_013770_, _013774_, _013776_);
  and g_106415_(_013769_, _013775_, _013777_);
  or g_106416_(_013768_, _013776_, _013778_);
  xor g_106417_(out[821], _009742_, _013779_);
  xor g_106418_(_001187_, _009742_, _013780_);
  or g_106419_(_013516_, _013677_, _013781_);
  not g_106420_(_013781_, _013783_);
  and g_106421_(_013520_, _013677_, _013784_);
  not g_106422_(_013784_, _013785_);
  and g_106423_(_013781_, _013785_, _013786_);
  or g_106424_(_013783_, _013784_, _013787_);
  and g_106425_(_013780_, _013786_, _013788_);
  or g_106426_(_013779_, _013787_, _013789_);
  and g_106427_(_013778_, _013789_, _013790_);
  or g_106428_(_013777_, _013788_, _013791_);
  and g_106429_(_013779_, _013787_, _013792_);
  not g_106430_(_013792_, _013794_);
  or g_106431_(_013769_, _013775_, _013795_);
  and g_106432_(_013794_, _013795_, _013796_);
  and g_106433_(_013790_, _013796_, _013797_);
  and g_106434_(_013764_, _013797_, _013798_);
  not g_106435_(_013798_, _013799_);
  and g_106436_(_013736_, _013798_, _013800_);
  or g_106437_(_013737_, _013799_, _013801_);
  xor g_106438_(out[819], _001338_, _013802_);
  xor g_106439_(_001242_, _001338_, _013803_);
  and g_106440_(_013598_, _013676_, _013805_);
  and g_106441_(_013602_, _013677_, _013806_);
  or g_106442_(_013805_, _013806_, _013807_);
  or g_106443_(_013803_, _013807_, _013808_);
  and g_106444_(_013607_, _013677_, _013809_);
  and g_106445_(_001211_, _013676_, _013810_);
  or g_106446_(_013809_, _013810_, _013811_);
  or g_106447_(_001340_, _013811_, _013812_);
  and g_106448_(_013808_, _013812_, _013813_);
  and g_106449_(_013803_, _013807_, _013814_);
  xor g_106450_(_013803_, _013807_, _013816_);
  xor g_106451_(_001340_, _013811_, _013817_);
  and g_106452_(_013816_, _013817_, _013818_);
  or g_106453_(_001077_, _013677_, _013819_);
  or g_106454_(_013625_, _013676_, _013820_);
  and g_106455_(_013819_, _013820_, _013821_);
  and g_106456_(out[817], _013821_, _013822_);
  or g_106457_(_001088_, _013677_, _013823_);
  or g_106458_(_013619_, _013676_, _013824_);
  and g_106459_(_013823_, _013824_, _013825_);
  and g_106460_(out[816], _013825_, _013827_);
  not g_106461_(_013827_, _013828_);
  xor g_106462_(out[817], _013821_, _013829_);
  xor g_106463_(_001209_, _013821_, _013830_);
  and g_106464_(_013828_, _013829_, _013831_);
  or g_106465_(_013827_, _013830_, _013832_);
  or g_106466_(_013822_, _013831_, _013833_);
  and g_106467_(_013818_, _013833_, _013834_);
  not g_106468_(_013834_, _013835_);
  or g_106469_(_013813_, _013814_, _013836_);
  not g_106470_(_013836_, _013838_);
  and g_106471_(_013835_, _013836_, _013839_);
  or g_106472_(_013834_, _013838_, _013840_);
  and g_106473_(_013800_, _013840_, _013841_);
  or g_106474_(_013801_, _013839_, _013842_);
  and g_106475_(_013791_, _013794_, _013843_);
  or g_106476_(_013790_, _013792_, _013844_);
  and g_106477_(_013764_, _013843_, _013845_);
  or g_106478_(_013765_, _013844_, _013846_);
  and g_106479_(_013756_, _013758_, _013847_);
  or g_106480_(_013755_, _013757_, _013849_);
  and g_106481_(_013748_, _013849_, _013850_);
  or g_106482_(_013747_, _013847_, _013851_);
  and g_106483_(_013846_, _013850_, _013852_);
  or g_106484_(_013845_, _013851_, _013853_);
  and g_106485_(_013736_, _013853_, _013854_);
  or g_106486_(_013737_, _013852_, _013855_);
  and g_106487_(_013714_, _013733_, _013856_);
  or g_106488_(_013715_, _013732_, _013857_);
  and g_106489_(_013692_, _013697_, _013858_);
  or g_106490_(_013691_, _013696_, _013860_);
  and g_106491_(_013857_, _013860_, _013861_);
  or g_106492_(_013856_, _013858_, _013862_);
  and g_106493_(_013855_, _013861_, _013863_);
  or g_106494_(_013854_, _013862_, _013864_);
  and g_106495_(_013842_, _013863_, _013865_);
  or g_106496_(_013841_, _013864_, _013866_);
  or g_106497_(out[816], _013825_, _013867_);
  and g_106498_(_013818_, _013867_, _013868_);
  not g_106499_(_013868_, _013869_);
  and g_106500_(_013831_, _013868_, _013871_);
  or g_106501_(_013832_, _013869_, _013872_);
  and g_106502_(_013800_, _013871_, _013873_);
  or g_106503_(_013801_, _013872_, _013874_);
  and g_106504_(_013866_, _013874_, _013875_);
  or g_106505_(_013865_, _013873_, _013876_);
  and g_106506_(_013684_, _013876_, _013877_);
  or g_106507_(_013682_, _013875_, _013878_);
  and g_106508_(_013685_, _013875_, _013879_);
  or g_106509_(_013686_, _013876_, _013880_);
  and g_106510_(_013878_, _013880_, _013882_);
  or g_106511_(_013877_, _013879_, _013883_);
  and g_106512_(_013811_, _013876_, _013884_);
  and g_106513_(_001339_, _013875_, _013885_);
  or g_106514_(_013884_, _013885_, _013886_);
  or g_106515_(_001516_, _013886_, _013887_);
  xor g_106516_(out[835], _001514_, _013888_);
  xor g_106517_(_001374_, _001514_, _013889_);
  and g_106518_(_013807_, _013876_, _013890_);
  and g_106519_(_013802_, _013875_, _013891_);
  or g_106520_(_013890_, _013891_, _013893_);
  or g_106521_(_013889_, _013893_, _013894_);
  and g_106522_(_013887_, _013894_, _013895_);
  and g_106523_(_013889_, _013893_, _013896_);
  xor g_106524_(_001516_, _013886_, _013897_);
  xor g_106525_(_001515_, _013886_, _013898_);
  xor g_106526_(_013889_, _013893_, _013899_);
  xor g_106527_(_013888_, _013893_, _013900_);
  and g_106528_(_013897_, _013899_, _013901_);
  or g_106529_(_013898_, _013900_, _013902_);
  or g_106530_(_001209_, _013876_, _013904_);
  or g_106531_(_013821_, _013875_, _013905_);
  and g_106532_(_013904_, _013905_, _013906_);
  and g_106533_(out[833], _013906_, _013907_);
  not g_106534_(_013907_, _013908_);
  and g_106535_(_013825_, _013876_, _013909_);
  not g_106536_(_013909_, _013910_);
  or g_106537_(out[816], _013876_, _013911_);
  not g_106538_(_013911_, _013912_);
  or g_106539_(_013909_, _013912_, _013913_);
  and g_106540_(_013910_, _013911_, _013915_);
  and g_106541_(out[832], _013913_, _013916_);
  or g_106542_(_001352_, _013915_, _013917_);
  xor g_106543_(out[833], _013906_, _013918_);
  xor g_106544_(_001341_, _013906_, _013919_);
  and g_106545_(_013917_, _013918_, _013920_);
  or g_106546_(_013916_, _013919_, _013921_);
  and g_106547_(_013908_, _013921_, _013922_);
  or g_106548_(_013907_, _013920_, _013923_);
  and g_106549_(_013901_, _013923_, _013924_);
  or g_106550_(_013902_, _013922_, _013926_);
  or g_106551_(_013895_, _013896_, _013927_);
  not g_106552_(_013927_, _013928_);
  and g_106553_(_013926_, _013927_, _013929_);
  or g_106554_(_013924_, _013928_, _013930_);
  and g_106555_(_009754_, _009769_, _013931_);
  or g_106556_(_009755_, _009768_, _013932_);
  xor g_106557_(out[842], _009765_, _013933_);
  not g_106558_(_013933_, _013934_);
  and g_106559_(_013882_, _013933_, _013935_);
  or g_106560_(_013883_, _013934_, _013937_);
  and g_106561_(_013932_, _013937_, _013938_);
  or g_106562_(_013931_, _013935_, _013939_);
  and g_106563_(_009755_, _009768_, _013940_);
  or g_106564_(_009754_, _009769_, _013941_);
  and g_106565_(_013883_, _013934_, _013942_);
  or g_106566_(_013882_, _013933_, _013943_);
  and g_106567_(_013941_, _013943_, _013944_);
  or g_106568_(_013940_, _013942_, _013945_);
  and g_106569_(_013938_, _013944_, _013946_);
  or g_106570_(_013939_, _013945_, _013948_);
  xor g_106571_(out[840], _009763_, _013949_);
  xor g_106572_(_001385_, _009763_, _013950_);
  and g_106573_(_013718_, _013875_, _013951_);
  and g_106574_(_013724_, _013876_, _013952_);
  or g_106575_(_013951_, _013952_, _013953_);
  or g_106576_(_013949_, _013953_, _013954_);
  not g_106577_(_013954_, _013955_);
  and g_106578_(out[841], _009764_, _013956_);
  xor g_106579_(out[841], _009764_, _013957_);
  xor g_106580_(_001396_, _009764_, _013959_);
  and g_106581_(_013707_, _013876_, _013960_);
  or g_106582_(_013706_, _013875_, _013961_);
  and g_106583_(_013700_, _013875_, _013962_);
  or g_106584_(_013699_, _013876_, _013963_);
  and g_106585_(_013961_, _013963_, _013964_);
  or g_106586_(_013960_, _013962_, _013965_);
  and g_106587_(_013957_, _013965_, _013966_);
  or g_106588_(_013959_, _013964_, _013967_);
  or g_106589_(_013955_, _013966_, _013968_);
  and g_106590_(_013949_, _013953_, _013970_);
  and g_106591_(_013959_, _013964_, _013971_);
  or g_106592_(_013957_, _013965_, _013972_);
  or g_106593_(_013970_, _013971_, _013973_);
  or g_106594_(_013968_, _013973_, _013974_);
  xor g_106595_(_013949_, _013953_, _013975_);
  and g_106596_(_013967_, _013972_, _013976_);
  and g_106597_(_013946_, _013976_, _013977_);
  and g_106598_(_013975_, _013977_, _013978_);
  or g_106599_(_013948_, _013974_, _013979_);
  xor g_106600_(out[839], _009762_, _013981_);
  xor g_106601_(_001297_, _009762_, _013982_);
  and g_106602_(_013739_, _013875_, _013983_);
  or g_106603_(_013740_, _013876_, _013984_);
  and g_106604_(_013746_, _013876_, _013985_);
  or g_106605_(_013745_, _013875_, _013986_);
  and g_106606_(_013984_, _013986_, _013987_);
  or g_106607_(_013983_, _013985_, _013988_);
  and g_106608_(_013981_, _013987_, _013989_);
  or g_106609_(_013982_, _013988_, _013990_);
  xor g_106610_(out[838], _009761_, _013992_);
  not g_106611_(_013992_, _013993_);
  and g_106612_(_013751_, _013875_, _013994_);
  and g_106613_(_013754_, _013876_, _013995_);
  or g_106614_(_013994_, _013995_, _013996_);
  or g_106615_(_013992_, _013996_, _013997_);
  not g_106616_(_013997_, _013998_);
  and g_106617_(_013982_, _013988_, _013999_);
  or g_106618_(_013981_, _013987_, _014000_);
  and g_106619_(_013990_, _014000_, _014001_);
  or g_106620_(_013989_, _013999_, _014003_);
  xor g_106621_(_013992_, _013996_, _014004_);
  xor g_106622_(_013993_, _013996_, _014005_);
  and g_106623_(_014001_, _014004_, _014006_);
  or g_106624_(_014003_, _014005_, _014007_);
  or g_106625_(_024914_, _001514_, _014008_);
  not g_106626_(_014008_, _014009_);
  and g_106627_(_009760_, _014008_, _014010_);
  or g_106628_(_009759_, _014009_, _014011_);
  and g_106629_(_013776_, _013876_, _014012_);
  not g_106630_(_014012_, _014014_);
  or g_106631_(_013768_, _013876_, _014015_);
  not g_106632_(_014015_, _014016_);
  and g_106633_(_014014_, _014015_, _014017_);
  or g_106634_(_014012_, _014016_, _014018_);
  and g_106635_(_014011_, _014017_, _014019_);
  or g_106636_(_014010_, _014018_, _014020_);
  xor g_106637_(out[837], _009759_, _014021_);
  xor g_106638_(_001319_, _009759_, _014022_);
  or g_106639_(_013779_, _013876_, _014023_);
  not g_106640_(_014023_, _014025_);
  and g_106641_(_013787_, _013876_, _014026_);
  not g_106642_(_014026_, _014027_);
  and g_106643_(_014023_, _014027_, _014028_);
  or g_106644_(_014025_, _014026_, _014029_);
  and g_106645_(_014022_, _014028_, _014030_);
  or g_106646_(_014021_, _014029_, _014031_);
  and g_106647_(_014020_, _014031_, _014032_);
  or g_106648_(_014019_, _014030_, _014033_);
  and g_106649_(_014021_, _014029_, _014034_);
  or g_106650_(_014022_, _014028_, _014036_);
  and g_106651_(_014010_, _014018_, _014037_);
  or g_106652_(_014011_, _014017_, _014038_);
  and g_106653_(_014036_, _014038_, _014039_);
  or g_106654_(_014034_, _014037_, _014040_);
  and g_106655_(_014032_, _014039_, _014041_);
  or g_106656_(_014033_, _014040_, _014042_);
  and g_106657_(_014006_, _014041_, _014043_);
  or g_106658_(_014007_, _014042_, _014044_);
  and g_106659_(_013978_, _014043_, _014045_);
  or g_106660_(_013979_, _014044_, _014047_);
  and g_106661_(_013930_, _014045_, _014048_);
  or g_106662_(_013929_, _014047_, _014049_);
  and g_106663_(_014006_, _014033_, _014050_);
  or g_106664_(_014007_, _014032_, _014051_);
  and g_106665_(_014036_, _014050_, _014052_);
  or g_106666_(_014034_, _014051_, _014053_);
  and g_106667_(_013998_, _014000_, _014054_);
  or g_106668_(_013997_, _013999_, _014055_);
  and g_106669_(_013990_, _014055_, _014056_);
  or g_106670_(_013989_, _014054_, _014058_);
  and g_106671_(_014053_, _014056_, _014059_);
  or g_106672_(_014052_, _014058_, _014060_);
  and g_106673_(_013978_, _014060_, _014061_);
  or g_106674_(_013979_, _014059_, _014062_);
  or g_106675_(_013954_, _013971_, _014063_);
  and g_106676_(_013967_, _014063_, _014064_);
  and g_106677_(_013939_, _013941_, _014065_);
  or g_106678_(_013938_, _013940_, _014066_);
  and g_106679_(_013946_, _013968_, _014067_);
  and g_106680_(_013972_, _014067_, _014069_);
  or g_106681_(_013948_, _014064_, _014070_);
  or g_106682_(_014065_, _014069_, _014071_);
  and g_106683_(_014066_, _014070_, _014072_);
  and g_106684_(_014062_, _014072_, _014073_);
  or g_106685_(_014061_, _014071_, _014074_);
  and g_106686_(_014049_, _014073_, _014075_);
  or g_106687_(_014048_, _014074_, _014076_);
  or g_106688_(out[832], _013913_, _014077_);
  not g_106689_(_014077_, _014078_);
  and g_106690_(_013901_, _014077_, _014080_);
  or g_106691_(_013902_, _014078_, _014081_);
  and g_106692_(_013920_, _014080_, _014082_);
  or g_106693_(_013921_, _014081_, _014083_);
  and g_106694_(_014045_, _014082_, _014084_);
  or g_106695_(_014047_, _014083_, _014085_);
  and g_106696_(_014076_, _014085_, _014086_);
  or g_106697_(_014075_, _014084_, _014087_);
  and g_106698_(_013883_, _014087_, _014088_);
  or g_106699_(_013882_, _014086_, _014089_);
  and g_106700_(_013933_, _014086_, _014091_);
  or g_106701_(_013934_, _014087_, _014092_);
  and g_106702_(_014089_, _014092_, _014093_);
  or g_106703_(_014088_, _014091_, _014094_);
  and g_106704_(_009771_, _009784_, _014095_);
  or g_106705_(_009770_, _009785_, _014096_);
  xor g_106706_(out[858], _009781_, _014097_);
  xor g_106707_(_001539_, _009781_, _014098_);
  and g_106708_(_014093_, _014097_, _014099_);
  or g_106709_(_014094_, _014098_, _014100_);
  and g_106710_(_009770_, _009785_, _014102_);
  or g_106711_(_009771_, _009784_, _014103_);
  and g_106712_(_014100_, _014103_, _014104_);
  or g_106713_(_014099_, _014102_, _014105_);
  and g_106714_(out[857], _009780_, _014106_);
  xor g_106715_(out[857], _009780_, _014107_);
  or g_106716_(_009782_, _014106_, _014108_);
  and g_106717_(_013965_, _014087_, _014109_);
  not g_106718_(_014109_, _014110_);
  or g_106719_(_013957_, _014087_, _014111_);
  not g_106720_(_014111_, _014113_);
  and g_106721_(_014110_, _014111_, _014114_);
  or g_106722_(_014109_, _014113_, _014115_);
  and g_106723_(_014107_, _014115_, _014116_);
  xor g_106724_(out[856], _009779_, _014117_);
  xor g_106725_(_001517_, _009779_, _014118_);
  or g_106726_(_013949_, _014087_, _014119_);
  not g_106727_(_014119_, _014120_);
  and g_106728_(_013953_, _014087_, _014121_);
  not g_106729_(_014121_, _014122_);
  and g_106730_(_014119_, _014122_, _014124_);
  or g_106731_(_014120_, _014121_, _014125_);
  and g_106732_(_014118_, _014124_, _014126_);
  or g_106733_(_014116_, _014126_, _014127_);
  and g_106734_(_014094_, _014098_, _014128_);
  or g_106735_(_014093_, _014097_, _014129_);
  and g_106736_(_014108_, _014114_, _014130_);
  or g_106737_(_014107_, _014115_, _014131_);
  and g_106738_(_014117_, _014125_, _014132_);
  xor g_106739_(_014108_, _014114_, _014133_);
  and g_106740_(_014096_, _014129_, _014135_);
  or g_106741_(_014095_, _014128_, _014136_);
  and g_106742_(_014104_, _014135_, _014137_);
  or g_106743_(_014105_, _014136_, _014138_);
  xor g_106744_(_014118_, _014124_, _014139_);
  and g_106745_(_014137_, _014139_, _014140_);
  or g_106746_(_014116_, _014132_, _014141_);
  or g_106747_(_014126_, _014130_, _014142_);
  or g_106748_(_014141_, _014142_, _014143_);
  and g_106749_(_014133_, _014140_, _014144_);
  or g_106750_(_014138_, _014143_, _014146_);
  xor g_106751_(out[855], _009777_, _014147_);
  xor g_106752_(_001429_, _009777_, _014148_);
  and g_106753_(_013981_, _014086_, _014149_);
  and g_106754_(_013988_, _014087_, _014150_);
  or g_106755_(_014149_, _014150_, _014151_);
  or g_106756_(_014148_, _014151_, _014152_);
  xor g_106757_(out[854], _009776_, _014153_);
  not g_106758_(_014153_, _014154_);
  and g_106759_(_013996_, _014087_, _014155_);
  and g_106760_(_013993_, _014086_, _014157_);
  or g_106761_(_014155_, _014157_, _014158_);
  or g_106762_(_014153_, _014158_, _014159_);
  and g_106763_(_014148_, _014151_, _014160_);
  xor g_106764_(_014148_, _014151_, _014161_);
  xor g_106765_(_014147_, _014151_, _014162_);
  xor g_106766_(_014153_, _014158_, _014163_);
  xor g_106767_(_014154_, _014158_, _014164_);
  and g_106768_(_014161_, _014163_, _014165_);
  or g_106769_(_014162_, _014164_, _014166_);
  xor g_106770_(out[853], _009774_, _014168_);
  xor g_106771_(_001451_, _009774_, _014169_);
  or g_106772_(_014021_, _014087_, _014170_);
  not g_106773_(_014170_, _014171_);
  and g_106774_(_014029_, _014087_, _014172_);
  not g_106775_(_014172_, _014173_);
  and g_106776_(_014170_, _014173_, _014174_);
  or g_106777_(_014171_, _014172_, _014175_);
  and g_106778_(_014168_, _014175_, _014176_);
  or g_106779_(_014169_, _014174_, _014177_);
  or g_106780_(_025068_, _001844_, _014179_);
  not g_106781_(_014179_, _014180_);
  and g_106782_(_009775_, _014179_, _014181_);
  or g_106783_(_009774_, _014180_, _014182_);
  and g_106784_(_014018_, _014087_, _014183_);
  not g_106785_(_014183_, _014184_);
  or g_106786_(_014010_, _014087_, _014185_);
  not g_106787_(_014185_, _014186_);
  and g_106788_(_014184_, _014185_, _014187_);
  or g_106789_(_014183_, _014186_, _014188_);
  and g_106790_(_014182_, _014187_, _014190_);
  or g_106791_(_014181_, _014188_, _014191_);
  and g_106792_(_014169_, _014174_, _014192_);
  or g_106793_(_014168_, _014175_, _014193_);
  and g_106794_(_014191_, _014193_, _014194_);
  or g_106795_(_014190_, _014192_, _014195_);
  and g_106796_(_014165_, _014195_, _014196_);
  or g_106797_(_014166_, _014194_, _014197_);
  and g_106798_(_014177_, _014196_, _014198_);
  or g_106799_(_014176_, _014197_, _014199_);
  or g_106800_(_014159_, _014160_, _014201_);
  and g_106801_(_014152_, _014201_, _014202_);
  not g_106802_(_014202_, _014203_);
  and g_106803_(_014199_, _014202_, _014204_);
  or g_106804_(_014198_, _014203_, _014205_);
  xor g_106805_(out[851], _001844_, _014206_);
  xor g_106806_(_001506_, _001844_, _014207_);
  and g_106807_(_013888_, _014086_, _014208_);
  and g_106808_(_013893_, _014087_, _014209_);
  or g_106809_(_014208_, _014209_, _014210_);
  not g_106810_(_014210_, _014212_);
  or g_106811_(_014207_, _014210_, _014213_);
  and g_106812_(_014207_, _014210_, _014214_);
  or g_106813_(_014206_, _014212_, _014215_);
  and g_106814_(_013886_, _014087_, _014216_);
  and g_106815_(_001515_, _014086_, _014217_);
  or g_106816_(_014216_, _014217_, _014218_);
  or g_106817_(_001846_, _014218_, _014219_);
  or g_106818_(_014214_, _014219_, _014220_);
  and g_106819_(_014213_, _014220_, _014221_);
  not g_106820_(_014221_, _014223_);
  or g_106821_(_001341_, _014087_, _014224_);
  or g_106822_(_013906_, _014086_, _014225_);
  and g_106823_(_014224_, _014225_, _014226_);
  and g_106824_(out[849], _014226_, _014227_);
  not g_106825_(_014227_, _014228_);
  or g_106826_(_001352_, _014087_, _014229_);
  not g_106827_(_014229_, _014230_);
  and g_106828_(_013915_, _014087_, _014231_);
  or g_106829_(_013913_, _014086_, _014232_);
  and g_106830_(_014229_, _014232_, _014234_);
  or g_106831_(_014230_, _014231_, _014235_);
  and g_106832_(out[848], _014234_, _014236_);
  or g_106833_(_001484_, _014235_, _014237_);
  xor g_106834_(out[849], _014226_, _014238_);
  xor g_106835_(_001473_, _014226_, _014239_);
  and g_106836_(_014237_, _014238_, _014240_);
  or g_106837_(_014236_, _014239_, _014241_);
  and g_106838_(_014228_, _014241_, _014242_);
  or g_106839_(_014227_, _014240_, _014243_);
  xor g_106840_(_001846_, _014218_, _014245_);
  xor g_106841_(_001845_, _014218_, _014246_);
  and g_106842_(_014215_, _014245_, _014247_);
  or g_106843_(_014214_, _014246_, _014248_);
  and g_106844_(_014243_, _014247_, _014249_);
  or g_106845_(_014242_, _014248_, _014250_);
  and g_106846_(_014221_, _014250_, _014251_);
  or g_106847_(_014223_, _014249_, _014252_);
  and g_106848_(_014181_, _014188_, _014253_);
  or g_106849_(_014182_, _014187_, _014254_);
  and g_106850_(_014177_, _014254_, _014256_);
  or g_106851_(_014176_, _014253_, _014257_);
  and g_106852_(_014194_, _014256_, _014258_);
  or g_106853_(_014195_, _014257_, _014259_);
  and g_106854_(_014165_, _014258_, _014260_);
  or g_106855_(_014166_, _014259_, _014261_);
  and g_106856_(_014144_, _014260_, _014262_);
  or g_106857_(_014146_, _014261_, _014263_);
  and g_106858_(_014252_, _014262_, _014264_);
  or g_106859_(_014251_, _014263_, _014265_);
  and g_106860_(_014127_, _014131_, _014267_);
  not g_106861_(_014267_, _014268_);
  and g_106862_(_014137_, _014267_, _014269_);
  or g_106863_(_014138_, _014268_, _014270_);
  and g_106864_(_014265_, _014270_, _014271_);
  or g_106865_(_014264_, _014269_, _014272_);
  and g_106866_(_014096_, _014105_, _014273_);
  or g_106867_(_014095_, _014104_, _014274_);
  and g_106868_(_014144_, _014205_, _014275_);
  or g_106869_(_014146_, _014204_, _014276_);
  and g_106870_(_014274_, _014276_, _014278_);
  or g_106871_(_014273_, _014275_, _014279_);
  and g_106872_(_014271_, _014278_, _014280_);
  or g_106873_(_014272_, _014279_, _014281_);
  or g_106874_(out[848], _014234_, _014282_);
  and g_106875_(_014213_, _014282_, _014283_);
  and g_106876_(_014247_, _014283_, _014284_);
  not g_106877_(_014284_, _014285_);
  or g_106878_(_014263_, _014285_, _014286_);
  or g_106879_(_014241_, _014286_, _014287_);
  not g_106880_(_014287_, _014289_);
  and g_106881_(_014281_, _014287_, _014290_);
  or g_106882_(_014280_, _014289_, _014291_);
  and g_106883_(_014094_, _014291_, _014292_);
  or g_106884_(_014093_, _014290_, _014293_);
  and g_106885_(_014097_, _014290_, _014294_);
  or g_106886_(_014098_, _014291_, _014295_);
  and g_106887_(_014293_, _014295_, _014296_);
  or g_106888_(_014292_, _014294_, _014297_);
  xor g_106889_(out[874], _009797_, _014298_);
  xor g_106890_(_001671_, _009797_, _014300_);
  and g_106891_(_014296_, _014298_, _014301_);
  or g_106892_(_014297_, _014300_, _014302_);
  and g_106893_(_009786_, _009802_, _014303_);
  or g_106894_(_009787_, _009801_, _014304_);
  and g_106895_(_014302_, _014304_, _014305_);
  or g_106896_(_014301_, _014303_, _014306_);
  and g_106897_(_009787_, _009801_, _014307_);
  and g_106898_(_014297_, _014300_, _014308_);
  or g_106899_(_014307_, _014308_, _014309_);
  not g_106900_(_014309_, _014311_);
  and g_106901_(_014305_, _014311_, _014312_);
  or g_106902_(_014306_, _014309_, _014313_);
  and g_106903_(out[873], _009796_, _014314_);
  xor g_106904_(out[873], _009796_, _014315_);
  or g_106905_(_009798_, _014314_, _014316_);
  and g_106906_(_014115_, _014291_, _014317_);
  and g_106907_(_014108_, _014290_, _014318_);
  or g_106908_(_014317_, _014318_, _014319_);
  or g_106909_(_014315_, _014319_, _014320_);
  xor g_106910_(out[872], _009795_, _014322_);
  xor g_106911_(_001649_, _009795_, _014323_);
  and g_106912_(_014118_, _014290_, _014324_);
  and g_106913_(_014125_, _014291_, _014325_);
  or g_106914_(_014324_, _014325_, _014326_);
  or g_106915_(_014322_, _014326_, _014327_);
  not g_106916_(_014327_, _014328_);
  and g_106917_(_014315_, _014319_, _014329_);
  xor g_106918_(_014315_, _014319_, _014330_);
  xor g_106919_(_014316_, _014319_, _014331_);
  xor g_106920_(_014322_, _014326_, _014333_);
  xor g_106921_(_014323_, _014326_, _014334_);
  and g_106922_(_014312_, _014333_, _014335_);
  or g_106923_(_014313_, _014334_, _014336_);
  and g_106924_(_014330_, _014335_, _014337_);
  or g_106925_(_014331_, _014336_, _014338_);
  xor g_106926_(out[871], _009794_, _014339_);
  xor g_106927_(_001561_, _009794_, _014340_);
  or g_106928_(_014148_, _014291_, _014341_);
  not g_106929_(_014341_, _014342_);
  and g_106930_(_014151_, _014291_, _014344_);
  not g_106931_(_014344_, _014345_);
  and g_106932_(_014341_, _014345_, _014346_);
  or g_106933_(_014342_, _014344_, _014347_);
  and g_106934_(_014339_, _014346_, _014348_);
  or g_106935_(_014339_, _014346_, _014349_);
  xor g_106936_(_014339_, _014346_, _014350_);
  xor g_106937_(_014340_, _014346_, _014351_);
  xor g_106938_(out[870], _009793_, _014352_);
  xor g_106939_(_001572_, _009793_, _014353_);
  or g_106940_(_014153_, _014291_, _014355_);
  and g_106941_(_014158_, _014291_, _014356_);
  not g_106942_(_014356_, _014357_);
  and g_106943_(_014355_, _014357_, _014358_);
  and g_106944_(_014353_, _014358_, _014359_);
  xor g_106945_(_014353_, _014358_, _014360_);
  xor g_106946_(_014352_, _014358_, _014361_);
  and g_106947_(_014350_, _014360_, _014362_);
  or g_106948_(_014351_, _014361_, _014363_);
  or g_106949_(_025222_, _002016_, _014364_);
  not g_106950_(_014364_, _014366_);
  and g_106951_(_009792_, _014364_, _014367_);
  or g_106952_(_009791_, _014366_, _014368_);
  and g_106953_(_014188_, _014291_, _014369_);
  and g_106954_(_014182_, _014290_, _014370_);
  or g_106955_(_014369_, _014370_, _014371_);
  or g_106956_(_014367_, _014371_, _014372_);
  not g_106957_(_014372_, _014373_);
  xor g_106958_(out[869], _009791_, _014374_);
  xor g_106959_(_001583_, _009791_, _014375_);
  and g_106960_(_014169_, _014290_, _014377_);
  and g_106961_(_014175_, _014291_, _014378_);
  or g_106962_(_014377_, _014378_, _014379_);
  or g_106963_(_014374_, _014379_, _014380_);
  not g_106964_(_014380_, _014381_);
  and g_106965_(_014372_, _014380_, _014382_);
  or g_106966_(_014373_, _014381_, _014383_);
  and g_106967_(_014374_, _014379_, _014384_);
  and g_106968_(_014367_, _014371_, _014385_);
  or g_106969_(_014384_, _014385_, _014386_);
  not g_106970_(_014386_, _014388_);
  and g_106971_(_014382_, _014388_, _014389_);
  or g_106972_(_014383_, _014386_, _014390_);
  and g_106973_(_014362_, _014389_, _014391_);
  or g_106974_(_014363_, _014390_, _014392_);
  and g_106975_(_014337_, _014391_, _014393_);
  or g_106976_(_014338_, _014392_, _014394_);
  and g_106977_(_014218_, _014291_, _014395_);
  and g_106978_(_001845_, _014290_, _014396_);
  or g_106979_(_014395_, _014396_, _014397_);
  xor g_106980_(out[867], _002016_, _014399_);
  xor g_106981_(_001638_, _002016_, _014400_);
  and g_106982_(_014210_, _014291_, _014401_);
  and g_106983_(_014206_, _014290_, _014402_);
  or g_106984_(_014401_, _014402_, _014403_);
  or g_106985_(_014400_, _014403_, _014404_);
  or g_106986_(_002017_, _014397_, _014405_);
  and g_106987_(_014400_, _014403_, _014406_);
  xor g_106988_(_002017_, _014397_, _014407_);
  xor g_106989_(_014400_, _014403_, _014408_);
  and g_106990_(_014407_, _014408_, _014410_);
  or g_106991_(_001473_, _014291_, _014411_);
  or g_106992_(_014226_, _014290_, _014412_);
  and g_106993_(_014411_, _014412_, _014413_);
  and g_106994_(out[865], _014413_, _014414_);
  or g_106995_(_001484_, _014291_, _014415_);
  or g_106996_(_014234_, _014290_, _014416_);
  and g_106997_(_014415_, _014416_, _014417_);
  and g_106998_(out[864], _014417_, _014418_);
  not g_106999_(_014418_, _014419_);
  xor g_107000_(out[865], _014413_, _014421_);
  and g_107001_(_014419_, _014421_, _014422_);
  or g_107002_(_014414_, _014422_, _014423_);
  and g_107003_(_014410_, _014423_, _014424_);
  not g_107004_(_014424_, _014425_);
  or g_107005_(_014405_, _014406_, _014426_);
  and g_107006_(_014404_, _014426_, _014427_);
  not g_107007_(_014427_, _014428_);
  and g_107008_(_014425_, _014427_, _014429_);
  or g_107009_(_014424_, _014428_, _014430_);
  and g_107010_(_014393_, _014430_, _014432_);
  or g_107011_(_014394_, _014429_, _014433_);
  or g_107012_(_014382_, _014384_, _014434_);
  or g_107013_(_014363_, _014434_, _014435_);
  not g_107014_(_014435_, _014436_);
  and g_107015_(_014349_, _014359_, _014437_);
  or g_107016_(_014348_, _014437_, _014438_);
  or g_107017_(_014436_, _014438_, _014439_);
  and g_107018_(_014337_, _014439_, _014440_);
  not g_107019_(_014440_, _014441_);
  or g_107020_(_014305_, _014307_, _014443_);
  not g_107021_(_014443_, _014444_);
  or g_107022_(_014328_, _014329_, _014445_);
  and g_107023_(_014320_, _014445_, _014446_);
  and g_107024_(_014312_, _014446_, _014447_);
  not g_107025_(_014447_, _014448_);
  and g_107026_(_014443_, _014448_, _014449_);
  or g_107027_(_014444_, _014447_, _014450_);
  and g_107028_(_014433_, _014449_, _014451_);
  or g_107029_(_014432_, _014450_, _014452_);
  and g_107030_(_014441_, _014451_, _014454_);
  or g_107031_(_014440_, _014452_, _014455_);
  or g_107032_(out[864], _014417_, _014456_);
  and g_107033_(_014410_, _014456_, _014457_);
  and g_107034_(_014422_, _014457_, _014458_);
  and g_107035_(_014393_, _014458_, _014459_);
  not g_107036_(_014459_, _014460_);
  and g_107037_(_014455_, _014460_, _014461_);
  or g_107038_(_014454_, _014459_, _014462_);
  and g_107039_(_014297_, _014462_, _014463_);
  not g_107040_(_014463_, _014465_);
  or g_107041_(_014300_, _014462_, _014466_);
  not g_107042_(_014466_, _014467_);
  and g_107043_(_014465_, _014466_, _014468_);
  or g_107044_(_014463_, _014467_, _014469_);
  xor g_107045_(out[890], _009814_, _014470_);
  xor g_107046_(_001803_, _009814_, _014471_);
  and g_107047_(_014468_, _014470_, _014472_);
  or g_107048_(_014469_, _014471_, _014473_);
  and g_107049_(_009803_, _009818_, _014474_);
  or g_107050_(_009804_, _009817_, _014476_);
  and g_107051_(_014473_, _014476_, _014477_);
  or g_107052_(_014472_, _014474_, _014478_);
  and g_107053_(_014469_, _014471_, _014479_);
  or g_107054_(_014468_, _014470_, _014480_);
  and g_107055_(_009804_, _009817_, _014481_);
  or g_107056_(_009803_, _009818_, _014482_);
  and g_107057_(out[889], _009813_, _014483_);
  xor g_107058_(out[889], _009813_, _014484_);
  or g_107059_(_009815_, _014483_, _014485_);
  and g_107060_(_014319_, _014462_, _014487_);
  not g_107061_(_014487_, _014488_);
  or g_107062_(_014315_, _014462_, _014489_);
  not g_107063_(_014489_, _014490_);
  and g_107064_(_014488_, _014489_, _014491_);
  or g_107065_(_014487_, _014490_, _014492_);
  and g_107066_(_014485_, _014491_, _014493_);
  or g_107067_(_014484_, _014492_, _014494_);
  and g_107068_(_014482_, _014494_, _014495_);
  or g_107069_(_014481_, _014493_, _014496_);
  and g_107070_(_014480_, _014495_, _014498_);
  or g_107071_(_014479_, _014496_, _014499_);
  and g_107072_(_014477_, _014498_, _014500_);
  or g_107073_(_014478_, _014499_, _014501_);
  xor g_107074_(out[888], _009812_, _014502_);
  xor g_107075_(_001781_, _009812_, _014503_);
  or g_107076_(_014322_, _014462_, _014504_);
  not g_107077_(_014504_, _014505_);
  and g_107078_(_014326_, _014462_, _014506_);
  not g_107079_(_014506_, _014507_);
  and g_107080_(_014504_, _014507_, _014509_);
  or g_107081_(_014505_, _014506_, _014510_);
  and g_107082_(_014502_, _014510_, _014511_);
  or g_107083_(_014503_, _014509_, _014512_);
  and g_107084_(_014484_, _014492_, _014513_);
  or g_107085_(_014485_, _014491_, _014514_);
  and g_107086_(_014503_, _014509_, _014515_);
  or g_107087_(_014502_, _014510_, _014516_);
  and g_107088_(_014514_, _014516_, _014517_);
  or g_107089_(_014513_, _014515_, _014518_);
  and g_107090_(_014512_, _014517_, _014520_);
  or g_107091_(_014511_, _014518_, _014521_);
  and g_107092_(_014500_, _014520_, _014522_);
  or g_107093_(_014501_, _014521_, _014523_);
  xor g_107094_(out[886], _009809_, _014524_);
  xor g_107095_(_001704_, _009809_, _014525_);
  or g_107096_(_014352_, _014462_, _014526_);
  or g_107097_(_014358_, _014461_, _014527_);
  and g_107098_(_014526_, _014527_, _014528_);
  not g_107099_(_014528_, _014529_);
  and g_107100_(_014525_, _014528_, _014531_);
  or g_107101_(_014524_, _014529_, _014532_);
  xor g_107102_(out[887], _009810_, _014533_);
  xor g_107103_(_001693_, _009810_, _014534_);
  and g_107104_(_014339_, _014461_, _014535_);
  or g_107105_(_014340_, _014462_, _014536_);
  and g_107106_(_014347_, _014462_, _014537_);
  or g_107107_(_014346_, _014461_, _014538_);
  and g_107108_(_014536_, _014538_, _014539_);
  or g_107109_(_014535_, _014537_, _014540_);
  and g_107110_(_014534_, _014540_, _014542_);
  or g_107111_(_014533_, _014539_, _014543_);
  and g_107112_(_014533_, _014539_, _014544_);
  or g_107113_(_014534_, _014540_, _014545_);
  xor g_107114_(_014525_, _014528_, _014546_);
  xor g_107115_(_014524_, _014528_, _014547_);
  and g_107116_(_014545_, _014546_, _014548_);
  or g_107117_(_014544_, _014547_, _014549_);
  and g_107118_(_014543_, _014548_, _014550_);
  or g_107119_(_014542_, _014549_, _014551_);
  or g_107120_(_025376_, _002075_, _014553_);
  not g_107121_(_014553_, _014554_);
  and g_107122_(_009808_, _014553_, _014555_);
  or g_107123_(_009807_, _014554_, _014556_);
  and g_107124_(_014371_, _014462_, _014557_);
  not g_107125_(_014557_, _014558_);
  or g_107126_(_014367_, _014462_, _014559_);
  not g_107127_(_014559_, _014560_);
  and g_107128_(_014558_, _014559_, _014561_);
  or g_107129_(_014557_, _014560_, _014562_);
  and g_107130_(_014556_, _014561_, _014564_);
  or g_107131_(_014555_, _014562_, _014565_);
  xor g_107132_(out[885], _009807_, _014566_);
  xor g_107133_(_001715_, _009807_, _014567_);
  or g_107134_(_014374_, _014462_, _014568_);
  not g_107135_(_014568_, _014569_);
  and g_107136_(_014379_, _014462_, _014570_);
  not g_107137_(_014570_, _014571_);
  and g_107138_(_014568_, _014571_, _014572_);
  or g_107139_(_014569_, _014570_, _014573_);
  and g_107140_(_014567_, _014572_, _014575_);
  or g_107141_(_014566_, _014573_, _014576_);
  and g_107142_(_014565_, _014576_, _014577_);
  or g_107143_(_014564_, _014575_, _014578_);
  and g_107144_(_014566_, _014573_, _014579_);
  or g_107145_(_014567_, _014572_, _014580_);
  and g_107146_(_014555_, _014562_, _014581_);
  or g_107147_(_014556_, _014561_, _014582_);
  and g_107148_(_014580_, _014582_, _014583_);
  or g_107149_(_014579_, _014581_, _014584_);
  and g_107150_(_014577_, _014583_, _014586_);
  or g_107151_(_014578_, _014584_, _014587_);
  and g_107152_(_014550_, _014586_, _014588_);
  or g_107153_(_014551_, _014587_, _014589_);
  and g_107154_(_014522_, _014588_, _014590_);
  or g_107155_(_014523_, _014589_, _014591_);
  or g_107156_(_001605_, _014462_, _014592_);
  or g_107157_(_014413_, _014461_, _014593_);
  and g_107158_(_014592_, _014593_, _014594_);
  or g_107159_(_001616_, _014462_, _014595_);
  or g_107160_(_014417_, _014461_, _014597_);
  and g_107161_(_014595_, _014597_, _014598_);
  and g_107162_(out[880], _014598_, _014599_);
  not g_107163_(_014599_, _014600_);
  and g_107164_(out[881], _014594_, _014601_);
  xor g_107165_(out[881], _014594_, _014602_);
  xor g_107166_(_001737_, _014594_, _014603_);
  and g_107167_(_014600_, _014602_, _014604_);
  or g_107168_(_014599_, _014603_, _014605_);
  or g_107169_(_002017_, _014462_, _014606_);
  not g_107170_(_014606_, _014608_);
  and g_107171_(_014397_, _014462_, _014609_);
  not g_107172_(_014609_, _014610_);
  and g_107173_(_014606_, _014610_, _014611_);
  or g_107174_(_014608_, _014609_, _014612_);
  and g_107175_(_002076_, _014611_, _014613_);
  or g_107176_(_002077_, _014612_, _014614_);
  xor g_107177_(out[883], _002075_, _014615_);
  xor g_107178_(_001770_, _002075_, _014616_);
  or g_107179_(_014400_, _014462_, _014617_);
  not g_107180_(_014617_, _014619_);
  and g_107181_(_014403_, _014462_, _014620_);
  not g_107182_(_014620_, _014621_);
  and g_107183_(_014617_, _014621_, _014622_);
  or g_107184_(_014619_, _014620_, _014623_);
  and g_107185_(_014616_, _014623_, _014624_);
  or g_107186_(_014615_, _014622_, _014625_);
  xor g_107187_(_002076_, _014611_, _014626_);
  xor g_107188_(_002077_, _014611_, _014627_);
  and g_107189_(_014625_, _014626_, _014628_);
  or g_107190_(_014624_, _014627_, _014630_);
  and g_107191_(_014615_, _014622_, _014631_);
  or g_107192_(_014616_, _014623_, _014632_);
  or g_107193_(out[880], _014598_, _014633_);
  not g_107194_(_014633_, _014634_);
  and g_107195_(_014632_, _014633_, _014635_);
  or g_107196_(_014631_, _014634_, _014636_);
  and g_107197_(_014628_, _014635_, _014637_);
  or g_107198_(_014630_, _014636_, _014638_);
  and g_107199_(_014604_, _014637_, _014639_);
  or g_107200_(_014605_, _014638_, _014641_);
  and g_107201_(_014590_, _014639_, _014642_);
  or g_107202_(_014591_, _014641_, _014643_);
  and g_107203_(_014613_, _014625_, _014644_);
  or g_107204_(_014614_, _014624_, _014645_);
  and g_107205_(_014632_, _014645_, _014646_);
  or g_107206_(_014631_, _014644_, _014647_);
  or g_107207_(_014601_, _014604_, _014648_);
  and g_107208_(_014628_, _014648_, _014649_);
  not g_107209_(_014649_, _014650_);
  and g_107210_(_014646_, _014650_, _014652_);
  or g_107211_(_014647_, _014649_, _014653_);
  and g_107212_(_014590_, _014653_, _014654_);
  or g_107213_(_014591_, _014652_, _014655_);
  and g_107214_(_014550_, _014578_, _014656_);
  or g_107215_(_014551_, _014577_, _014657_);
  and g_107216_(_014580_, _014656_, _014658_);
  or g_107217_(_014579_, _014657_, _014659_);
  and g_107218_(_014531_, _014543_, _014660_);
  or g_107219_(_014532_, _014542_, _014661_);
  and g_107220_(_014545_, _014661_, _014663_);
  or g_107221_(_014544_, _014660_, _014664_);
  and g_107222_(_014659_, _014663_, _014665_);
  or g_107223_(_014658_, _014664_, _014666_);
  and g_107224_(_014522_, _014666_, _014667_);
  or g_107225_(_014523_, _014665_, _014668_);
  and g_107226_(_014500_, _014518_, _014669_);
  or g_107227_(_014501_, _014517_, _014670_);
  and g_107228_(_014478_, _014482_, _014671_);
  or g_107229_(_014477_, _014481_, _014672_);
  and g_107230_(_014670_, _014672_, _014674_);
  or g_107231_(_014669_, _014671_, _014675_);
  and g_107232_(_014668_, _014674_, _014676_);
  or g_107233_(_014667_, _014675_, _014677_);
  and g_107234_(_014655_, _014676_, _014678_);
  or g_107235_(_014654_, _014677_, _014679_);
  and g_107236_(_014643_, _014679_, _014680_);
  or g_107237_(_014642_, _014678_, _014681_);
  and g_107238_(_014469_, _014681_, _014682_);
  or g_107239_(_014468_, _014680_, _014683_);
  and g_107240_(_014470_, _014680_, _014685_);
  or g_107241_(_014471_, _014681_, _014686_);
  and g_107242_(_014683_, _014686_, _014687_);
  or g_107243_(_014682_, _014685_, _014688_);
  xor g_107244_(out[906], _009830_, _014689_);
  xor g_107245_(_001935_, _009830_, _014690_);
  and g_107246_(_014687_, _014689_, _014691_);
  or g_107247_(_014688_, _014690_, _014692_);
  and g_107248_(_009819_, _009835_, _014693_);
  or g_107249_(_009820_, _009834_, _014694_);
  and g_107250_(_014692_, _014694_, _014696_);
  or g_107251_(_014691_, _014693_, _014697_);
  and g_107252_(_009820_, _009834_, _014698_);
  or g_107253_(_009819_, _009835_, _014699_);
  and g_107254_(_014688_, _014690_, _014700_);
  or g_107255_(_014687_, _014689_, _014701_);
  and g_107256_(_014699_, _014701_, _014702_);
  or g_107257_(_014698_, _014700_, _014703_);
  and g_107258_(out[905], _009829_, _014704_);
  xor g_107259_(out[905], _009829_, _014705_);
  or g_107260_(_009831_, _014704_, _014707_);
  and g_107261_(_014492_, _014681_, _014708_);
  and g_107262_(_014485_, _014680_, _014709_);
  or g_107263_(_014708_, _014709_, _014710_);
  or g_107264_(_014705_, _014710_, _014711_);
  xor g_107265_(out[904], _009828_, _014712_);
  xor g_107266_(_001913_, _009828_, _014713_);
  and g_107267_(_014503_, _014680_, _014714_);
  not g_107268_(_014714_, _014715_);
  or g_107269_(_014509_, _014680_, _014716_);
  not g_107270_(_014716_, _014718_);
  and g_107271_(_014715_, _014716_, _014719_);
  or g_107272_(_014714_, _014718_, _014720_);
  and g_107273_(_014705_, _014710_, _014721_);
  and g_107274_(_014713_, _014719_, _014722_);
  or g_107275_(_014721_, _014722_, _014723_);
  xor g_107276_(_014713_, _014719_, _014724_);
  xor g_107277_(_014712_, _014719_, _014725_);
  and g_107278_(_014696_, _014702_, _014726_);
  or g_107279_(_014697_, _014703_, _014727_);
  xor g_107280_(_014705_, _014710_, _014729_);
  xor g_107281_(_014707_, _014710_, _014730_);
  and g_107282_(_014726_, _014729_, _014731_);
  or g_107283_(_014727_, _014730_, _014732_);
  and g_107284_(_014724_, _014731_, _014733_);
  or g_107285_(_014725_, _014732_, _014734_);
  xor g_107286_(out[903], _009827_, _014735_);
  xor g_107287_(_001825_, _009827_, _014736_);
  and g_107288_(_014533_, _014680_, _014737_);
  not g_107289_(_014737_, _014738_);
  or g_107290_(_014539_, _014680_, _014740_);
  not g_107291_(_014740_, _014741_);
  and g_107292_(_014738_, _014740_, _014742_);
  or g_107293_(_014737_, _014741_, _014743_);
  and g_107294_(_014736_, _014743_, _014744_);
  or g_107295_(_014735_, _014742_, _014745_);
  xor g_107296_(out[902], _009826_, _014746_);
  and g_107297_(_014525_, _014680_, _014747_);
  and g_107298_(_014529_, _014681_, _014748_);
  or g_107299_(_014747_, _014748_, _014749_);
  or g_107300_(_014746_, _014749_, _014751_);
  not g_107301_(_014751_, _014752_);
  or g_107302_(_014744_, _014752_, _014753_);
  and g_107303_(_014735_, _014742_, _014754_);
  or g_107304_(_014736_, _014743_, _014755_);
  and g_107305_(_014746_, _014749_, _014756_);
  or g_107306_(_014754_, _014756_, _014757_);
  and g_107307_(_014745_, _014755_, _014758_);
  xor g_107308_(_014746_, _014749_, _014759_);
  and g_107309_(_014758_, _014759_, _014760_);
  or g_107310_(_014753_, _014757_, _014762_);
  or g_107311_(_025530_, _002332_, _014763_);
  not g_107312_(_014763_, _014764_);
  and g_107313_(_009825_, _014763_, _014765_);
  or g_107314_(_009824_, _014764_, _014766_);
  and g_107315_(_014562_, _014681_, _014767_);
  and g_107316_(_014556_, _014680_, _014768_);
  or g_107317_(_014767_, _014768_, _014769_);
  or g_107318_(_014765_, _014769_, _014770_);
  not g_107319_(_014770_, _014771_);
  xor g_107320_(out[901], _009824_, _014773_);
  xor g_107321_(_001847_, _009824_, _014774_);
  and g_107322_(_014567_, _014680_, _014775_);
  not g_107323_(_014775_, _014776_);
  or g_107324_(_014572_, _014680_, _014777_);
  not g_107325_(_014777_, _014778_);
  and g_107326_(_014776_, _014777_, _014779_);
  or g_107327_(_014775_, _014778_, _014780_);
  and g_107328_(_014774_, _014779_, _014781_);
  or g_107329_(_014773_, _014780_, _014782_);
  and g_107330_(_014770_, _014782_, _014784_);
  or g_107331_(_014771_, _014781_, _014785_);
  and g_107332_(_014773_, _014780_, _014786_);
  or g_107333_(_014774_, _014779_, _014787_);
  and g_107334_(_014765_, _014769_, _014788_);
  or g_107335_(_014786_, _014788_, _014789_);
  not g_107336_(_014789_, _014790_);
  and g_107337_(_014784_, _014790_, _014791_);
  or g_107338_(_014785_, _014789_, _014792_);
  or g_107339_(_014762_, _014792_, _014793_);
  and g_107340_(_014733_, _014791_, _014795_);
  and g_107341_(_014760_, _014795_, _014796_);
  or g_107342_(_014734_, _014793_, _014797_);
  xor g_107343_(out[899], _002332_, _014798_);
  xor g_107344_(_001902_, _002332_, _014799_);
  and g_107345_(_014615_, _014680_, _014800_);
  and g_107346_(_014623_, _014681_, _014801_);
  or g_107347_(_014800_, _014801_, _014802_);
  not g_107348_(_014802_, _014803_);
  and g_107349_(_014798_, _014803_, _014804_);
  or g_107350_(_014799_, _014802_, _014806_);
  or g_107351_(_014611_, _014680_, _014807_);
  or g_107352_(_002077_, _014681_, _014808_);
  and g_107353_(_014807_, _014808_, _014809_);
  not g_107354_(_014809_, _014810_);
  and g_107355_(_002333_, _014809_, _014811_);
  or g_107356_(_002334_, _014810_, _014812_);
  and g_107357_(_014806_, _014812_, _014813_);
  or g_107358_(_014804_, _014811_, _014814_);
  and g_107359_(_014799_, _014802_, _014815_);
  or g_107360_(_014798_, _014803_, _014817_);
  and g_107361_(_002334_, _014810_, _014818_);
  or g_107362_(_002333_, _014809_, _014819_);
  and g_107363_(_014817_, _014819_, _014820_);
  or g_107364_(_014815_, _014818_, _014821_);
  and g_107365_(_014813_, _014820_, _014822_);
  or g_107366_(_014814_, _014821_, _014823_);
  and g_107367_(out[881], _014680_, _014824_);
  not g_107368_(_014824_, _014825_);
  or g_107369_(_014594_, _014680_, _014826_);
  not g_107370_(_014826_, _014828_);
  and g_107371_(_014825_, _014826_, _014829_);
  or g_107372_(_014824_, _014828_, _014830_);
  and g_107373_(out[897], _014829_, _014831_);
  or g_107374_(_001869_, _014830_, _014832_);
  and g_107375_(out[880], _014680_, _014833_);
  not g_107376_(_014833_, _014834_);
  or g_107377_(_014598_, _014680_, _014835_);
  not g_107378_(_014835_, _014836_);
  and g_107379_(_014834_, _014835_, _014837_);
  or g_107380_(_014833_, _014836_, _014839_);
  and g_107381_(out[896], _014837_, _014840_);
  or g_107382_(_001880_, _014839_, _014841_);
  xor g_107383_(out[897], _014829_, _014842_);
  xor g_107384_(_001869_, _014829_, _014843_);
  and g_107385_(_014841_, _014842_, _014844_);
  or g_107386_(_014840_, _014843_, _014845_);
  and g_107387_(_014832_, _014845_, _014846_);
  or g_107388_(_014831_, _014844_, _014847_);
  and g_107389_(_014822_, _014847_, _014848_);
  or g_107390_(_014823_, _014846_, _014850_);
  and g_107391_(_014814_, _014817_, _014851_);
  or g_107392_(_014813_, _014815_, _014852_);
  and g_107393_(_014850_, _014852_, _014853_);
  or g_107394_(_014848_, _014851_, _014854_);
  and g_107395_(_014796_, _014854_, _014855_);
  or g_107396_(_014797_, _014853_, _014856_);
  and g_107397_(_014785_, _014787_, _014857_);
  or g_107398_(_014784_, _014786_, _014858_);
  and g_107399_(_014760_, _014857_, _014859_);
  or g_107400_(_014762_, _014858_, _014861_);
  and g_107401_(_014745_, _014752_, _014862_);
  or g_107402_(_014744_, _014751_, _014863_);
  and g_107403_(_014755_, _014863_, _014864_);
  or g_107404_(_014754_, _014862_, _014865_);
  and g_107405_(_014861_, _014864_, _014866_);
  or g_107406_(_014859_, _014865_, _014867_);
  and g_107407_(_014733_, _014867_, _014868_);
  or g_107408_(_014734_, _014866_, _014869_);
  and g_107409_(_014697_, _014699_, _014870_);
  or g_107410_(_014696_, _014698_, _014872_);
  and g_107411_(_014723_, _014726_, _014873_);
  and g_107412_(_014711_, _014873_, _014874_);
  not g_107413_(_014874_, _014875_);
  and g_107414_(_014872_, _014875_, _014876_);
  or g_107415_(_014870_, _014874_, _014877_);
  and g_107416_(_014869_, _014876_, _014878_);
  or g_107417_(_014868_, _014877_, _014879_);
  and g_107418_(_014856_, _014878_, _014880_);
  or g_107419_(_014855_, _014879_, _014881_);
  or g_107420_(out[896], _014837_, _014883_);
  and g_107421_(_014796_, _014883_, _014884_);
  not g_107422_(_014884_, _014885_);
  and g_107423_(_014844_, _014884_, _014886_);
  or g_107424_(_014845_, _014885_, _014887_);
  and g_107425_(_014822_, _014886_, _014888_);
  or g_107426_(_014823_, _014887_, _014889_);
  and g_107427_(_014881_, _014889_, _014890_);
  or g_107428_(_014880_, _014888_, _014891_);
  and g_107429_(_014688_, _014891_, _014892_);
  or g_107430_(_014687_, _014890_, _014894_);
  and g_107431_(_014689_, _014890_, _014895_);
  or g_107432_(_014690_, _014891_, _014896_);
  and g_107433_(_014894_, _014896_, _014897_);
  or g_107434_(_014892_, _014895_, _014898_);
  xor g_107435_(out[915], _002528_, _014899_);
  xor g_107436_(_002034_, _002528_, _014900_);
  and g_107437_(_014798_, _014890_, _014901_);
  and g_107438_(_014802_, _014891_, _014902_);
  or g_107439_(_014901_, _014902_, _014903_);
  and g_107440_(_014900_, _014903_, _014905_);
  or g_107441_(_014900_, _014903_, _014906_);
  xor g_107442_(_014900_, _014903_, _014907_);
  xor g_107443_(_014899_, _014903_, _014908_);
  and g_107444_(_014810_, _014891_, _014909_);
  and g_107445_(_002333_, _014890_, _014910_);
  or g_107446_(_014909_, _014910_, _014911_);
  or g_107447_(_002531_, _014911_, _014912_);
  xor g_107448_(_002531_, _014911_, _014913_);
  xor g_107449_(_002530_, _014911_, _014914_);
  and g_107450_(_014907_, _014913_, _014916_);
  or g_107451_(_014908_, _014914_, _014917_);
  or g_107452_(_001869_, _014891_, _014918_);
  or g_107453_(_014829_, _014890_, _014919_);
  and g_107454_(_014918_, _014919_, _014920_);
  and g_107455_(out[913], _014920_, _014921_);
  not g_107456_(_014921_, _014922_);
  or g_107457_(_001880_, _014891_, _014923_);
  not g_107458_(_014923_, _014924_);
  and g_107459_(_014839_, _014891_, _014925_);
  or g_107460_(_014837_, _014890_, _014927_);
  and g_107461_(_014923_, _014927_, _014928_);
  or g_107462_(_014924_, _014925_, _014929_);
  and g_107463_(out[912], _014928_, _014930_);
  or g_107464_(_002012_, _014929_, _014931_);
  xor g_107465_(out[913], _014920_, _014932_);
  xor g_107466_(_002001_, _014920_, _014933_);
  and g_107467_(_014931_, _014932_, _014934_);
  or g_107468_(_014930_, _014933_, _014935_);
  and g_107469_(_014922_, _014935_, _014936_);
  or g_107470_(_014921_, _014934_, _014938_);
  and g_107471_(_014916_, _014938_, _014939_);
  or g_107472_(_014917_, _014936_, _014940_);
  and g_107473_(_014906_, _014912_, _014941_);
  or g_107474_(_014905_, _014941_, _014942_);
  not g_107475_(_014942_, _014943_);
  and g_107476_(_014940_, _014942_, _014944_);
  or g_107477_(_014939_, _014943_, _014945_);
  xor g_107478_(out[922], _009847_, _014946_);
  xor g_107479_(_002067_, _009847_, _014947_);
  and g_107480_(_014897_, _014946_, _014949_);
  or g_107481_(_014898_, _014947_, _014950_);
  and g_107482_(_009836_, _009851_, _014951_);
  or g_107483_(_009837_, _009850_, _014952_);
  and g_107484_(_014950_, _014952_, _014953_);
  or g_107485_(_014949_, _014951_, _014954_);
  and g_107486_(_009837_, _009850_, _014955_);
  or g_107487_(_009836_, _009851_, _014956_);
  and g_107488_(_014898_, _014947_, _014957_);
  or g_107489_(_014897_, _014946_, _014958_);
  and g_107490_(_014956_, _014958_, _014960_);
  or g_107491_(_014955_, _014957_, _014961_);
  and g_107492_(out[921], _009846_, _014962_);
  xor g_107493_(out[921], _009846_, _014963_);
  or g_107494_(_009848_, _014962_, _014964_);
  and g_107495_(_014710_, _014891_, _014965_);
  and g_107496_(_014707_, _014890_, _014966_);
  or g_107497_(_014965_, _014966_, _014967_);
  or g_107498_(_014963_, _014967_, _014968_);
  not g_107499_(_014968_, _014969_);
  xor g_107500_(out[920], _009845_, _014971_);
  xor g_107501_(_002045_, _009845_, _014972_);
  and g_107502_(_014713_, _014890_, _014973_);
  and g_107503_(_014720_, _014891_, _014974_);
  or g_107504_(_014973_, _014974_, _014975_);
  and g_107505_(_014963_, _014967_, _014976_);
  not g_107506_(_014976_, _014977_);
  or g_107507_(_014971_, _014975_, _014978_);
  and g_107508_(_014977_, _014978_, _014979_);
  xor g_107509_(_014971_, _014975_, _014980_);
  xor g_107510_(_014972_, _014975_, _014982_);
  and g_107511_(_014953_, _014960_, _014983_);
  or g_107512_(_014954_, _014961_, _014984_);
  and g_107513_(_014968_, _014977_, _014985_);
  or g_107514_(_014969_, _014976_, _014986_);
  and g_107515_(_014983_, _014985_, _014987_);
  or g_107516_(_014984_, _014986_, _014988_);
  and g_107517_(_014980_, _014987_, _014989_);
  or g_107518_(_014982_, _014988_, _014990_);
  xor g_107519_(out[919], _009843_, _014991_);
  xor g_107520_(_001957_, _009843_, _014993_);
  and g_107521_(_014735_, _014890_, _014994_);
  or g_107522_(_014736_, _014891_, _014995_);
  and g_107523_(_014743_, _014891_, _014996_);
  or g_107524_(_014742_, _014890_, _014997_);
  and g_107525_(_014995_, _014997_, _014998_);
  or g_107526_(_014994_, _014996_, _014999_);
  and g_107527_(_014991_, _014998_, _015000_);
  or g_107528_(_014993_, _014999_, _015001_);
  xor g_107529_(out[918], _009842_, _015002_);
  not g_107530_(_015002_, _015004_);
  or g_107531_(_014746_, _014891_, _015005_);
  not g_107532_(_015005_, _015006_);
  and g_107533_(_014749_, _014891_, _015007_);
  not g_107534_(_015007_, _015008_);
  and g_107535_(_015005_, _015008_, _015009_);
  or g_107536_(_015006_, _015007_, _015010_);
  and g_107537_(_015002_, _015010_, _015011_);
  or g_107538_(_015004_, _015009_, _015012_);
  and g_107539_(_015001_, _015012_, _015013_);
  or g_107540_(_015000_, _015011_, _015015_);
  and g_107541_(_015004_, _015009_, _015016_);
  or g_107542_(_015002_, _015010_, _015017_);
  xor g_107543_(out[917], _009840_, _015018_);
  xor g_107544_(_001979_, _009840_, _015019_);
  and g_107545_(_014780_, _014891_, _015020_);
  or g_107546_(_014779_, _014890_, _015021_);
  and g_107547_(_014774_, _014890_, _015022_);
  or g_107548_(_014773_, _014891_, _015023_);
  and g_107549_(_015021_, _015023_, _015024_);
  or g_107550_(_015020_, _015022_, _015026_);
  and g_107551_(_015018_, _015026_, _015027_);
  or g_107552_(_015019_, _015024_, _015028_);
  and g_107553_(_014993_, _014999_, _015029_);
  or g_107554_(_014991_, _014998_, _015030_);
  and g_107555_(_015028_, _015030_, _015031_);
  or g_107556_(_015027_, _015029_, _015032_);
  and g_107557_(_015017_, _015031_, _015033_);
  or g_107558_(_015016_, _015032_, _015034_);
  and g_107559_(_015013_, _015033_, _015035_);
  or g_107560_(_015015_, _015034_, _015037_);
  or g_107561_(_025684_, _002528_, _015038_);
  not g_107562_(_015038_, _015039_);
  and g_107563_(_009841_, _015038_, _015040_);
  or g_107564_(_009840_, _015039_, _015041_);
  and g_107565_(_014769_, _014891_, _015042_);
  not g_107566_(_015042_, _015043_);
  or g_107567_(_014765_, _014891_, _015044_);
  not g_107568_(_015044_, _015045_);
  and g_107569_(_015043_, _015044_, _015046_);
  or g_107570_(_015042_, _015045_, _015048_);
  and g_107571_(_015041_, _015046_, _015049_);
  or g_107572_(_015040_, _015048_, _015050_);
  or g_107573_(_015018_, _015026_, _015051_);
  not g_107574_(_015051_, _015052_);
  and g_107575_(_015050_, _015051_, _015053_);
  or g_107576_(_015049_, _015052_, _015054_);
  and g_107577_(_015040_, _015048_, _015055_);
  not g_107578_(_015055_, _015056_);
  and g_107579_(_015053_, _015056_, _015057_);
  or g_107580_(_015054_, _015055_, _015059_);
  and g_107581_(_015035_, _015057_, _015060_);
  or g_107582_(_015037_, _015059_, _015061_);
  and g_107583_(_014989_, _015060_, _015062_);
  or g_107584_(_014990_, _015061_, _015063_);
  and g_107585_(_014945_, _015062_, _015064_);
  or g_107586_(_014944_, _015063_, _015065_);
  and g_107587_(_015035_, _015054_, _015066_);
  or g_107588_(_015037_, _015053_, _015067_);
  or g_107589_(_015017_, _015029_, _015068_);
  not g_107590_(_015068_, _015070_);
  and g_107591_(_015001_, _015068_, _015071_);
  or g_107592_(_015000_, _015070_, _015072_);
  and g_107593_(_015067_, _015071_, _015073_);
  or g_107594_(_015066_, _015072_, _015074_);
  and g_107595_(_014989_, _015074_, _015075_);
  or g_107596_(_014990_, _015073_, _015076_);
  or g_107597_(_014953_, _014955_, _015077_);
  not g_107598_(_015077_, _015078_);
  or g_107599_(_014979_, _014984_, _015079_);
  not g_107600_(_015079_, _015081_);
  and g_107601_(_014968_, _015081_, _015082_);
  or g_107602_(_014969_, _015079_, _015083_);
  and g_107603_(_015077_, _015083_, _015084_);
  or g_107604_(_015078_, _015082_, _015085_);
  and g_107605_(_015076_, _015084_, _015086_);
  or g_107606_(_015075_, _015085_, _015087_);
  and g_107607_(_015065_, _015086_, _015088_);
  or g_107608_(_015064_, _015087_, _015089_);
  or g_107609_(out[912], _014928_, _015090_);
  not g_107610_(_015090_, _015092_);
  or g_107611_(_014917_, _014935_, _015093_);
  or g_107612_(_015063_, _015093_, _015094_);
  not g_107613_(_015094_, _015095_);
  and g_107614_(_015090_, _015095_, _015096_);
  or g_107615_(_015092_, _015094_, _015097_);
  and g_107616_(_015089_, _015097_, _015098_);
  or g_107617_(_015088_, _015096_, _015099_);
  and g_107618_(_014898_, _015099_, _015100_);
  not g_107619_(_015100_, _015101_);
  or g_107620_(_014947_, _015099_, _015103_);
  not g_107621_(_015103_, _015104_);
  and g_107622_(_015101_, _015103_, _015105_);
  or g_107623_(_015100_, _015104_, _015106_);
  and g_107624_(_009857_, _015105_, _015107_);
  or g_107625_(_009858_, _015106_, _015108_);
  and g_107626_(_009854_, _015108_, _015109_);
  or g_107627_(_009856_, _015107_, _015110_);
  and g_107628_(_009409_, _009853_, _015111_);
  or g_107629_(_009410_, _009852_, _015112_);
  and g_107630_(_009858_, _015106_, _015114_);
  or g_107631_(_009857_, _015105_, _015115_);
  and g_107632_(_015112_, _015115_, _015116_);
  or g_107633_(_015111_, _015114_, _015117_);
  and g_107634_(out[937], _009406_, _015118_);
  xor g_107635_(out[937], _009406_, _015119_);
  xor g_107636_(_002166_, _009406_, _015120_);
  and g_107637_(_014967_, _015099_, _015121_);
  not g_107638_(_015121_, _015122_);
  or g_107639_(_014963_, _015099_, _015123_);
  and g_107640_(_015122_, _015123_, _015125_);
  not g_107641_(_015125_, _015126_);
  or g_107642_(_015119_, _015126_, _015127_);
  xor g_107643_(out[936], _009405_, _015128_);
  xor g_107644_(_002155_, _009405_, _015129_);
  or g_107645_(_014971_, _015099_, _015130_);
  and g_107646_(_014975_, _015099_, _015131_);
  not g_107647_(_015131_, _015132_);
  and g_107648_(_015130_, _015132_, _015133_);
  and g_107649_(_015119_, _015126_, _015134_);
  and g_107650_(_015129_, _015133_, _015136_);
  or g_107651_(_015134_, _015136_, _015137_);
  xor g_107652_(_015129_, _015133_, _015138_);
  xor g_107653_(_015128_, _015133_, _015139_);
  and g_107654_(_015109_, _015116_, _015140_);
  or g_107655_(_015110_, _015117_, _015141_);
  xor g_107656_(_015120_, _015125_, _015142_);
  xor g_107657_(_015119_, _015125_, _015143_);
  and g_107658_(_015140_, _015142_, _015144_);
  or g_107659_(_015141_, _015143_, _015145_);
  and g_107660_(_015138_, _015144_, _015147_);
  or g_107661_(_015139_, _015145_, _015148_);
  xor g_107662_(out[935], _009403_, _015149_);
  xor g_107663_(_002078_, _009403_, _015150_);
  or g_107664_(_014993_, _015099_, _015151_);
  or g_107665_(_014998_, _015098_, _015152_);
  and g_107666_(_015151_, _015152_, _015153_);
  or g_107667_(_015149_, _015153_, _015154_);
  xor g_107668_(out[934], _009402_, _015155_);
  not g_107669_(_015155_, _015156_);
  or g_107670_(_015002_, _015099_, _015158_);
  or g_107671_(_015009_, _015098_, _015159_);
  and g_107672_(_015158_, _015159_, _015160_);
  and g_107673_(_015156_, _015160_, _015161_);
  and g_107674_(_015149_, _015153_, _015162_);
  xor g_107675_(_015149_, _015153_, _015163_);
  xor g_107676_(_015150_, _015153_, _015164_);
  xor g_107677_(_015156_, _015160_, _015165_);
  xor g_107678_(_015155_, _015160_, _015166_);
  and g_107679_(_015163_, _015165_, _015167_);
  or g_107680_(_015164_, _015166_, _015169_);
  or g_107681_(_025838_, _002719_, _015170_);
  not g_107682_(_015170_, _015171_);
  and g_107683_(_009401_, _015170_, _015172_);
  or g_107684_(_009400_, _015171_, _015173_);
  or g_107685_(_015046_, _015098_, _015174_);
  or g_107686_(_015040_, _015099_, _015175_);
  and g_107687_(_015174_, _015175_, _015176_);
  and g_107688_(_015173_, _015176_, _015177_);
  xor g_107689_(out[933], _009400_, _015178_);
  xor g_107690_(_002089_, _009400_, _015180_);
  or g_107691_(_015018_, _015099_, _015181_);
  or g_107692_(_015024_, _015098_, _015182_);
  and g_107693_(_015181_, _015182_, _015183_);
  and g_107694_(_015180_, _015183_, _015184_);
  or g_107695_(_015177_, _015184_, _015185_);
  or g_107696_(_015180_, _015183_, _015186_);
  or g_107697_(_015173_, _015176_, _015187_);
  and g_107698_(_015186_, _015187_, _015188_);
  not g_107699_(_015188_, _015189_);
  or g_107700_(_015185_, _015189_, _015191_);
  or g_107701_(_015169_, _015191_, _015192_);
  not g_107702_(_015192_, _015193_);
  and g_107703_(_015147_, _015193_, _015194_);
  or g_107704_(_015148_, _015192_, _015195_);
  xor g_107705_(out[931], _002719_, _015196_);
  xor g_107706_(_002144_, _002719_, _015197_);
  and g_107707_(_014899_, _015098_, _015198_);
  and g_107708_(_014903_, _015099_, _015199_);
  or g_107709_(_015198_, _015199_, _015200_);
  not g_107710_(_015200_, _015202_);
  and g_107711_(_015197_, _015200_, _015203_);
  or g_107712_(_015196_, _015202_, _015204_);
  and g_107713_(_014911_, _015099_, _015205_);
  not g_107714_(_015205_, _015206_);
  or g_107715_(_002531_, _015099_, _015207_);
  and g_107716_(_015206_, _015207_, _015208_);
  and g_107717_(_002720_, _015208_, _015209_);
  not g_107718_(_015209_, _015210_);
  and g_107719_(_015196_, _015202_, _015211_);
  or g_107720_(_015197_, _015200_, _015213_);
  and g_107721_(_015210_, _015213_, _015214_);
  or g_107722_(_015209_, _015211_, _015215_);
  or g_107723_(_002001_, _015099_, _015216_);
  or g_107724_(_014920_, _015098_, _015217_);
  and g_107725_(_015216_, _015217_, _015218_);
  and g_107726_(out[929], _015218_, _015219_);
  not g_107727_(_015219_, _015220_);
  or g_107728_(_002012_, _015099_, _015221_);
  or g_107729_(_014928_, _015098_, _015222_);
  and g_107730_(_015221_, _015222_, _015224_);
  and g_107731_(out[928], _015224_, _015225_);
  not g_107732_(_015225_, _015226_);
  xor g_107733_(out[929], _015218_, _015227_);
  xor g_107734_(_002111_, _015218_, _015228_);
  and g_107735_(_015226_, _015227_, _015229_);
  or g_107736_(_015225_, _015228_, _015230_);
  and g_107737_(_015220_, _015230_, _015231_);
  or g_107738_(_015219_, _015229_, _015232_);
  xor g_107739_(_002721_, _015208_, _015233_);
  or g_107740_(_015231_, _015233_, _015235_);
  and g_107741_(_015214_, _015235_, _015236_);
  or g_107742_(_015203_, _015211_, _015237_);
  or g_107743_(_015233_, _015237_, _015238_);
  not g_107744_(_015238_, _015239_);
  and g_107745_(_015232_, _015239_, _015240_);
  and g_107746_(_015204_, _015215_, _015241_);
  or g_107747_(_015240_, _015241_, _015242_);
  or g_107748_(_015203_, _015236_, _015243_);
  and g_107749_(_015194_, _015242_, _015244_);
  or g_107750_(_015195_, _015243_, _015246_);
  and g_107751_(_015167_, _015185_, _015247_);
  and g_107752_(_015186_, _015247_, _015248_);
  and g_107753_(_015154_, _015161_, _015249_);
  or g_107754_(_015162_, _015249_, _015250_);
  or g_107755_(_015248_, _015250_, _015251_);
  and g_107756_(_015147_, _015251_, _015252_);
  and g_107757_(_015137_, _015140_, _015253_);
  and g_107758_(_015127_, _015253_, _015254_);
  and g_107759_(_015110_, _015112_, _015255_);
  or g_107760_(_015254_, _015255_, _015257_);
  or g_107761_(_015252_, _015257_, _015258_);
  not g_107762_(_015258_, _015259_);
  and g_107763_(_015246_, _015259_, _015260_);
  or g_107764_(_015244_, _015258_, _015261_);
  or g_107765_(out[928], _015224_, _015262_);
  not g_107766_(_015262_, _015263_);
  and g_107767_(_015194_, _015262_, _015264_);
  or g_107768_(_015195_, _015263_, _015265_);
  and g_107769_(_015229_, _015264_, _015266_);
  or g_107770_(_015230_, _015265_, _015268_);
  and g_107771_(_015239_, _015266_, _015269_);
  or g_107772_(_015238_, _015268_, _015270_);
  and g_107773_(_015261_, _015270_, _015271_);
  or g_107774_(_015260_, _015269_, _015272_);
  and g_107775_(_009409_, _015271_, _015273_);
  or g_107776_(_009853_, _015271_, _015274_);
  not g_107777_(_015274_, _015275_);
  or g_107778_(_015273_, _015275_, _015276_);
  not g_107779_(_015276_, _015277_);
  and g_107780_(_009396_, _015277_, _015279_);
  xor g_107781_(out[954], _009392_, _015280_);
  xor g_107782_(_002287_, _009392_, _015281_);
  and g_107783_(_015106_, _015272_, _015282_);
  and g_107784_(_009857_, _015271_, _015283_);
  or g_107785_(_015282_, _015283_, _015284_);
  not g_107786_(_015284_, _015285_);
  and g_107787_(_015281_, _015284_, _015286_);
  or g_107788_(_015279_, _015286_, _015287_);
  and g_107789_(_015280_, _015285_, _015288_);
  or g_107790_(_015281_, _015284_, _015290_);
  and g_107791_(_009397_, _015276_, _015291_);
  or g_107792_(_009396_, _015277_, _015292_);
  and g_107793_(_015290_, _015292_, _015293_);
  or g_107794_(_015288_, _015291_, _015294_);
  or g_107795_(_015287_, _015294_, _015295_);
  xor g_107796_(out[952], _009388_, _015296_);
  xor g_107797_(_002265_, _009388_, _015297_);
  or g_107798_(_015128_, _015272_, _015298_);
  or g_107799_(_015133_, _015271_, _015299_);
  and g_107800_(_015298_, _015299_, _015301_);
  and g_107801_(_015297_, _015301_, _015302_);
  and g_107802_(out[953], _009391_, _015303_);
  xor g_107803_(out[953], _009391_, _015304_);
  or g_107804_(_009394_, _015303_, _015305_);
  and g_107805_(_015126_, _015272_, _015306_);
  and g_107806_(_015120_, _015271_, _015307_);
  or g_107807_(_015306_, _015307_, _015308_);
  and g_107808_(_015304_, _015308_, _015309_);
  or g_107809_(_015302_, _015309_, _015310_);
  not g_107810_(_015310_, _015312_);
  or g_107811_(_015304_, _015308_, _015313_);
  or g_107812_(_015297_, _015301_, _015314_);
  and g_107813_(_015313_, _015314_, _015315_);
  not g_107814_(_015315_, _015316_);
  and g_107815_(_015312_, _015315_, _015317_);
  or g_107816_(_015310_, _015316_, _015318_);
  xor g_107817_(out[950], _009386_, _015319_);
  xor g_107818_(_002199_, _009386_, _015320_);
  or g_107819_(_015155_, _015272_, _015321_);
  or g_107820_(_015160_, _015271_, _015323_);
  and g_107821_(_015321_, _015323_, _015324_);
  and g_107822_(_015320_, _015324_, _015325_);
  or g_107823_(_015150_, _015272_, _015326_);
  or g_107824_(_015153_, _015271_, _015327_);
  and g_107825_(_015326_, _015327_, _015328_);
  and g_107826_(_009389_, _015328_, _015329_);
  or g_107827_(_015325_, _015329_, _015330_);
  or g_107828_(_009389_, _015328_, _015331_);
  or g_107829_(_015320_, _015324_, _015332_);
  and g_107830_(_015331_, _015332_, _015334_);
  not g_107831_(_015334_, _015335_);
  or g_107832_(_015330_, _015335_, _015336_);
  xor g_107833_(out[948], _009384_, _015337_);
  xor g_107834_(_002221_, _009384_, _015338_);
  or g_107835_(_015176_, _015271_, _015339_);
  not g_107836_(_015339_, _015340_);
  and g_107837_(_015173_, _015271_, _015341_);
  or g_107838_(_015340_, _015341_, _015342_);
  or g_107839_(_015337_, _015342_, _015343_);
  xor g_107840_(out[949], _009385_, _015345_);
  xor g_107841_(_002210_, _009385_, _015346_);
  and g_107842_(_015180_, _015271_, _015347_);
  or g_107843_(_015183_, _015271_, _015348_);
  not g_107844_(_015348_, _015349_);
  or g_107845_(_015347_, _015349_, _015350_);
  or g_107846_(_015345_, _015350_, _015351_);
  and g_107847_(_015343_, _015351_, _015352_);
  not g_107848_(_015352_, _015353_);
  and g_107849_(_015345_, _015350_, _015354_);
  and g_107850_(_015337_, _015342_, _015356_);
  or g_107851_(_015354_, _015356_, _015357_);
  or g_107852_(_015336_, _015357_, _015358_);
  or g_107853_(_015353_, _015358_, _015359_);
  xor g_107854_(out[947], _002904_, _015360_);
  xor g_107855_(_002254_, _002904_, _015361_);
  and g_107856_(_015196_, _015271_, _015362_);
  and g_107857_(_015200_, _015272_, _015363_);
  or g_107858_(_015362_, _015363_, _015364_);
  or g_107859_(_015361_, _015364_, _015365_);
  or g_107860_(_015208_, _015271_, _015367_);
  not g_107861_(_015367_, _015368_);
  and g_107862_(_002720_, _015271_, _015369_);
  or g_107863_(_015368_, _015369_, _015370_);
  and g_107864_(_015361_, _015364_, _015371_);
  or g_107865_(_002906_, _015370_, _015372_);
  xor g_107866_(_015361_, _015364_, _015373_);
  xor g_107867_(_015360_, _015364_, _015374_);
  xor g_107868_(_002906_, _015370_, _015375_);
  xor g_107869_(_002905_, _015370_, _015376_);
  and g_107870_(_015373_, _015375_, _015378_);
  or g_107871_(_015374_, _015376_, _015379_);
  or g_107872_(_002111_, _015272_, _015380_);
  or g_107873_(_015218_, _015271_, _015381_);
  and g_107874_(_015380_, _015381_, _015382_);
  and g_107875_(out[945], _015382_, _015383_);
  and g_107876_(_015378_, _015383_, _015384_);
  not g_107877_(_015384_, _015385_);
  or g_107878_(_015371_, _015372_, _015386_);
  and g_107879_(_015365_, _015386_, _015387_);
  and g_107880_(out[928], _015271_, _015389_);
  or g_107881_(_015224_, _015271_, _015390_);
  not g_107882_(_015390_, _015391_);
  or g_107883_(_015389_, _015391_, _015392_);
  not g_107884_(_015392_, _015393_);
  and g_107885_(out[944], _015393_, _015394_);
  or g_107886_(_002232_, _015392_, _015395_);
  xor g_107887_(out[945], _015382_, _015396_);
  xor g_107888_(_054336_, _015382_, _015397_);
  and g_107889_(_015395_, _015396_, _015398_);
  or g_107890_(_015394_, _015397_, _015400_);
  and g_107891_(_015378_, _015398_, _015401_);
  or g_107892_(_015379_, _015400_, _015402_);
  and g_107893_(_015387_, _015402_, _015403_);
  and g_107894_(_015385_, _015403_, _015404_);
  or g_107895_(_015359_, _015404_, _015405_);
  and g_107896_(_015330_, _015331_, _015406_);
  not g_107897_(_015406_, _015407_);
  or g_107898_(_015352_, _015354_, _015408_);
  or g_107899_(_015336_, _015408_, _015409_);
  and g_107900_(_015407_, _015409_, _015411_);
  and g_107901_(_015405_, _015411_, _015412_);
  or g_107902_(_015318_, _015412_, _015413_);
  and g_107903_(_015302_, _015313_, _015414_);
  or g_107904_(_015309_, _015414_, _015415_);
  not g_107905_(_015415_, _015416_);
  and g_107906_(_015413_, _015416_, _015417_);
  or g_107907_(_015295_, _015417_, _015418_);
  or g_107908_(_015279_, _015293_, _015419_);
  and g_107909_(_015418_, _015419_, _015420_);
  or g_107910_(out[944], _015393_, _015422_);
  or g_107911_(_015295_, _015359_, _015423_);
  not g_107912_(_015423_, _015424_);
  and g_107913_(_015401_, _015422_, _015425_);
  and g_107914_(_015317_, _015424_, _015426_);
  and g_107915_(_015425_, _015426_, _015427_);
  or g_107916_(_015420_, _015427_, _015428_);
  not g_107917_(_015428_, _015429_);
  or g_107918_(_009390_, _015428_, _015430_);
  or g_107919_(_015328_, _015429_, _015431_);
  and g_107920_(_015430_, _015431_, _015433_);
  or g_107921_(_009383_, _015433_, _015434_);
  and g_107922_(_009181_, _009183_, _015435_);
  and g_107923_(_009396_, _015276_, _015436_);
  xor g_107924_(_015435_, _015436_, _015437_);
  or g_107925_(_009233_, _009379_, _015438_);
  or g_107926_(_009236_, _009378_, _015439_);
  and g_107927_(_015438_, _015439_, _015440_);
  or g_107928_(_015324_, _015429_, _015441_);
  or g_107929_(_015319_, _015428_, _015442_);
  and g_107930_(_015441_, _015442_, _015444_);
  and g_107931_(out[465], _009378_, _015445_);
  and g_107932_(_009320_, _009379_, _015446_);
  or g_107933_(_015445_, _015446_, _015447_);
  or g_107934_(_054336_, _015428_, _015448_);
  or g_107935_(_015382_, _015429_, _015449_);
  and g_107936_(_015448_, _015449_, _015450_);
  or g_107937_(_015447_, _015450_, _015451_);
  or g_107938_(_009204_, _009379_, _015452_);
  or g_107939_(_009209_, _009378_, _015453_);
  and g_107940_(_015452_, _015453_, _015455_);
  and g_107941_(_015301_, _015428_, _015456_);
  and g_107942_(_015296_, _015429_, _015457_);
  or g_107943_(_015456_, _015457_, _015458_);
  xor g_107944_(_015455_, _015458_, _015459_);
  and g_107945_(_009271_, _009379_, _015460_);
  or g_107946_(_009270_, _009378_, _015461_);
  and g_107947_(_009265_, _009378_, _015462_);
  or g_107948_(_009264_, _009379_, _015463_);
  and g_107949_(_015461_, _015463_, _015464_);
  or g_107950_(_015460_, _015462_, _015466_);
  or g_107951_(_015345_, _015428_, _015467_);
  not g_107952_(_015467_, _015468_);
  and g_107953_(_015350_, _015428_, _015469_);
  not g_107954_(_015469_, _015470_);
  and g_107955_(_015467_, _015470_, _015471_);
  or g_107956_(_015468_, _015469_, _015472_);
  and g_107957_(_009199_, _009379_, _015473_);
  or g_107958_(_009198_, _009378_, _015474_);
  and g_107959_(_009192_, _009378_, _015475_);
  or g_107960_(_009191_, _009379_, _015477_);
  and g_107961_(_015474_, _015477_, _015478_);
  or g_107962_(_015473_, _015475_, _015479_);
  and g_107963_(_015308_, _015428_, _015480_);
  not g_107964_(_015480_, _015481_);
  or g_107965_(_015304_, _015428_, _015482_);
  not g_107966_(_015482_, _015483_);
  and g_107967_(_015481_, _015482_, _015484_);
  or g_107968_(_015480_, _015483_, _015485_);
  or g_107969_(_015478_, _015485_, _015486_);
  or g_107970_(_009178_, _009378_, _015488_);
  or g_107971_(_003136_, _009379_, _015489_);
  and g_107972_(_015488_, _015489_, _015490_);
  or g_107973_(_015281_, _015428_, _015491_);
  or g_107974_(_015285_, _015429_, _015492_);
  and g_107975_(_015491_, _015492_, _015493_);
  or g_107976_(_015479_, _015484_, _015494_);
  and g_107977_(_015338_, _015429_, _015495_);
  and g_107978_(_015342_, _015428_, _015496_);
  or g_107979_(_015495_, _015496_, _015497_);
  and g_107980_(_009254_, _009378_, _015499_);
  and g_107981_(_009259_, _009379_, _015500_);
  or g_107982_(_015499_, _015500_, _015501_);
  and g_107983_(_015497_, _015501_, _015502_);
  or g_107984_(_009291_, _009379_, _015503_);
  or g_107985_(_009296_, _009378_, _015504_);
  and g_107986_(_015503_, _015504_, _015505_);
  and g_107987_(_015360_, _015429_, _015506_);
  and g_107988_(_015364_, _015428_, _015507_);
  or g_107989_(_015506_, _015507_, _015508_);
  or g_107990_(_015505_, _015508_, _015510_);
  and g_107991_(_009383_, _015433_, _015511_);
  and g_107992_(_015505_, _015508_, _015512_);
  or g_107993_(_009328_, _009378_, _015513_);
  or g_107994_(out[464], _009379_, _015514_);
  and g_107995_(_015513_, _015514_, _015515_);
  or g_107996_(_015392_, _015429_, _015516_);
  or g_107997_(out[944], _015428_, _015517_);
  and g_107998_(_015516_, _015517_, _015518_);
  and g_107999_(_009302_, _009379_, _015519_);
  and g_108000_(_053881_, _009378_, _015521_);
  or g_108001_(_015519_, _015521_, _015522_);
  and g_108002_(_015370_, _015428_, _015523_);
  and g_108003_(_002905_, _015429_, _015524_);
  or g_108004_(_015523_, _015524_, _015525_);
  or g_108005_(_015497_, _015501_, _015526_);
  and g_108006_(_015447_, _015450_, _015527_);
  or g_108007_(_015466_, _015471_, _015528_);
  or g_108008_(_015464_, _015472_, _015529_);
  and g_108009_(_015486_, _015510_, _015530_);
  and g_108010_(_015529_, _015530_, _015532_);
  and g_108011_(_015494_, _015526_, _015533_);
  and g_108012_(_015434_, _015451_, _015534_);
  and g_108013_(_015533_, _015534_, _015535_);
  and g_108014_(_015532_, _015535_, _015536_);
  and g_108015_(_015528_, _015536_, _015537_);
  xor g_108016_(_015490_, _015493_, _015538_);
  or g_108017_(_015459_, _015538_, _015539_);
  xor g_108018_(_015515_, _015518_, _015540_);
  xor g_108019_(_015440_, _015444_, _015541_);
  or g_108020_(_015540_, _015541_, _015543_);
  or g_108021_(_015539_, _015543_, _015544_);
  or g_108022_(_015437_, _015527_, _015545_);
  xor g_108023_(_015522_, _015525_, _015546_);
  or g_108024_(_015502_, _015512_, _015547_);
  or g_108025_(_015546_, _015547_, _015548_);
  or g_108026_(_015511_, _015548_, _015549_);
  or g_108027_(_015545_, _015549_, _015550_);
  or g_108028_(_015544_, _015550_, _015551_);
  not g_108029_(_015551_, _015552_);
  and g_108030_(_015537_, _015552_, _015554_);
  not g_108031_(_015554_, _015555_);
  and g_108032_(out[4], out[3], _015556_);
  not g_108033_(_015556_, _015557_);
  or g_108034_(out[5], _015556_, _015558_);
  or g_108035_(out[6], _015558_, _015559_);
  or g_108036_(out[7], _015559_, _015560_);
  or g_108037_(out[8], _015560_, _015561_);
  and g_108038_(out[9], _015561_, _015562_);
  or g_108039_(out[10], _015562_, _015563_);
  xor g_108040_(out[11], _015563_, _015565_);
  xor g_108041_(_002298_, _015563_, _015566_);
  and g_108042_(out[20], out[19], _015567_);
  not g_108043_(_015567_, _015568_);
  or g_108044_(out[21], _015567_, _015569_);
  or g_108045_(out[22], _015569_, _015570_);
  or g_108046_(out[23], _015570_, _015571_);
  or g_108047_(out[24], _015571_, _015572_);
  and g_108048_(out[25], _015572_, _015573_);
  or g_108049_(out[26], _015573_, _015574_);
  xor g_108050_(out[27], _015574_, _015576_);
  xor g_108051_(_002430_, _015574_, _015577_);
  and g_108052_(_015566_, _015576_, _015578_);
  or g_108053_(_015565_, _015577_, _015579_);
  xor g_108054_(out[24], _015571_, _015580_);
  xor g_108055_(_002529_, _015571_, _015581_);
  xor g_108056_(out[8], _015560_, _015582_);
  xor g_108057_(_002397_, _015560_, _015583_);
  and g_108058_(_015581_, _015582_, _015584_);
  or g_108059_(_015580_, _015583_, _015585_);
  xor g_108060_(out[7], _015559_, _015587_);
  not g_108061_(_015587_, _015588_);
  xor g_108062_(out[23], _015570_, _015589_);
  not g_108063_(_015589_, _015590_);
  and g_108064_(_015588_, _015589_, _015591_);
  or g_108065_(_015587_, _015590_, _015592_);
  and g_108066_(_015587_, _015590_, _015593_);
  or g_108067_(_015588_, _015589_, _015594_);
  and g_108068_(_002375_, out[18], _015595_);
  or g_108069_(out[2], _002507_, _015596_);
  and g_108070_(_002386_, out[19], _015598_);
  or g_108071_(out[3], _002518_, _015599_);
  and g_108072_(out[2], _002507_, _015600_);
  or g_108073_(_002375_, out[18], _015601_);
  and g_108074_(_006016_, _015601_, _015602_);
  or g_108075_(_006005_, _015600_, _015603_);
  and g_108076_(_006082_, _015602_, _015604_);
  or g_108077_(_006071_, _015603_, _015605_);
  and g_108078_(_015596_, _015605_, _015606_);
  or g_108079_(_015595_, _015604_, _015607_);
  and g_108080_(_015599_, _015607_, _015609_);
  or g_108081_(_015598_, _015606_, _015610_);
  and g_108082_(out[3], _002518_, _015611_);
  or g_108083_(_002386_, out[19], _015612_);
  and g_108084_(_005301_, _015557_, _015613_);
  or g_108085_(_005312_, _015556_, _015614_);
  and g_108086_(_005466_, _015568_, _015615_);
  or g_108087_(_005477_, _015567_, _015616_);
  and g_108088_(_015614_, _015615_, _015617_);
  or g_108089_(_015613_, _015616_, _015618_);
  and g_108090_(_015612_, _015618_, _015620_);
  or g_108091_(_015611_, _015617_, _015621_);
  and g_108092_(_006324_, _015620_, _015622_);
  or g_108093_(_006313_, _015621_, _015623_);
  and g_108094_(_015610_, _015622_, _015624_);
  or g_108095_(_015609_, _015623_, _015625_);
  and g_108096_(_015613_, _015616_, _015626_);
  or g_108097_(_015614_, _015615_, _015627_);
  and g_108098_(out[5], _015556_, _015628_);
  xor g_108099_(out[5], _015556_, _015629_);
  xor g_108100_(_002331_, _015556_, _015631_);
  and g_108101_(out[21], _015567_, _015632_);
  xor g_108102_(out[21], _015567_, _015633_);
  xor g_108103_(_002463_, _015567_, _015634_);
  and g_108104_(_015631_, _015633_, _015635_);
  or g_108105_(_015629_, _015634_, _015636_);
  and g_108106_(_015627_, _015636_, _015637_);
  or g_108107_(_015626_, _015635_, _015638_);
  and g_108108_(_015625_, _015637_, _015639_);
  or g_108109_(_015624_, _015638_, _015640_);
  and g_108110_(_015629_, _015634_, _015642_);
  or g_108111_(_015631_, _015633_, _015643_);
  xor g_108112_(out[6], _015558_, _015644_);
  xor g_108113_(_002320_, _015558_, _015645_);
  xor g_108114_(out[22], _015569_, _015646_);
  xor g_108115_(_002452_, _015569_, _015647_);
  and g_108116_(_015644_, _015647_, _015648_);
  or g_108117_(_015645_, _015646_, _015649_);
  and g_108118_(_015643_, _015649_, _015650_);
  or g_108119_(_015642_, _015648_, _015651_);
  and g_108120_(_015640_, _015650_, _015653_);
  or g_108121_(_015639_, _015651_, _015654_);
  and g_108122_(_015645_, _015646_, _015655_);
  or g_108123_(_015644_, _015647_, _015656_);
  and g_108124_(_015592_, _015656_, _015657_);
  or g_108125_(_015591_, _015655_, _015658_);
  and g_108126_(_015654_, _015657_, _015659_);
  or g_108127_(_015653_, _015658_, _015660_);
  and g_108128_(_015585_, _015594_, _015661_);
  or g_108129_(_015584_, _015593_, _015662_);
  and g_108130_(_015660_, _015661_, _015664_);
  or g_108131_(_015659_, _015662_, _015665_);
  and g_108132_(_015580_, _015583_, _015666_);
  or g_108133_(_015581_, _015582_, _015667_);
  xor g_108134_(out[9], _015561_, _015668_);
  xor g_108135_(_002408_, _015561_, _015669_);
  xor g_108136_(out[25], _015572_, _015670_);
  xor g_108137_(_002540_, _015572_, _015671_);
  and g_108138_(_015668_, _015671_, _015672_);
  or g_108139_(_015669_, _015670_, _015673_);
  and g_108140_(_015667_, _015673_, _015675_);
  or g_108141_(_015666_, _015672_, _015676_);
  and g_108142_(_015665_, _015675_, _015677_);
  or g_108143_(_015664_, _015676_, _015678_);
  xor g_108144_(out[10], _015562_, _015679_);
  xor g_108145_(_002419_, _015562_, _015680_);
  xor g_108146_(out[26], _015573_, _015681_);
  xor g_108147_(_002551_, _015573_, _015682_);
  and g_108148_(_015679_, _015682_, _015683_);
  or g_108149_(_015680_, _015681_, _015684_);
  and g_108150_(_015669_, _015670_, _015686_);
  or g_108151_(_015668_, _015671_, _015687_);
  and g_108152_(_015684_, _015687_, _015688_);
  or g_108153_(_015683_, _015686_, _015689_);
  and g_108154_(_015678_, _015688_, _015690_);
  or g_108155_(_015677_, _015689_, _015691_);
  and g_108156_(_015565_, _015577_, _015692_);
  or g_108157_(_015566_, _015576_, _015693_);
  and g_108158_(_015680_, _015681_, _015694_);
  or g_108159_(_015679_, _015682_, _015695_);
  and g_108160_(_015693_, _015695_, _015697_);
  or g_108161_(_015692_, _015694_, _015698_);
  and g_108162_(_015691_, _015697_, _015699_);
  or g_108163_(_015690_, _015698_, _015700_);
  and g_108164_(_015579_, _015700_, _015701_);
  or g_108165_(_015578_, _015699_, _015702_);
  or g_108166_(out[1], _015701_, _015703_);
  or g_108167_(out[17], _015702_, _015704_);
  and g_108168_(_015703_, _015704_, _015705_);
  not g_108169_(_015705_, _015706_);
  and g_108170_(out[36], out[35], _015708_);
  or g_108171_(out[37], _015708_, _015709_);
  or g_108172_(out[38], _015709_, _015710_);
  or g_108173_(out[39], _015710_, _015711_);
  xor g_108174_(out[39], _015710_, _015712_);
  xor g_108175_(_002573_, _015710_, _015713_);
  or g_108176_(_015589_, _015702_, _015714_);
  or g_108177_(_015587_, _015701_, _015715_);
  and g_108178_(_015714_, _015715_, _015716_);
  not g_108179_(_015716_, _015717_);
  and g_108180_(_015713_, _015716_, _015719_);
  or g_108181_(_015712_, _015717_, _015720_);
  xor g_108182_(out[37], _015708_, _015721_);
  xor g_108183_(_002595_, _015708_, _015722_);
  and g_108184_(_015634_, _015701_, _015723_);
  or g_108185_(_015633_, _015702_, _015724_);
  and g_108186_(_015631_, _015702_, _015725_);
  or g_108187_(_015629_, _015701_, _015726_);
  and g_108188_(_015724_, _015726_, _015727_);
  or g_108189_(_015723_, _015725_, _015728_);
  and g_108190_(_015722_, _015727_, _015730_);
  or g_108191_(_015721_, _015728_, _015731_);
  xor g_108192_(out[38], _015709_, _015732_);
  not g_108193_(_015732_, _015733_);
  or g_108194_(_015647_, _015702_, _015734_);
  or g_108195_(_015645_, _015701_, _015735_);
  and g_108196_(_015734_, _015735_, _015736_);
  not g_108197_(_015736_, _015737_);
  and g_108198_(_015732_, _015736_, _015738_);
  not g_108199_(_015738_, _015739_);
  and g_108200_(_015712_, _015717_, _015741_);
  or g_108201_(_015713_, _015716_, _015742_);
  and g_108202_(_015739_, _015742_, _015743_);
  or g_108203_(_015738_, _015741_, _015744_);
  and g_108204_(_015681_, _015701_, _015745_);
  or g_108205_(_015682_, _015702_, _015746_);
  and g_108206_(_015679_, _015702_, _015747_);
  or g_108207_(_015680_, _015701_, _015748_);
  and g_108208_(_015746_, _015748_, _015749_);
  or g_108209_(_015745_, _015747_, _015750_);
  or g_108210_(out[40], _015711_, _015752_);
  and g_108211_(out[41], _015752_, _015753_);
  or g_108212_(out[42], _015753_, _015754_);
  xor g_108213_(out[42], _015753_, _015755_);
  not g_108214_(_015755_, _015756_);
  and g_108215_(_015749_, _015755_, _015757_);
  or g_108216_(_015750_, _015756_, _015758_);
  and g_108217_(_015565_, _015576_, _015759_);
  or g_108218_(_015566_, _015577_, _015760_);
  xor g_108219_(out[43], _015754_, _015761_);
  xor g_108220_(_002562_, _015754_, _015763_);
  and g_108221_(_015759_, _015763_, _015764_);
  or g_108222_(_015760_, _015761_, _015765_);
  and g_108223_(_015760_, _015761_, _015766_);
  or g_108224_(_015759_, _015763_, _015767_);
  and g_108225_(_015765_, _015767_, _015768_);
  or g_108226_(_015764_, _015766_, _015769_);
  xor g_108227_(_015749_, _015755_, _015770_);
  xor g_108228_(_015750_, _015755_, _015771_);
  and g_108229_(_015768_, _015770_, _015772_);
  or g_108230_(_015769_, _015771_, _015774_);
  xor g_108231_(out[40], _015711_, _015775_);
  xor g_108232_(_002661_, _015711_, _015776_);
  and g_108233_(_015581_, _015701_, _015777_);
  or g_108234_(_015580_, _015702_, _015778_);
  and g_108235_(_015583_, _015702_, _015779_);
  or g_108236_(_015582_, _015701_, _015780_);
  and g_108237_(_015778_, _015780_, _015781_);
  or g_108238_(_015777_, _015779_, _015782_);
  and g_108239_(_015776_, _015781_, _015783_);
  or g_108240_(_015775_, _015782_, _015785_);
  xor g_108241_(out[41], _015752_, _015786_);
  xor g_108242_(_002672_, _015752_, _015787_);
  and g_108243_(_015670_, _015701_, _015788_);
  or g_108244_(_015671_, _015702_, _015789_);
  and g_108245_(_015668_, _015702_, _015790_);
  or g_108246_(_015669_, _015701_, _015791_);
  and g_108247_(_015789_, _015791_, _015792_);
  or g_108248_(_015788_, _015790_, _015793_);
  and g_108249_(_015786_, _015792_, _015794_);
  or g_108250_(_015787_, _015793_, _015796_);
  and g_108251_(_015785_, _015796_, _015797_);
  or g_108252_(_015783_, _015794_, _015798_);
  and g_108253_(_015787_, _015793_, _015799_);
  or g_108254_(_015786_, _015792_, _015800_);
  and g_108255_(_015775_, _015782_, _015801_);
  or g_108256_(_015776_, _015781_, _015802_);
  and g_108257_(_015800_, _015802_, _015803_);
  or g_108258_(_015799_, _015801_, _015804_);
  and g_108259_(_015797_, _015803_, _015805_);
  or g_108260_(_015798_, _015804_, _015807_);
  and g_108261_(_015772_, _015805_, _015808_);
  or g_108262_(_015774_, _015807_, _015809_);
  and g_108263_(_015721_, _015728_, _015810_);
  or g_108264_(_015722_, _015727_, _015811_);
  xor g_108265_(out[36], out[35], _015812_);
  xor g_108266_(_002606_, out[35], _015813_);
  and g_108267_(_015615_, _015701_, _015814_);
  or g_108268_(_015616_, _015702_, _015815_);
  and g_108269_(_015613_, _015702_, _015816_);
  or g_108270_(_015614_, _015701_, _015818_);
  and g_108271_(_015815_, _015818_, _015819_);
  or g_108272_(_015814_, _015816_, _015820_);
  and g_108273_(_015813_, _015820_, _015821_);
  or g_108274_(_015812_, _015819_, _015822_);
  and g_108275_(_015811_, _015822_, _015823_);
  or g_108276_(_015810_, _015821_, _015824_);
  and g_108277_(_015812_, _015819_, _015825_);
  or g_108278_(_015813_, _015820_, _015826_);
  xor g_108279_(_015732_, _015736_, _015827_);
  xor g_108280_(_015733_, _015736_, _015829_);
  and g_108281_(_015720_, _015742_, _015830_);
  or g_108282_(_015719_, _015741_, _015831_);
  and g_108283_(_015827_, _015830_, _015832_);
  or g_108284_(_015829_, _015831_, _015833_);
  and g_108285_(_015731_, _015826_, _015834_);
  or g_108286_(_015730_, _015825_, _015835_);
  and g_108287_(_015823_, _015834_, _015836_);
  or g_108288_(_015824_, _015835_, _015837_);
  and g_108289_(_015808_, _015836_, _015838_);
  or g_108290_(_015809_, _015837_, _015840_);
  and g_108291_(_015832_, _015838_, _015841_);
  or g_108292_(_015833_, _015840_, _015842_);
  and g_108293_(out[19], _015701_, _015843_);
  and g_108294_(out[3], _015702_, _015844_);
  or g_108295_(_015843_, _015844_, _015845_);
  not g_108296_(_015845_, _015846_);
  or g_108297_(_002650_, _015845_, _015847_);
  not g_108298_(_015847_, _015848_);
  or g_108299_(out[2], _015701_, _015849_);
  or g_108300_(out[18], _015702_, _015851_);
  and g_108301_(_015849_, _015851_, _015852_);
  not g_108302_(_015852_, _015853_);
  and g_108303_(out[34], _015853_, _015854_);
  or g_108304_(_015848_, _015854_, _015855_);
  or g_108305_(out[35], _015846_, _015856_);
  not g_108306_(_015856_, _015857_);
  and g_108307_(_002639_, _015852_, _015858_);
  or g_108308_(out[34], _015853_, _015859_);
  or g_108309_(_015857_, _015858_, _015860_);
  or g_108310_(_015855_, _015860_, _015862_);
  not g_108311_(_015862_, _015863_);
  and g_108312_(_002364_, _015702_, _015864_);
  or g_108313_(out[0], _015701_, _015865_);
  and g_108314_(_002496_, _015701_, _015866_);
  or g_108315_(out[16], _015702_, _015867_);
  and g_108316_(_015865_, _015867_, _015868_);
  or g_108317_(_015864_, _015866_, _015869_);
  and g_108318_(out[32], _015869_, _015870_);
  or g_108319_(_002628_, _015868_, _015871_);
  and g_108320_(_002617_, _015705_, _015873_);
  or g_108321_(out[33], _015706_, _015874_);
  xor g_108322_(_002617_, _015705_, _015875_);
  xor g_108323_(out[33], _015705_, _015876_);
  and g_108324_(_015871_, _015875_, _015877_);
  or g_108325_(_015870_, _015876_, _015878_);
  and g_108326_(_002628_, _015868_, _015879_);
  or g_108327_(_015878_, _015879_, _015880_);
  or g_108328_(_015862_, _015880_, _015881_);
  not g_108329_(_015881_, _015882_);
  and g_108330_(_015841_, _015882_, _015884_);
  or g_108331_(_015842_, _015881_, _015885_);
  and g_108332_(_015874_, _015878_, _015886_);
  or g_108333_(_015873_, _015877_, _015887_);
  and g_108334_(_015863_, _015887_, _015888_);
  or g_108335_(_015862_, _015886_, _015889_);
  and g_108336_(_015856_, _015858_, _015890_);
  or g_108337_(_015857_, _015859_, _015891_);
  and g_108338_(_015847_, _015891_, _015892_);
  or g_108339_(_015848_, _015890_, _015893_);
  and g_108340_(_015889_, _015892_, _015895_);
  or g_108341_(_015888_, _015893_, _015896_);
  and g_108342_(_015841_, _015896_, _015897_);
  or g_108343_(_015842_, _015895_, _015898_);
  and g_108344_(_015824_, _015832_, _015899_);
  or g_108345_(_015823_, _015833_, _015900_);
  and g_108346_(_015731_, _015899_, _015901_);
  or g_108347_(_015730_, _015900_, _015902_);
  and g_108348_(_015720_, _015744_, _015903_);
  or g_108349_(_015719_, _015743_, _015904_);
  and g_108350_(_015902_, _015904_, _015906_);
  or g_108351_(_015901_, _015903_, _015907_);
  and g_108352_(_015808_, _015907_, _015908_);
  or g_108353_(_015809_, _015906_, _015909_);
  and g_108354_(_015757_, _015767_, _015910_);
  or g_108355_(_015758_, _015766_, _015911_);
  and g_108356_(_015765_, _015911_, _015912_);
  or g_108357_(_015764_, _015910_, _015913_);
  and g_108358_(_015772_, _015804_, _015914_);
  or g_108359_(_015774_, _015803_, _015915_);
  and g_108360_(_015796_, _015914_, _015917_);
  or g_108361_(_015794_, _015915_, _015918_);
  and g_108362_(_015912_, _015918_, _015919_);
  or g_108363_(_015913_, _015917_, _015920_);
  and g_108364_(_015909_, _015919_, _015921_);
  or g_108365_(_015908_, _015920_, _015922_);
  and g_108366_(_015898_, _015921_, _015923_);
  or g_108367_(_015897_, _015922_, _015924_);
  and g_108368_(_015885_, _015924_, _015925_);
  or g_108369_(_015884_, _015923_, _015926_);
  or g_108370_(_015705_, _015925_, _015928_);
  or g_108371_(out[33], _015926_, _015929_);
  and g_108372_(_015928_, _015929_, _015930_);
  not g_108373_(_015930_, _015931_);
  or g_108374_(_015852_, _015925_, _015932_);
  or g_108375_(out[34], _015926_, _015933_);
  and g_108376_(_015932_, _015933_, _015934_);
  not g_108377_(_015934_, _015935_);
  and g_108378_(_002771_, _015934_, _015936_);
  or g_108379_(out[50], _015935_, _015937_);
  and g_108380_(out[35], _015925_, _015939_);
  or g_108381_(_002650_, _015926_, _015940_);
  and g_108382_(_015845_, _015926_, _015941_);
  or g_108383_(_015846_, _015925_, _015942_);
  and g_108384_(_015940_, _015942_, _015943_);
  or g_108385_(_015939_, _015941_, _015944_);
  or g_108386_(_002782_, _015944_, _015945_);
  not g_108387_(_015945_, _015946_);
  and g_108388_(_015937_, _015945_, _015947_);
  or g_108389_(_015936_, _015946_, _015948_);
  and g_108390_(out[50], _015935_, _015950_);
  or g_108391_(out[51], _015943_, _015951_);
  not g_108392_(_015951_, _015952_);
  or g_108393_(_015950_, _015952_, _015953_);
  or g_108394_(_015948_, _015953_, _015954_);
  not g_108395_(_015954_, _015955_);
  and g_108396_(_002749_, _015930_, _015956_);
  or g_108397_(out[49], _015931_, _015957_);
  and g_108398_(_015869_, _015926_, _015958_);
  or g_108399_(_015868_, _015925_, _015959_);
  and g_108400_(_002628_, _015925_, _015961_);
  or g_108401_(out[32], _015926_, _015962_);
  and g_108402_(_015959_, _015962_, _015963_);
  or g_108403_(_015958_, _015961_, _015964_);
  and g_108404_(out[48], _015964_, _015965_);
  or g_108405_(_002760_, _015963_, _015966_);
  xor g_108406_(_002749_, _015930_, _015967_);
  xor g_108407_(out[49], _015930_, _015968_);
  and g_108408_(_015966_, _015967_, _015969_);
  or g_108409_(_015965_, _015968_, _015970_);
  and g_108410_(_015957_, _015970_, _015972_);
  or g_108411_(_015956_, _015969_, _015973_);
  and g_108412_(_015955_, _015973_, _015974_);
  or g_108413_(_015954_, _015972_, _015975_);
  and g_108414_(_015948_, _015951_, _015976_);
  or g_108415_(_015947_, _015952_, _015977_);
  and g_108416_(_015975_, _015977_, _015978_);
  or g_108417_(_015974_, _015976_, _015979_);
  and g_108418_(_015755_, _015925_, _015980_);
  or g_108419_(_015756_, _015926_, _015981_);
  and g_108420_(_015750_, _015926_, _015983_);
  or g_108421_(_015749_, _015925_, _015984_);
  and g_108422_(_015981_, _015984_, _015985_);
  or g_108423_(_015980_, _015983_, _015986_);
  and g_108424_(out[52], out[51], _015987_);
  or g_108425_(out[53], _015987_, _015988_);
  or g_108426_(out[54], _015988_, _015989_);
  or g_108427_(out[55], _015989_, _015990_);
  or g_108428_(out[56], _015990_, _015991_);
  and g_108429_(out[57], _015991_, _015992_);
  or g_108430_(out[58], _015992_, _015994_);
  xor g_108431_(out[58], _015992_, _015995_);
  xor g_108432_(_002815_, _015992_, _015996_);
  and g_108433_(_015985_, _015995_, _015997_);
  or g_108434_(_015986_, _015996_, _015998_);
  and g_108435_(_015759_, _015761_, _015999_);
  or g_108436_(_015760_, _015763_, _016000_);
  xor g_108437_(out[59], _015994_, _016001_);
  xor g_108438_(_002694_, _015994_, _016002_);
  and g_108439_(_015999_, _016002_, _016003_);
  or g_108440_(_016000_, _016001_, _016005_);
  and g_108441_(_015998_, _016005_, _016006_);
  or g_108442_(_015997_, _016003_, _016007_);
  and g_108443_(_016000_, _016001_, _016008_);
  or g_108444_(_015999_, _016002_, _016009_);
  and g_108445_(_015986_, _015996_, _016010_);
  or g_108446_(_015985_, _015995_, _016011_);
  and g_108447_(_016009_, _016011_, _016012_);
  or g_108448_(_016008_, _016010_, _016013_);
  xor g_108449_(out[57], _015991_, _016014_);
  xor g_108450_(_002804_, _015991_, _016016_);
  and g_108451_(_015786_, _015925_, _016017_);
  or g_108452_(_015787_, _015926_, _016018_);
  and g_108453_(_015793_, _015926_, _016019_);
  or g_108454_(_015792_, _015925_, _016020_);
  and g_108455_(_016018_, _016020_, _016021_);
  or g_108456_(_016017_, _016019_, _016022_);
  and g_108457_(_016014_, _016021_, _016023_);
  or g_108458_(_016016_, _016022_, _016024_);
  xor g_108459_(out[56], _015990_, _016025_);
  xor g_108460_(_002793_, _015990_, _016027_);
  and g_108461_(_015776_, _015925_, _016028_);
  or g_108462_(_015775_, _015926_, _016029_);
  and g_108463_(_015782_, _015926_, _016030_);
  or g_108464_(_015781_, _015925_, _016031_);
  and g_108465_(_016029_, _016031_, _016032_);
  or g_108466_(_016028_, _016030_, _016033_);
  and g_108467_(_016025_, _016033_, _016034_);
  or g_108468_(_016027_, _016032_, _016035_);
  and g_108469_(_016016_, _016022_, _016036_);
  or g_108470_(_016014_, _016021_, _016038_);
  and g_108471_(_016035_, _016038_, _016039_);
  or g_108472_(_016034_, _016036_, _016040_);
  and g_108473_(_016027_, _016032_, _016041_);
  or g_108474_(_016025_, _016033_, _016042_);
  and g_108475_(_016006_, _016012_, _016043_);
  or g_108476_(_016007_, _016013_, _016044_);
  and g_108477_(_016024_, _016042_, _016045_);
  or g_108478_(_016023_, _016041_, _016046_);
  and g_108479_(_016039_, _016045_, _016047_);
  or g_108480_(_016040_, _016046_, _016049_);
  and g_108481_(_016043_, _016047_, _016050_);
  or g_108482_(_016044_, _016049_, _016051_);
  xor g_108483_(out[55], _015989_, _016052_);
  not g_108484_(_016052_, _016053_);
  and g_108485_(_015713_, _015925_, _016054_);
  or g_108486_(_015712_, _015926_, _016055_);
  and g_108487_(_015717_, _015926_, _016056_);
  or g_108488_(_015716_, _015925_, _016057_);
  and g_108489_(_016055_, _016057_, _016058_);
  or g_108490_(_016054_, _016056_, _016060_);
  and g_108491_(_016052_, _016060_, _016061_);
  or g_108492_(_016053_, _016058_, _016062_);
  xor g_108493_(out[54], _015988_, _016063_);
  xor g_108494_(_002716_, _015988_, _016064_);
  and g_108495_(_015732_, _015925_, _016065_);
  or g_108496_(_015733_, _015926_, _016066_);
  and g_108497_(_015737_, _015926_, _016067_);
  or g_108498_(_015736_, _015925_, _016068_);
  and g_108499_(_016066_, _016068_, _016069_);
  or g_108500_(_016065_, _016067_, _016071_);
  and g_108501_(_016063_, _016069_, _016072_);
  or g_108502_(_016064_, _016071_, _016073_);
  and g_108503_(_016062_, _016073_, _016074_);
  or g_108504_(_016061_, _016072_, _016075_);
  and g_108505_(_016053_, _016058_, _016076_);
  or g_108506_(_016052_, _016060_, _016077_);
  and g_108507_(_016064_, _016071_, _016078_);
  or g_108508_(_016063_, _016069_, _016079_);
  and g_108509_(_016077_, _016079_, _016080_);
  or g_108510_(_016076_, _016078_, _016082_);
  and g_108511_(_016074_, _016080_, _016083_);
  or g_108512_(_016075_, _016082_, _016084_);
  xor g_108513_(out[52], out[51], _016085_);
  xor g_108514_(_002738_, out[51], _016086_);
  and g_108515_(_015812_, _015925_, _016087_);
  or g_108516_(_015813_, _015926_, _016088_);
  and g_108517_(_015820_, _015926_, _016089_);
  or g_108518_(_015819_, _015925_, _016090_);
  and g_108519_(_016088_, _016090_, _016091_);
  or g_108520_(_016087_, _016089_, _016093_);
  and g_108521_(_016086_, _016093_, _016094_);
  or g_108522_(_016085_, _016091_, _016095_);
  xor g_108523_(out[53], _015987_, _016096_);
  xor g_108524_(_002727_, _015987_, _016097_);
  and g_108525_(_015722_, _015925_, _016098_);
  or g_108526_(_015721_, _015926_, _016099_);
  and g_108527_(_015728_, _015926_, _016100_);
  or g_108528_(_015727_, _015925_, _016101_);
  and g_108529_(_016099_, _016101_, _016102_);
  or g_108530_(_016098_, _016100_, _016104_);
  and g_108531_(_016096_, _016104_, _016105_);
  or g_108532_(_016097_, _016102_, _016106_);
  and g_108533_(_016095_, _016106_, _016107_);
  or g_108534_(_016094_, _016105_, _016108_);
  and g_108535_(_016097_, _016102_, _016109_);
  or g_108536_(_016096_, _016104_, _016110_);
  and g_108537_(_016085_, _016091_, _016111_);
  or g_108538_(_016086_, _016093_, _016112_);
  and g_108539_(_016110_, _016112_, _016113_);
  or g_108540_(_016109_, _016111_, _016115_);
  and g_108541_(_016107_, _016113_, _016116_);
  or g_108542_(_016108_, _016115_, _016117_);
  and g_108543_(_016083_, _016116_, _016118_);
  or g_108544_(_016084_, _016117_, _016119_);
  and g_108545_(_016050_, _016118_, _016120_);
  or g_108546_(_016051_, _016119_, _016121_);
  and g_108547_(_015979_, _016120_, _016122_);
  or g_108548_(_015978_, _016121_, _016123_);
  and g_108549_(_016108_, _016110_, _016124_);
  or g_108550_(_016107_, _016109_, _016126_);
  and g_108551_(_016083_, _016124_, _016127_);
  or g_108552_(_016084_, _016126_, _016128_);
  or g_108553_(_016074_, _016076_, _016129_);
  not g_108554_(_016129_, _016130_);
  and g_108555_(_016128_, _016129_, _016131_);
  or g_108556_(_016127_, _016130_, _016132_);
  and g_108557_(_016050_, _016132_, _016133_);
  or g_108558_(_016051_, _016131_, _016134_);
  and g_108559_(_016007_, _016009_, _016135_);
  or g_108560_(_016006_, _016008_, _016137_);
  and g_108561_(_016024_, _016040_, _016138_);
  or g_108562_(_016023_, _016039_, _016139_);
  and g_108563_(_016043_, _016138_, _016140_);
  or g_108564_(_016044_, _016139_, _016141_);
  and g_108565_(_016137_, _016141_, _016142_);
  or g_108566_(_016135_, _016140_, _016143_);
  and g_108567_(_016134_, _016142_, _016144_);
  or g_108568_(_016133_, _016143_, _016145_);
  and g_108569_(_016123_, _016144_, _016146_);
  or g_108570_(_016122_, _016145_, _016148_);
  and g_108571_(_002760_, _015963_, _016149_);
  or g_108572_(_015954_, _015970_, _016150_);
  or g_108573_(_016149_, _016150_, _016151_);
  not g_108574_(_016151_, _016152_);
  and g_108575_(_016120_, _016152_, _016153_);
  or g_108576_(_016121_, _016151_, _016154_);
  and g_108577_(_016148_, _016154_, _016155_);
  or g_108578_(_016146_, _016153_, _016156_);
  and g_108579_(_015931_, _016156_, _016157_);
  or g_108580_(_015930_, _016155_, _016159_);
  and g_108581_(_002749_, _016155_, _016160_);
  or g_108582_(out[49], _016156_, _016161_);
  and g_108583_(_016159_, _016161_, _016162_);
  or g_108584_(_016157_, _016160_, _016163_);
  and g_108585_(out[68], out[67], _016164_);
  or g_108586_(out[69], _016164_, _016165_);
  or g_108587_(out[70], _016165_, _016166_);
  or g_108588_(out[71], _016166_, _016167_);
  or g_108589_(out[72], _016167_, _016168_);
  and g_108590_(out[73], _016168_, _016170_);
  or g_108591_(out[74], _016170_, _016171_);
  xor g_108592_(out[74], _016170_, _016172_);
  xor g_108593_(_002947_, _016170_, _016173_);
  and g_108594_(_015995_, _016155_, _016174_);
  or g_108595_(_015996_, _016156_, _016175_);
  and g_108596_(_015986_, _016156_, _016176_);
  not g_108597_(_016176_, _016177_);
  and g_108598_(_016175_, _016177_, _016178_);
  or g_108599_(_016174_, _016176_, _016179_);
  and g_108600_(_016172_, _016178_, _016181_);
  or g_108601_(_016173_, _016179_, _016182_);
  and g_108602_(_015999_, _016001_, _016183_);
  or g_108603_(_016000_, _016002_, _016184_);
  xor g_108604_(out[75], _016171_, _016185_);
  xor g_108605_(_002826_, _016171_, _016186_);
  and g_108606_(_016183_, _016186_, _016187_);
  or g_108607_(_016184_, _016185_, _016188_);
  and g_108608_(_016182_, _016188_, _016189_);
  or g_108609_(_016181_, _016187_, _016190_);
  and g_108610_(_016184_, _016185_, _016192_);
  or g_108611_(_016183_, _016186_, _016193_);
  and g_108612_(_016190_, _016193_, _016194_);
  or g_108613_(_016189_, _016192_, _016195_);
  xor g_108614_(out[73], _016168_, _016196_);
  xor g_108615_(_002936_, _016168_, _016197_);
  and g_108616_(_016014_, _016155_, _016198_);
  or g_108617_(_016016_, _016156_, _016199_);
  and g_108618_(_016022_, _016156_, _016200_);
  or g_108619_(_016021_, _016155_, _016201_);
  and g_108620_(_016199_, _016201_, _016203_);
  or g_108621_(_016198_, _016200_, _016204_);
  and g_108622_(_016197_, _016204_, _016205_);
  or g_108623_(_016196_, _016203_, _016206_);
  or g_108624_(_016025_, _016156_, _016207_);
  not g_108625_(_016207_, _016208_);
  and g_108626_(_016033_, _016156_, _016209_);
  or g_108627_(_016032_, _016155_, _016210_);
  and g_108628_(_016207_, _016210_, _016211_);
  or g_108629_(_016208_, _016209_, _016212_);
  xor g_108630_(out[72], _016167_, _016214_);
  xor g_108631_(_002925_, _016167_, _016215_);
  and g_108632_(_016212_, _016214_, _016216_);
  or g_108633_(_016211_, _016215_, _016217_);
  and g_108634_(_016206_, _016217_, _016218_);
  or g_108635_(_016205_, _016216_, _016219_);
  xor g_108636_(out[70], _016165_, _016220_);
  not g_108637_(_016220_, _016221_);
  and g_108638_(_016063_, _016155_, _016222_);
  or g_108639_(_016064_, _016156_, _016223_);
  and g_108640_(_016071_, _016156_, _016225_);
  or g_108641_(_016069_, _016155_, _016226_);
  and g_108642_(_016223_, _016226_, _016227_);
  or g_108643_(_016222_, _016225_, _016228_);
  and g_108644_(_016220_, _016227_, _016229_);
  not g_108645_(_016229_, _016230_);
  xor g_108646_(out[71], _016166_, _016231_);
  xor g_108647_(_002837_, _016166_, _016232_);
  or g_108648_(_016052_, _016156_, _016233_);
  or g_108649_(_016058_, _016155_, _016234_);
  and g_108650_(_016233_, _016234_, _016236_);
  or g_108651_(_016232_, _016236_, _016237_);
  and g_108652_(_016230_, _016237_, _016238_);
  and g_108653_(_016221_, _016228_, _016239_);
  xor g_108654_(out[69], _016164_, _016240_);
  xor g_108655_(_002859_, _016164_, _016241_);
  or g_108656_(_016096_, _016156_, _016242_);
  not g_108657_(_016242_, _016243_);
  and g_108658_(_016104_, _016156_, _016244_);
  or g_108659_(_016102_, _016155_, _016245_);
  and g_108660_(_016242_, _016245_, _016247_);
  or g_108661_(_016243_, _016244_, _016248_);
  and g_108662_(_016241_, _016247_, _016249_);
  or g_108663_(_016240_, _016248_, _016250_);
  or g_108664_(_016239_, _016249_, _016251_);
  and g_108665_(_016240_, _016248_, _016252_);
  or g_108666_(_016241_, _016247_, _016253_);
  xor g_108667_(out[68], out[67], _016254_);
  xor g_108668_(_002870_, out[67], _016255_);
  and g_108669_(_016085_, _016155_, _016256_);
  or g_108670_(_016086_, _016156_, _016258_);
  and g_108671_(_016093_, _016156_, _016259_);
  or g_108672_(_016091_, _016155_, _016260_);
  and g_108673_(_016258_, _016260_, _016261_);
  or g_108674_(_016256_, _016259_, _016262_);
  and g_108675_(_016255_, _016262_, _016263_);
  or g_108676_(_016254_, _016261_, _016264_);
  and g_108677_(_016253_, _016264_, _016265_);
  or g_108678_(_016252_, _016263_, _016266_);
  or g_108679_(_002782_, _016156_, _016267_);
  or g_108680_(_015943_, _016155_, _016269_);
  and g_108681_(_016267_, _016269_, _016270_);
  or g_108682_(out[67], _016270_, _016271_);
  and g_108683_(out[67], _016270_, _016272_);
  xor g_108684_(out[67], _016270_, _016273_);
  xor g_108685_(_002914_, _016270_, _016274_);
  or g_108686_(_015934_, _016155_, _016275_);
  or g_108687_(out[50], _016156_, _016276_);
  and g_108688_(_016275_, _016276_, _016277_);
  and g_108689_(_002903_, _016277_, _016278_);
  xor g_108690_(_002903_, _016277_, _016280_);
  xor g_108691_(out[66], _016277_, _016281_);
  and g_108692_(_016273_, _016280_, _016282_);
  or g_108693_(_016274_, _016281_, _016283_);
  or g_108694_(out[65], _016163_, _016284_);
  not g_108695_(_016284_, _016285_);
  and g_108696_(_015964_, _016156_, _016286_);
  or g_108697_(_015963_, _016155_, _016287_);
  and g_108698_(_002760_, _016155_, _016288_);
  or g_108699_(out[48], _016156_, _016289_);
  and g_108700_(_016287_, _016289_, _016291_);
  or g_108701_(_016286_, _016288_, _016292_);
  and g_108702_(out[64], _016292_, _016293_);
  or g_108703_(_002892_, _016291_, _016294_);
  and g_108704_(out[65], _016163_, _016295_);
  or g_108705_(_002881_, _016162_, _016296_);
  and g_108706_(_016294_, _016296_, _016297_);
  or g_108707_(_016293_, _016295_, _016298_);
  and g_108708_(_016284_, _016298_, _016299_);
  or g_108709_(_016285_, _016297_, _016300_);
  and g_108710_(_016282_, _016300_, _016302_);
  or g_108711_(_016283_, _016299_, _016303_);
  and g_108712_(_016271_, _016278_, _016304_);
  or g_108713_(_016272_, _016304_, _016305_);
  not g_108714_(_016305_, _016306_);
  and g_108715_(_016303_, _016306_, _016307_);
  or g_108716_(_016302_, _016305_, _016308_);
  and g_108717_(_016254_, _016261_, _016309_);
  or g_108718_(_016255_, _016262_, _016310_);
  or g_108719_(_016307_, _016309_, _016311_);
  and g_108720_(_016265_, _016311_, _016313_);
  or g_108721_(_016251_, _016313_, _016314_);
  and g_108722_(_016238_, _016314_, _016315_);
  and g_108723_(_016232_, _016236_, _016316_);
  and g_108724_(_016211_, _016215_, _016317_);
  or g_108725_(_016212_, _016214_, _016318_);
  or g_108726_(_016316_, _016317_, _016319_);
  or g_108727_(_016315_, _016319_, _016320_);
  xor g_108728_(_016220_, _016227_, _016321_);
  xor g_108729_(_016232_, _016236_, _016322_);
  and g_108730_(_016321_, _016322_, _016324_);
  and g_108731_(_016250_, _016310_, _016325_);
  and g_108732_(_016265_, _016325_, _016326_);
  and g_108733_(_016324_, _016326_, _016327_);
  and g_108734_(_016308_, _016327_, _016328_);
  and g_108735_(_016266_, _016324_, _016329_);
  and g_108736_(_016250_, _016329_, _016330_);
  or g_108737_(_016238_, _016316_, _016331_);
  not g_108738_(_016331_, _016332_);
  or g_108739_(_016330_, _016332_, _016333_);
  or g_108740_(_016328_, _016333_, _016335_);
  and g_108741_(_016218_, _016318_, _016336_);
  and g_108742_(_016335_, _016336_, _016337_);
  and g_108743_(_016218_, _016320_, _016338_);
  or g_108744_(_016219_, _016337_, _016339_);
  and g_108745_(_016173_, _016179_, _016340_);
  or g_108746_(_016172_, _016178_, _016341_);
  and g_108747_(_016193_, _016341_, _016342_);
  or g_108748_(_016192_, _016340_, _016343_);
  and g_108749_(_016189_, _016342_, _016344_);
  or g_108750_(_016190_, _016343_, _016346_);
  and g_108751_(_016196_, _016203_, _016347_);
  or g_108752_(_016197_, _016204_, _016348_);
  and g_108753_(_016344_, _016348_, _016349_);
  or g_108754_(_016346_, _016347_, _016350_);
  and g_108755_(_016339_, _016349_, _016351_);
  or g_108756_(_016338_, _016350_, _016352_);
  and g_108757_(_016195_, _016352_, _016353_);
  or g_108758_(_016194_, _016351_, _016354_);
  or g_108759_(out[64], _016292_, _016355_);
  and g_108760_(_016344_, _016355_, _016357_);
  and g_108761_(_016282_, _016348_, _016358_);
  and g_108762_(_016284_, _016297_, _016359_);
  and g_108763_(_016336_, _016359_, _016360_);
  and g_108764_(_016358_, _016360_, _016361_);
  and g_108765_(_016357_, _016361_, _016362_);
  and g_108766_(_016327_, _016362_, _016363_);
  not g_108767_(_016363_, _016364_);
  and g_108768_(_016354_, _016364_, _016365_);
  or g_108769_(_016353_, _016363_, _016366_);
  and g_108770_(_016163_, _016366_, _016368_);
  not g_108771_(_016368_, _016369_);
  or g_108772_(out[65], _016366_, _016370_);
  not g_108773_(_016370_, _016371_);
  and g_108774_(_016369_, _016370_, _016372_);
  or g_108775_(_016368_, _016371_, _016373_);
  and g_108776_(_016179_, _016366_, _016374_);
  or g_108777_(_016178_, _016365_, _016375_);
  and g_108778_(_016172_, _016365_, _016376_);
  or g_108779_(_016173_, _016366_, _016377_);
  and g_108780_(_016375_, _016377_, _016379_);
  or g_108781_(_016374_, _016376_, _016380_);
  and g_108782_(out[84], out[83], _016381_);
  or g_108783_(out[85], _016381_, _016382_);
  or g_108784_(out[86], _016382_, _016383_);
  or g_108785_(out[87], _016383_, _016384_);
  or g_108786_(out[88], _016384_, _016385_);
  and g_108787_(out[89], _016385_, _016386_);
  or g_108788_(out[90], _016386_, _016387_);
  xor g_108789_(out[90], _016386_, _016388_);
  xor g_108790_(_003079_, _016386_, _016390_);
  and g_108791_(_016379_, _016388_, _016391_);
  or g_108792_(_016380_, _016390_, _016392_);
  and g_108793_(_016183_, _016185_, _016393_);
  or g_108794_(_016184_, _016186_, _016394_);
  xor g_108795_(out[91], _016387_, _016395_);
  xor g_108796_(_002958_, _016387_, _016396_);
  and g_108797_(_016393_, _016396_, _016397_);
  or g_108798_(_016394_, _016395_, _016398_);
  and g_108799_(_016392_, _016398_, _016399_);
  or g_108800_(_016391_, _016397_, _016401_);
  and g_108801_(_016380_, _016390_, _016402_);
  or g_108802_(_016379_, _016388_, _016403_);
  and g_108803_(_016394_, _016395_, _016404_);
  or g_108804_(_016393_, _016396_, _016405_);
  xor g_108805_(out[89], _016385_, _016406_);
  xor g_108806_(_003068_, _016385_, _016407_);
  and g_108807_(_016204_, _016366_, _016408_);
  or g_108808_(_016203_, _016365_, _016409_);
  and g_108809_(_016196_, _016365_, _016410_);
  or g_108810_(_016197_, _016366_, _016412_);
  and g_108811_(_016409_, _016412_, _016413_);
  or g_108812_(_016408_, _016410_, _016414_);
  and g_108813_(_016406_, _016413_, _016415_);
  or g_108814_(_016407_, _016414_, _016416_);
  xor g_108815_(out[88], _016384_, _016417_);
  xor g_108816_(_003057_, _016384_, _016418_);
  and g_108817_(_016212_, _016366_, _016419_);
  or g_108818_(_016211_, _016365_, _016420_);
  and g_108819_(_016215_, _016365_, _016421_);
  or g_108820_(_016214_, _016366_, _016423_);
  and g_108821_(_016420_, _016423_, _016424_);
  or g_108822_(_016419_, _016421_, _016425_);
  and g_108823_(_016417_, _016425_, _016426_);
  or g_108824_(_016418_, _016424_, _016427_);
  and g_108825_(_016407_, _016414_, _016428_);
  or g_108826_(_016406_, _016413_, _016429_);
  and g_108827_(_016427_, _016429_, _016430_);
  or g_108828_(_016426_, _016428_, _016431_);
  and g_108829_(_016418_, _016424_, _016432_);
  or g_108830_(_016417_, _016425_, _016434_);
  and g_108831_(_016403_, _016405_, _016435_);
  or g_108832_(_016402_, _016404_, _016436_);
  and g_108833_(_016399_, _016435_, _016437_);
  or g_108834_(_016401_, _016436_, _016438_);
  and g_108835_(_016416_, _016434_, _016439_);
  or g_108836_(_016415_, _016432_, _016440_);
  and g_108837_(_016430_, _016439_, _016441_);
  or g_108838_(_016431_, _016440_, _016442_);
  and g_108839_(_016437_, _016441_, _016443_);
  or g_108840_(_016438_, _016442_, _016445_);
  xor g_108841_(out[86], _016382_, _016446_);
  not g_108842_(_016446_, _016447_);
  or g_108843_(_016227_, _016365_, _016448_);
  or g_108844_(_016221_, _016366_, _016449_);
  and g_108845_(_016448_, _016449_, _016450_);
  not g_108846_(_016450_, _016451_);
  and g_108847_(_016446_, _016450_, _016452_);
  not g_108848_(_016452_, _016453_);
  xor g_108849_(out[87], _016383_, _016454_);
  xor g_108850_(_002969_, _016383_, _016456_);
  or g_108851_(_016236_, _016365_, _016457_);
  or g_108852_(_016231_, _016366_, _016458_);
  and g_108853_(_016457_, _016458_, _016459_);
  not g_108854_(_016459_, _016460_);
  and g_108855_(_016454_, _016460_, _016461_);
  or g_108856_(_016456_, _016459_, _016462_);
  and g_108857_(_016453_, _016462_, _016463_);
  or g_108858_(_016452_, _016461_, _016464_);
  and g_108859_(_016447_, _016451_, _016465_);
  or g_108860_(_016446_, _016450_, _016467_);
  and g_108861_(_016456_, _016459_, _016468_);
  or g_108862_(_016454_, _016460_, _016469_);
  and g_108863_(_016467_, _016469_, _016470_);
  or g_108864_(_016465_, _016468_, _016471_);
  and g_108865_(_016463_, _016470_, _016472_);
  or g_108866_(_016464_, _016471_, _016473_);
  xor g_108867_(out[85], _016381_, _016474_);
  xor g_108868_(_002991_, _016381_, _016475_);
  and g_108869_(_016248_, _016366_, _016476_);
  or g_108870_(_016247_, _016365_, _016478_);
  and g_108871_(_016241_, _016365_, _016479_);
  or g_108872_(_016240_, _016366_, _016480_);
  and g_108873_(_016478_, _016480_, _016481_);
  or g_108874_(_016476_, _016479_, _016482_);
  and g_108875_(_016475_, _016481_, _016483_);
  or g_108876_(_016474_, _016482_, _016484_);
  xor g_108877_(out[84], out[83], _016485_);
  xor g_108878_(_003002_, out[83], _016486_);
  and g_108879_(_016254_, _016365_, _016487_);
  or g_108880_(_016255_, _016366_, _016489_);
  and g_108881_(_016262_, _016366_, _016490_);
  or g_108882_(_016261_, _016365_, _016491_);
  and g_108883_(_016489_, _016491_, _016492_);
  or g_108884_(_016487_, _016490_, _016493_);
  and g_108885_(_016485_, _016492_, _016494_);
  or g_108886_(_016486_, _016493_, _016495_);
  and g_108887_(_016484_, _016495_, _016496_);
  or g_108888_(_016483_, _016494_, _016497_);
  and g_108889_(_016474_, _016482_, _016498_);
  or g_108890_(_016475_, _016481_, _016500_);
  and g_108891_(_016486_, _016493_, _016501_);
  or g_108892_(_016485_, _016492_, _016502_);
  and g_108893_(_016500_, _016502_, _016503_);
  or g_108894_(_016498_, _016501_, _016504_);
  and g_108895_(_016472_, _016503_, _016505_);
  or g_108896_(_016473_, _016504_, _016506_);
  and g_108897_(_016443_, _016505_, _016507_);
  or g_108898_(_016445_, _016506_, _016508_);
  and g_108899_(_016496_, _016507_, _016509_);
  or g_108900_(_016497_, _016508_, _016511_);
  or g_108901_(_002914_, _016366_, _016512_);
  or g_108902_(_016270_, _016365_, _016513_);
  and g_108903_(_016512_, _016513_, _016514_);
  not g_108904_(_016514_, _016515_);
  and g_108905_(out[83], _016514_, _016516_);
  or g_108906_(_016277_, _016365_, _016517_);
  or g_108907_(out[66], _016366_, _016518_);
  and g_108908_(_016517_, _016518_, _016519_);
  not g_108909_(_016519_, _016520_);
  and g_108910_(_003035_, _016519_, _016522_);
  or g_108911_(out[83], _016514_, _016523_);
  xor g_108912_(out[83], _016514_, _016524_);
  xor g_108913_(_003046_, _016514_, _016525_);
  xor g_108914_(_003035_, _016519_, _016526_);
  xor g_108915_(out[82], _016519_, _016527_);
  and g_108916_(_016524_, _016526_, _016528_);
  or g_108917_(_016525_, _016527_, _016529_);
  and g_108918_(_003013_, _016372_, _016530_);
  or g_108919_(out[81], _016373_, _016531_);
  and g_108920_(_016522_, _016523_, _016533_);
  or g_108921_(_016516_, _016533_, _016534_);
  not g_108922_(_016534_, _016535_);
  and g_108923_(_016292_, _016366_, _016536_);
  not g_108924_(_016536_, _016537_);
  or g_108925_(out[64], _016366_, _016538_);
  not g_108926_(_016538_, _016539_);
  and g_108927_(_016537_, _016538_, _016540_);
  or g_108928_(_016536_, _016539_, _016541_);
  and g_108929_(out[80], _016541_, _016542_);
  or g_108930_(_003024_, _016540_, _016544_);
  xor g_108931_(_003013_, _016372_, _016545_);
  xor g_108932_(out[81], _016372_, _016546_);
  and g_108933_(_016544_, _016545_, _016547_);
  or g_108934_(_016542_, _016546_, _016548_);
  and g_108935_(_016528_, _016547_, _016549_);
  or g_108936_(_016529_, _016548_, _016550_);
  and g_108937_(_016531_, _016548_, _016551_);
  or g_108938_(_016530_, _016547_, _016552_);
  and g_108939_(_016528_, _016552_, _016553_);
  or g_108940_(_016529_, _016551_, _016555_);
  and g_108941_(_016535_, _016555_, _016556_);
  or g_108942_(_016534_, _016553_, _016557_);
  and g_108943_(_016509_, _016557_, _016558_);
  or g_108944_(_016511_, _016556_, _016559_);
  and g_108945_(_016464_, _016469_, _016560_);
  or g_108946_(_016463_, _016468_, _016561_);
  and g_108947_(_016484_, _016504_, _016562_);
  or g_108948_(_016483_, _016503_, _016563_);
  and g_108949_(_016472_, _016562_, _016564_);
  or g_108950_(_016473_, _016563_, _016566_);
  and g_108951_(_016561_, _016566_, _016567_);
  or g_108952_(_016560_, _016564_, _016568_);
  and g_108953_(_016443_, _016568_, _016569_);
  or g_108954_(_016445_, _016567_, _016570_);
  and g_108955_(_016416_, _016431_, _016571_);
  or g_108956_(_016415_, _016430_, _016572_);
  and g_108957_(_016437_, _016571_, _016573_);
  or g_108958_(_016438_, _016572_, _016574_);
  and g_108959_(_016401_, _016405_, _016575_);
  or g_108960_(_016399_, _016404_, _016577_);
  and g_108961_(_016574_, _016577_, _016578_);
  or g_108962_(_016573_, _016575_, _016579_);
  and g_108963_(_016570_, _016578_, _016580_);
  or g_108964_(_016569_, _016579_, _016581_);
  and g_108965_(_016559_, _016580_, _016582_);
  or g_108966_(_016558_, _016581_, _016583_);
  and g_108967_(_003024_, _016540_, _016584_);
  or g_108968_(out[80], _016541_, _016585_);
  and g_108969_(_016549_, _016585_, _016586_);
  or g_108970_(_016550_, _016584_, _016588_);
  and g_108971_(_016509_, _016586_, _016589_);
  or g_108972_(_016511_, _016588_, _016590_);
  and g_108973_(_016583_, _016590_, _016591_);
  or g_108974_(_016582_, _016589_, _016592_);
  and g_108975_(_016373_, _016592_, _016593_);
  or g_108976_(_016372_, _016591_, _016594_);
  and g_108977_(_003013_, _016591_, _016595_);
  or g_108978_(out[81], _016592_, _016596_);
  and g_108979_(_016594_, _016596_, _016597_);
  or g_108980_(_016593_, _016595_, _016599_);
  and g_108981_(_016393_, _016395_, _016600_);
  or g_108982_(_016394_, _016396_, _016601_);
  and g_108983_(out[100], out[99], _016602_);
  or g_108984_(out[101], _016602_, _016603_);
  or g_108985_(out[102], _016603_, _016604_);
  or g_108986_(out[103], _016604_, _016605_);
  or g_108987_(out[104], _016605_, _016606_);
  and g_108988_(out[105], _016606_, _016607_);
  or g_108989_(out[106], _016607_, _016608_);
  xor g_108990_(out[107], _016608_, _016610_);
  xor g_108991_(_003090_, _016608_, _016611_);
  and g_108992_(_016600_, _016611_, _016612_);
  or g_108993_(_016601_, _016610_, _016613_);
  xor g_108994_(out[106], _016607_, _016614_);
  xor g_108995_(_003211_, _016607_, _016615_);
  or g_108996_(_016390_, _016592_, _016616_);
  not g_108997_(_016616_, _016617_);
  and g_108998_(_016380_, _016592_, _016618_);
  not g_108999_(_016618_, _016619_);
  and g_109000_(_016616_, _016619_, _016621_);
  or g_109001_(_016617_, _016618_, _016622_);
  and g_109002_(_016614_, _016621_, _016623_);
  or g_109003_(_016615_, _016622_, _016624_);
  and g_109004_(_016613_, _016624_, _016625_);
  or g_109005_(_016612_, _016623_, _016626_);
  and g_109006_(_016601_, _016610_, _016627_);
  or g_109007_(_016600_, _016611_, _016628_);
  and g_109008_(_016615_, _016622_, _016629_);
  or g_109009_(_016614_, _016621_, _016630_);
  and g_109010_(_016628_, _016630_, _016632_);
  or g_109011_(_016627_, _016629_, _016633_);
  and g_109012_(_016625_, _016632_, _016634_);
  or g_109013_(_016626_, _016633_, _016635_);
  xor g_109014_(out[105], _016606_, _016636_);
  xor g_109015_(_003200_, _016606_, _016637_);
  or g_109016_(_016407_, _016592_, _016638_);
  not g_109017_(_016638_, _016639_);
  and g_109018_(_016414_, _016592_, _016640_);
  not g_109019_(_016640_, _016641_);
  and g_109020_(_016638_, _016641_, _016643_);
  or g_109021_(_016639_, _016640_, _016644_);
  and g_109022_(_016637_, _016644_, _016645_);
  or g_109023_(_016636_, _016643_, _016646_);
  xor g_109024_(out[104], _016605_, _016647_);
  xor g_109025_(_003189_, _016605_, _016648_);
  or g_109026_(_016417_, _016592_, _016649_);
  not g_109027_(_016649_, _016650_);
  and g_109028_(_016425_, _016592_, _016651_);
  not g_109029_(_016651_, _016652_);
  and g_109030_(_016649_, _016652_, _016654_);
  or g_109031_(_016650_, _016651_, _016655_);
  and g_109032_(_016647_, _016655_, _016656_);
  or g_109033_(_016648_, _016654_, _016657_);
  and g_109034_(_016646_, _016657_, _016658_);
  or g_109035_(_016645_, _016656_, _016659_);
  and g_109036_(_016636_, _016643_, _016660_);
  or g_109037_(_016637_, _016644_, _016661_);
  and g_109038_(_016648_, _016654_, _016662_);
  or g_109039_(_016647_, _016655_, _016663_);
  and g_109040_(_016661_, _016663_, _016665_);
  or g_109041_(_016660_, _016662_, _016666_);
  and g_109042_(_016658_, _016665_, _016667_);
  or g_109043_(_016659_, _016666_, _016668_);
  and g_109044_(_016634_, _016667_, _016669_);
  or g_109045_(_016635_, _016668_, _016670_);
  xor g_109046_(out[102], _016603_, _016671_);
  xor g_109047_(_003112_, _016603_, _016672_);
  and g_109048_(_016446_, _016591_, _016673_);
  or g_109049_(_016447_, _016592_, _016674_);
  and g_109050_(_016451_, _016592_, _016676_);
  or g_109051_(_016450_, _016591_, _016677_);
  and g_109052_(_016674_, _016677_, _016678_);
  or g_109053_(_016673_, _016676_, _016679_);
  and g_109054_(_016671_, _016678_, _016680_);
  or g_109055_(_016672_, _016679_, _016681_);
  xor g_109056_(out[103], _016604_, _016682_);
  xor g_109057_(_003101_, _016604_, _016683_);
  and g_109058_(_016456_, _016591_, _016684_);
  or g_109059_(_016454_, _016592_, _016685_);
  and g_109060_(_016460_, _016592_, _016687_);
  or g_109061_(_016459_, _016591_, _016688_);
  and g_109062_(_016685_, _016688_, _016689_);
  or g_109063_(_016684_, _016687_, _016690_);
  and g_109064_(_016682_, _016690_, _016691_);
  or g_109065_(_016683_, _016689_, _016692_);
  and g_109066_(_016681_, _016692_, _016693_);
  or g_109067_(_016680_, _016691_, _016694_);
  xor g_109068_(out[101], _016602_, _016695_);
  xor g_109069_(_003123_, _016602_, _016696_);
  or g_109070_(_016474_, _016592_, _016698_);
  not g_109071_(_016698_, _016699_);
  and g_109072_(_016482_, _016592_, _016700_);
  not g_109073_(_016700_, _016701_);
  and g_109074_(_016698_, _016701_, _016702_);
  or g_109075_(_016699_, _016700_, _016703_);
  and g_109076_(_016696_, _016702_, _016704_);
  or g_109077_(_016695_, _016703_, _016705_);
  and g_109078_(_016683_, _016689_, _016706_);
  or g_109079_(_016682_, _016690_, _016707_);
  and g_109080_(_016672_, _016679_, _016709_);
  or g_109081_(_016671_, _016678_, _016710_);
  xor g_109082_(out[100], out[99], _016711_);
  xor g_109083_(_003134_, out[99], _016712_);
  or g_109084_(_016486_, _016592_, _016713_);
  not g_109085_(_016713_, _016714_);
  and g_109086_(_016493_, _016592_, _016715_);
  not g_109087_(_016715_, _016716_);
  and g_109088_(_016713_, _016716_, _016717_);
  or g_109089_(_016714_, _016715_, _016718_);
  and g_109090_(_016712_, _016718_, _016720_);
  or g_109091_(_016711_, _016717_, _016721_);
  and g_109092_(_016695_, _016703_, _016722_);
  or g_109093_(_016696_, _016702_, _016723_);
  and g_109094_(_016721_, _016723_, _016724_);
  or g_109095_(_016720_, _016722_, _016725_);
  and g_109096_(_016711_, _016717_, _016726_);
  or g_109097_(_016712_, _016718_, _016727_);
  and g_109098_(_016681_, _016707_, _016728_);
  or g_109099_(_016680_, _016706_, _016729_);
  and g_109100_(_016692_, _016710_, _016731_);
  or g_109101_(_016691_, _016709_, _016732_);
  and g_109102_(_016728_, _016731_, _016733_);
  or g_109103_(_016729_, _016732_, _016734_);
  and g_109104_(_016705_, _016727_, _016735_);
  or g_109105_(_016704_, _016726_, _016736_);
  and g_109106_(_016724_, _016735_, _016737_);
  or g_109107_(_016725_, _016736_, _016738_);
  and g_109108_(_016733_, _016737_, _016739_);
  or g_109109_(_016734_, _016738_, _016740_);
  and g_109110_(out[83], _016591_, _016742_);
  or g_109111_(_003046_, _016592_, _016743_);
  and g_109112_(_016515_, _016592_, _016744_);
  or g_109113_(_016514_, _016591_, _016745_);
  and g_109114_(_016743_, _016745_, _016746_);
  or g_109115_(_016742_, _016744_, _016747_);
  or g_109116_(out[99], _016746_, _016748_);
  not g_109117_(_016748_, _016749_);
  or g_109118_(_003178_, _016747_, _016750_);
  not g_109119_(_016750_, _016751_);
  and g_109120_(_016748_, _016750_, _016753_);
  or g_109121_(_016749_, _016751_, _016754_);
  and g_109122_(_016520_, _016592_, _016755_);
  or g_109123_(_016519_, _016591_, _016756_);
  or g_109124_(out[82], _016592_, _016757_);
  not g_109125_(_016757_, _016758_);
  and g_109126_(_016756_, _016757_, _016759_);
  or g_109127_(_016755_, _016758_, _016760_);
  and g_109128_(_003167_, _016759_, _016761_);
  or g_109129_(out[98], _016760_, _016762_);
  xor g_109130_(_003167_, _016759_, _016764_);
  xor g_109131_(out[98], _016759_, _016765_);
  and g_109132_(_016753_, _016764_, _016766_);
  or g_109133_(_016754_, _016765_, _016767_);
  and g_109134_(_003145_, _016597_, _016768_);
  not g_109135_(_016768_, _016769_);
  and g_109136_(_016541_, _016592_, _016770_);
  or g_109137_(_016540_, _016591_, _016771_);
  and g_109138_(_003024_, _016591_, _016772_);
  or g_109139_(out[80], _016592_, _016773_);
  and g_109140_(_016771_, _016773_, _016775_);
  or g_109141_(_016770_, _016772_, _016776_);
  and g_109142_(out[96], _016776_, _016777_);
  or g_109143_(_003156_, _016775_, _016778_);
  and g_109144_(out[97], _016599_, _016779_);
  or g_109145_(_003145_, _016597_, _016780_);
  and g_109146_(_016778_, _016780_, _016781_);
  or g_109147_(_016777_, _016779_, _016782_);
  and g_109148_(_016769_, _016782_, _016783_);
  or g_109149_(_016768_, _016781_, _016784_);
  and g_109150_(_016766_, _016784_, _016786_);
  or g_109151_(_016767_, _016783_, _016787_);
  and g_109152_(_016748_, _016761_, _016788_);
  or g_109153_(_016749_, _016762_, _016789_);
  and g_109154_(_016750_, _016789_, _016790_);
  or g_109155_(_016751_, _016788_, _016791_);
  and g_109156_(_016787_, _016790_, _016792_);
  or g_109157_(_016786_, _016791_, _016793_);
  and g_109158_(_016739_, _016793_, _016794_);
  or g_109159_(_016740_, _016792_, _016795_);
  and g_109160_(_016725_, _016733_, _016797_);
  or g_109161_(_016724_, _016734_, _016798_);
  and g_109162_(_016705_, _016797_, _016799_);
  or g_109163_(_016704_, _016798_, _016800_);
  and g_109164_(_016694_, _016707_, _016801_);
  or g_109165_(_016693_, _016706_, _016802_);
  and g_109166_(_016800_, _016802_, _016803_);
  or g_109167_(_016799_, _016801_, _016804_);
  and g_109168_(_016795_, _016803_, _016805_);
  or g_109169_(_016794_, _016804_, _016806_);
  and g_109170_(_016669_, _016806_, _016808_);
  or g_109171_(_016670_, _016805_, _016809_);
  and g_109172_(_016626_, _016628_, _016810_);
  or g_109173_(_016625_, _016627_, _016811_);
  and g_109174_(_016659_, _016661_, _016812_);
  or g_109175_(_016658_, _016660_, _016813_);
  and g_109176_(_016634_, _016812_, _016814_);
  or g_109177_(_016635_, _016813_, _016815_);
  and g_109178_(_016811_, _016815_, _016816_);
  or g_109179_(_016810_, _016814_, _016817_);
  and g_109180_(_016809_, _016816_, _016819_);
  or g_109181_(_016808_, _016817_, _016820_);
  and g_109182_(_003156_, _016775_, _016821_);
  or g_109183_(out[96], _016776_, _016822_);
  and g_109184_(_016769_, _016822_, _016823_);
  or g_109185_(_016768_, _016821_, _016824_);
  and g_109186_(_016766_, _016781_, _016825_);
  not g_109187_(_016825_, _016826_);
  and g_109188_(_016823_, _016825_, _016827_);
  or g_109189_(_016824_, _016826_, _016828_);
  and g_109190_(_016669_, _016827_, _016830_);
  or g_109191_(_016670_, _016828_, _016831_);
  and g_109192_(_016739_, _016830_, _016832_);
  or g_109193_(_016740_, _016831_, _016833_);
  and g_109194_(_016820_, _016833_, _016834_);
  or g_109195_(_016819_, _016832_, _016835_);
  or g_109196_(_016597_, _016834_, _016836_);
  or g_109197_(out[97], _016835_, _016837_);
  and g_109198_(_016836_, _016837_, _016838_);
  not g_109199_(_016838_, _016839_);
  and g_109200_(_016614_, _016834_, _016841_);
  not g_109201_(_016841_, _016842_);
  or g_109202_(_016621_, _016834_, _016843_);
  not g_109203_(_016843_, _016844_);
  and g_109204_(_016842_, _016843_, _016845_);
  or g_109205_(_016841_, _016844_, _016846_);
  and g_109206_(out[116], out[115], _016847_);
  or g_109207_(out[117], _016847_, _016848_);
  or g_109208_(out[118], _016848_, _016849_);
  or g_109209_(out[119], _016849_, _016850_);
  or g_109210_(out[120], _016850_, _016852_);
  and g_109211_(out[121], _016852_, _016853_);
  or g_109212_(out[122], _016853_, _016854_);
  xor g_109213_(out[122], _016853_, _016855_);
  xor g_109214_(_003343_, _016853_, _016856_);
  and g_109215_(_016845_, _016855_, _016857_);
  or g_109216_(_016846_, _016856_, _016858_);
  and g_109217_(_016600_, _016610_, _016859_);
  or g_109218_(_016601_, _016611_, _016860_);
  xor g_109219_(out[123], _016854_, _016861_);
  xor g_109220_(_003222_, _016854_, _016863_);
  and g_109221_(_016859_, _016863_, _016864_);
  or g_109222_(_016860_, _016861_, _016865_);
  and g_109223_(_016858_, _016865_, _016866_);
  or g_109224_(_016857_, _016864_, _016867_);
  and g_109225_(_016860_, _016861_, _016868_);
  or g_109226_(_016859_, _016863_, _016869_);
  and g_109227_(_016846_, _016856_, _016870_);
  or g_109228_(_016845_, _016855_, _016871_);
  and g_109229_(_016869_, _016871_, _016872_);
  or g_109230_(_016868_, _016870_, _016874_);
  xor g_109231_(out[121], _016852_, _016875_);
  xor g_109232_(_003332_, _016852_, _016876_);
  and g_109233_(_016636_, _016834_, _016877_);
  not g_109234_(_016877_, _016878_);
  or g_109235_(_016643_, _016834_, _016879_);
  not g_109236_(_016879_, _016880_);
  and g_109237_(_016878_, _016879_, _016881_);
  or g_109238_(_016877_, _016880_, _016882_);
  and g_109239_(_016875_, _016881_, _016883_);
  or g_109240_(_016876_, _016882_, _016885_);
  and g_109241_(_016866_, _016872_, _016886_);
  or g_109242_(_016867_, _016874_, _016887_);
  and g_109243_(_016885_, _016886_, _016888_);
  or g_109244_(_016883_, _016887_, _016889_);
  and g_109245_(_016876_, _016882_, _016890_);
  or g_109246_(_016875_, _016881_, _016891_);
  xor g_109247_(out[120], _016850_, _016892_);
  xor g_109248_(_003321_, _016850_, _016893_);
  and g_109249_(_016648_, _016834_, _016894_);
  not g_109250_(_016894_, _016896_);
  or g_109251_(_016654_, _016834_, _016897_);
  not g_109252_(_016897_, _016898_);
  and g_109253_(_016896_, _016897_, _016899_);
  or g_109254_(_016894_, _016898_, _016900_);
  and g_109255_(_016892_, _016900_, _016901_);
  or g_109256_(_016893_, _016899_, _016902_);
  and g_109257_(_016891_, _016902_, _016903_);
  or g_109258_(_016890_, _016901_, _016904_);
  and g_109259_(_016893_, _016899_, _016905_);
  or g_109260_(_016892_, _016900_, _016907_);
  and g_109261_(_016903_, _016907_, _016908_);
  or g_109262_(_016904_, _016905_, _016909_);
  and g_109263_(_016888_, _016908_, _016910_);
  or g_109264_(_016889_, _016909_, _016911_);
  xor g_109265_(out[119], _016849_, _016912_);
  xor g_109266_(_003233_, _016849_, _016913_);
  and g_109267_(_016683_, _016834_, _016914_);
  or g_109268_(_016682_, _016835_, _016915_);
  and g_109269_(_016690_, _016835_, _016916_);
  or g_109270_(_016689_, _016834_, _016918_);
  and g_109271_(_016915_, _016918_, _016919_);
  or g_109272_(_016914_, _016916_, _016920_);
  and g_109273_(_016912_, _016920_, _016921_);
  or g_109274_(_016913_, _016919_, _016922_);
  xor g_109275_(out[118], _016848_, _016923_);
  xor g_109276_(_003244_, _016848_, _016924_);
  and g_109277_(_016671_, _016834_, _016925_);
  or g_109278_(_016672_, _016835_, _016926_);
  and g_109279_(_016679_, _016835_, _016927_);
  or g_109280_(_016678_, _016834_, _016929_);
  and g_109281_(_016926_, _016929_, _016930_);
  or g_109282_(_016925_, _016927_, _016931_);
  and g_109283_(_016923_, _016930_, _016932_);
  or g_109284_(_016924_, _016931_, _016933_);
  and g_109285_(_016922_, _016933_, _016934_);
  or g_109286_(_016921_, _016932_, _016935_);
  and g_109287_(_016913_, _016919_, _016936_);
  or g_109288_(_016912_, _016920_, _016937_);
  and g_109289_(_016924_, _016931_, _016938_);
  or g_109290_(_016923_, _016930_, _016940_);
  and g_109291_(_016937_, _016940_, _016941_);
  or g_109292_(_016936_, _016938_, _016942_);
  and g_109293_(_016934_, _016941_, _016943_);
  or g_109294_(_016935_, _016942_, _016944_);
  xor g_109295_(out[116], out[115], _016945_);
  xor g_109296_(_003266_, out[115], _016946_);
  and g_109297_(_016711_, _016834_, _016947_);
  not g_109298_(_016947_, _016948_);
  or g_109299_(_016717_, _016834_, _016949_);
  not g_109300_(_016949_, _016951_);
  and g_109301_(_016948_, _016949_, _016952_);
  or g_109302_(_016947_, _016951_, _016953_);
  and g_109303_(_016946_, _016953_, _016954_);
  or g_109304_(_016945_, _016952_, _016955_);
  xor g_109305_(out[117], _016847_, _016956_);
  xor g_109306_(_003255_, _016847_, _016957_);
  and g_109307_(_016696_, _016834_, _016958_);
  not g_109308_(_016958_, _016959_);
  or g_109309_(_016702_, _016834_, _016960_);
  not g_109310_(_016960_, _016962_);
  and g_109311_(_016959_, _016960_, _016963_);
  or g_109312_(_016958_, _016962_, _016964_);
  and g_109313_(_016956_, _016964_, _016965_);
  or g_109314_(_016957_, _016963_, _016966_);
  and g_109315_(_016955_, _016966_, _016967_);
  or g_109316_(_016954_, _016965_, _016968_);
  and g_109317_(_016957_, _016963_, _016969_);
  or g_109318_(_016956_, _016964_, _016970_);
  and g_109319_(_016945_, _016952_, _016971_);
  or g_109320_(_016946_, _016953_, _016973_);
  and g_109321_(_016970_, _016973_, _016974_);
  or g_109322_(_016969_, _016971_, _016975_);
  and g_109323_(_016967_, _016974_, _016976_);
  or g_109324_(_016968_, _016975_, _016977_);
  and g_109325_(_016943_, _016976_, _016978_);
  or g_109326_(_016944_, _016977_, _016979_);
  and g_109327_(out[99], _016834_, _016980_);
  not g_109328_(_016980_, _016981_);
  and g_109329_(_016747_, _016835_, _016982_);
  not g_109330_(_016982_, _016984_);
  and g_109331_(_016981_, _016984_, _016985_);
  or g_109332_(_016980_, _016982_, _016986_);
  and g_109333_(out[115], _016985_, _016987_);
  or g_109334_(_003310_, _016986_, _016988_);
  or g_109335_(_016759_, _016834_, _016989_);
  not g_109336_(_016989_, _016990_);
  and g_109337_(_003167_, _016834_, _016991_);
  not g_109338_(_016991_, _016992_);
  and g_109339_(_016989_, _016992_, _016993_);
  or g_109340_(_016990_, _016991_, _016995_);
  and g_109341_(out[114], _016995_, _016996_);
  or g_109342_(_003299_, _016993_, _016997_);
  and g_109343_(_016988_, _016997_, _016998_);
  or g_109344_(_016987_, _016996_, _016999_);
  and g_109345_(_003310_, _016986_, _017000_);
  or g_109346_(out[115], _016985_, _017001_);
  and g_109347_(_003299_, _016993_, _017002_);
  or g_109348_(out[114], _016995_, _017003_);
  and g_109349_(_017001_, _017003_, _017004_);
  or g_109350_(_017000_, _017002_, _017006_);
  and g_109351_(_016998_, _017004_, _017007_);
  or g_109352_(_016999_, _017006_, _017008_);
  and g_109353_(_003277_, _016838_, _017009_);
  or g_109354_(out[113], _016839_, _017010_);
  and g_109355_(_016776_, _016835_, _017011_);
  or g_109356_(_016775_, _016834_, _017012_);
  and g_109357_(_003156_, _016834_, _017013_);
  or g_109358_(out[96], _016835_, _017014_);
  and g_109359_(_017012_, _017014_, _017015_);
  or g_109360_(_017011_, _017013_, _017017_);
  and g_109361_(out[112], _017017_, _017018_);
  or g_109362_(_003288_, _017015_, _017019_);
  xor g_109363_(_003277_, _016838_, _017020_);
  xor g_109364_(out[113], _016838_, _017021_);
  and g_109365_(_017019_, _017020_, _017022_);
  or g_109366_(_017018_, _017021_, _017023_);
  and g_109367_(_017010_, _017023_, _017024_);
  or g_109368_(_017009_, _017022_, _017025_);
  and g_109369_(_017007_, _017025_, _017026_);
  or g_109370_(_017008_, _017024_, _017028_);
  and g_109371_(_017001_, _017002_, _017029_);
  or g_109372_(_017000_, _017003_, _017030_);
  and g_109373_(_016988_, _017030_, _017031_);
  or g_109374_(_016987_, _017029_, _017032_);
  and g_109375_(_017028_, _017031_, _017033_);
  or g_109376_(_017026_, _017032_, _017034_);
  and g_109377_(_016978_, _017034_, _017035_);
  or g_109378_(_016979_, _017033_, _017036_);
  and g_109379_(_016968_, _016970_, _017037_);
  or g_109380_(_016967_, _016969_, _017039_);
  and g_109381_(_016943_, _017037_, _017040_);
  or g_109382_(_016944_, _017039_, _017041_);
  and g_109383_(_016935_, _016937_, _017042_);
  or g_109384_(_016934_, _016936_, _017043_);
  and g_109385_(_017041_, _017043_, _017044_);
  or g_109386_(_017040_, _017042_, _017045_);
  and g_109387_(_017036_, _017044_, _017046_);
  or g_109388_(_017035_, _017045_, _017047_);
  and g_109389_(_016910_, _017047_, _017048_);
  or g_109390_(_016911_, _017046_, _017050_);
  and g_109391_(_016867_, _016869_, _017051_);
  or g_109392_(_016866_, _016868_, _017052_);
  and g_109393_(_016888_, _016904_, _017053_);
  or g_109394_(_016889_, _016903_, _017054_);
  and g_109395_(_017052_, _017054_, _017055_);
  or g_109396_(_017051_, _017053_, _017056_);
  and g_109397_(_017050_, _017055_, _017057_);
  or g_109398_(_017048_, _017056_, _017058_);
  and g_109399_(_003288_, _017015_, _017059_);
  or g_109400_(out[112], _017017_, _017061_);
  or g_109401_(_017008_, _017023_, _017062_);
  not g_109402_(_017062_, _017063_);
  and g_109403_(_016910_, _017063_, _017064_);
  or g_109404_(_016911_, _017062_, _017065_);
  and g_109405_(_016978_, _017064_, _017066_);
  or g_109406_(_016979_, _017065_, _017067_);
  and g_109407_(_017061_, _017066_, _017068_);
  or g_109408_(_017059_, _017067_, _017069_);
  and g_109409_(_017058_, _017069_, _017070_);
  or g_109410_(_017057_, _017068_, _017072_);
  or g_109411_(_016838_, _017070_, _017073_);
  or g_109412_(out[113], _017072_, _017074_);
  and g_109413_(_017073_, _017074_, _017075_);
  not g_109414_(_017075_, _017076_);
  and g_109415_(_016846_, _017072_, _017077_);
  not g_109416_(_017077_, _017078_);
  or g_109417_(_016856_, _017072_, _017079_);
  not g_109418_(_017079_, _017080_);
  and g_109419_(_017078_, _017079_, _017081_);
  or g_109420_(_017077_, _017080_, _017083_);
  and g_109421_(out[132], out[131], _017084_);
  or g_109422_(out[133], _017084_, _017085_);
  or g_109423_(out[134], _017085_, _017086_);
  or g_109424_(out[135], _017086_, _017087_);
  or g_109425_(out[136], _017087_, _017088_);
  and g_109426_(out[137], _017088_, _017089_);
  or g_109427_(out[138], _017089_, _017090_);
  xor g_109428_(out[138], _017089_, _017091_);
  xor g_109429_(_003475_, _017089_, _017092_);
  and g_109430_(_017081_, _017091_, _017094_);
  or g_109431_(_017083_, _017092_, _017095_);
  and g_109432_(_016859_, _016861_, _017096_);
  or g_109433_(_016860_, _016863_, _017097_);
  xor g_109434_(out[139], _017090_, _017098_);
  xor g_109435_(_003354_, _017090_, _017099_);
  and g_109436_(_017096_, _017099_, _017100_);
  or g_109437_(_017097_, _017098_, _017101_);
  and g_109438_(_017095_, _017101_, _017102_);
  or g_109439_(_017094_, _017100_, _017103_);
  and g_109440_(_017097_, _017098_, _017105_);
  or g_109441_(_017096_, _017099_, _017106_);
  and g_109442_(_017083_, _017092_, _017107_);
  or g_109443_(_017081_, _017091_, _017108_);
  and g_109444_(_017106_, _017108_, _017109_);
  or g_109445_(_017105_, _017107_, _017110_);
  xor g_109446_(out[137], _017088_, _017111_);
  xor g_109447_(_003464_, _017088_, _017112_);
  and g_109448_(_016882_, _017072_, _017113_);
  not g_109449_(_017113_, _017114_);
  or g_109450_(_016876_, _017072_, _017116_);
  not g_109451_(_017116_, _017117_);
  and g_109452_(_017114_, _017116_, _017118_);
  or g_109453_(_017113_, _017117_, _017119_);
  and g_109454_(_017111_, _017118_, _017120_);
  or g_109455_(_017112_, _017119_, _017121_);
  and g_109456_(_017102_, _017109_, _017122_);
  or g_109457_(_017103_, _017110_, _017123_);
  and g_109458_(_017121_, _017122_, _017124_);
  or g_109459_(_017120_, _017123_, _017125_);
  and g_109460_(_017112_, _017119_, _017127_);
  or g_109461_(_017111_, _017118_, _017128_);
  xor g_109462_(out[136], _017087_, _017129_);
  xor g_109463_(_003453_, _017087_, _017130_);
  and g_109464_(_016900_, _017072_, _017131_);
  not g_109465_(_017131_, _017132_);
  or g_109466_(_016892_, _017072_, _017133_);
  not g_109467_(_017133_, _017134_);
  and g_109468_(_017132_, _017133_, _017135_);
  or g_109469_(_017131_, _017134_, _017136_);
  and g_109470_(_017129_, _017136_, _017138_);
  or g_109471_(_017130_, _017135_, _017139_);
  and g_109472_(_017128_, _017139_, _017140_);
  or g_109473_(_017127_, _017138_, _017141_);
  and g_109474_(_017130_, _017135_, _017142_);
  or g_109475_(_017129_, _017136_, _017143_);
  and g_109476_(_017140_, _017143_, _017144_);
  or g_109477_(_017141_, _017142_, _017145_);
  and g_109478_(_017124_, _017144_, _017146_);
  or g_109479_(_017125_, _017145_, _017147_);
  xor g_109480_(out[134], _017085_, _017149_);
  xor g_109481_(_003376_, _017085_, _017150_);
  and g_109482_(_016931_, _017072_, _017151_);
  or g_109483_(_016930_, _017070_, _017152_);
  and g_109484_(_016923_, _017070_, _017153_);
  or g_109485_(_016924_, _017072_, _017154_);
  and g_109486_(_017152_, _017154_, _017155_);
  or g_109487_(_017151_, _017153_, _017156_);
  and g_109488_(_017149_, _017155_, _017157_);
  or g_109489_(_017150_, _017156_, _017158_);
  xor g_109490_(out[135], _017086_, _017160_);
  not g_109491_(_017160_, _017161_);
  and g_109492_(_016920_, _017072_, _017162_);
  or g_109493_(_016919_, _017070_, _017163_);
  and g_109494_(_016913_, _017070_, _017164_);
  or g_109495_(_016912_, _017072_, _017165_);
  and g_109496_(_017163_, _017165_, _017166_);
  or g_109497_(_017162_, _017164_, _017167_);
  and g_109498_(_017160_, _017167_, _017168_);
  or g_109499_(_017161_, _017166_, _017169_);
  and g_109500_(_017158_, _017169_, _017171_);
  or g_109501_(_017157_, _017168_, _017172_);
  or g_109502_(_017149_, _017155_, _017173_);
  not g_109503_(_017173_, _017174_);
  and g_109504_(_017161_, _017166_, _017175_);
  or g_109505_(_017160_, _017167_, _017176_);
  xor g_109506_(out[133], _017084_, _017177_);
  xor g_109507_(_003387_, _017084_, _017178_);
  and g_109508_(_016964_, _017072_, _017179_);
  or g_109509_(_016963_, _017070_, _017180_);
  and g_109510_(_016957_, _017070_, _017182_);
  or g_109511_(_016956_, _017072_, _017183_);
  and g_109512_(_017180_, _017183_, _017184_);
  or g_109513_(_017179_, _017182_, _017185_);
  and g_109514_(_017178_, _017184_, _017186_);
  or g_109515_(_017177_, _017185_, _017187_);
  xor g_109516_(out[132], out[131], _017188_);
  xor g_109517_(_003398_, out[131], _017189_);
  and g_109518_(_016945_, _017070_, _017190_);
  or g_109519_(_016946_, _017072_, _017191_);
  and g_109520_(_016953_, _017072_, _017193_);
  or g_109521_(_016952_, _017070_, _017194_);
  and g_109522_(_017191_, _017194_, _017195_);
  or g_109523_(_017190_, _017193_, _017196_);
  and g_109524_(_017188_, _017195_, _017197_);
  or g_109525_(_017189_, _017196_, _017198_);
  and g_109526_(_017189_, _017196_, _017199_);
  or g_109527_(_017188_, _017195_, _017200_);
  and g_109528_(_017177_, _017185_, _017201_);
  or g_109529_(_017178_, _017184_, _017202_);
  and g_109530_(_017200_, _017202_, _017204_);
  or g_109531_(_017199_, _017201_, _017205_);
  and g_109532_(_017187_, _017204_, _017206_);
  or g_109533_(_017186_, _017205_, _017207_);
  and g_109534_(_017171_, _017173_, _017208_);
  or g_109535_(_017172_, _017174_, _017209_);
  and g_109536_(_017176_, _017208_, _017210_);
  or g_109537_(_017175_, _017209_, _017211_);
  and g_109538_(_017198_, _017206_, _017212_);
  or g_109539_(_017197_, _017207_, _017213_);
  and g_109540_(_017210_, _017212_, _017215_);
  or g_109541_(_017211_, _017213_, _017216_);
  and g_109542_(_016995_, _017072_, _017217_);
  not g_109543_(_017217_, _017218_);
  or g_109544_(out[114], _017072_, _017219_);
  not g_109545_(_017219_, _017220_);
  and g_109546_(_017218_, _017219_, _017221_);
  or g_109547_(_017217_, _017220_, _017222_);
  and g_109548_(_003431_, _017221_, _017223_);
  or g_109549_(out[130], _017222_, _017224_);
  or g_109550_(_003310_, _017072_, _017226_);
  not g_109551_(_017226_, _017227_);
  and g_109552_(_016986_, _017072_, _017228_);
  not g_109553_(_017228_, _017229_);
  and g_109554_(_017226_, _017229_, _017230_);
  or g_109555_(_017227_, _017228_, _017231_);
  and g_109556_(out[131], _017230_, _017232_);
  or g_109557_(_003442_, _017231_, _017233_);
  and g_109558_(_017224_, _017233_, _017234_);
  or g_109559_(_017223_, _017232_, _017235_);
  and g_109560_(_003442_, _017231_, _017237_);
  or g_109561_(out[131], _017230_, _017238_);
  and g_109562_(out[130], _017222_, _017239_);
  or g_109563_(_003431_, _017221_, _017240_);
  and g_109564_(_017238_, _017240_, _017241_);
  or g_109565_(_017237_, _017239_, _017242_);
  and g_109566_(_017234_, _017241_, _017243_);
  or g_109567_(_017235_, _017242_, _017244_);
  and g_109568_(_003409_, _017075_, _017245_);
  or g_109569_(out[129], _017076_, _017246_);
  and g_109570_(_017017_, _017072_, _017248_);
  or g_109571_(_017015_, _017070_, _017249_);
  and g_109572_(_003288_, _017070_, _017250_);
  or g_109573_(out[112], _017072_, _017251_);
  and g_109574_(_017249_, _017251_, _017252_);
  or g_109575_(_017248_, _017250_, _017253_);
  and g_109576_(out[128], _017253_, _017254_);
  or g_109577_(_003420_, _017252_, _017255_);
  xor g_109578_(_003409_, _017075_, _017256_);
  xor g_109579_(out[129], _017075_, _017257_);
  and g_109580_(_017255_, _017256_, _017259_);
  or g_109581_(_017254_, _017257_, _017260_);
  and g_109582_(_017246_, _017260_, _017261_);
  or g_109583_(_017245_, _017259_, _017262_);
  and g_109584_(_017243_, _017262_, _017263_);
  or g_109585_(_017244_, _017261_, _017264_);
  and g_109586_(_017223_, _017238_, _017265_);
  or g_109587_(_017224_, _017237_, _017266_);
  and g_109588_(_017233_, _017266_, _017267_);
  or g_109589_(_017232_, _017265_, _017268_);
  and g_109590_(_017264_, _017267_, _017270_);
  or g_109591_(_017263_, _017268_, _017271_);
  and g_109592_(_017215_, _017271_, _017272_);
  or g_109593_(_017216_, _017270_, _017273_);
  and g_109594_(_017205_, _017210_, _017274_);
  or g_109595_(_017204_, _017211_, _017275_);
  and g_109596_(_017187_, _017274_, _017276_);
  or g_109597_(_017186_, _017275_, _017277_);
  or g_109598_(_017171_, _017175_, _017278_);
  not g_109599_(_017278_, _017279_);
  and g_109600_(_017277_, _017278_, _017281_);
  or g_109601_(_017276_, _017279_, _017282_);
  and g_109602_(_017273_, _017281_, _017283_);
  or g_109603_(_017272_, _017282_, _017284_);
  and g_109604_(_017146_, _017284_, _017285_);
  or g_109605_(_017147_, _017283_, _017286_);
  and g_109606_(_017103_, _017106_, _017287_);
  or g_109607_(_017102_, _017105_, _017288_);
  and g_109608_(_017124_, _017141_, _017289_);
  or g_109609_(_017125_, _017140_, _017290_);
  and g_109610_(_017288_, _017290_, _017292_);
  or g_109611_(_017287_, _017289_, _017293_);
  and g_109612_(_017286_, _017292_, _017294_);
  or g_109613_(_017285_, _017293_, _017295_);
  and g_109614_(_003420_, _017252_, _017296_);
  or g_109615_(_017244_, _017260_, _017297_);
  or g_109616_(_017296_, _017297_, _017298_);
  or g_109617_(_017216_, _017298_, _017299_);
  not g_109618_(_017299_, _017300_);
  and g_109619_(_017146_, _017300_, _017301_);
  or g_109620_(_017147_, _017299_, _017303_);
  and g_109621_(_017295_, _017303_, _017304_);
  or g_109622_(_017294_, _017301_, _017305_);
  and g_109623_(_017076_, _017305_, _017306_);
  and g_109624_(_003409_, _017304_, _017307_);
  or g_109625_(_017306_, _017307_, _017308_);
  and g_109626_(_017091_, _017304_, _017309_);
  or g_109627_(_017092_, _017305_, _017310_);
  and g_109628_(_017083_, _017305_, _017311_);
  or g_109629_(_017081_, _017304_, _017312_);
  and g_109630_(_017310_, _017312_, _017314_);
  or g_109631_(_017309_, _017311_, _017315_);
  and g_109632_(out[148], out[147], _017316_);
  or g_109633_(out[149], _017316_, _017317_);
  or g_109634_(out[150], _017317_, _017318_);
  or g_109635_(out[151], _017318_, _017319_);
  or g_109636_(out[152], _017319_, _017320_);
  and g_109637_(out[153], _017320_, _017321_);
  or g_109638_(out[154], _017321_, _017322_);
  xor g_109639_(out[154], _017321_, _017323_);
  xor g_109640_(_003607_, _017321_, _017325_);
  and g_109641_(_017314_, _017323_, _017326_);
  or g_109642_(_017315_, _017325_, _017327_);
  and g_109643_(_017096_, _017098_, _017328_);
  or g_109644_(_017097_, _017099_, _017329_);
  xor g_109645_(out[155], _017322_, _017330_);
  xor g_109646_(_003486_, _017322_, _017331_);
  and g_109647_(_017328_, _017331_, _017332_);
  or g_109648_(_017329_, _017330_, _017333_);
  and g_109649_(_017327_, _017333_, _017334_);
  or g_109650_(_017326_, _017332_, _017336_);
  and g_109651_(_017329_, _017330_, _017337_);
  or g_109652_(_017328_, _017331_, _017338_);
  and g_109653_(_017315_, _017325_, _017339_);
  or g_109654_(_017314_, _017323_, _017340_);
  and g_109655_(_017338_, _017340_, _017341_);
  or g_109656_(_017337_, _017339_, _017342_);
  and g_109657_(_017334_, _017341_, _017343_);
  or g_109658_(_017336_, _017342_, _017344_);
  xor g_109659_(out[153], _017320_, _017345_);
  xor g_109660_(_003596_, _017320_, _017347_);
  and g_109661_(_017111_, _017304_, _017348_);
  or g_109662_(_017112_, _017305_, _017349_);
  and g_109663_(_017119_, _017305_, _017350_);
  or g_109664_(_017118_, _017304_, _017351_);
  and g_109665_(_017349_, _017351_, _017352_);
  or g_109666_(_017348_, _017350_, _017353_);
  and g_109667_(_017347_, _017353_, _017354_);
  or g_109668_(_017345_, _017352_, _017355_);
  xor g_109669_(out[152], _017319_, _017356_);
  not g_109670_(_017356_, _017358_);
  and g_109671_(_017130_, _017304_, _017359_);
  or g_109672_(_017129_, _017305_, _017360_);
  and g_109673_(_017136_, _017305_, _017361_);
  or g_109674_(_017135_, _017304_, _017362_);
  and g_109675_(_017360_, _017362_, _017363_);
  or g_109676_(_017359_, _017361_, _017364_);
  and g_109677_(_017356_, _017364_, _017365_);
  or g_109678_(_017358_, _017363_, _017366_);
  and g_109679_(_017355_, _017366_, _017367_);
  or g_109680_(_017354_, _017365_, _017369_);
  and g_109681_(_017345_, _017352_, _017370_);
  or g_109682_(_017347_, _017353_, _017371_);
  and g_109683_(_017358_, _017363_, _017372_);
  or g_109684_(_017356_, _017364_, _017373_);
  and g_109685_(_017371_, _017373_, _017374_);
  or g_109686_(_017370_, _017372_, _017375_);
  and g_109687_(_017367_, _017374_, _017376_);
  or g_109688_(_017369_, _017375_, _017377_);
  and g_109689_(_017343_, _017376_, _017378_);
  or g_109690_(_017344_, _017377_, _017380_);
  xor g_109691_(out[150], _017317_, _017381_);
  xor g_109692_(_003508_, _017317_, _017382_);
  or g_109693_(_017150_, _017305_, _017383_);
  or g_109694_(_017155_, _017304_, _017384_);
  and g_109695_(_017383_, _017384_, _017385_);
  not g_109696_(_017385_, _017386_);
  and g_109697_(_017381_, _017385_, _017387_);
  xor g_109698_(out[151], _017318_, _017388_);
  xor g_109699_(_003497_, _017318_, _017389_);
  or g_109700_(_017160_, _017305_, _017391_);
  or g_109701_(_017166_, _017304_, _017392_);
  and g_109702_(_017391_, _017392_, _017393_);
  not g_109703_(_017393_, _017394_);
  and g_109704_(_017388_, _017394_, _017395_);
  or g_109705_(_017387_, _017395_, _017396_);
  and g_109706_(_017382_, _017386_, _017397_);
  and g_109707_(_017389_, _017393_, _017398_);
  or g_109708_(_017388_, _017394_, _017399_);
  or g_109709_(_017397_, _017398_, _017400_);
  xor g_109710_(_017381_, _017385_, _017402_);
  xor g_109711_(_017389_, _017393_, _017403_);
  and g_109712_(_017402_, _017403_, _017404_);
  or g_109713_(_017396_, _017400_, _017405_);
  xor g_109714_(out[149], _017316_, _017406_);
  xor g_109715_(_003519_, _017316_, _017407_);
  and g_109716_(_017178_, _017304_, _017408_);
  or g_109717_(_017177_, _017305_, _017409_);
  and g_109718_(_017185_, _017305_, _017410_);
  or g_109719_(_017184_, _017304_, _017411_);
  and g_109720_(_017409_, _017411_, _017413_);
  or g_109721_(_017408_, _017410_, _017414_);
  or g_109722_(_017406_, _017414_, _017415_);
  xor g_109723_(out[148], out[147], _017416_);
  xor g_109724_(_003530_, out[147], _017417_);
  and g_109725_(_017188_, _017304_, _017418_);
  or g_109726_(_017189_, _017305_, _017419_);
  and g_109727_(_017196_, _017305_, _017420_);
  or g_109728_(_017195_, _017304_, _017421_);
  and g_109729_(_017419_, _017421_, _017422_);
  or g_109730_(_017418_, _017420_, _017424_);
  or g_109731_(_017417_, _017424_, _017425_);
  and g_109732_(_017415_, _017425_, _017426_);
  not g_109733_(_017426_, _017427_);
  and g_109734_(_017406_, _017414_, _017428_);
  or g_109735_(_017407_, _017413_, _017429_);
  and g_109736_(_017417_, _017424_, _017430_);
  or g_109737_(_017416_, _017422_, _017431_);
  and g_109738_(_017429_, _017431_, _017432_);
  or g_109739_(_017428_, _017430_, _017433_);
  and g_109740_(_017426_, _017432_, _017435_);
  or g_109741_(_017427_, _017433_, _017436_);
  and g_109742_(_017404_, _017435_, _017437_);
  or g_109743_(_017380_, _017436_, _017438_);
  and g_109744_(_017378_, _017437_, _017439_);
  or g_109745_(_017405_, _017438_, _017440_);
  and g_109746_(out[131], _017304_, _017441_);
  and g_109747_(_017231_, _017305_, _017442_);
  or g_109748_(_017441_, _017442_, _017443_);
  not g_109749_(_017443_, _017444_);
  and g_109750_(out[147], _017444_, _017446_);
  or g_109751_(_003574_, _017443_, _017447_);
  and g_109752_(_017222_, _017305_, _017448_);
  and g_109753_(_003431_, _017304_, _017449_);
  or g_109754_(_017448_, _017449_, _017450_);
  not g_109755_(_017450_, _017451_);
  and g_109756_(out[146], _017450_, _017452_);
  or g_109757_(_003563_, _017451_, _017453_);
  and g_109758_(_017447_, _017453_, _017454_);
  or g_109759_(_017446_, _017452_, _017455_);
  and g_109760_(_003574_, _017443_, _017457_);
  or g_109761_(out[147], _017444_, _017458_);
  or g_109762_(out[146], _017450_, _017459_);
  not g_109763_(_017459_, _017460_);
  and g_109764_(_017458_, _017459_, _017461_);
  or g_109765_(_017457_, _017460_, _017462_);
  and g_109766_(_017454_, _017461_, _017463_);
  or g_109767_(_017455_, _017462_, _017464_);
  or g_109768_(out[145], _017308_, _017465_);
  not g_109769_(_017465_, _017466_);
  or g_109770_(_017252_, _017304_, _017468_);
  not g_109771_(_017468_, _017469_);
  and g_109772_(_003420_, _017304_, _017470_);
  not g_109773_(_017470_, _017471_);
  and g_109774_(_017468_, _017471_, _017472_);
  or g_109775_(_017469_, _017470_, _017473_);
  and g_109776_(out[144], _017473_, _017474_);
  or g_109777_(_003552_, _017472_, _017475_);
  xor g_109778_(out[145], _017308_, _017476_);
  xor g_109779_(_003541_, _017308_, _017477_);
  and g_109780_(_017475_, _017476_, _017479_);
  or g_109781_(_017474_, _017477_, _017480_);
  and g_109782_(_017465_, _017480_, _017481_);
  or g_109783_(_017466_, _017479_, _017482_);
  and g_109784_(_017463_, _017482_, _017483_);
  or g_109785_(_017464_, _017481_, _017484_);
  and g_109786_(_017458_, _017460_, _017485_);
  or g_109787_(_017457_, _017459_, _017486_);
  and g_109788_(_017447_, _017486_, _017487_);
  or g_109789_(_017446_, _017485_, _017488_);
  and g_109790_(_017484_, _017487_, _017490_);
  or g_109791_(_017483_, _017488_, _017491_);
  and g_109792_(_017439_, _017491_, _017492_);
  or g_109793_(_017440_, _017490_, _017493_);
  and g_109794_(_017396_, _017399_, _017494_);
  and g_109795_(_017404_, _017433_, _017495_);
  and g_109796_(_017415_, _017495_, _017496_);
  or g_109797_(_017494_, _017496_, _017497_);
  and g_109798_(_017378_, _017497_, _017498_);
  and g_109799_(_017336_, _017338_, _017499_);
  and g_109800_(_017369_, _017371_, _017501_);
  and g_109801_(_017343_, _017501_, _017502_);
  or g_109802_(_017499_, _017502_, _017503_);
  or g_109803_(_017498_, _017503_, _017504_);
  not g_109804_(_017504_, _017505_);
  and g_109805_(_017493_, _017505_, _017506_);
  or g_109806_(_017492_, _017504_, _017507_);
  or g_109807_(out[144], _017473_, _017508_);
  not g_109808_(_017508_, _017509_);
  or g_109809_(_017464_, _017509_, _017510_);
  or g_109810_(_017480_, _017510_, _017512_);
  or g_109811_(_017440_, _017512_, _017513_);
  not g_109812_(_017513_, _017514_);
  and g_109813_(_017507_, _017513_, _017515_);
  or g_109814_(_017506_, _017514_, _017516_);
  and g_109815_(_017308_, _017516_, _017517_);
  and g_109816_(_003541_, _017515_, _017518_);
  or g_109817_(_017517_, _017518_, _017519_);
  and g_109818_(_017323_, _017515_, _017520_);
  or g_109819_(_017325_, _017516_, _017521_);
  and g_109820_(_017315_, _017516_, _017523_);
  or g_109821_(_017314_, _017515_, _017524_);
  and g_109822_(_017521_, _017524_, _017525_);
  or g_109823_(_017520_, _017523_, _017526_);
  and g_109824_(out[164], out[163], _017527_);
  or g_109825_(out[165], _017527_, _017528_);
  or g_109826_(out[166], _017528_, _017529_);
  or g_109827_(out[167], _017529_, _017530_);
  or g_109828_(out[168], _017530_, _017531_);
  and g_109829_(out[169], _017531_, _017532_);
  or g_109830_(out[170], _017532_, _017534_);
  xor g_109831_(out[170], _017532_, _017535_);
  xor g_109832_(_003739_, _017532_, _017536_);
  and g_109833_(_017525_, _017535_, _017537_);
  or g_109834_(_017526_, _017536_, _017538_);
  and g_109835_(_017328_, _017330_, _017539_);
  or g_109836_(_017329_, _017331_, _017540_);
  xor g_109837_(out[171], _017534_, _017541_);
  xor g_109838_(_003618_, _017534_, _017542_);
  and g_109839_(_017539_, _017542_, _017543_);
  or g_109840_(_017540_, _017541_, _017545_);
  and g_109841_(_017538_, _017545_, _017546_);
  or g_109842_(_017537_, _017543_, _017547_);
  and g_109843_(_017540_, _017541_, _017548_);
  or g_109844_(_017539_, _017542_, _017549_);
  and g_109845_(_017526_, _017536_, _017550_);
  or g_109846_(_017525_, _017535_, _017551_);
  and g_109847_(_017549_, _017551_, _017552_);
  or g_109848_(_017548_, _017550_, _017553_);
  xor g_109849_(out[169], _017531_, _017554_);
  xor g_109850_(_003728_, _017531_, _017556_);
  or g_109851_(_017347_, _017516_, _017557_);
  not g_109852_(_017557_, _017558_);
  and g_109853_(_017353_, _017516_, _017559_);
  not g_109854_(_017559_, _017560_);
  and g_109855_(_017557_, _017560_, _017561_);
  or g_109856_(_017558_, _017559_, _017562_);
  and g_109857_(_017554_, _017561_, _017563_);
  or g_109858_(_017556_, _017562_, _017564_);
  and g_109859_(_017546_, _017552_, _017565_);
  or g_109860_(_017547_, _017553_, _017567_);
  and g_109861_(_017564_, _017565_, _017568_);
  or g_109862_(_017563_, _017567_, _017569_);
  and g_109863_(_017556_, _017562_, _017570_);
  or g_109864_(_017554_, _017561_, _017571_);
  xor g_109865_(out[168], _017530_, _017572_);
  xor g_109866_(_003717_, _017530_, _017573_);
  or g_109867_(_017356_, _017516_, _017574_);
  not g_109868_(_017574_, _017575_);
  and g_109869_(_017364_, _017516_, _017576_);
  not g_109870_(_017576_, _017578_);
  and g_109871_(_017574_, _017578_, _017579_);
  or g_109872_(_017575_, _017576_, _017580_);
  and g_109873_(_017572_, _017580_, _017581_);
  or g_109874_(_017573_, _017579_, _017582_);
  and g_109875_(_017571_, _017582_, _017583_);
  or g_109876_(_017570_, _017581_, _017584_);
  and g_109877_(_017573_, _017579_, _017585_);
  or g_109878_(_017572_, _017580_, _017586_);
  and g_109879_(_017583_, _017586_, _017587_);
  or g_109880_(_017584_, _017585_, _017589_);
  and g_109881_(_017568_, _017587_, _017590_);
  or g_109882_(_017569_, _017589_, _017591_);
  xor g_109883_(out[167], _017529_, _017592_);
  xor g_109884_(_003629_, _017529_, _017593_);
  or g_109885_(_017388_, _017516_, _017594_);
  not g_109886_(_017594_, _017595_);
  and g_109887_(_017394_, _017516_, _017596_);
  not g_109888_(_017596_, _017597_);
  and g_109889_(_017594_, _017597_, _017598_);
  or g_109890_(_017595_, _017596_, _017600_);
  and g_109891_(_017592_, _017600_, _017601_);
  or g_109892_(_017593_, _017598_, _017602_);
  xor g_109893_(out[166], _017528_, _017603_);
  xor g_109894_(_003640_, _017528_, _017604_);
  or g_109895_(_017382_, _017516_, _017605_);
  not g_109896_(_017605_, _017606_);
  and g_109897_(_017386_, _017516_, _017607_);
  not g_109898_(_017607_, _017608_);
  and g_109899_(_017605_, _017608_, _017609_);
  or g_109900_(_017606_, _017607_, _017611_);
  and g_109901_(_017603_, _017609_, _017612_);
  or g_109902_(_017604_, _017611_, _017613_);
  and g_109903_(_017602_, _017613_, _017614_);
  or g_109904_(_017601_, _017612_, _017615_);
  and g_109905_(_017593_, _017598_, _017616_);
  or g_109906_(_017592_, _017600_, _017617_);
  and g_109907_(_017604_, _017611_, _017618_);
  or g_109908_(_017603_, _017609_, _017619_);
  and g_109909_(_017617_, _017619_, _017620_);
  or g_109910_(_017616_, _017618_, _017622_);
  and g_109911_(_017614_, _017620_, _017623_);
  or g_109912_(_017615_, _017622_, _017624_);
  xor g_109913_(out[164], out[163], _017625_);
  xor g_109914_(_003662_, out[163], _017626_);
  or g_109915_(_017417_, _017516_, _017627_);
  not g_109916_(_017627_, _017628_);
  and g_109917_(_017424_, _017516_, _017629_);
  not g_109918_(_017629_, _017630_);
  and g_109919_(_017627_, _017630_, _017631_);
  or g_109920_(_017628_, _017629_, _017633_);
  and g_109921_(_017626_, _017633_, _017634_);
  or g_109922_(_017625_, _017631_, _017635_);
  xor g_109923_(out[165], _017527_, _017636_);
  xor g_109924_(_003651_, _017527_, _017637_);
  or g_109925_(_017406_, _017516_, _017638_);
  not g_109926_(_017638_, _017639_);
  and g_109927_(_017414_, _017516_, _017640_);
  not g_109928_(_017640_, _017641_);
  and g_109929_(_017638_, _017641_, _017642_);
  or g_109930_(_017639_, _017640_, _017644_);
  and g_109931_(_017636_, _017644_, _017645_);
  or g_109932_(_017637_, _017642_, _017646_);
  and g_109933_(_017635_, _017646_, _017647_);
  or g_109934_(_017634_, _017645_, _017648_);
  and g_109935_(_017637_, _017642_, _017649_);
  or g_109936_(_017636_, _017644_, _017650_);
  and g_109937_(_017625_, _017631_, _017651_);
  or g_109938_(_017626_, _017633_, _017652_);
  and g_109939_(_017650_, _017652_, _017653_);
  or g_109940_(_017649_, _017651_, _017655_);
  and g_109941_(_017647_, _017653_, _017656_);
  or g_109942_(_017648_, _017655_, _017657_);
  and g_109943_(_017623_, _017656_, _017658_);
  or g_109944_(_017624_, _017657_, _017659_);
  and g_109945_(_017590_, _017658_, _017660_);
  or g_109946_(_017591_, _017659_, _017661_);
  or g_109947_(_003574_, _017516_, _017662_);
  not g_109948_(_017662_, _017663_);
  and g_109949_(_017443_, _017516_, _017664_);
  not g_109950_(_017664_, _017666_);
  and g_109951_(_017662_, _017666_, _017667_);
  or g_109952_(_017663_, _017664_, _017668_);
  and g_109953_(out[163], _017667_, _017669_);
  or g_109954_(_003706_, _017668_, _017670_);
  and g_109955_(_017450_, _017516_, _017671_);
  not g_109956_(_017671_, _017672_);
  or g_109957_(out[146], _017516_, _017673_);
  not g_109958_(_017673_, _017674_);
  and g_109959_(_017672_, _017673_, _017675_);
  or g_109960_(_017671_, _017674_, _017677_);
  and g_109961_(out[162], _017677_, _017678_);
  or g_109962_(_003695_, _017675_, _017679_);
  and g_109963_(_017670_, _017679_, _017680_);
  or g_109964_(_017669_, _017678_, _017681_);
  and g_109965_(_003706_, _017668_, _017682_);
  or g_109966_(out[163], _017667_, _017683_);
  and g_109967_(_003695_, _017675_, _017684_);
  or g_109968_(out[162], _017677_, _017685_);
  and g_109969_(_017683_, _017685_, _017686_);
  or g_109970_(_017682_, _017684_, _017688_);
  and g_109971_(_017680_, _017686_, _017689_);
  or g_109972_(_017681_, _017688_, _017690_);
  or g_109973_(out[161], _017519_, _017691_);
  and g_109974_(_017473_, _017516_, _017692_);
  not g_109975_(_017692_, _017693_);
  or g_109976_(out[144], _017516_, _017694_);
  not g_109977_(_017694_, _017695_);
  and g_109978_(_017693_, _017694_, _017696_);
  or g_109979_(_017692_, _017695_, _017697_);
  and g_109980_(out[160], _017697_, _017699_);
  xor g_109981_(_003673_, _017519_, _017700_);
  or g_109982_(_017699_, _017700_, _017701_);
  not g_109983_(_017701_, _017702_);
  and g_109984_(_017691_, _017701_, _017703_);
  not g_109985_(_017703_, _017704_);
  and g_109986_(_017689_, _017704_, _017705_);
  or g_109987_(_017690_, _017703_, _017706_);
  and g_109988_(_017683_, _017684_, _017707_);
  or g_109989_(_017682_, _017685_, _017708_);
  and g_109990_(_017670_, _017708_, _017710_);
  or g_109991_(_017669_, _017707_, _017711_);
  and g_109992_(_017706_, _017710_, _017712_);
  or g_109993_(_017705_, _017711_, _017713_);
  and g_109994_(_017660_, _017713_, _017714_);
  or g_109995_(_017661_, _017712_, _017715_);
  and g_109996_(_017648_, _017650_, _017716_);
  or g_109997_(_017647_, _017649_, _017717_);
  and g_109998_(_017623_, _017716_, _017718_);
  or g_109999_(_017624_, _017717_, _017719_);
  and g_110000_(_017615_, _017617_, _017721_);
  or g_110001_(_017614_, _017616_, _017722_);
  and g_110002_(_017719_, _017722_, _017723_);
  or g_110003_(_017718_, _017721_, _017724_);
  and g_110004_(_017590_, _017724_, _017725_);
  or g_110005_(_017591_, _017723_, _017726_);
  and g_110006_(_017568_, _017584_, _017727_);
  or g_110007_(_017569_, _017583_, _017728_);
  and g_110008_(_017547_, _017549_, _017729_);
  or g_110009_(_017546_, _017548_, _017730_);
  and g_110010_(_017728_, _017730_, _017732_);
  or g_110011_(_017727_, _017729_, _017733_);
  or g_110012_(_017725_, _017733_, _017734_);
  and g_110013_(_017715_, _017732_, _017735_);
  and g_110014_(_017726_, _017735_, _017736_);
  or g_110015_(_017714_, _017734_, _017737_);
  and g_110016_(_003684_, _017696_, _017738_);
  or g_110017_(out[160], _017697_, _017739_);
  and g_110018_(_017689_, _017739_, _017740_);
  or g_110019_(_017690_, _017738_, _017741_);
  and g_110020_(_017702_, _017740_, _017743_);
  or g_110021_(_017701_, _017741_, _017744_);
  and g_110022_(_017660_, _017743_, _017745_);
  or g_110023_(_017661_, _017744_, _017746_);
  and g_110024_(_017737_, _017746_, _017747_);
  or g_110025_(_017736_, _017745_, _017748_);
  and g_110026_(_017519_, _017748_, _017749_);
  and g_110027_(_003673_, _017747_, _017750_);
  or g_110028_(_017749_, _017750_, _017751_);
  and g_110029_(_017539_, _017541_, _017752_);
  or g_110030_(_017540_, _017542_, _017754_);
  and g_110031_(out[180], out[179], _017755_);
  or g_110032_(out[181], _017755_, _017756_);
  or g_110033_(out[182], _017756_, _017757_);
  or g_110034_(out[183], _017757_, _017758_);
  or g_110035_(out[184], _017758_, _017759_);
  and g_110036_(out[185], _017759_, _017760_);
  or g_110037_(out[186], _017760_, _017761_);
  xor g_110038_(out[187], _017761_, _017762_);
  xor g_110039_(_003750_, _017761_, _017763_);
  and g_110040_(_017752_, _017763_, _017765_);
  or g_110041_(_017754_, _017762_, _017766_);
  and g_110042_(_017535_, _017747_, _017767_);
  and g_110043_(_017526_, _017748_, _017768_);
  or g_110044_(_017767_, _017768_, _017769_);
  xor g_110045_(_003871_, _017760_, _017770_);
  or g_110046_(_017769_, _017770_, _017771_);
  not g_110047_(_017771_, _017772_);
  and g_110048_(_017766_, _017771_, _017773_);
  or g_110049_(_017765_, _017772_, _017774_);
  and g_110050_(_017769_, _017770_, _017776_);
  not g_110051_(_017776_, _017777_);
  and g_110052_(_017754_, _017762_, _017778_);
  or g_110053_(_017752_, _017763_, _017779_);
  xor g_110054_(_003860_, _017759_, _017780_);
  and g_110055_(_017554_, _017747_, _017781_);
  and g_110056_(_017562_, _017748_, _017782_);
  or g_110057_(_017781_, _017782_, _017783_);
  or g_110058_(_017780_, _017783_, _017784_);
  not g_110059_(_017784_, _017785_);
  and g_110060_(_017779_, _017784_, _017787_);
  or g_110061_(_017778_, _017785_, _017788_);
  and g_110062_(_017777_, _017787_, _017789_);
  or g_110063_(_017776_, _017788_, _017790_);
  and g_110064_(_017773_, _017789_, _017791_);
  or g_110065_(_017774_, _017790_, _017792_);
  xor g_110066_(out[184], _017758_, _017793_);
  and g_110067_(_017573_, _017747_, _017794_);
  and g_110068_(_017580_, _017748_, _017795_);
  or g_110069_(_017794_, _017795_, _017796_);
  and g_110070_(_017793_, _017796_, _017798_);
  not g_110071_(_017798_, _017799_);
  and g_110072_(_017780_, _017783_, _017800_);
  not g_110073_(_017800_, _017801_);
  and g_110074_(_017799_, _017801_, _017802_);
  or g_110075_(_017798_, _017800_, _017803_);
  or g_110076_(_017793_, _017796_, _017804_);
  not g_110077_(_017804_, _017805_);
  and g_110078_(_017802_, _017804_, _017806_);
  or g_110079_(_017803_, _017805_, _017807_);
  and g_110080_(_017791_, _017806_, _017809_);
  or g_110081_(_017792_, _017807_, _017810_);
  xor g_110082_(out[182], _017756_, _017811_);
  xor g_110083_(_003772_, _017756_, _017812_);
  and g_110084_(_017603_, _017747_, _017813_);
  or g_110085_(_017604_, _017748_, _017814_);
  and g_110086_(_017611_, _017748_, _017815_);
  or g_110087_(_017609_, _017747_, _017816_);
  and g_110088_(_017814_, _017816_, _017817_);
  or g_110089_(_017813_, _017815_, _017818_);
  and g_110090_(_017811_, _017817_, _017820_);
  or g_110091_(_017812_, _017818_, _017821_);
  xor g_110092_(out[183], _017757_, _017822_);
  xor g_110093_(_003761_, _017757_, _017823_);
  and g_110094_(_017593_, _017747_, _017824_);
  or g_110095_(_017592_, _017748_, _017825_);
  and g_110096_(_017600_, _017748_, _017826_);
  or g_110097_(_017598_, _017747_, _017827_);
  and g_110098_(_017825_, _017827_, _017828_);
  or g_110099_(_017824_, _017826_, _017829_);
  and g_110100_(_017822_, _017829_, _017831_);
  or g_110101_(_017823_, _017828_, _017832_);
  and g_110102_(_017821_, _017832_, _017833_);
  or g_110103_(_017820_, _017831_, _017834_);
  and g_110104_(_017823_, _017828_, _017835_);
  or g_110105_(_017822_, _017829_, _017836_);
  and g_110106_(_017812_, _017818_, _017837_);
  or g_110107_(_017811_, _017817_, _017838_);
  and g_110108_(_017836_, _017838_, _017839_);
  or g_110109_(_017835_, _017837_, _017840_);
  and g_110110_(_017833_, _017839_, _017842_);
  or g_110111_(_017834_, _017840_, _017843_);
  xor g_110112_(out[180], out[179], _017844_);
  xor g_110113_(_003794_, out[179], _017845_);
  and g_110114_(_017625_, _017747_, _017846_);
  or g_110115_(_017626_, _017748_, _017847_);
  and g_110116_(_017633_, _017748_, _017848_);
  or g_110117_(_017631_, _017747_, _017849_);
  and g_110118_(_017847_, _017849_, _017850_);
  or g_110119_(_017846_, _017848_, _017851_);
  and g_110120_(_017845_, _017851_, _017853_);
  or g_110121_(_017844_, _017850_, _017854_);
  xor g_110122_(out[181], _017755_, _017855_);
  xor g_110123_(_003783_, _017755_, _017856_);
  and g_110124_(_017637_, _017747_, _017857_);
  or g_110125_(_017636_, _017748_, _017858_);
  and g_110126_(_017644_, _017748_, _017859_);
  or g_110127_(_017642_, _017747_, _017860_);
  and g_110128_(_017858_, _017860_, _017861_);
  or g_110129_(_017857_, _017859_, _017862_);
  and g_110130_(_017855_, _017862_, _017864_);
  or g_110131_(_017856_, _017861_, _017865_);
  and g_110132_(_017854_, _017865_, _017866_);
  or g_110133_(_017853_, _017864_, _017867_);
  or g_110134_(_017855_, _017862_, _017868_);
  or g_110135_(_017845_, _017851_, _017869_);
  and g_110136_(_017868_, _017869_, _017870_);
  not g_110137_(_017870_, _017871_);
  and g_110138_(_017866_, _017870_, _017872_);
  or g_110139_(_017867_, _017871_, _017873_);
  and g_110140_(_017842_, _017872_, _017875_);
  or g_110141_(_017843_, _017873_, _017876_);
  and g_110142_(out[163], _017747_, _017877_);
  or g_110143_(_003706_, _017748_, _017878_);
  and g_110144_(_017668_, _017748_, _017879_);
  or g_110145_(_017667_, _017747_, _017880_);
  and g_110146_(_017878_, _017880_, _017881_);
  or g_110147_(_017877_, _017879_, _017882_);
  and g_110148_(out[179], _017881_, _017883_);
  or g_110149_(_003838_, _017882_, _017884_);
  and g_110150_(_017677_, _017748_, _017886_);
  not g_110151_(_017886_, _017887_);
  or g_110152_(out[162], _017748_, _017888_);
  not g_110153_(_017888_, _017889_);
  and g_110154_(_017887_, _017888_, _017890_);
  or g_110155_(_017886_, _017889_, _017891_);
  and g_110156_(out[178], _017891_, _017892_);
  or g_110157_(_003827_, _017890_, _017893_);
  and g_110158_(_017884_, _017893_, _017894_);
  or g_110159_(_017883_, _017892_, _017895_);
  and g_110160_(_003838_, _017882_, _017897_);
  or g_110161_(out[179], _017881_, _017898_);
  and g_110162_(_003827_, _017890_, _017899_);
  or g_110163_(out[178], _017891_, _017900_);
  and g_110164_(_017898_, _017900_, _017901_);
  or g_110165_(_017897_, _017899_, _017902_);
  and g_110166_(_017894_, _017901_, _017903_);
  or g_110167_(_017895_, _017902_, _017904_);
  or g_110168_(out[177], _017751_, _017905_);
  not g_110169_(_017905_, _017906_);
  and g_110170_(_017697_, _017748_, _017908_);
  or g_110171_(_017696_, _017747_, _017909_);
  and g_110172_(_003684_, _017747_, _017910_);
  or g_110173_(out[160], _017748_, _017911_);
  and g_110174_(_017909_, _017911_, _017912_);
  or g_110175_(_017908_, _017910_, _017913_);
  and g_110176_(out[176], _017913_, _017914_);
  or g_110177_(_003816_, _017912_, _017915_);
  xor g_110178_(out[177], _017751_, _017916_);
  xor g_110179_(_003805_, _017751_, _017917_);
  and g_110180_(_017915_, _017916_, _017919_);
  or g_110181_(_017914_, _017917_, _017920_);
  and g_110182_(_017905_, _017920_, _017921_);
  or g_110183_(_017906_, _017919_, _017922_);
  and g_110184_(_017903_, _017922_, _017923_);
  or g_110185_(_017904_, _017921_, _017924_);
  and g_110186_(_017898_, _017899_, _017925_);
  or g_110187_(_017897_, _017900_, _017926_);
  and g_110188_(_017884_, _017926_, _017927_);
  or g_110189_(_017883_, _017925_, _017928_);
  and g_110190_(_017924_, _017927_, _017930_);
  or g_110191_(_017923_, _017928_, _017931_);
  and g_110192_(_017875_, _017931_, _017932_);
  or g_110193_(_017876_, _017930_, _017933_);
  and g_110194_(_017867_, _017868_, _017934_);
  and g_110195_(_017842_, _017934_, _017935_);
  not g_110196_(_017935_, _017936_);
  and g_110197_(_017834_, _017836_, _017937_);
  or g_110198_(_017833_, _017835_, _017938_);
  and g_110199_(_017936_, _017938_, _017939_);
  or g_110200_(_017935_, _017937_, _017941_);
  and g_110201_(_017933_, _017939_, _017942_);
  or g_110202_(_017932_, _017941_, _017943_);
  and g_110203_(_017809_, _017943_, _017944_);
  or g_110204_(_017810_, _017942_, _017945_);
  and g_110205_(_017774_, _017779_, _017946_);
  or g_110206_(_017773_, _017778_, _017947_);
  and g_110207_(_017791_, _017803_, _017948_);
  not g_110208_(_017948_, _017949_);
  and g_110209_(_017947_, _017949_, _017950_);
  or g_110210_(_017946_, _017948_, _017952_);
  and g_110211_(_017945_, _017950_, _017953_);
  or g_110212_(_017944_, _017952_, _017954_);
  and g_110213_(_003816_, _017912_, _017955_);
  or g_110214_(_017904_, _017920_, _017956_);
  or g_110215_(_017955_, _017956_, _017957_);
  or g_110216_(_017876_, _017957_, _017958_);
  not g_110217_(_017958_, _017959_);
  and g_110218_(_017809_, _017959_, _017960_);
  or g_110219_(_017810_, _017958_, _017961_);
  and g_110220_(_017954_, _017961_, _017963_);
  or g_110221_(_017953_, _017960_, _017964_);
  and g_110222_(_017751_, _017964_, _017965_);
  and g_110223_(_003805_, _017963_, _017966_);
  or g_110224_(_017965_, _017966_, _017967_);
  and g_110225_(out[196], out[195], _017968_);
  or g_110226_(out[197], _017968_, _017969_);
  or g_110227_(out[198], _017969_, _017970_);
  or g_110228_(out[199], _017970_, _017971_);
  or g_110229_(out[200], _017971_, _017972_);
  and g_110230_(out[201], _017972_, _017974_);
  or g_110231_(out[202], _017974_, _017975_);
  xor g_110232_(out[202], _017974_, _017976_);
  not g_110233_(_017976_, _017977_);
  and g_110234_(_017769_, _017964_, _017978_);
  not g_110235_(_017978_, _017979_);
  or g_110236_(_017770_, _017964_, _017980_);
  not g_110237_(_017980_, _017981_);
  and g_110238_(_017979_, _017980_, _017982_);
  or g_110239_(_017978_, _017981_, _017983_);
  and g_110240_(_017976_, _017982_, _017985_);
  or g_110241_(_017977_, _017983_, _017986_);
  and g_110242_(_017752_, _017762_, _017987_);
  or g_110243_(_017754_, _017763_, _017988_);
  xor g_110244_(out[203], _017975_, _017989_);
  xor g_110245_(_003882_, _017975_, _017990_);
  and g_110246_(_017987_, _017990_, _017991_);
  or g_110247_(_017988_, _017989_, _017992_);
  and g_110248_(_017986_, _017992_, _017993_);
  or g_110249_(_017985_, _017991_, _017994_);
  or g_110250_(_017976_, _017982_, _017996_);
  not g_110251_(_017996_, _017997_);
  and g_110252_(_017988_, _017989_, _017998_);
  or g_110253_(_017987_, _017990_, _017999_);
  and g_110254_(_017783_, _017964_, _018000_);
  not g_110255_(_018000_, _018001_);
  or g_110256_(_017780_, _017964_, _018002_);
  and g_110257_(_018001_, _018002_, _018003_);
  xor g_110258_(out[201], _017972_, _018004_);
  and g_110259_(_018003_, _018004_, _018005_);
  not g_110260_(_018005_, _018007_);
  or g_110261_(_017998_, _018005_, _018008_);
  or g_110262_(_017997_, _018008_, _018009_);
  and g_110263_(_017996_, _017999_, _018010_);
  and g_110264_(_017993_, _018010_, _018011_);
  and g_110265_(_018007_, _018011_, _018012_);
  or g_110266_(_017994_, _018009_, _018013_);
  or g_110267_(_018003_, _018004_, _018014_);
  not g_110268_(_018014_, _018015_);
  xor g_110269_(_003981_, _017971_, _018016_);
  and g_110270_(_017796_, _017964_, _018018_);
  not g_110271_(_018018_, _018019_);
  or g_110272_(_017793_, _017964_, _018020_);
  and g_110273_(_018019_, _018020_, _018021_);
  or g_110274_(_018016_, _018021_, _018022_);
  not g_110275_(_018022_, _018023_);
  and g_110276_(_018014_, _018022_, _018024_);
  or g_110277_(_018015_, _018023_, _018025_);
  and g_110278_(_018016_, _018021_, _018026_);
  not g_110279_(_018026_, _018027_);
  and g_110280_(_018024_, _018027_, _018029_);
  or g_110281_(_018025_, _018026_, _018030_);
  and g_110282_(_018012_, _018029_, _018031_);
  or g_110283_(_018013_, _018030_, _018032_);
  xor g_110284_(out[199], _017970_, _018033_);
  xor g_110285_(_003893_, _017970_, _018034_);
  and g_110286_(_017829_, _017964_, _018035_);
  or g_110287_(_017828_, _017963_, _018036_);
  and g_110288_(_017823_, _017963_, _018037_);
  or g_110289_(_017822_, _017964_, _018038_);
  and g_110290_(_018036_, _018038_, _018040_);
  or g_110291_(_018035_, _018037_, _018041_);
  and g_110292_(_018034_, _018040_, _018042_);
  or g_110293_(_018033_, _018041_, _018043_);
  xor g_110294_(out[198], _017969_, _018044_);
  not g_110295_(_018044_, _018045_);
  and g_110296_(_017818_, _017964_, _018046_);
  or g_110297_(_017817_, _017963_, _018047_);
  and g_110298_(_017811_, _017963_, _018048_);
  or g_110299_(_017812_, _017964_, _018049_);
  and g_110300_(_018047_, _018049_, _018051_);
  or g_110301_(_018046_, _018048_, _018052_);
  and g_110302_(_018044_, _018051_, _018053_);
  or g_110303_(_018045_, _018052_, _018054_);
  and g_110304_(_018033_, _018041_, _018055_);
  or g_110305_(_018034_, _018040_, _018056_);
  and g_110306_(_018054_, _018056_, _018057_);
  or g_110307_(_018053_, _018055_, _018058_);
  and g_110308_(_018043_, _018058_, _018059_);
  not g_110309_(_018059_, _018060_);
  xor g_110310_(_003915_, _017968_, _018062_);
  or g_110311_(_017861_, _017963_, _018063_);
  or g_110312_(_017855_, _017964_, _018064_);
  and g_110313_(_018063_, _018064_, _018065_);
  and g_110314_(_018062_, _018065_, _018066_);
  not g_110315_(_018066_, _018067_);
  or g_110316_(_018044_, _018051_, _018068_);
  not g_110317_(_018068_, _018069_);
  and g_110318_(_018043_, _018068_, _018070_);
  and g_110319_(_018067_, _018070_, _018071_);
  or g_110320_(_018058_, _018069_, _018073_);
  or g_110321_(_018042_, _018073_, _018074_);
  and g_110322_(_018057_, _018071_, _018075_);
  or g_110323_(_018066_, _018074_, _018076_);
  or g_110324_(_018062_, _018065_, _018077_);
  not g_110325_(_018077_, _018078_);
  xor g_110326_(out[196], out[195], _018079_);
  or g_110327_(_017845_, _017964_, _018080_);
  or g_110328_(_017850_, _017963_, _018081_);
  and g_110329_(_018080_, _018081_, _018082_);
  or g_110330_(_018079_, _018082_, _018084_);
  not g_110331_(_018084_, _018085_);
  and g_110332_(_018077_, _018084_, _018086_);
  or g_110333_(_018078_, _018085_, _018087_);
  and g_110334_(_018075_, _018087_, _018088_);
  or g_110335_(_018076_, _018086_, _018089_);
  and g_110336_(_018060_, _018089_, _018090_);
  or g_110337_(_018059_, _018088_, _018091_);
  and g_110338_(_018031_, _018091_, _018092_);
  or g_110339_(_018032_, _018090_, _018093_);
  and g_110340_(_018079_, _018082_, _018095_);
  or g_110341_(_018087_, _018095_, _018096_);
  or g_110342_(_018076_, _018096_, _018097_);
  not g_110343_(_018097_, _018098_);
  and g_110344_(_018031_, _018098_, _018099_);
  or g_110345_(_018032_, _018097_, _018100_);
  or g_110346_(_003838_, _017964_, _018101_);
  not g_110347_(_018101_, _018102_);
  and g_110348_(_017882_, _017964_, _018103_);
  or g_110349_(_017881_, _017963_, _018104_);
  and g_110350_(_018101_, _018104_, _018106_);
  or g_110351_(_018102_, _018103_, _018107_);
  and g_110352_(out[195], _018106_, _018108_);
  not g_110353_(_018108_, _018109_);
  and g_110354_(_017891_, _017964_, _018110_);
  and g_110355_(_003827_, _017963_, _018111_);
  or g_110356_(_018110_, _018111_, _018112_);
  or g_110357_(out[194], _018112_, _018113_);
  and g_110358_(_003970_, _018107_, _018114_);
  xor g_110359_(_003959_, _018112_, _018115_);
  or g_110360_(_018114_, _018115_, _018117_);
  or g_110361_(_018108_, _018117_, _018118_);
  or g_110362_(out[193], _017967_, _018119_);
  and g_110363_(_017913_, _017964_, _018120_);
  or g_110364_(_017912_, _017963_, _018121_);
  or g_110365_(out[176], _017964_, _018122_);
  not g_110366_(_018122_, _018123_);
  and g_110367_(_018121_, _018122_, _018124_);
  or g_110368_(_018120_, _018123_, _018125_);
  and g_110369_(out[192], _018125_, _018126_);
  xor g_110370_(_003937_, _017967_, _018128_);
  or g_110371_(_018126_, _018128_, _018129_);
  and g_110372_(_018119_, _018129_, _018130_);
  or g_110373_(_018118_, _018130_, _018131_);
  or g_110374_(_018113_, _018114_, _018132_);
  and g_110375_(_018131_, _018132_, _018133_);
  not g_110376_(_018133_, _018134_);
  and g_110377_(_018109_, _018133_, _018135_);
  or g_110378_(_018108_, _018134_, _018136_);
  and g_110379_(_018099_, _018136_, _018137_);
  or g_110380_(_018100_, _018135_, _018139_);
  and g_110381_(_017994_, _017999_, _018140_);
  not g_110382_(_018140_, _018141_);
  or g_110383_(_018013_, _018024_, _018142_);
  not g_110384_(_018142_, _018143_);
  and g_110385_(_018141_, _018142_, _018144_);
  and g_110386_(_018139_, _018144_, _018145_);
  or g_110387_(_018092_, _018143_, _018146_);
  or g_110388_(_018137_, _018146_, _018147_);
  and g_110389_(_018093_, _018145_, _018148_);
  or g_110390_(_018140_, _018147_, _018150_);
  or g_110391_(out[192], _018125_, _018151_);
  not g_110392_(_018151_, _018152_);
  or g_110393_(_018118_, _018129_, _018153_);
  or g_110394_(_018100_, _018153_, _018154_);
  not g_110395_(_018154_, _018155_);
  and g_110396_(_018151_, _018155_, _018156_);
  or g_110397_(_018152_, _018154_, _018157_);
  and g_110398_(_018150_, _018157_, _018158_);
  or g_110399_(_018148_, _018156_, _018159_);
  and g_110400_(_017967_, _018159_, _018161_);
  and g_110401_(_003937_, _018158_, _018162_);
  or g_110402_(_018161_, _018162_, _018163_);
  and g_110403_(out[212], out[211], _018164_);
  or g_110404_(out[213], _018164_, _018165_);
  or g_110405_(out[214], _018165_, _018166_);
  or g_110406_(out[215], _018166_, _018167_);
  or g_110407_(out[216], _018167_, _018168_);
  and g_110408_(out[217], _018168_, _018169_);
  or g_110409_(out[218], _018169_, _018170_);
  xor g_110410_(out[218], _018169_, _018172_);
  not g_110411_(_018172_, _018173_);
  and g_110412_(_017976_, _018158_, _018174_);
  not g_110413_(_018174_, _018175_);
  or g_110414_(_017982_, _018158_, _018176_);
  not g_110415_(_018176_, _018177_);
  and g_110416_(_018175_, _018176_, _018178_);
  or g_110417_(_018174_, _018177_, _018179_);
  and g_110418_(_018172_, _018178_, _018180_);
  or g_110419_(_018173_, _018179_, _018181_);
  and g_110420_(_017987_, _017989_, _018183_);
  or g_110421_(_017988_, _017990_, _018184_);
  xor g_110422_(out[219], _018170_, _018185_);
  xor g_110423_(_003992_, _018170_, _018186_);
  and g_110424_(_018183_, _018186_, _018187_);
  or g_110425_(_018184_, _018185_, _018188_);
  and g_110426_(_018181_, _018188_, _018189_);
  or g_110427_(_018180_, _018187_, _018190_);
  and g_110428_(_018184_, _018185_, _018191_);
  and g_110429_(_018173_, _018179_, _018192_);
  or g_110430_(_018191_, _018192_, _018194_);
  or g_110431_(_018190_, _018194_, _018195_);
  xor g_110432_(out[216], _018167_, _018196_);
  not g_110433_(_018196_, _018197_);
  and g_110434_(_018016_, _018158_, _018198_);
  not g_110435_(_018198_, _018199_);
  or g_110436_(_018021_, _018158_, _018200_);
  not g_110437_(_018200_, _018201_);
  and g_110438_(_018199_, _018200_, _018202_);
  or g_110439_(_018198_, _018201_, _018203_);
  or g_110440_(_018197_, _018202_, _018205_);
  and g_110441_(_018004_, _018158_, _018206_);
  not g_110442_(_018206_, _018207_);
  or g_110443_(_018003_, _018158_, _018208_);
  not g_110444_(_018208_, _018209_);
  and g_110445_(_018207_, _018208_, _018210_);
  or g_110446_(_018206_, _018209_, _018211_);
  xor g_110447_(out[217], _018168_, _018212_);
  or g_110448_(_018210_, _018212_, _018213_);
  and g_110449_(_018205_, _018213_, _018214_);
  not g_110450_(_018214_, _018216_);
  and g_110451_(_018210_, _018212_, _018217_);
  and g_110452_(_018197_, _018202_, _018218_);
  or g_110453_(_018217_, _018218_, _018219_);
  or g_110454_(_018216_, _018219_, _018220_);
  or g_110455_(_018195_, _018220_, _018221_);
  xor g_110456_(out[215], _018166_, _018222_);
  not g_110457_(_018222_, _018223_);
  and g_110458_(_018034_, _018158_, _018224_);
  or g_110459_(_018033_, _018159_, _018225_);
  and g_110460_(_018041_, _018159_, _018227_);
  or g_110461_(_018040_, _018158_, _018228_);
  and g_110462_(_018225_, _018228_, _018229_);
  or g_110463_(_018224_, _018227_, _018230_);
  or g_110464_(_018223_, _018229_, _018231_);
  and g_110465_(_018223_, _018229_, _018232_);
  xor g_110466_(_018222_, _018229_, _018233_);
  xor g_110467_(out[214], _018165_, _018234_);
  not g_110468_(_018234_, _018235_);
  and g_110469_(_018044_, _018158_, _018236_);
  and g_110470_(_018052_, _018159_, _018238_);
  or g_110471_(_018236_, _018238_, _018239_);
  or g_110472_(_018235_, _018239_, _018240_);
  xor g_110473_(_018234_, _018239_, _018241_);
  or g_110474_(_018233_, _018241_, _018242_);
  xor g_110475_(out[212], out[211], _018243_);
  and g_110476_(_018079_, _018158_, _018244_);
  not g_110477_(_018244_, _018245_);
  or g_110478_(_018082_, _018158_, _018246_);
  not g_110479_(_018246_, _018247_);
  and g_110480_(_018245_, _018246_, _018249_);
  or g_110481_(_018244_, _018247_, _018250_);
  or g_110482_(_018243_, _018249_, _018251_);
  xor g_110483_(out[213], _018164_, _018252_);
  xor g_110484_(_004025_, _018164_, _018253_);
  and g_110485_(_018062_, _018158_, _018254_);
  not g_110486_(_018254_, _018255_);
  or g_110487_(_018065_, _018158_, _018256_);
  not g_110488_(_018256_, _018257_);
  and g_110489_(_018255_, _018256_, _018258_);
  or g_110490_(_018254_, _018257_, _018260_);
  or g_110491_(_018253_, _018258_, _018261_);
  and g_110492_(_018251_, _018261_, _018262_);
  not g_110493_(_018262_, _018263_);
  and g_110494_(_018253_, _018258_, _018264_);
  and g_110495_(_018243_, _018249_, _018265_);
  or g_110496_(_018264_, _018265_, _018266_);
  or g_110497_(_018242_, _018263_, _018267_);
  or g_110498_(_018266_, _018267_, _018268_);
  or g_110499_(_018221_, _018268_, _018269_);
  and g_110500_(_018112_, _018159_, _018271_);
  and g_110501_(_003959_, _018158_, _018272_);
  or g_110502_(_018271_, _018272_, _018273_);
  or g_110503_(out[210], _018273_, _018274_);
  and g_110504_(out[195], _018158_, _018275_);
  not g_110505_(_018275_, _018276_);
  or g_110506_(_018106_, _018158_, _018277_);
  not g_110507_(_018277_, _018278_);
  and g_110508_(_018276_, _018277_, _018279_);
  or g_110509_(_018275_, _018278_, _018280_);
  or g_110510_(_004080_, _018280_, _018282_);
  and g_110511_(_018274_, _018282_, _018283_);
  and g_110512_(_004080_, _018280_, _018284_);
  xor g_110513_(_004069_, _018273_, _018285_);
  xor g_110514_(_004080_, _018279_, _018286_);
  or g_110515_(_018285_, _018286_, _018287_);
  or g_110516_(out[209], _018163_, _018288_);
  and g_110517_(out[192], _018158_, _018289_);
  not g_110518_(_018289_, _018290_);
  and g_110519_(_018124_, _018159_, _018291_);
  or g_110520_(_018125_, _018158_, _018293_);
  or g_110521_(_018289_, _018291_, _018294_);
  and g_110522_(_018290_, _018293_, _018295_);
  and g_110523_(out[208], _018295_, _018296_);
  xor g_110524_(_004047_, _018163_, _018297_);
  or g_110525_(_018296_, _018297_, _018298_);
  and g_110526_(_018288_, _018298_, _018299_);
  or g_110527_(_018287_, _018299_, _018300_);
  or g_110528_(_018283_, _018284_, _018301_);
  and g_110529_(_018300_, _018301_, _018302_);
  or g_110530_(_018269_, _018302_, _018304_);
  or g_110531_(_018242_, _018262_, _018305_);
  or g_110532_(_018264_, _018305_, _018306_);
  and g_110533_(_018231_, _018240_, _018307_);
  or g_110534_(_018232_, _018307_, _018308_);
  and g_110535_(_018306_, _018308_, _018309_);
  or g_110536_(_018221_, _018309_, _018310_);
  or g_110537_(_018214_, _018217_, _018311_);
  or g_110538_(_018195_, _018311_, _018312_);
  or g_110539_(_018189_, _018191_, _018313_);
  and g_110540_(_018312_, _018313_, _018315_);
  and g_110541_(_018310_, _018315_, _018316_);
  and g_110542_(_018304_, _018316_, _018317_);
  and g_110543_(_004058_, _018294_, _018318_);
  or g_110544_(_018287_, _018298_, _018319_);
  or g_110545_(_018318_, _018319_, _018320_);
  or g_110546_(_018269_, _018320_, _018321_);
  not g_110547_(_018321_, _018322_);
  or g_110548_(_018317_, _018322_, _018323_);
  not g_110549_(_018323_, _018324_);
  and g_110550_(_018163_, _018323_, _018326_);
  and g_110551_(_004047_, _018324_, _018327_);
  or g_110552_(_018326_, _018327_, _018328_);
  and g_110553_(_018172_, _018324_, _018329_);
  or g_110554_(_018173_, _018323_, _018330_);
  and g_110555_(_018179_, _018323_, _018331_);
  or g_110556_(_018178_, _018324_, _018332_);
  and g_110557_(_018330_, _018332_, _018333_);
  or g_110558_(_018329_, _018331_, _018334_);
  and g_110559_(out[228], out[227], _018335_);
  or g_110560_(out[229], _018335_, _018337_);
  or g_110561_(out[230], _018337_, _018338_);
  or g_110562_(out[231], _018338_, _018339_);
  or g_110563_(out[232], _018339_, _018340_);
  and g_110564_(out[233], _018340_, _018341_);
  or g_110565_(out[234], _018341_, _018342_);
  xor g_110566_(out[234], _018341_, _018343_);
  not g_110567_(_018343_, _018344_);
  or g_110568_(_018334_, _018344_, _018345_);
  and g_110569_(_018183_, _018185_, _018346_);
  or g_110570_(_018184_, _018186_, _018348_);
  xor g_110571_(out[235], _018342_, _018349_);
  xor g_110572_(_004124_, _018342_, _018350_);
  or g_110573_(_018348_, _018349_, _018351_);
  and g_110574_(_018345_, _018351_, _018352_);
  or g_110575_(_018333_, _018343_, _018353_);
  and g_110576_(_018348_, _018349_, _018354_);
  and g_110577_(_018210_, _018323_, _018355_);
  or g_110578_(_018211_, _018324_, _018356_);
  or g_110579_(_018212_, _018323_, _018357_);
  not g_110580_(_018357_, _018359_);
  or g_110581_(_018355_, _018359_, _018360_);
  and g_110582_(_018356_, _018357_, _018361_);
  xor g_110583_(out[233], _018340_, _018362_);
  and g_110584_(_018360_, _018362_, _018363_);
  not g_110585_(_018363_, _018364_);
  xor g_110586_(out[232], _018339_, _018365_);
  not g_110587_(_018365_, _018366_);
  or g_110588_(_018196_, _018323_, _018367_);
  not g_110589_(_018367_, _018368_);
  and g_110590_(_018203_, _018323_, _018370_);
  or g_110591_(_018202_, _018324_, _018371_);
  and g_110592_(_018367_, _018371_, _018372_);
  or g_110593_(_018368_, _018370_, _018373_);
  or g_110594_(_018366_, _018372_, _018374_);
  or g_110595_(_018360_, _018362_, _018375_);
  and g_110596_(_018374_, _018375_, _018376_);
  not g_110597_(_018376_, _018377_);
  and g_110598_(_018366_, _018372_, _018378_);
  or g_110599_(_018365_, _018373_, _018379_);
  and g_110600_(_018352_, _018353_, _018381_);
  not g_110601_(_018381_, _018382_);
  or g_110602_(_018354_, _018382_, _018383_);
  not g_110603_(_018383_, _018384_);
  and g_110604_(_018364_, _018379_, _018385_);
  or g_110605_(_018363_, _018378_, _018386_);
  and g_110606_(_018376_, _018385_, _018387_);
  or g_110607_(_018377_, _018386_, _018388_);
  and g_110608_(_018384_, _018387_, _018389_);
  or g_110609_(_018383_, _018388_, _018390_);
  xor g_110610_(out[230], _018337_, _018392_);
  not g_110611_(_018392_, _018393_);
  and g_110612_(_018234_, _018324_, _018394_);
  or g_110613_(_018235_, _018323_, _018395_);
  and g_110614_(_018239_, _018323_, _018396_);
  not g_110615_(_018396_, _018397_);
  and g_110616_(_018395_, _018397_, _018398_);
  or g_110617_(_018394_, _018396_, _018399_);
  and g_110618_(_018392_, _018398_, _018400_);
  or g_110619_(_018393_, _018399_, _018401_);
  xor g_110620_(out[231], _018338_, _018403_);
  not g_110621_(_018403_, _018404_);
  or g_110622_(_018222_, _018323_, _018405_);
  not g_110623_(_018405_, _018406_);
  and g_110624_(_018230_, _018323_, _018407_);
  or g_110625_(_018229_, _018324_, _018408_);
  and g_110626_(_018405_, _018408_, _018409_);
  or g_110627_(_018406_, _018407_, _018410_);
  and g_110628_(_018403_, _018410_, _018411_);
  or g_110629_(_018404_, _018409_, _018412_);
  and g_110630_(_018401_, _018412_, _018414_);
  or g_110631_(_018400_, _018411_, _018415_);
  and g_110632_(_018404_, _018409_, _018416_);
  and g_110633_(_018393_, _018399_, _018417_);
  or g_110634_(_018416_, _018417_, _018418_);
  or g_110635_(_018415_, _018418_, _018419_);
  xor g_110636_(out[229], _018335_, _018420_);
  xor g_110637_(_004157_, _018335_, _018421_);
  or g_110638_(_018252_, _018323_, _018422_);
  not g_110639_(_018422_, _018423_);
  and g_110640_(_018260_, _018323_, _018425_);
  or g_110641_(_018258_, _018324_, _018426_);
  and g_110642_(_018422_, _018426_, _018427_);
  or g_110643_(_018423_, _018425_, _018428_);
  or g_110644_(_018421_, _018427_, _018429_);
  xor g_110645_(out[228], out[227], _018430_);
  and g_110646_(_018249_, _018323_, _018431_);
  or g_110647_(_018250_, _018324_, _018432_);
  or g_110648_(_018243_, _018323_, _018433_);
  not g_110649_(_018433_, _018434_);
  or g_110650_(_018431_, _018434_, _018436_);
  and g_110651_(_018432_, _018433_, _018437_);
  or g_110652_(_018430_, _018436_, _018438_);
  and g_110653_(_018429_, _018438_, _018439_);
  not g_110654_(_018439_, _018440_);
  and g_110655_(_018421_, _018427_, _018441_);
  not g_110656_(_018441_, _018442_);
  and g_110657_(_018430_, _018436_, _018443_);
  and g_110658_(_018439_, _018442_, _018444_);
  or g_110659_(_018440_, _018441_, _018445_);
  or g_110660_(_018419_, _018443_, _018447_);
  not g_110661_(_018447_, _018448_);
  and g_110662_(_018444_, _018448_, _018449_);
  or g_110663_(_018445_, _018447_, _018450_);
  and g_110664_(_018295_, _018323_, _018451_);
  and g_110665_(_004058_, _018324_, _018452_);
  or g_110666_(_018451_, _018452_, _018453_);
  and g_110667_(out[224], _018453_, _018454_);
  not g_110668_(_018454_, _018455_);
  or g_110669_(out[225], _018328_, _018456_);
  xor g_110670_(out[225], _018328_, _018458_);
  xor g_110671_(_004179_, _018328_, _018459_);
  and g_110672_(_018455_, _018458_, _018460_);
  or g_110673_(_018454_, _018459_, _018461_);
  or g_110674_(out[224], _018453_, _018462_);
  and g_110675_(out[211], _018324_, _018463_);
  or g_110676_(_004080_, _018323_, _018464_);
  and g_110677_(_018280_, _018323_, _018465_);
  or g_110678_(_018279_, _018324_, _018466_);
  and g_110679_(_018464_, _018466_, _018467_);
  or g_110680_(_018463_, _018465_, _018469_);
  or g_110681_(_004212_, _018469_, _018470_);
  and g_110682_(_018273_, _018323_, _018471_);
  and g_110683_(_004069_, _018324_, _018472_);
  or g_110684_(_018471_, _018472_, _018473_);
  and g_110685_(_004212_, _018469_, _018474_);
  or g_110686_(out[226], _018473_, _018475_);
  xor g_110687_(out[227], _018467_, _018476_);
  xor g_110688_(_004212_, _018467_, _018477_);
  xor g_110689_(out[226], _018473_, _018478_);
  xor g_110690_(_004201_, _018473_, _018480_);
  and g_110691_(_018476_, _018478_, _018481_);
  or g_110692_(_018477_, _018480_, _018482_);
  and g_110693_(_018462_, _018481_, _018483_);
  and g_110694_(_018460_, _018483_, _018484_);
  and g_110695_(_018449_, _018484_, _018485_);
  and g_110696_(_018389_, _018485_, _018486_);
  and g_110697_(_018456_, _018461_, _018487_);
  or g_110698_(_018482_, _018487_, _018488_);
  or g_110699_(_018474_, _018475_, _018489_);
  and g_110700_(_018470_, _018489_, _018491_);
  and g_110701_(_018488_, _018491_, _018492_);
  or g_110702_(_018450_, _018492_, _018493_);
  or g_110703_(_018414_, _018416_, _018494_);
  or g_110704_(_018439_, _018441_, _018495_);
  or g_110705_(_018419_, _018495_, _018496_);
  and g_110706_(_018494_, _018496_, _018497_);
  and g_110707_(_018493_, _018497_, _018498_);
  or g_110708_(_018390_, _018498_, _018499_);
  or g_110709_(_018363_, _018376_, _018500_);
  or g_110710_(_018383_, _018500_, _018502_);
  or g_110711_(_018352_, _018354_, _018503_);
  and g_110712_(_018502_, _018503_, _018504_);
  and g_110713_(_018499_, _018504_, _018505_);
  or g_110714_(_018486_, _018505_, _018506_);
  not g_110715_(_018506_, _018507_);
  and g_110716_(_018328_, _018506_, _018508_);
  not g_110717_(_018508_, _018509_);
  or g_110718_(out[225], _018506_, _018510_);
  not g_110719_(_018510_, _018511_);
  and g_110720_(_018509_, _018510_, _018513_);
  or g_110721_(_018508_, _018511_, _018514_);
  and g_110722_(_018346_, _018349_, _018515_);
  or g_110723_(_018348_, _018350_, _018516_);
  and g_110724_(out[244], out[243], _018517_);
  or g_110725_(out[245], _018517_, _018518_);
  or g_110726_(out[246], _018518_, _018519_);
  or g_110727_(out[247], _018519_, _018520_);
  or g_110728_(out[248], _018520_, _018521_);
  and g_110729_(out[249], _018521_, _018522_);
  or g_110730_(out[250], _018522_, _018524_);
  xor g_110731_(out[251], _018524_, _018525_);
  xor g_110732_(_004245_, _018524_, _018526_);
  and g_110733_(_018515_, _018526_, _018527_);
  or g_110734_(_018516_, _018525_, _018528_);
  and g_110735_(_018334_, _018506_, _018529_);
  or g_110736_(_018333_, _018507_, _018530_);
  and g_110737_(_018343_, _018507_, _018531_);
  or g_110738_(_018344_, _018506_, _018532_);
  and g_110739_(_018530_, _018532_, _018533_);
  or g_110740_(_018529_, _018531_, _018535_);
  xor g_110741_(out[250], _018522_, _018536_);
  xor g_110742_(_004355_, _018522_, _018537_);
  and g_110743_(_018533_, _018536_, _018538_);
  or g_110744_(_018535_, _018537_, _018539_);
  and g_110745_(_018528_, _018539_, _018540_);
  or g_110746_(_018527_, _018538_, _018541_);
  and g_110747_(_018535_, _018537_, _018542_);
  or g_110748_(_018533_, _018536_, _018543_);
  and g_110749_(_018516_, _018525_, _018544_);
  or g_110750_(_018515_, _018526_, _018546_);
  and g_110751_(_018360_, _018506_, _018547_);
  or g_110752_(_018361_, _018507_, _018548_);
  or g_110753_(_018362_, _018506_, _018549_);
  not g_110754_(_018549_, _018550_);
  or g_110755_(_018547_, _018550_, _018551_);
  and g_110756_(_018548_, _018549_, _018552_);
  xor g_110757_(out[249], _018521_, _018553_);
  xor g_110758_(_004344_, _018521_, _018554_);
  and g_110759_(_018551_, _018553_, _018555_);
  or g_110760_(_018552_, _018554_, _018557_);
  xor g_110761_(out[248], _018520_, _018558_);
  xor g_110762_(_004333_, _018520_, _018559_);
  and g_110763_(_018373_, _018506_, _018560_);
  or g_110764_(_018372_, _018507_, _018561_);
  or g_110765_(_018365_, _018506_, _018562_);
  not g_110766_(_018562_, _018563_);
  and g_110767_(_018561_, _018562_, _018564_);
  or g_110768_(_018560_, _018563_, _018565_);
  and g_110769_(_018558_, _018565_, _018566_);
  or g_110770_(_018559_, _018564_, _018568_);
  and g_110771_(_018552_, _018554_, _018569_);
  or g_110772_(_018551_, _018553_, _018570_);
  and g_110773_(_018568_, _018570_, _018571_);
  or g_110774_(_018566_, _018569_, _018572_);
  and g_110775_(_018559_, _018564_, _018573_);
  or g_110776_(_018558_, _018565_, _018574_);
  and g_110777_(_018543_, _018546_, _018575_);
  or g_110778_(_018542_, _018544_, _018576_);
  and g_110779_(_018540_, _018575_, _018577_);
  or g_110780_(_018541_, _018576_, _018579_);
  and g_110781_(_018557_, _018574_, _018580_);
  or g_110782_(_018555_, _018573_, _018581_);
  and g_110783_(_018571_, _018580_, _018582_);
  or g_110784_(_018572_, _018581_, _018583_);
  and g_110785_(_018577_, _018582_, _018584_);
  or g_110786_(_018579_, _018583_, _018585_);
  xor g_110787_(out[247], _018519_, _018586_);
  xor g_110788_(_004256_, _018519_, _018587_);
  and g_110789_(_018410_, _018506_, _018588_);
  or g_110790_(_018409_, _018507_, _018590_);
  or g_110791_(_018403_, _018506_, _018591_);
  not g_110792_(_018591_, _018592_);
  and g_110793_(_018590_, _018591_, _018593_);
  or g_110794_(_018588_, _018592_, _018594_);
  and g_110795_(_018586_, _018594_, _018595_);
  xor g_110796_(out[246], _018518_, _018596_);
  not g_110797_(_018596_, _018597_);
  and g_110798_(_018399_, _018506_, _018598_);
  or g_110799_(_018398_, _018507_, _018599_);
  and g_110800_(_018392_, _018507_, _018601_);
  or g_110801_(_018393_, _018506_, _018602_);
  and g_110802_(_018599_, _018602_, _018603_);
  or g_110803_(_018598_, _018601_, _018604_);
  and g_110804_(_018596_, _018603_, _018605_);
  or g_110805_(_018595_, _018605_, _018606_);
  and g_110806_(_018597_, _018604_, _018607_);
  and g_110807_(_018587_, _018593_, _018608_);
  or g_110808_(_018586_, _018594_, _018609_);
  or g_110809_(_018607_, _018608_, _018610_);
  xor g_110810_(_018596_, _018603_, _018612_);
  xor g_110811_(_018587_, _018593_, _018613_);
  and g_110812_(_018612_, _018613_, _018614_);
  or g_110813_(_018606_, _018610_, _018615_);
  xor g_110814_(out[244], out[243], _018616_);
  xor g_110815_(_004289_, out[243], _018617_);
  and g_110816_(_018436_, _018506_, _018618_);
  or g_110817_(_018437_, _018507_, _018619_);
  or g_110818_(_018430_, _018506_, _018620_);
  not g_110819_(_018620_, _018621_);
  or g_110820_(_018618_, _018621_, _018623_);
  and g_110821_(_018619_, _018620_, _018624_);
  and g_110822_(_018617_, _018624_, _018625_);
  or g_110823_(_018616_, _018623_, _018626_);
  xor g_110824_(out[245], _018517_, _018627_);
  xor g_110825_(_004278_, _018517_, _018628_);
  and g_110826_(_018428_, _018506_, _018629_);
  or g_110827_(_018427_, _018507_, _018630_);
  or g_110828_(_018420_, _018506_, _018631_);
  not g_110829_(_018631_, _018632_);
  and g_110830_(_018630_, _018631_, _018634_);
  or g_110831_(_018629_, _018632_, _018635_);
  and g_110832_(_018627_, _018635_, _018636_);
  or g_110833_(_018628_, _018634_, _018637_);
  and g_110834_(_018626_, _018637_, _018638_);
  or g_110835_(_018625_, _018636_, _018639_);
  and g_110836_(_018628_, _018634_, _018640_);
  or g_110837_(_018627_, _018635_, _018641_);
  and g_110838_(_018616_, _018623_, _018642_);
  or g_110839_(_018617_, _018624_, _018643_);
  and g_110840_(_018641_, _018643_, _018645_);
  or g_110841_(_018640_, _018642_, _018646_);
  and g_110842_(_018638_, _018645_, _018647_);
  or g_110843_(_018639_, _018646_, _018648_);
  and g_110844_(_018614_, _018647_, _018649_);
  or g_110845_(_018615_, _018648_, _018650_);
  and g_110846_(_018584_, _018649_, _018651_);
  or g_110847_(_018585_, _018650_, _018652_);
  and g_110848_(_018469_, _018506_, _018653_);
  or g_110849_(_018467_, _018507_, _018654_);
  and g_110850_(out[227], _018507_, _018656_);
  or g_110851_(_004212_, _018506_, _018657_);
  and g_110852_(_018654_, _018657_, _018658_);
  or g_110853_(_018653_, _018656_, _018659_);
  and g_110854_(out[243], _018658_, _018660_);
  or g_110855_(_004322_, _018659_, _018661_);
  and g_110856_(_018473_, _018506_, _018662_);
  not g_110857_(_018662_, _018663_);
  or g_110858_(out[226], _018506_, _018664_);
  not g_110859_(_018664_, _018665_);
  and g_110860_(_018663_, _018664_, _018667_);
  or g_110861_(_018662_, _018665_, _018668_);
  and g_110862_(out[242], _018668_, _018669_);
  or g_110863_(_004311_, _018667_, _018670_);
  and g_110864_(_018661_, _018670_, _018671_);
  or g_110865_(_018660_, _018669_, _018672_);
  and g_110866_(_004322_, _018659_, _018673_);
  or g_110867_(out[243], _018658_, _018674_);
  and g_110868_(_004311_, _018667_, _018675_);
  or g_110869_(out[242], _018668_, _018676_);
  and g_110870_(_018674_, _018676_, _018678_);
  or g_110871_(_018673_, _018675_, _018679_);
  and g_110872_(_018671_, _018678_, _018680_);
  or g_110873_(_018672_, _018679_, _018681_);
  or g_110874_(out[241], _018514_, _018682_);
  and g_110875_(_018453_, _018506_, _018683_);
  not g_110876_(_018683_, _018684_);
  or g_110877_(out[224], _018506_, _018685_);
  not g_110878_(_018685_, _018686_);
  and g_110879_(_018684_, _018685_, _018687_);
  or g_110880_(_018683_, _018686_, _018689_);
  and g_110881_(out[240], _018689_, _018690_);
  xor g_110882_(out[241], _018513_, _018691_);
  or g_110883_(_018690_, _018691_, _018692_);
  not g_110884_(_018692_, _018693_);
  and g_110885_(_018682_, _018692_, _018694_);
  not g_110886_(_018694_, _018695_);
  and g_110887_(_018680_, _018695_, _018696_);
  or g_110888_(_018681_, _018694_, _018697_);
  and g_110889_(_018674_, _018675_, _018698_);
  or g_110890_(_018673_, _018676_, _018700_);
  and g_110891_(_018661_, _018700_, _018701_);
  or g_110892_(_018660_, _018698_, _018702_);
  and g_110893_(_018697_, _018701_, _018703_);
  or g_110894_(_018696_, _018702_, _018704_);
  and g_110895_(_018651_, _018704_, _018705_);
  or g_110896_(_018652_, _018703_, _018706_);
  or g_110897_(_018638_, _018640_, _018707_);
  and g_110898_(_018614_, _018639_, _018708_);
  and g_110899_(_018641_, _018708_, _018709_);
  or g_110900_(_018615_, _018707_, _018711_);
  and g_110901_(_018606_, _018609_, _018712_);
  not g_110902_(_018712_, _018713_);
  and g_110903_(_018711_, _018713_, _018714_);
  or g_110904_(_018709_, _018712_, _018715_);
  and g_110905_(_018584_, _018715_, _018716_);
  or g_110906_(_018585_, _018714_, _018717_);
  and g_110907_(_018557_, _018572_, _018718_);
  or g_110908_(_018555_, _018571_, _018719_);
  and g_110909_(_018577_, _018718_, _018720_);
  or g_110910_(_018579_, _018719_, _018722_);
  and g_110911_(_018541_, _018546_, _018723_);
  or g_110912_(_018540_, _018544_, _018724_);
  and g_110913_(_018722_, _018724_, _018725_);
  or g_110914_(_018720_, _018723_, _018726_);
  or g_110915_(_018716_, _018726_, _018727_);
  and g_110916_(_018706_, _018725_, _018728_);
  and g_110917_(_018717_, _018728_, _018729_);
  or g_110918_(_018705_, _018727_, _018730_);
  and g_110919_(_004300_, _018687_, _018731_);
  or g_110920_(out[240], _018689_, _018733_);
  and g_110921_(_018680_, _018733_, _018734_);
  or g_110922_(_018681_, _018731_, _018735_);
  and g_110923_(_018693_, _018734_, _018736_);
  or g_110924_(_018692_, _018735_, _018737_);
  and g_110925_(_018651_, _018736_, _018738_);
  or g_110926_(_018652_, _018737_, _018739_);
  and g_110927_(_018730_, _018739_, _018740_);
  or g_110928_(_018729_, _018738_, _018741_);
  and g_110929_(_018514_, _018741_, _018742_);
  or g_110930_(_018513_, _018740_, _018744_);
  and g_110931_(_053038_, _018740_, _018745_);
  or g_110932_(out[241], _018741_, _018746_);
  and g_110933_(_018744_, _018746_, _018747_);
  or g_110934_(_018742_, _018745_, _018748_);
  and g_110935_(out[260], out[259], _018749_);
  or g_110936_(out[261], _018749_, _018750_);
  or g_110937_(out[262], _018750_, _018751_);
  xor g_110938_(out[262], _018750_, _018752_);
  xor g_110939_(_052983_, _018750_, _018753_);
  and g_110940_(_018604_, _018741_, _018755_);
  or g_110941_(_018603_, _018740_, _018756_);
  and g_110942_(_018596_, _018740_, _018757_);
  or g_110943_(_018597_, _018741_, _018758_);
  and g_110944_(_018756_, _018758_, _018759_);
  or g_110945_(_018755_, _018757_, _018760_);
  and g_110946_(_018752_, _018759_, _018761_);
  or g_110947_(_018753_, _018760_, _018762_);
  or g_110948_(out[263], _018751_, _018763_);
  xor g_110949_(out[263], _018751_, _018764_);
  xor g_110950_(_004377_, _018751_, _018766_);
  and g_110951_(_018594_, _018741_, _018767_);
  or g_110952_(_018593_, _018740_, _018768_);
  and g_110953_(_018587_, _018740_, _018769_);
  or g_110954_(_018586_, _018741_, _018770_);
  and g_110955_(_018768_, _018770_, _018771_);
  or g_110956_(_018767_, _018769_, _018772_);
  and g_110957_(_018764_, _018772_, _018773_);
  or g_110958_(_018766_, _018771_, _018774_);
  and g_110959_(_018762_, _018774_, _018775_);
  or g_110960_(_018761_, _018773_, _018777_);
  and g_110961_(_018659_, _018741_, _018778_);
  or g_110962_(_018658_, _018740_, _018779_);
  and g_110963_(out[243], _018740_, _018780_);
  or g_110964_(_004322_, _018741_, _018781_);
  and g_110965_(_018779_, _018781_, _018782_);
  or g_110966_(_018778_, _018780_, _018783_);
  and g_110967_(out[259], _018782_, _018784_);
  or g_110968_(_053005_, _018783_, _018785_);
  and g_110969_(_018668_, _018741_, _018786_);
  or g_110970_(_018667_, _018740_, _018788_);
  and g_110971_(_004311_, _018740_, _018789_);
  or g_110972_(out[242], _018741_, _018790_);
  and g_110973_(_018788_, _018790_, _018791_);
  or g_110974_(_018786_, _018789_, _018792_);
  and g_110975_(out[258], _018792_, _018793_);
  or g_110976_(_053016_, _018791_, _018794_);
  and g_110977_(_018689_, _018741_, _018795_);
  or g_110978_(_018687_, _018740_, _018796_);
  and g_110979_(_004300_, _018740_, _018797_);
  or g_110980_(out[240], _018741_, _018799_);
  and g_110981_(_018796_, _018799_, _018800_);
  or g_110982_(_018795_, _018797_, _018801_);
  and g_110983_(out[256], _018801_, _018802_);
  or g_110984_(_004388_, _018800_, _018803_);
  and g_110985_(out[257], _018748_, _018804_);
  or g_110986_(_053027_, _018747_, _018805_);
  and g_110987_(_018803_, _018805_, _018806_);
  or g_110988_(_018802_, _018804_, _018807_);
  and g_110989_(_053016_, _018791_, _018808_);
  or g_110990_(out[258], _018792_, _018810_);
  and g_110991_(_053027_, _018747_, _018811_);
  or g_110992_(out[257], _018748_, _018812_);
  and g_110993_(_018810_, _018812_, _018813_);
  or g_110994_(_018808_, _018811_, _018814_);
  and g_110995_(_018807_, _018813_, _018815_);
  or g_110996_(_018806_, _018814_, _018816_);
  and g_110997_(_018794_, _018816_, _018817_);
  or g_110998_(_018793_, _018815_, _018818_);
  and g_110999_(_018785_, _018818_, _018819_);
  or g_111000_(_018784_, _018817_, _018821_);
  xor g_111001_(out[260], out[259], _018822_);
  xor g_111002_(_052994_, out[259], _018823_);
  and g_111003_(_018616_, _018740_, _018824_);
  and g_111004_(_018624_, _018741_, _018825_);
  or g_111005_(_018824_, _018825_, _018826_);
  not g_111006_(_018826_, _018827_);
  and g_111007_(_018822_, _018827_, _018828_);
  or g_111008_(_018823_, _018826_, _018829_);
  and g_111009_(_053005_, _018783_, _018830_);
  or g_111010_(out[259], _018782_, _018832_);
  and g_111011_(_018829_, _018832_, _018833_);
  or g_111012_(_018828_, _018830_, _018834_);
  and g_111013_(_018821_, _018833_, _018835_);
  or g_111014_(_018819_, _018834_, _018836_);
  xor g_111015_(out[261], _018749_, _018837_);
  and g_111016_(_018635_, _018741_, _018838_);
  and g_111017_(_018628_, _018740_, _018839_);
  or g_111018_(_018838_, _018839_, _018840_);
  and g_111019_(_018837_, _018840_, _018841_);
  not g_111020_(_018841_, _018843_);
  and g_111021_(_018823_, _018826_, _018844_);
  or g_111022_(_018822_, _018827_, _018845_);
  and g_111023_(_018843_, _018845_, _018846_);
  or g_111024_(_018841_, _018844_, _018847_);
  and g_111025_(_018836_, _018846_, _018848_);
  or g_111026_(_018835_, _018847_, _018849_);
  or g_111027_(_018837_, _018840_, _018850_);
  not g_111028_(_018850_, _018851_);
  and g_111029_(_018753_, _018760_, _018852_);
  or g_111030_(_018752_, _018759_, _018854_);
  and g_111031_(_018850_, _018854_, _018855_);
  or g_111032_(_018851_, _018852_, _018856_);
  and g_111033_(_018849_, _018855_, _018857_);
  or g_111034_(_018848_, _018856_, _018858_);
  and g_111035_(_018775_, _018858_, _018859_);
  or g_111036_(_018777_, _018857_, _018860_);
  or g_111037_(out[264], _018763_, _018861_);
  and g_111038_(out[265], _018861_, _018862_);
  or g_111039_(out[266], _018862_, _018863_);
  xor g_111040_(out[266], _018862_, _018865_);
  xor g_111041_(_004421_, _018862_, _018866_);
  and g_111042_(_018535_, _018741_, _018867_);
  and g_111043_(_018536_, _018740_, _018868_);
  or g_111044_(_018867_, _018868_, _018869_);
  not g_111045_(_018869_, _018870_);
  and g_111046_(_018865_, _018870_, _018871_);
  or g_111047_(_018866_, _018869_, _018872_);
  and g_111048_(_018515_, _018525_, _018873_);
  or g_111049_(_018516_, _018526_, _018874_);
  xor g_111050_(out[267], _018863_, _018876_);
  xor g_111051_(_004366_, _018863_, _018877_);
  and g_111052_(_018873_, _018877_, _018878_);
  or g_111053_(_018874_, _018876_, _018879_);
  and g_111054_(_018872_, _018879_, _018880_);
  or g_111055_(_018871_, _018878_, _018881_);
  and g_111056_(_018874_, _018876_, _018882_);
  or g_111057_(_018873_, _018877_, _018883_);
  and g_111058_(_018866_, _018869_, _018884_);
  or g_111059_(_018865_, _018870_, _018885_);
  or g_111060_(_018882_, _018884_, _018887_);
  and g_111061_(_018880_, _018885_, _018888_);
  and g_111062_(_018883_, _018888_, _018889_);
  or g_111063_(_018881_, _018887_, _018890_);
  xor g_111064_(out[264], _018763_, _018891_);
  not g_111065_(_018891_, _018892_);
  and g_111066_(_018565_, _018741_, _018893_);
  or g_111067_(_018564_, _018740_, _018894_);
  and g_111068_(_018559_, _018740_, _018895_);
  or g_111069_(_018558_, _018741_, _018896_);
  and g_111070_(_018894_, _018896_, _018898_);
  or g_111071_(_018893_, _018895_, _018899_);
  and g_111072_(_018891_, _018899_, _018900_);
  or g_111073_(_018892_, _018898_, _018901_);
  and g_111074_(_018552_, _018741_, _018902_);
  and g_111075_(_018553_, _018740_, _018903_);
  or g_111076_(_018902_, _018903_, _018904_);
  not g_111077_(_018904_, _018905_);
  xor g_111078_(out[265], _018861_, _018906_);
  xor g_111079_(_004410_, _018861_, _018907_);
  and g_111080_(_018904_, _018907_, _018909_);
  or g_111081_(_018905_, _018906_, _018910_);
  and g_111082_(_018901_, _018910_, _018911_);
  or g_111083_(_018900_, _018909_, _018912_);
  or g_111084_(_018904_, _018907_, _018913_);
  or g_111085_(_018891_, _018899_, _018914_);
  and g_111086_(_018913_, _018914_, _018915_);
  or g_111087_(_018764_, _018772_, _018916_);
  and g_111088_(_018915_, _018916_, _018917_);
  not g_111089_(_018917_, _018918_);
  and g_111090_(_018911_, _018917_, _018920_);
  or g_111091_(_018912_, _018918_, _018921_);
  and g_111092_(_018889_, _018920_, _018922_);
  or g_111093_(_018890_, _018921_, _018923_);
  and g_111094_(_018860_, _018922_, _018924_);
  or g_111095_(_018859_, _018923_, _018925_);
  and g_111096_(_018881_, _018883_, _018926_);
  or g_111097_(_018880_, _018882_, _018927_);
  and g_111098_(_018912_, _018913_, _018928_);
  not g_111099_(_018928_, _018929_);
  and g_111100_(_018889_, _018928_, _018931_);
  or g_111101_(_018890_, _018929_, _018932_);
  and g_111102_(_018927_, _018932_, _018933_);
  or g_111103_(_018926_, _018931_, _018934_);
  and g_111104_(_018925_, _018933_, _018935_);
  or g_111105_(_018924_, _018934_, _018936_);
  and g_111106_(_018813_, _018833_, _018937_);
  not g_111107_(_018937_, _018938_);
  and g_111108_(_018846_, _018855_, _018939_);
  or g_111109_(_018847_, _018856_, _018940_);
  and g_111110_(_018937_, _018939_, _018942_);
  or g_111111_(_018938_, _018940_, _018943_);
  and g_111112_(_004388_, _018800_, _018944_);
  or g_111113_(_018784_, _018793_, _018945_);
  or g_111114_(_018944_, _018945_, _018946_);
  or g_111115_(_018777_, _018807_, _018947_);
  or g_111116_(_018946_, _018947_, _018948_);
  not g_111117_(_018948_, _018949_);
  and g_111118_(_018942_, _018949_, _018950_);
  or g_111119_(_018943_, _018948_, _018951_);
  and g_111120_(_018922_, _018950_, _018953_);
  or g_111121_(_018923_, _018951_, _018954_);
  and g_111122_(_018936_, _018954_, _018955_);
  or g_111123_(_018935_, _018953_, _018956_);
  and g_111124_(_018748_, _018956_, _018957_);
  and g_111125_(_053027_, _018955_, _018958_);
  or g_111126_(_018957_, _018958_, _018959_);
  and g_111127_(out[275], out[276], _018960_);
  or g_111128_(out[277], _018960_, _018961_);
  or g_111129_(out[278], _018961_, _018962_);
  or g_111130_(out[279], _018962_, _018964_);
  or g_111131_(out[280], _018964_, _018965_);
  and g_111132_(out[281], _018965_, _018966_);
  or g_111133_(out[282], _018966_, _018967_);
  xor g_111134_(out[282], _018966_, _018968_);
  xor g_111135_(_004454_, _018966_, _018969_);
  or g_111136_(_018866_, _018956_, _018970_);
  not g_111137_(_018970_, _018971_);
  and g_111138_(_018869_, _018956_, _018972_);
  not g_111139_(_018972_, _018973_);
  and g_111140_(_018970_, _018973_, _018975_);
  or g_111141_(_018971_, _018972_, _018976_);
  and g_111142_(_018968_, _018975_, _018977_);
  or g_111143_(_018969_, _018976_, _018978_);
  and g_111144_(_018873_, _018876_, _018979_);
  or g_111145_(_018874_, _018877_, _018980_);
  xor g_111146_(out[283], _018967_, _018981_);
  xor g_111147_(_004432_, _018967_, _018982_);
  and g_111148_(_018979_, _018982_, _018983_);
  or g_111149_(_018980_, _018981_, _018984_);
  and g_111150_(_018978_, _018984_, _018986_);
  or g_111151_(_018977_, _018983_, _018987_);
  and g_111152_(_018980_, _018981_, _018988_);
  or g_111153_(_018979_, _018982_, _018989_);
  and g_111154_(_018969_, _018976_, _018990_);
  or g_111155_(_018968_, _018975_, _018991_);
  and g_111156_(_018989_, _018991_, _018992_);
  or g_111157_(_018988_, _018990_, _018993_);
  and g_111158_(_018986_, _018992_, _018994_);
  or g_111159_(_018987_, _018993_, _018995_);
  or g_111160_(_018891_, _018956_, _018997_);
  not g_111161_(_018997_, _018998_);
  and g_111162_(_018899_, _018956_, _018999_);
  not g_111163_(_018999_, _019000_);
  and g_111164_(_018997_, _019000_, _019001_);
  or g_111165_(_018998_, _018999_, _019002_);
  xor g_111166_(out[280], _018964_, _019003_);
  xor g_111167_(_053060_, _018964_, _019004_);
  and g_111168_(_019002_, _019003_, _019005_);
  or g_111169_(_019001_, _019004_, _019006_);
  or g_111170_(_018907_, _018956_, _019008_);
  not g_111171_(_019008_, _019009_);
  and g_111172_(_018904_, _018956_, _019010_);
  not g_111173_(_019010_, _019011_);
  and g_111174_(_019008_, _019011_, _019012_);
  or g_111175_(_019009_, _019010_, _019013_);
  xor g_111176_(out[281], _018965_, _019014_);
  xor g_111177_(_053137_, _018965_, _019015_);
  and g_111178_(_019013_, _019015_, _019016_);
  or g_111179_(_019012_, _019014_, _019017_);
  and g_111180_(_019006_, _019017_, _019019_);
  or g_111181_(_019005_, _019016_, _019020_);
  and g_111182_(_019012_, _019014_, _019021_);
  or g_111183_(_019013_, _019015_, _019022_);
  and g_111184_(_019001_, _019004_, _019023_);
  or g_111185_(_019002_, _019003_, _019024_);
  and g_111186_(_019022_, _019024_, _019025_);
  or g_111187_(_019021_, _019023_, _019026_);
  and g_111188_(_019019_, _019025_, _019027_);
  or g_111189_(_019020_, _019026_, _019028_);
  and g_111190_(_018994_, _019027_, _019030_);
  or g_111191_(_018995_, _019028_, _019031_);
  xor g_111192_(out[278], _018961_, _019032_);
  xor g_111193_(_053082_, _018961_, _019033_);
  and g_111194_(_018752_, _018955_, _019034_);
  or g_111195_(_018753_, _018956_, _019035_);
  and g_111196_(_018760_, _018956_, _019036_);
  or g_111197_(_018759_, _018955_, _019037_);
  and g_111198_(_019035_, _019037_, _019038_);
  or g_111199_(_019034_, _019036_, _019039_);
  and g_111200_(_019032_, _019038_, _019041_);
  or g_111201_(_019033_, _019039_, _019042_);
  xor g_111202_(out[279], _018962_, _019043_);
  xor g_111203_(_053049_, _018962_, _019044_);
  and g_111204_(_018766_, _018955_, _019045_);
  or g_111205_(_018764_, _018956_, _019046_);
  and g_111206_(_018772_, _018956_, _019047_);
  or g_111207_(_018771_, _018955_, _019048_);
  and g_111208_(_019046_, _019048_, _019049_);
  or g_111209_(_019045_, _019047_, _019050_);
  and g_111210_(_019043_, _019050_, _019052_);
  or g_111211_(_019044_, _019049_, _019053_);
  and g_111212_(_019042_, _019053_, _019054_);
  or g_111213_(_019041_, _019052_, _019055_);
  and g_111214_(_019044_, _019049_, _019056_);
  or g_111215_(_019043_, _019050_, _019057_);
  and g_111216_(_019033_, _019039_, _019058_);
  or g_111217_(_019032_, _019038_, _019059_);
  and g_111218_(_019057_, _019059_, _019060_);
  or g_111219_(_019056_, _019058_, _019061_);
  and g_111220_(_019054_, _019060_, _019063_);
  or g_111221_(_019055_, _019061_, _019064_);
  xor g_111222_(out[277], _018960_, _019065_);
  xor g_111223_(_053071_, _018960_, _019066_);
  or g_111224_(_018837_, _018956_, _019067_);
  not g_111225_(_019067_, _019068_);
  and g_111226_(_018840_, _018956_, _019069_);
  not g_111227_(_019069_, _019070_);
  and g_111228_(_019067_, _019070_, _019071_);
  or g_111229_(_019068_, _019069_, _019072_);
  and g_111230_(_019065_, _019072_, _019074_);
  or g_111231_(_019066_, _019071_, _019075_);
  xor g_111232_(out[275], out[276], _019076_);
  xor g_111233_(_053093_, out[276], _019077_);
  or g_111234_(_018823_, _018956_, _019078_);
  not g_111235_(_019078_, _019079_);
  and g_111236_(_018826_, _018956_, _019080_);
  not g_111237_(_019080_, _019081_);
  and g_111238_(_019078_, _019081_, _019082_);
  or g_111239_(_019079_, _019080_, _019083_);
  and g_111240_(_019077_, _019083_, _019085_);
  or g_111241_(_019076_, _019082_, _019086_);
  and g_111242_(_019075_, _019086_, _019087_);
  or g_111243_(_019074_, _019085_, _019088_);
  and g_111244_(_019076_, _019082_, _019089_);
  or g_111245_(_019077_, _019083_, _019090_);
  and g_111246_(_019066_, _019071_, _019091_);
  or g_111247_(_019065_, _019072_, _019092_);
  and g_111248_(_019090_, _019092_, _019093_);
  or g_111249_(_019089_, _019091_, _019094_);
  and g_111250_(_019087_, _019093_, _019096_);
  or g_111251_(_019088_, _019094_, _019097_);
  and g_111252_(_019063_, _019096_, _019098_);
  or g_111253_(_019064_, _019097_, _019099_);
  and g_111254_(_018792_, _018956_, _019100_);
  not g_111255_(_019100_, _019101_);
  or g_111256_(out[258], _018956_, _019102_);
  not g_111257_(_019102_, _019103_);
  and g_111258_(_019101_, _019102_, _019104_);
  or g_111259_(_019100_, _019103_, _019105_);
  and g_111260_(_053115_, _019104_, _019107_);
  or g_111261_(out[274], _019105_, _019108_);
  and g_111262_(out[259], _018955_, _019109_);
  or g_111263_(_053005_, _018956_, _019110_);
  and g_111264_(_018783_, _018956_, _019111_);
  or g_111265_(_018782_, _018955_, _019112_);
  and g_111266_(_019110_, _019112_, _019113_);
  or g_111267_(_019109_, _019111_, _019114_);
  and g_111268_(out[275], _019113_, _019115_);
  or g_111269_(_053093_, _019114_, _019116_);
  or g_111270_(_019107_, _019115_, _019118_);
  and g_111271_(_053093_, _019114_, _019119_);
  or g_111272_(out[275], _019113_, _019120_);
  and g_111273_(out[274], _019105_, _019121_);
  or g_111274_(_019119_, _019121_, _019122_);
  and g_111275_(_019116_, _019120_, _019123_);
  xor g_111276_(_053115_, _019104_, _019124_);
  and g_111277_(_019123_, _019124_, _019125_);
  or g_111278_(_019118_, _019122_, _019126_);
  or g_111279_(out[273], _018959_, _019127_);
  not g_111280_(_019127_, _019129_);
  and g_111281_(_018801_, _018956_, _019130_);
  or g_111282_(_018800_, _018955_, _019131_);
  and g_111283_(_004388_, _018955_, _019132_);
  or g_111284_(out[256], _018956_, _019133_);
  and g_111285_(_019131_, _019133_, _019134_);
  or g_111286_(_019130_, _019132_, _019135_);
  and g_111287_(out[272], _019135_, _019136_);
  or g_111288_(_004443_, _019134_, _019137_);
  xor g_111289_(out[273], _018959_, _019138_);
  xor g_111290_(_053126_, _018959_, _019140_);
  and g_111291_(_019137_, _019138_, _019141_);
  or g_111292_(_019136_, _019140_, _019142_);
  and g_111293_(_019127_, _019142_, _019143_);
  or g_111294_(_019129_, _019141_, _019144_);
  and g_111295_(_019125_, _019144_, _019145_);
  or g_111296_(_019126_, _019143_, _019146_);
  and g_111297_(_019107_, _019120_, _019147_);
  or g_111298_(_019108_, _019119_, _019148_);
  and g_111299_(_019116_, _019148_, _019149_);
  or g_111300_(_019115_, _019147_, _019151_);
  and g_111301_(_019146_, _019149_, _019152_);
  or g_111302_(_019145_, _019151_, _019153_);
  and g_111303_(_019098_, _019153_, _019154_);
  or g_111304_(_019099_, _019152_, _019155_);
  and g_111305_(_019055_, _019057_, _019156_);
  or g_111306_(_019054_, _019056_, _019157_);
  and g_111307_(_019063_, _019088_, _019158_);
  or g_111308_(_019064_, _019087_, _019159_);
  and g_111309_(_019092_, _019158_, _019160_);
  or g_111310_(_019091_, _019159_, _019162_);
  and g_111311_(_019157_, _019162_, _019163_);
  or g_111312_(_019156_, _019160_, _019164_);
  and g_111313_(_019155_, _019163_, _019165_);
  or g_111314_(_019154_, _019164_, _019166_);
  and g_111315_(_019030_, _019166_, _019167_);
  or g_111316_(_019031_, _019165_, _019168_);
  and g_111317_(_018987_, _018989_, _019169_);
  or g_111318_(_018986_, _018988_, _019170_);
  and g_111319_(_019020_, _019022_, _019171_);
  or g_111320_(_019019_, _019021_, _019173_);
  and g_111321_(_018994_, _019171_, _019174_);
  or g_111322_(_018995_, _019173_, _019175_);
  and g_111323_(_019170_, _019175_, _019176_);
  or g_111324_(_019169_, _019174_, _019177_);
  and g_111325_(_019168_, _019176_, _019178_);
  or g_111326_(_019167_, _019177_, _019179_);
  and g_111327_(_004443_, _019134_, _019180_);
  or g_111328_(out[272], _019135_, _019181_);
  and g_111329_(_019125_, _019141_, _019182_);
  or g_111330_(_019126_, _019142_, _019184_);
  and g_111331_(_019181_, _019182_, _019185_);
  or g_111332_(_019180_, _019184_, _019186_);
  or g_111333_(_019031_, _019099_, _019187_);
  and g_111334_(_019098_, _019185_, _019188_);
  and g_111335_(_019030_, _019188_, _019189_);
  or g_111336_(_019186_, _019187_, _019190_);
  and g_111337_(_019179_, _019190_, _019191_);
  or g_111338_(_019178_, _019189_, _019192_);
  and g_111339_(_018959_, _019192_, _019193_);
  and g_111340_(_053126_, _019191_, _019195_);
  or g_111341_(_019193_, _019195_, _019196_);
  and g_111342_(_018979_, _018981_, _019197_);
  or g_111343_(_018980_, _018982_, _019198_);
  and g_111344_(out[291], out[292], _019199_);
  or g_111345_(out[293], _019199_, _019200_);
  or g_111346_(out[294], _019200_, _019201_);
  or g_111347_(out[295], _019201_, _019202_);
  or g_111348_(out[296], _019202_, _019203_);
  and g_111349_(out[297], _019203_, _019204_);
  or g_111350_(out[298], _019204_, _019206_);
  xor g_111351_(out[299], _019206_, _019207_);
  xor g_111352_(_004465_, _019206_, _019208_);
  or g_111353_(_019198_, _019207_, _019209_);
  xor g_111354_(out[298], _019204_, _019210_);
  not g_111355_(_019210_, _019211_);
  and g_111356_(_018976_, _019192_, _019212_);
  not g_111357_(_019212_, _019213_);
  or g_111358_(_018969_, _019192_, _019214_);
  not g_111359_(_019214_, _019215_);
  and g_111360_(_019213_, _019214_, _019217_);
  or g_111361_(_019212_, _019215_, _019218_);
  or g_111362_(_019211_, _019218_, _019219_);
  and g_111363_(_019209_, _019219_, _019220_);
  not g_111364_(_019220_, _019221_);
  and g_111365_(_019211_, _019218_, _019222_);
  and g_111366_(_019198_, _019207_, _019223_);
  and g_111367_(_019013_, _019192_, _019224_);
  not g_111368_(_019224_, _019225_);
  or g_111369_(_019015_, _019192_, _019226_);
  not g_111370_(_019226_, _019228_);
  and g_111371_(_019225_, _019226_, _019229_);
  or g_111372_(_019224_, _019228_, _019230_);
  xor g_111373_(out[297], _019203_, _019231_);
  and g_111374_(_019229_, _019231_, _019232_);
  or g_111375_(_019223_, _019232_, _019233_);
  or g_111376_(_019222_, _019233_, _019234_);
  or g_111377_(_019221_, _019234_, _019235_);
  not g_111378_(_019235_, _019236_);
  and g_111379_(_019002_, _019192_, _019237_);
  not g_111380_(_019237_, _019239_);
  or g_111381_(_019003_, _019192_, _019240_);
  not g_111382_(_019240_, _019241_);
  and g_111383_(_019239_, _019240_, _019242_);
  or g_111384_(_019237_, _019241_, _019243_);
  xor g_111385_(out[296], _019202_, _019244_);
  not g_111386_(_019244_, _019245_);
  or g_111387_(_019242_, _019245_, _019246_);
  or g_111388_(_019229_, _019231_, _019247_);
  and g_111389_(_019246_, _019247_, _019248_);
  or g_111390_(_019243_, _019244_, _019250_);
  and g_111391_(_019248_, _019250_, _019251_);
  not g_111392_(_019251_, _019252_);
  and g_111393_(_019236_, _019251_, _019253_);
  or g_111394_(_019235_, _019252_, _019254_);
  xor g_111395_(out[294], _019200_, _019255_);
  not g_111396_(_019255_, _019256_);
  and g_111397_(_019039_, _019192_, _019257_);
  and g_111398_(_019032_, _019191_, _019258_);
  or g_111399_(_019257_, _019258_, _019259_);
  or g_111400_(_019256_, _019259_, _019261_);
  xor g_111401_(out[295], _019201_, _019262_);
  not g_111402_(_019262_, _019263_);
  or g_111403_(_019049_, _019191_, _019264_);
  or g_111404_(_019043_, _019192_, _019265_);
  and g_111405_(_019264_, _019265_, _019266_);
  not g_111406_(_019266_, _019267_);
  or g_111407_(_019263_, _019266_, _019268_);
  and g_111408_(_019261_, _019268_, _019269_);
  and g_111409_(_019263_, _019266_, _019270_);
  xor g_111410_(out[293], _019199_, _019272_);
  xor g_111411_(_053170_, _019199_, _019273_);
  and g_111412_(_019072_, _019192_, _019274_);
  not g_111413_(_019274_, _019275_);
  or g_111414_(_019065_, _019192_, _019276_);
  not g_111415_(_019276_, _019277_);
  and g_111416_(_019275_, _019276_, _019278_);
  or g_111417_(_019274_, _019277_, _019279_);
  and g_111418_(_019273_, _019278_, _019280_);
  xor g_111419_(_019255_, _019259_, _019281_);
  xor g_111420_(_019262_, _019266_, _019283_);
  or g_111421_(_019281_, _019283_, _019284_);
  or g_111422_(_019280_, _019284_, _019285_);
  not g_111423_(_019285_, _019286_);
  and g_111424_(_019272_, _019279_, _019287_);
  or g_111425_(_019273_, _019278_, _019288_);
  xor g_111426_(out[291], out[292], _019289_);
  not g_111427_(_019289_, _019290_);
  or g_111428_(_019077_, _019192_, _019291_);
  not g_111429_(_019291_, _019292_);
  and g_111430_(_019083_, _019192_, _019294_);
  not g_111431_(_019294_, _019295_);
  and g_111432_(_019291_, _019295_, _019296_);
  or g_111433_(_019292_, _019294_, _019297_);
  and g_111434_(_019290_, _019297_, _019298_);
  or g_111435_(_019289_, _019296_, _019299_);
  and g_111436_(_019288_, _019299_, _019300_);
  or g_111437_(_019287_, _019298_, _019301_);
  and g_111438_(_019289_, _019296_, _019302_);
  or g_111439_(_019290_, _019297_, _019303_);
  and g_111440_(_019300_, _019303_, _019305_);
  or g_111441_(_019301_, _019302_, _019306_);
  and g_111442_(_019286_, _019305_, _019307_);
  or g_111443_(_019285_, _019306_, _019308_);
  and g_111444_(out[275], _019191_, _019309_);
  or g_111445_(_053093_, _019192_, _019310_);
  and g_111446_(_019114_, _019192_, _019311_);
  or g_111447_(_019113_, _019191_, _019312_);
  and g_111448_(_019310_, _019312_, _019313_);
  or g_111449_(_019309_, _019311_, _019314_);
  or g_111450_(_053192_, _019314_, _019316_);
  and g_111451_(_019105_, _019192_, _019317_);
  and g_111452_(_053115_, _019191_, _019318_);
  or g_111453_(_019317_, _019318_, _019319_);
  and g_111454_(_053192_, _019314_, _019320_);
  or g_111455_(out[290], _019319_, _019321_);
  xor g_111456_(out[291], _019313_, _019322_);
  xor g_111457_(_053192_, _019313_, _019323_);
  xor g_111458_(out[290], _019319_, _019324_);
  xor g_111459_(_053214_, _019319_, _019325_);
  and g_111460_(_019322_, _019324_, _019327_);
  or g_111461_(_019323_, _019325_, _019328_);
  or g_111462_(out[289], _019196_, _019329_);
  and g_111463_(_019135_, _019192_, _019330_);
  and g_111464_(_004443_, _019191_, _019331_);
  or g_111465_(_019330_, _019331_, _019332_);
  and g_111466_(out[288], _019332_, _019333_);
  not g_111467_(_019333_, _019334_);
  xor g_111468_(out[289], _019196_, _019335_);
  xor g_111469_(_053225_, _019196_, _019336_);
  and g_111470_(_019334_, _019335_, _019338_);
  or g_111471_(_019333_, _019336_, _019339_);
  and g_111472_(_019329_, _019339_, _019340_);
  or g_111473_(_019328_, _019340_, _019341_);
  or g_111474_(_019320_, _019321_, _019342_);
  and g_111475_(_019316_, _019342_, _019343_);
  and g_111476_(_019341_, _019343_, _019344_);
  or g_111477_(_019308_, _019344_, _019345_);
  or g_111478_(_019285_, _019300_, _019346_);
  or g_111479_(_019269_, _019270_, _019347_);
  and g_111480_(_019346_, _019347_, _019349_);
  and g_111481_(_019345_, _019349_, _019350_);
  or g_111482_(_019254_, _019350_, _019351_);
  or g_111483_(_019220_, _019223_, _019352_);
  or g_111484_(_019235_, _019248_, _019353_);
  and g_111485_(_019352_, _019353_, _019354_);
  and g_111486_(_019351_, _019354_, _019355_);
  or g_111487_(out[288], _019332_, _019356_);
  and g_111488_(_019327_, _019356_, _019357_);
  and g_111489_(_019338_, _019357_, _019358_);
  and g_111490_(_019307_, _019358_, _019360_);
  and g_111491_(_019253_, _019360_, _019361_);
  or g_111492_(_019355_, _019361_, _019362_);
  not g_111493_(_019362_, _019363_);
  and g_111494_(_019196_, _019362_, _019364_);
  not g_111495_(_019364_, _019365_);
  or g_111496_(out[289], _019362_, _019366_);
  not g_111497_(_019366_, _019367_);
  and g_111498_(_019365_, _019366_, _019368_);
  or g_111499_(_019364_, _019367_, _019369_);
  and g_111500_(out[308], out[307], _019371_);
  or g_111501_(out[309], _019371_, _019372_);
  or g_111502_(out[310], _019372_, _019373_);
  or g_111503_(out[311], _019373_, _019374_);
  or g_111504_(out[312], _019374_, _019375_);
  and g_111505_(out[313], _019375_, _019376_);
  or g_111506_(out[314], _019376_, _019377_);
  xor g_111507_(out[314], _019376_, _019378_);
  xor g_111508_(_004520_, _019376_, _019379_);
  and g_111509_(_019218_, _019362_, _019380_);
  or g_111510_(_019217_, _019363_, _019382_);
  and g_111511_(_019210_, _019363_, _019383_);
  or g_111512_(_019211_, _019362_, _019384_);
  and g_111513_(_019382_, _019384_, _019385_);
  or g_111514_(_019380_, _019383_, _019386_);
  and g_111515_(_019378_, _019385_, _019387_);
  or g_111516_(_019379_, _019386_, _019388_);
  and g_111517_(_019197_, _019207_, _019389_);
  or g_111518_(_019198_, _019208_, _019390_);
  xor g_111519_(out[315], _019377_, _019391_);
  xor g_111520_(_004498_, _019377_, _019393_);
  and g_111521_(_019389_, _019393_, _019394_);
  or g_111522_(_019390_, _019391_, _019395_);
  and g_111523_(_019388_, _019395_, _019396_);
  or g_111524_(_019387_, _019394_, _019397_);
  and g_111525_(_019390_, _019391_, _019398_);
  or g_111526_(_019389_, _019393_, _019399_);
  and g_111527_(_019379_, _019386_, _019400_);
  or g_111528_(_019378_, _019385_, _019401_);
  and g_111529_(_019399_, _019401_, _019402_);
  or g_111530_(_019398_, _019400_, _019404_);
  and g_111531_(_019229_, _019362_, _019405_);
  or g_111532_(_019230_, _019363_, _019406_);
  or g_111533_(_019231_, _019362_, _019407_);
  not g_111534_(_019407_, _019408_);
  or g_111535_(_019405_, _019408_, _019409_);
  and g_111536_(_019406_, _019407_, _019410_);
  xor g_111537_(out[313], _019375_, _019411_);
  xor g_111538_(_053335_, _019375_, _019412_);
  and g_111539_(_019409_, _019411_, _019413_);
  or g_111540_(_019410_, _019412_, _019415_);
  and g_111541_(_019243_, _019362_, _019416_);
  or g_111542_(_019242_, _019363_, _019417_);
  or g_111543_(_019244_, _019362_, _019418_);
  not g_111544_(_019418_, _019419_);
  and g_111545_(_019417_, _019418_, _019420_);
  or g_111546_(_019416_, _019419_, _019421_);
  xor g_111547_(out[312], _019374_, _019422_);
  xor g_111548_(_053258_, _019374_, _019423_);
  and g_111549_(_019421_, _019422_, _019424_);
  or g_111550_(_019420_, _019423_, _019426_);
  and g_111551_(_019410_, _019412_, _019427_);
  or g_111552_(_019409_, _019411_, _019428_);
  and g_111553_(_019426_, _019428_, _019429_);
  or g_111554_(_019424_, _019427_, _019430_);
  and g_111555_(_019420_, _019423_, _019431_);
  or g_111556_(_019421_, _019422_, _019432_);
  and g_111557_(_019396_, _019402_, _019433_);
  or g_111558_(_019397_, _019404_, _019434_);
  and g_111559_(_019415_, _019432_, _019435_);
  or g_111560_(_019413_, _019431_, _019437_);
  and g_111561_(_019429_, _019435_, _019438_);
  or g_111562_(_019430_, _019437_, _019439_);
  and g_111563_(_019433_, _019438_, _019440_);
  or g_111564_(_019434_, _019439_, _019441_);
  xor g_111565_(out[311], _019373_, _019442_);
  xor g_111566_(_053247_, _019373_, _019443_);
  and g_111567_(_019267_, _019362_, _019444_);
  or g_111568_(_019266_, _019363_, _019445_);
  or g_111569_(_019262_, _019362_, _019446_);
  not g_111570_(_019446_, _019448_);
  and g_111571_(_019445_, _019446_, _019449_);
  or g_111572_(_019444_, _019448_, _019450_);
  and g_111573_(_019442_, _019450_, _019451_);
  or g_111574_(_019443_, _019449_, _019452_);
  xor g_111575_(out[310], _019372_, _019453_);
  xor g_111576_(_053280_, _019372_, _019454_);
  and g_111577_(_019259_, _019362_, _019455_);
  not g_111578_(_019455_, _019456_);
  and g_111579_(_019255_, _019363_, _019457_);
  or g_111580_(_019256_, _019362_, _019459_);
  and g_111581_(_019456_, _019459_, _019460_);
  or g_111582_(_019455_, _019457_, _019461_);
  and g_111583_(_019453_, _019460_, _019462_);
  or g_111584_(_019454_, _019461_, _019463_);
  and g_111585_(_019452_, _019463_, _019464_);
  or g_111586_(_019451_, _019462_, _019465_);
  xor g_111587_(out[309], _019371_, _019466_);
  xor g_111588_(_053269_, _019371_, _019467_);
  and g_111589_(_019279_, _019362_, _019468_);
  or g_111590_(_019278_, _019363_, _019470_);
  or g_111591_(_019272_, _019362_, _019471_);
  not g_111592_(_019471_, _019472_);
  and g_111593_(_019470_, _019471_, _019473_);
  or g_111594_(_019468_, _019472_, _019474_);
  and g_111595_(_019467_, _019473_, _019475_);
  or g_111596_(_019466_, _019474_, _019476_);
  and g_111597_(_019443_, _019449_, _019477_);
  or g_111598_(_019442_, _019450_, _019478_);
  and g_111599_(_019454_, _019461_, _019479_);
  or g_111600_(_019453_, _019460_, _019481_);
  and g_111601_(_019478_, _019481_, _019482_);
  or g_111602_(_019477_, _019479_, _019483_);
  and g_111603_(_019476_, _019482_, _019484_);
  or g_111604_(_019475_, _019483_, _019485_);
  and g_111605_(_019464_, _019484_, _019486_);
  or g_111606_(_019465_, _019485_, _019487_);
  and g_111607_(_019466_, _019474_, _019488_);
  or g_111608_(_019467_, _019473_, _019489_);
  xor g_111609_(out[308], out[307], _019490_);
  xor g_111610_(_053291_, out[307], _019492_);
  and g_111611_(_019289_, _019363_, _019493_);
  or g_111612_(_019290_, _019362_, _019494_);
  and g_111613_(_019297_, _019362_, _019495_);
  or g_111614_(_019296_, _019363_, _019496_);
  and g_111615_(_019494_, _019496_, _019497_);
  or g_111616_(_019493_, _019495_, _019498_);
  and g_111617_(_019492_, _019498_, _019499_);
  or g_111618_(_019490_, _019497_, _019500_);
  and g_111619_(_019489_, _019500_, _019501_);
  or g_111620_(_019488_, _019499_, _019503_);
  and g_111621_(_019490_, _019497_, _019504_);
  or g_111622_(_019492_, _019498_, _019505_);
  and g_111623_(_019501_, _019505_, _019506_);
  or g_111624_(_019503_, _019504_, _019507_);
  and g_111625_(_019486_, _019506_, _019508_);
  or g_111626_(_019487_, _019507_, _019509_);
  and g_111627_(out[291], _019363_, _019510_);
  or g_111628_(_053192_, _019362_, _019511_);
  and g_111629_(_019314_, _019362_, _019512_);
  or g_111630_(_019313_, _019363_, _019514_);
  and g_111631_(_019511_, _019514_, _019515_);
  or g_111632_(_019510_, _019512_, _019516_);
  and g_111633_(out[307], _019515_, _019517_);
  or g_111634_(_053302_, _019516_, _019518_);
  and g_111635_(_019319_, _019362_, _019519_);
  not g_111636_(_019519_, _019520_);
  or g_111637_(out[290], _019362_, _019521_);
  not g_111638_(_019521_, _019522_);
  and g_111639_(_019520_, _019521_, _019523_);
  or g_111640_(_019519_, _019522_, _019525_);
  and g_111641_(_053313_, _019523_, _019526_);
  or g_111642_(out[306], _019525_, _019527_);
  or g_111643_(_019517_, _019526_, _019528_);
  and g_111644_(_053302_, _019516_, _019529_);
  or g_111645_(out[307], _019515_, _019530_);
  and g_111646_(out[306], _019525_, _019531_);
  or g_111647_(_019529_, _019531_, _019532_);
  and g_111648_(_019518_, _019530_, _019533_);
  xor g_111649_(_053313_, _019523_, _019534_);
  and g_111650_(_019533_, _019534_, _019536_);
  or g_111651_(_019528_, _019532_, _019537_);
  and g_111652_(_019332_, _019362_, _019538_);
  not g_111653_(_019538_, _019539_);
  or g_111654_(out[288], _019362_, _019540_);
  not g_111655_(_019540_, _019541_);
  and g_111656_(_019539_, _019540_, _019542_);
  or g_111657_(_019538_, _019541_, _019543_);
  and g_111658_(out[304], _019543_, _019544_);
  or g_111659_(_004509_, _019542_, _019545_);
  and g_111660_(_053324_, _019368_, _019547_);
  or g_111661_(out[305], _019369_, _019548_);
  xor g_111662_(_053324_, _019368_, _019549_);
  xor g_111663_(out[305], _019368_, _019550_);
  and g_111664_(_019545_, _019549_, _019551_);
  or g_111665_(_019544_, _019550_, _019552_);
  and g_111666_(_004509_, _019542_, _019553_);
  or g_111667_(out[304], _019543_, _019554_);
  and g_111668_(_019551_, _019554_, _019555_);
  or g_111669_(_019552_, _019553_, _019556_);
  and g_111670_(_019536_, _019555_, _019558_);
  or g_111671_(_019537_, _019556_, _019559_);
  or g_111672_(_019509_, _019559_, _019560_);
  and g_111673_(_019440_, _019558_, _019561_);
  and g_111674_(_019508_, _019561_, _019562_);
  or g_111675_(_019441_, _019560_, _019563_);
  and g_111676_(_019548_, _019552_, _019564_);
  or g_111677_(_019547_, _019551_, _019565_);
  and g_111678_(_019536_, _019565_, _019566_);
  or g_111679_(_019537_, _019564_, _019567_);
  and g_111680_(_019526_, _019530_, _019569_);
  or g_111681_(_019527_, _019529_, _019570_);
  and g_111682_(_019518_, _019570_, _019571_);
  or g_111683_(_019517_, _019569_, _019572_);
  and g_111684_(_019567_, _019571_, _019573_);
  or g_111685_(_019566_, _019572_, _019574_);
  and g_111686_(_019508_, _019574_, _019575_);
  or g_111687_(_019509_, _019573_, _019576_);
  and g_111688_(_019486_, _019503_, _019577_);
  or g_111689_(_019487_, _019501_, _019578_);
  and g_111690_(_019465_, _019478_, _019580_);
  or g_111691_(_019464_, _019477_, _019581_);
  and g_111692_(_019578_, _019581_, _019582_);
  or g_111693_(_019577_, _019580_, _019583_);
  and g_111694_(_019576_, _019582_, _019584_);
  or g_111695_(_019575_, _019583_, _019585_);
  and g_111696_(_019440_, _019585_, _019586_);
  or g_111697_(_019441_, _019584_, _019587_);
  and g_111698_(_019397_, _019399_, _019588_);
  or g_111699_(_019396_, _019398_, _019589_);
  and g_111700_(_019415_, _019430_, _019591_);
  or g_111701_(_019413_, _019429_, _019592_);
  and g_111702_(_019433_, _019591_, _019593_);
  or g_111703_(_019434_, _019592_, _019594_);
  and g_111704_(_019589_, _019594_, _019595_);
  or g_111705_(_019588_, _019593_, _019596_);
  and g_111706_(_019587_, _019595_, _019597_);
  or g_111707_(_019586_, _019596_, _019598_);
  and g_111708_(_019563_, _019598_, _019599_);
  or g_111709_(_019562_, _019597_, _019600_);
  or g_111710_(_019368_, _019599_, _019602_);
  or g_111711_(out[305], _019600_, _019603_);
  and g_111712_(_019602_, _019603_, _019604_);
  and g_111713_(out[323], out[324], _019605_);
  or g_111714_(out[325], _019605_, _019606_);
  or g_111715_(out[326], _019606_, _019607_);
  or g_111716_(out[327], _019607_, _019608_);
  or g_111717_(out[328], _019608_, _019609_);
  and g_111718_(out[329], _019609_, _019610_);
  or g_111719_(out[330], _019610_, _019611_);
  xor g_111720_(out[330], _019610_, _019613_);
  not g_111721_(_019613_, _019614_);
  and g_111722_(_019386_, _019600_, _019615_);
  not g_111723_(_019615_, _019616_);
  and g_111724_(_019378_, _019599_, _019617_);
  or g_111725_(_019379_, _019600_, _019618_);
  and g_111726_(_019616_, _019618_, _019619_);
  or g_111727_(_019615_, _019617_, _019620_);
  and g_111728_(_019613_, _019619_, _019621_);
  or g_111729_(_019614_, _019620_, _019622_);
  and g_111730_(_019389_, _019391_, _019624_);
  or g_111731_(_019390_, _019393_, _019625_);
  xor g_111732_(out[331], _019611_, _019626_);
  xor g_111733_(_004531_, _019611_, _019627_);
  and g_111734_(_019624_, _019627_, _019628_);
  or g_111735_(_019625_, _019626_, _019629_);
  and g_111736_(_019622_, _019629_, _019630_);
  or g_111737_(_019621_, _019628_, _019631_);
  or g_111738_(_019613_, _019619_, _019632_);
  or g_111739_(_019624_, _019627_, _019633_);
  and g_111740_(_019410_, _019600_, _019635_);
  not g_111741_(_019635_, _019636_);
  or g_111742_(_019412_, _019600_, _019637_);
  not g_111743_(_019637_, _019638_);
  and g_111744_(_019636_, _019637_, _019639_);
  or g_111745_(_019635_, _019638_, _019640_);
  xor g_111746_(out[329], _019609_, _019641_);
  not g_111747_(_019641_, _019642_);
  or g_111748_(_019640_, _019642_, _019643_);
  xor g_111749_(out[328], _019608_, _019644_);
  not g_111750_(_019644_, _019646_);
  and g_111751_(_019421_, _019600_, _019647_);
  not g_111752_(_019647_, _019648_);
  or g_111753_(_019422_, _019600_, _019649_);
  not g_111754_(_019649_, _019650_);
  and g_111755_(_019648_, _019649_, _019651_);
  or g_111756_(_019647_, _019650_, _019652_);
  and g_111757_(_019644_, _019652_, _019653_);
  or g_111758_(_019646_, _019651_, _019654_);
  and g_111759_(_019640_, _019642_, _019655_);
  or g_111760_(_019639_, _019641_, _019657_);
  and g_111761_(_019654_, _019657_, _019658_);
  or g_111762_(_019653_, _019655_, _019659_);
  or g_111763_(_019644_, _019652_, _019660_);
  and g_111764_(_019630_, _019632_, _019661_);
  and g_111765_(_019633_, _019661_, _019662_);
  and g_111766_(_019643_, _019660_, _019663_);
  and g_111767_(_019658_, _019663_, _019664_);
  and g_111768_(_019662_, _019664_, _019665_);
  not g_111769_(_019665_, _019666_);
  xor g_111770_(out[327], _019607_, _019668_);
  and g_111771_(_019450_, _019600_, _019669_);
  not g_111772_(_019669_, _019670_);
  or g_111773_(_019442_, _019600_, _019671_);
  not g_111774_(_019671_, _019672_);
  and g_111775_(_019670_, _019671_, _019673_);
  or g_111776_(_019669_, _019672_, _019674_);
  and g_111777_(_019668_, _019674_, _019675_);
  xor g_111778_(out[326], _019606_, _019676_);
  and g_111779_(_019461_, _019600_, _019677_);
  not g_111780_(_019677_, _019679_);
  or g_111781_(_019454_, _019600_, _019680_);
  not g_111782_(_019680_, _019681_);
  and g_111783_(_019679_, _019680_, _019682_);
  or g_111784_(_019677_, _019681_, _019683_);
  and g_111785_(_019676_, _019682_, _019684_);
  or g_111786_(_019675_, _019684_, _019685_);
  not g_111787_(_019685_, _019686_);
  or g_111788_(_019668_, _019674_, _019687_);
  or g_111789_(_019676_, _019682_, _019688_);
  and g_111790_(_019687_, _019688_, _019690_);
  and g_111791_(_019686_, _019690_, _019691_);
  not g_111792_(_019691_, _019692_);
  xor g_111793_(out[323], out[324], _019693_);
  not g_111794_(_019693_, _019694_);
  or g_111795_(_019492_, _019600_, _019695_);
  not g_111796_(_019695_, _019696_);
  and g_111797_(_019498_, _019600_, _019697_);
  not g_111798_(_019697_, _019698_);
  and g_111799_(_019695_, _019698_, _019699_);
  or g_111800_(_019696_, _019697_, _019701_);
  and g_111801_(_019694_, _019701_, _019702_);
  xor g_111802_(out[325], _019605_, _019703_);
  and g_111803_(_019474_, _019600_, _019704_);
  not g_111804_(_019704_, _019705_);
  or g_111805_(_019466_, _019600_, _019706_);
  not g_111806_(_019706_, _019707_);
  and g_111807_(_019705_, _019706_, _019708_);
  or g_111808_(_019704_, _019707_, _019709_);
  and g_111809_(_019703_, _019709_, _019710_);
  or g_111810_(_019702_, _019710_, _019712_);
  not g_111811_(_019712_, _019713_);
  or g_111812_(_019703_, _019709_, _019714_);
  not g_111813_(_019714_, _019715_);
  and g_111814_(_019693_, _019699_, _019716_);
  or g_111815_(_019694_, _019701_, _019717_);
  and g_111816_(_019714_, _019717_, _019718_);
  or g_111817_(_019715_, _019716_, _019719_);
  and g_111818_(_019713_, _019718_, _019720_);
  or g_111819_(_019712_, _019719_, _019721_);
  and g_111820_(_019665_, _019720_, _019723_);
  or g_111821_(_019666_, _019721_, _019724_);
  and g_111822_(_019691_, _019723_, _019725_);
  or g_111823_(_019692_, _019724_, _019726_);
  or g_111824_(_053302_, _019600_, _019727_);
  not g_111825_(_019727_, _019728_);
  and g_111826_(_019516_, _019600_, _019729_);
  not g_111827_(_019729_, _019730_);
  and g_111828_(_019727_, _019730_, _019731_);
  or g_111829_(_019728_, _019729_, _019732_);
  and g_111830_(out[323], _019731_, _019734_);
  or g_111831_(_019523_, _019599_, _019735_);
  or g_111832_(out[306], _019600_, _019736_);
  and g_111833_(_019735_, _019736_, _019737_);
  and g_111834_(_053412_, _019737_, _019738_);
  or g_111835_(out[323], _019731_, _019739_);
  xor g_111836_(out[323], _019731_, _019740_);
  xor g_111837_(_053390_, _019731_, _019741_);
  xor g_111838_(_053412_, _019737_, _019742_);
  xor g_111839_(out[322], _019737_, _019743_);
  and g_111840_(_019740_, _019742_, _019745_);
  or g_111841_(_019741_, _019743_, _019746_);
  and g_111842_(_053423_, _019604_, _019747_);
  or g_111843_(_019542_, _019599_, _019748_);
  or g_111844_(out[304], _019600_, _019749_);
  and g_111845_(_019748_, _019749_, _019750_);
  not g_111846_(_019750_, _019751_);
  and g_111847_(out[320], _019751_, _019752_);
  or g_111848_(_004542_, _019750_, _019753_);
  xor g_111849_(_053423_, _019604_, _019754_);
  xor g_111850_(out[321], _019604_, _019756_);
  and g_111851_(_019753_, _019754_, _019757_);
  or g_111852_(_019752_, _019756_, _019758_);
  or g_111853_(_019747_, _019757_, _019759_);
  and g_111854_(_019745_, _019759_, _019760_);
  and g_111855_(_019738_, _019739_, _019761_);
  or g_111856_(_019734_, _019761_, _019762_);
  or g_111857_(_019760_, _019762_, _019763_);
  and g_111858_(_019725_, _019763_, _019764_);
  and g_111859_(_019712_, _019714_, _019765_);
  and g_111860_(_019691_, _019765_, _019767_);
  and g_111861_(_019685_, _019687_, _019768_);
  or g_111862_(_019767_, _019768_, _019769_);
  and g_111863_(_019665_, _019769_, _019770_);
  and g_111864_(_019643_, _019659_, _019771_);
  and g_111865_(_019662_, _019771_, _019772_);
  and g_111866_(_019631_, _019633_, _019773_);
  or g_111867_(_019772_, _019773_, _019774_);
  or g_111868_(_019764_, _019774_, _019775_);
  or g_111869_(_019770_, _019775_, _019776_);
  and g_111870_(_004542_, _019750_, _019778_);
  or g_111871_(_019746_, _019778_, _019779_);
  or g_111872_(_019758_, _019779_, _019780_);
  or g_111873_(_019726_, _019780_, _019781_);
  and g_111874_(_019776_, _019781_, _019782_);
  not g_111875_(_019782_, _019783_);
  or g_111876_(_019604_, _019782_, _019784_);
  not g_111877_(_019784_, _019785_);
  and g_111878_(_053423_, _019782_, _019786_);
  or g_111879_(_019785_, _019786_, _019787_);
  and g_111880_(_019624_, _019626_, _019789_);
  or g_111881_(_019625_, _019627_, _019790_);
  and g_111882_(out[339], out[340], _019791_);
  or g_111883_(out[341], _019791_, _019792_);
  or g_111884_(out[342], _019792_, _019793_);
  or g_111885_(out[343], _019793_, _019794_);
  or g_111886_(out[344], _019794_, _019795_);
  and g_111887_(out[345], _019795_, _019796_);
  or g_111888_(out[346], _019796_, _019797_);
  xor g_111889_(out[347], _019797_, _019798_);
  xor g_111890_(_004564_, _019797_, _019800_);
  or g_111891_(_019790_, _019798_, _019801_);
  xor g_111892_(out[346], _019796_, _019802_);
  not g_111893_(_019802_, _019803_);
  and g_111894_(_019613_, _019782_, _019804_);
  not g_111895_(_019804_, _019805_);
  or g_111896_(_019619_, _019782_, _019806_);
  not g_111897_(_019806_, _019807_);
  and g_111898_(_019805_, _019806_, _019808_);
  or g_111899_(_019804_, _019807_, _019809_);
  or g_111900_(_019803_, _019809_, _019811_);
  and g_111901_(_019801_, _019811_, _019812_);
  not g_111902_(_019812_, _019813_);
  and g_111903_(_019803_, _019809_, _019814_);
  and g_111904_(_019641_, _019782_, _019815_);
  not g_111905_(_019815_, _019816_);
  and g_111906_(_019640_, _019783_, _019817_);
  or g_111907_(_019639_, _019782_, _019818_);
  and g_111908_(_019816_, _019818_, _019819_);
  or g_111909_(_019815_, _019817_, _019820_);
  xor g_111910_(out[345], _019795_, _019822_);
  and g_111911_(_019819_, _019822_, _019823_);
  not g_111912_(_019823_, _019824_);
  and g_111913_(_019790_, _019798_, _019825_);
  xor g_111914_(out[344], _019794_, _019826_);
  not g_111915_(_019826_, _019827_);
  and g_111916_(_019651_, _019783_, _019828_);
  or g_111917_(_019652_, _019782_, _019829_);
  and g_111918_(_019644_, _019782_, _019830_);
  not g_111919_(_019830_, _019831_);
  or g_111920_(_019828_, _019830_, _019833_);
  and g_111921_(_019829_, _019831_, _019834_);
  or g_111922_(_019827_, _019833_, _019835_);
  or g_111923_(_019819_, _019822_, _019836_);
  and g_111924_(_019835_, _019836_, _019837_);
  not g_111925_(_019837_, _019838_);
  and g_111926_(_019827_, _019833_, _019839_);
  or g_111927_(_019826_, _019834_, _019840_);
  or g_111928_(_019814_, _019825_, _019841_);
  or g_111929_(_019813_, _019841_, _019842_);
  not g_111930_(_019842_, _019844_);
  and g_111931_(_019824_, _019840_, _019845_);
  or g_111932_(_019823_, _019839_, _019846_);
  and g_111933_(_019837_, _019845_, _019847_);
  or g_111934_(_019838_, _019846_, _019848_);
  and g_111935_(_019844_, _019847_, _019849_);
  or g_111936_(_019842_, _019848_, _019850_);
  xor g_111937_(out[342], _019792_, _019851_);
  not g_111938_(_019851_, _019852_);
  and g_111939_(_019676_, _019782_, _019853_);
  and g_111940_(_019683_, _019783_, _019855_);
  or g_111941_(_019853_, _019855_, _019856_);
  or g_111942_(_019852_, _019856_, _019857_);
  xor g_111943_(out[343], _019793_, _019858_);
  not g_111944_(_019858_, _019859_);
  or g_111945_(_019668_, _019783_, _019860_);
  or g_111946_(_019673_, _019782_, _019861_);
  and g_111947_(_019860_, _019861_, _019862_);
  or g_111948_(_019859_, _019862_, _019863_);
  and g_111949_(_019857_, _019863_, _019864_);
  and g_111950_(_019859_, _019862_, _019866_);
  xor g_111951_(_019851_, _019856_, _019867_);
  xor g_111952_(_019858_, _019862_, _019868_);
  or g_111953_(_019867_, _019868_, _019869_);
  not g_111954_(_019869_, _019870_);
  xor g_111955_(out[339], out[340], _019871_);
  and g_111956_(_019693_, _019782_, _019872_);
  not g_111957_(_019872_, _019873_);
  and g_111958_(_019701_, _019783_, _019874_);
  or g_111959_(_019699_, _019782_, _019875_);
  and g_111960_(_019873_, _019875_, _019877_);
  or g_111961_(_019872_, _019874_, _019878_);
  or g_111962_(_019871_, _019877_, _019879_);
  xor g_111963_(out[341], _019791_, _019880_);
  xor g_111964_(_053467_, _019791_, _019881_);
  and g_111965_(_019708_, _019783_, _019882_);
  or g_111966_(_019709_, _019782_, _019883_);
  and g_111967_(_019703_, _019782_, _019884_);
  not g_111968_(_019884_, _019885_);
  or g_111969_(_019882_, _019884_, _019886_);
  and g_111970_(_019883_, _019885_, _019888_);
  or g_111971_(_019881_, _019886_, _019889_);
  and g_111972_(_019879_, _019889_, _019890_);
  not g_111973_(_019890_, _019891_);
  and g_111974_(_019881_, _019886_, _019892_);
  and g_111975_(_019871_, _019877_, _019893_);
  or g_111976_(_019892_, _019893_, _019894_);
  not g_111977_(_019894_, _019895_);
  and g_111978_(_019890_, _019895_, _019896_);
  or g_111979_(_019891_, _019894_, _019897_);
  and g_111980_(_019870_, _019896_, _019899_);
  or g_111981_(_019869_, _019897_, _019900_);
  and g_111982_(out[323], _019782_, _019901_);
  not g_111983_(_019901_, _019902_);
  and g_111984_(_019732_, _019783_, _019903_);
  or g_111985_(_019731_, _019782_, _019904_);
  and g_111986_(_019902_, _019904_, _019905_);
  or g_111987_(_019901_, _019903_, _019906_);
  or g_111988_(_053489_, _019906_, _019907_);
  or g_111989_(_019737_, _019782_, _019908_);
  not g_111990_(_019908_, _019910_);
  and g_111991_(_053412_, _019782_, _019911_);
  or g_111992_(_019910_, _019911_, _019912_);
  and g_111993_(_053489_, _019906_, _019913_);
  or g_111994_(out[338], _019912_, _019914_);
  xor g_111995_(out[339], _019905_, _019915_);
  xor g_111996_(_053489_, _019905_, _019916_);
  xor g_111997_(out[338], _019912_, _019917_);
  xor g_111998_(_053511_, _019912_, _019918_);
  and g_111999_(_019915_, _019917_, _019919_);
  or g_112000_(_019916_, _019918_, _019921_);
  or g_112001_(out[337], _019787_, _019922_);
  and g_112002_(_019751_, _019783_, _019923_);
  and g_112003_(_004542_, _019782_, _019924_);
  or g_112004_(_019923_, _019924_, _019925_);
  and g_112005_(out[336], _019925_, _019926_);
  not g_112006_(_019926_, _019927_);
  xor g_112007_(out[337], _019787_, _019928_);
  xor g_112008_(_053522_, _019787_, _019929_);
  and g_112009_(_019927_, _019928_, _019930_);
  or g_112010_(_019926_, _019929_, _019932_);
  and g_112011_(_019922_, _019932_, _019933_);
  or g_112012_(_019921_, _019933_, _019934_);
  or g_112013_(_019913_, _019914_, _019935_);
  and g_112014_(_019907_, _019935_, _019936_);
  and g_112015_(_019934_, _019936_, _019937_);
  or g_112016_(_019900_, _019937_, _019938_);
  or g_112017_(_019869_, _019890_, _019939_);
  or g_112018_(_019892_, _019939_, _019940_);
  or g_112019_(_019864_, _019866_, _019941_);
  and g_112020_(_019940_, _019941_, _019943_);
  and g_112021_(_019938_, _019943_, _019944_);
  or g_112022_(_019850_, _019944_, _019945_);
  or g_112023_(_019823_, _019837_, _019946_);
  or g_112024_(_019842_, _019946_, _019947_);
  or g_112025_(_019812_, _019825_, _019948_);
  and g_112026_(_019947_, _019948_, _019949_);
  and g_112027_(_019945_, _019949_, _019950_);
  or g_112028_(out[336], _019925_, _019951_);
  and g_112029_(_019919_, _019951_, _019952_);
  and g_112030_(_019930_, _019952_, _019954_);
  and g_112031_(_019899_, _019954_, _019955_);
  and g_112032_(_019849_, _019955_, _019956_);
  or g_112033_(_019950_, _019956_, _019957_);
  not g_112034_(_019957_, _019958_);
  and g_112035_(_019787_, _019957_, _019959_);
  and g_112036_(_053522_, _019958_, _019960_);
  or g_112037_(_019959_, _019960_, _019961_);
  and g_112038_(out[355], out[356], _019962_);
  or g_112039_(out[357], _019962_, _019963_);
  or g_112040_(out[358], _019963_, _019965_);
  or g_112041_(out[359], _019965_, _019966_);
  or g_112042_(out[360], _019966_, _019967_);
  and g_112043_(out[361], _019967_, _019968_);
  or g_112044_(out[362], _019968_, _019969_);
  xor g_112045_(out[362], _019968_, _019970_);
  not g_112046_(_019970_, _019971_);
  and g_112047_(_019802_, _019958_, _019972_);
  or g_112048_(_019803_, _019957_, _019973_);
  and g_112049_(_019809_, _019957_, _019974_);
  or g_112050_(_019808_, _019958_, _019976_);
  and g_112051_(_019973_, _019976_, _019977_);
  or g_112052_(_019972_, _019974_, _019978_);
  or g_112053_(_019971_, _019978_, _019979_);
  and g_112054_(_019789_, _019798_, _019980_);
  or g_112055_(_019790_, _019800_, _019981_);
  xor g_112056_(out[363], _019969_, _019982_);
  xor g_112057_(_004597_, _019969_, _019983_);
  or g_112058_(_019981_, _019982_, _019984_);
  and g_112059_(_019979_, _019984_, _019985_);
  not g_112060_(_019985_, _019987_);
  and g_112061_(_019971_, _019978_, _019988_);
  and g_112062_(_019819_, _019957_, _019989_);
  or g_112063_(_019820_, _019958_, _019990_);
  or g_112064_(_019822_, _019957_, _019991_);
  not g_112065_(_019991_, _019992_);
  or g_112066_(_019989_, _019992_, _019993_);
  and g_112067_(_019990_, _019991_, _019994_);
  xor g_112068_(out[361], _019967_, _019995_);
  and g_112069_(_019993_, _019995_, _019996_);
  not g_112070_(_019996_, _019998_);
  and g_112071_(_019981_, _019982_, _019999_);
  xor g_112072_(out[360], _019966_, _020000_);
  not g_112073_(_020000_, _020001_);
  or g_112074_(_019826_, _019957_, _020002_);
  not g_112075_(_020002_, _020003_);
  and g_112076_(_019834_, _019957_, _020004_);
  or g_112077_(_019833_, _019958_, _020005_);
  and g_112078_(_020002_, _020005_, _020006_);
  or g_112079_(_020003_, _020004_, _020007_);
  or g_112080_(_020001_, _020006_, _020009_);
  or g_112081_(_019993_, _019995_, _020010_);
  and g_112082_(_020009_, _020010_, _020011_);
  not g_112083_(_020011_, _020012_);
  and g_112084_(_020001_, _020006_, _020013_);
  or g_112085_(_020000_, _020007_, _020014_);
  or g_112086_(_019988_, _019999_, _020015_);
  or g_112087_(_019987_, _020015_, _020016_);
  not g_112088_(_020016_, _020017_);
  and g_112089_(_019998_, _020014_, _020018_);
  or g_112090_(_019996_, _020013_, _020020_);
  and g_112091_(_020011_, _020018_, _020021_);
  or g_112092_(_020012_, _020020_, _020022_);
  and g_112093_(_020017_, _020021_, _020023_);
  or g_112094_(_020016_, _020022_, _020024_);
  xor g_112095_(out[359], _019965_, _020025_);
  not g_112096_(_020025_, _020026_);
  or g_112097_(_019858_, _019957_, _020027_);
  or g_112098_(_019862_, _019958_, _020028_);
  and g_112099_(_020027_, _020028_, _020029_);
  not g_112100_(_020029_, _020031_);
  or g_112101_(_020026_, _020029_, _020032_);
  xor g_112102_(out[358], _019963_, _020033_);
  not g_112103_(_020033_, _020034_);
  and g_112104_(_019851_, _019958_, _020035_);
  and g_112105_(_019856_, _019957_, _020036_);
  or g_112106_(_020035_, _020036_, _020037_);
  or g_112107_(_020034_, _020037_, _020038_);
  and g_112108_(_020032_, _020038_, _020039_);
  and g_112109_(_020026_, _020029_, _020040_);
  xor g_112110_(_020025_, _020029_, _020042_);
  xor g_112111_(_020033_, _020037_, _020043_);
  or g_112112_(_020042_, _020043_, _020044_);
  not g_112113_(_020044_, _020045_);
  xor g_112114_(out[357], _019962_, _020046_);
  xor g_112115_(_053566_, _019962_, _020047_);
  or g_112116_(_019880_, _019957_, _020048_);
  not g_112117_(_020048_, _020049_);
  and g_112118_(_019888_, _019957_, _020050_);
  or g_112119_(_019886_, _019958_, _020051_);
  and g_112120_(_020048_, _020051_, _020053_);
  or g_112121_(_020049_, _020050_, _020054_);
  or g_112122_(_020047_, _020053_, _020055_);
  xor g_112123_(out[355], out[356], _020056_);
  and g_112124_(_019877_, _019957_, _020057_);
  or g_112125_(_019878_, _019958_, _020058_);
  or g_112126_(_019871_, _019957_, _020059_);
  not g_112127_(_020059_, _020060_);
  or g_112128_(_020057_, _020060_, _020061_);
  and g_112129_(_020058_, _020059_, _020062_);
  or g_112130_(_020056_, _020061_, _020064_);
  and g_112131_(_020055_, _020064_, _020065_);
  not g_112132_(_020065_, _020066_);
  and g_112133_(_020047_, _020053_, _020067_);
  and g_112134_(_020056_, _020061_, _020068_);
  or g_112135_(_020067_, _020068_, _020069_);
  not g_112136_(_020069_, _020070_);
  and g_112137_(_020065_, _020070_, _020071_);
  or g_112138_(_020066_, _020069_, _020072_);
  and g_112139_(_020045_, _020071_, _020073_);
  or g_112140_(_020044_, _020072_, _020075_);
  and g_112141_(out[339], _019958_, _020076_);
  or g_112142_(_053489_, _019957_, _020077_);
  and g_112143_(_019906_, _019957_, _020078_);
  or g_112144_(_019905_, _019958_, _020079_);
  and g_112145_(_020077_, _020079_, _020080_);
  or g_112146_(_020076_, _020078_, _020081_);
  or g_112147_(_053588_, _020081_, _020082_);
  and g_112148_(_019912_, _019957_, _020083_);
  and g_112149_(_053511_, _019958_, _020084_);
  or g_112150_(_020083_, _020084_, _020086_);
  or g_112151_(out[354], _020086_, _020087_);
  and g_112152_(_053588_, _020081_, _020088_);
  xor g_112153_(_053588_, _020080_, _020089_);
  xor g_112154_(_053610_, _020086_, _020090_);
  or g_112155_(_020089_, _020090_, _020091_);
  not g_112156_(_020091_, _020092_);
  or g_112157_(out[353], _019961_, _020093_);
  or g_112158_(_020087_, _020088_, _020094_);
  and g_112159_(_020082_, _020094_, _020095_);
  and g_112160_(_019925_, _019957_, _020097_);
  and g_112161_(_004575_, _019958_, _020098_);
  or g_112162_(_020097_, _020098_, _020099_);
  and g_112163_(out[352], _020099_, _020100_);
  not g_112164_(_020100_, _020101_);
  xor g_112165_(out[353], _019961_, _020102_);
  xor g_112166_(_053621_, _019961_, _020103_);
  and g_112167_(_020101_, _020102_, _020104_);
  or g_112168_(_020100_, _020103_, _020105_);
  and g_112169_(_020092_, _020104_, _020106_);
  and g_112170_(_020093_, _020105_, _020108_);
  or g_112171_(_020091_, _020108_, _020109_);
  and g_112172_(_020095_, _020109_, _020110_);
  or g_112173_(_020075_, _020110_, _020111_);
  or g_112174_(_020039_, _020040_, _020112_);
  or g_112175_(_020065_, _020067_, _020113_);
  or g_112176_(_020044_, _020113_, _020114_);
  and g_112177_(_020112_, _020114_, _020115_);
  and g_112178_(_020111_, _020115_, _020116_);
  or g_112179_(_020024_, _020116_, _020117_);
  or g_112180_(_019996_, _020011_, _020119_);
  or g_112181_(_020016_, _020119_, _020120_);
  or g_112182_(_019985_, _019999_, _020121_);
  and g_112183_(_020120_, _020121_, _020122_);
  and g_112184_(_020117_, _020122_, _020123_);
  or g_112185_(out[352], _020099_, _020124_);
  and g_112186_(_020106_, _020124_, _020125_);
  and g_112187_(_020023_, _020125_, _020126_);
  and g_112188_(_020073_, _020126_, _020127_);
  or g_112189_(_020123_, _020127_, _020128_);
  not g_112190_(_020128_, _020130_);
  and g_112191_(_019961_, _020128_, _020131_);
  and g_112192_(_053621_, _020130_, _020132_);
  or g_112193_(_020131_, _020132_, _020133_);
  and g_112194_(out[371], out[372], _020134_);
  or g_112195_(out[373], _020134_, _020135_);
  or g_112196_(out[374], _020135_, _020136_);
  or g_112197_(out[375], _020136_, _020137_);
  or g_112198_(out[376], _020137_, _020138_);
  and g_112199_(out[377], _020138_, _020139_);
  or g_112200_(out[378], _020139_, _020141_);
  xor g_112201_(out[378], _020139_, _020142_);
  not g_112202_(_020142_, _020143_);
  and g_112203_(_019970_, _020130_, _020144_);
  or g_112204_(_019971_, _020128_, _020145_);
  and g_112205_(_019978_, _020128_, _020146_);
  or g_112206_(_019977_, _020130_, _020147_);
  and g_112207_(_020145_, _020147_, _020148_);
  or g_112208_(_020144_, _020146_, _020149_);
  and g_112209_(_020142_, _020148_, _020150_);
  or g_112210_(_020143_, _020149_, _020152_);
  and g_112211_(_019980_, _019982_, _020153_);
  or g_112212_(_019981_, _019983_, _020154_);
  xor g_112213_(out[379], _020141_, _020155_);
  xor g_112214_(_004630_, _020141_, _020156_);
  and g_112215_(_020153_, _020156_, _020157_);
  or g_112216_(_020154_, _020155_, _020158_);
  and g_112217_(_020152_, _020158_, _020159_);
  or g_112218_(_020150_, _020157_, _020160_);
  and g_112219_(_020143_, _020149_, _020161_);
  and g_112220_(_020154_, _020155_, _020163_);
  and g_112221_(_019993_, _020128_, _020164_);
  or g_112222_(_019994_, _020130_, _020165_);
  or g_112223_(_019995_, _020128_, _020166_);
  not g_112224_(_020166_, _020167_);
  or g_112225_(_020164_, _020167_, _020168_);
  and g_112226_(_020165_, _020166_, _020169_);
  xor g_112227_(out[377], _020138_, _020170_);
  and g_112228_(_020168_, _020170_, _020171_);
  or g_112229_(_020161_, _020163_, _020172_);
  or g_112230_(_020160_, _020172_, _020174_);
  or g_112231_(_020171_, _020174_, _020175_);
  or g_112232_(_020168_, _020170_, _020176_);
  xor g_112233_(out[376], _020137_, _020177_);
  not g_112234_(_020177_, _020178_);
  or g_112235_(_020000_, _020128_, _020179_);
  not g_112236_(_020179_, _020180_);
  and g_112237_(_020007_, _020128_, _020181_);
  or g_112238_(_020006_, _020130_, _020182_);
  and g_112239_(_020179_, _020182_, _020183_);
  or g_112240_(_020180_, _020181_, _020185_);
  or g_112241_(_020178_, _020183_, _020186_);
  and g_112242_(_020176_, _020186_, _020187_);
  or g_112243_(_020177_, _020185_, _020188_);
  and g_112244_(_020187_, _020188_, _020189_);
  not g_112245_(_020189_, _020190_);
  or g_112246_(_020175_, _020190_, _020191_);
  xor g_112247_(out[374], _020135_, _020192_);
  not g_112248_(_020192_, _020193_);
  and g_112249_(_020033_, _020130_, _020194_);
  or g_112250_(_020034_, _020128_, _020196_);
  and g_112251_(_020037_, _020128_, _020197_);
  not g_112252_(_020197_, _020198_);
  and g_112253_(_020196_, _020198_, _020199_);
  or g_112254_(_020194_, _020197_, _020200_);
  or g_112255_(_020193_, _020200_, _020201_);
  xor g_112256_(out[375], _020136_, _020202_);
  not g_112257_(_020202_, _020203_);
  or g_112258_(_020025_, _020128_, _020204_);
  not g_112259_(_020204_, _020205_);
  and g_112260_(_020031_, _020128_, _020207_);
  or g_112261_(_020029_, _020130_, _020208_);
  and g_112262_(_020204_, _020208_, _020209_);
  or g_112263_(_020205_, _020207_, _020210_);
  or g_112264_(_020203_, _020209_, _020211_);
  and g_112265_(_020201_, _020211_, _020212_);
  and g_112266_(_020203_, _020209_, _020213_);
  or g_112267_(_020192_, _020199_, _020214_);
  and g_112268_(_020212_, _020214_, _020215_);
  not g_112269_(_020215_, _020216_);
  or g_112270_(_020213_, _020216_, _020218_);
  xor g_112271_(out[373], _020134_, _020219_);
  xor g_112272_(_053665_, _020134_, _020220_);
  or g_112273_(_020046_, _020128_, _020221_);
  not g_112274_(_020221_, _020222_);
  and g_112275_(_020054_, _020128_, _020223_);
  or g_112276_(_020053_, _020130_, _020224_);
  and g_112277_(_020221_, _020224_, _020225_);
  or g_112278_(_020222_, _020223_, _020226_);
  or g_112279_(_020220_, _020225_, _020227_);
  xor g_112280_(out[371], out[372], _020229_);
  and g_112281_(_020061_, _020128_, _020230_);
  or g_112282_(_020062_, _020130_, _020231_);
  or g_112283_(_020056_, _020128_, _020232_);
  not g_112284_(_020232_, _020233_);
  or g_112285_(_020230_, _020233_, _020234_);
  and g_112286_(_020231_, _020232_, _020235_);
  or g_112287_(_020229_, _020234_, _020236_);
  and g_112288_(_020227_, _020236_, _020237_);
  not g_112289_(_020237_, _020238_);
  and g_112290_(_020229_, _020234_, _020240_);
  and g_112291_(out[355], _020130_, _020241_);
  or g_112292_(_053588_, _020128_, _020242_);
  and g_112293_(_020081_, _020128_, _020243_);
  or g_112294_(_020080_, _020130_, _020244_);
  and g_112295_(_020242_, _020244_, _020245_);
  or g_112296_(_020241_, _020243_, _020246_);
  and g_112297_(_053687_, _020246_, _020247_);
  and g_112298_(_020220_, _020225_, _020248_);
  and g_112299_(_020086_, _020128_, _020249_);
  and g_112300_(_053610_, _020130_, _020251_);
  or g_112301_(_020249_, _020251_, _020252_);
  or g_112302_(out[370], _020252_, _020253_);
  or g_112303_(_053687_, _020246_, _020254_);
  xor g_112304_(out[370], _020252_, _020255_);
  xor g_112305_(_053709_, _020252_, _020256_);
  xor g_112306_(out[371], _020245_, _020257_);
  xor g_112307_(_053687_, _020245_, _020258_);
  and g_112308_(_020255_, _020257_, _020259_);
  or g_112309_(_020256_, _020258_, _020260_);
  or g_112310_(_020238_, _020248_, _020262_);
  or g_112311_(_020240_, _020262_, _020263_);
  or g_112312_(_020191_, _020263_, _020264_);
  or g_112313_(_020218_, _020264_, _020265_);
  and g_112314_(_020099_, _020128_, _020266_);
  and g_112315_(_004608_, _020130_, _020267_);
  or g_112316_(_020266_, _020267_, _020268_);
  and g_112317_(out[368], _020268_, _020269_);
  not g_112318_(_020269_, _020270_);
  or g_112319_(out[369], _020133_, _020271_);
  xor g_112320_(out[369], _020133_, _020273_);
  xor g_112321_(_053720_, _020133_, _020274_);
  and g_112322_(_020270_, _020273_, _020275_);
  or g_112323_(_020269_, _020274_, _020276_);
  or g_112324_(out[368], _020268_, _020277_);
  not g_112325_(_020277_, _020278_);
  and g_112326_(_020259_, _020275_, _020279_);
  or g_112327_(_020265_, _020278_, _020280_);
  not g_112328_(_020280_, _020281_);
  and g_112329_(_020279_, _020281_, _020282_);
  and g_112330_(_020271_, _020276_, _020284_);
  or g_112331_(_020212_, _020213_, _020285_);
  or g_112332_(_020237_, _020248_, _020286_);
  or g_112333_(_020218_, _020286_, _020287_);
  and g_112334_(_020285_, _020287_, _020288_);
  or g_112335_(_020191_, _020288_, _020289_);
  or g_112336_(_020175_, _020187_, _020290_);
  or g_112337_(_020159_, _020163_, _020291_);
  or g_112338_(_020247_, _020253_, _020292_);
  and g_112339_(_020254_, _020292_, _020293_);
  or g_112340_(_020260_, _020284_, _020295_);
  and g_112341_(_020293_, _020295_, _020296_);
  or g_112342_(_020265_, _020296_, _020297_);
  and g_112343_(_020290_, _020297_, _020298_);
  and g_112344_(_020289_, _020291_, _020299_);
  and g_112345_(_020298_, _020299_, _020300_);
  or g_112346_(_020282_, _020300_, _020301_);
  not g_112347_(_020301_, _020302_);
  and g_112348_(_020133_, _020301_, _020303_);
  and g_112349_(_053720_, _020302_, _020304_);
  or g_112350_(_020303_, _020304_, _020306_);
  and g_112351_(out[371], _020302_, _020307_);
  or g_112352_(_053687_, _020301_, _020308_);
  and g_112353_(_020246_, _020301_, _020309_);
  or g_112354_(_020245_, _020302_, _020310_);
  and g_112355_(_020308_, _020310_, _020311_);
  or g_112356_(_020307_, _020309_, _020312_);
  and g_112357_(out[387], _020311_, _020313_);
  or g_112358_(_053786_, _020312_, _020314_);
  and g_112359_(_020252_, _020301_, _020315_);
  not g_112360_(_020315_, _020317_);
  or g_112361_(out[370], _020301_, _020318_);
  not g_112362_(_020318_, _020319_);
  and g_112363_(_020317_, _020318_, _020320_);
  or g_112364_(_020315_, _020319_, _020321_);
  and g_112365_(out[386], _020321_, _020322_);
  or g_112366_(_020313_, _020322_, _020323_);
  and g_112367_(_053786_, _020312_, _020324_);
  or g_112368_(out[387], _020311_, _020325_);
  and g_112369_(_053808_, _020320_, _020326_);
  or g_112370_(out[386], _020321_, _020328_);
  or g_112371_(_020324_, _020326_, _020329_);
  or g_112372_(_020323_, _020329_, _020330_);
  or g_112373_(out[385], _020306_, _020331_);
  and g_112374_(_020268_, _020301_, _020332_);
  not g_112375_(_020332_, _020333_);
  or g_112376_(out[368], _020301_, _020334_);
  not g_112377_(_020334_, _020335_);
  and g_112378_(_020333_, _020334_, _020336_);
  or g_112379_(_020332_, _020335_, _020337_);
  and g_112380_(out[384], _020337_, _020339_);
  xor g_112381_(_053819_, _020306_, _020340_);
  or g_112382_(_020339_, _020340_, _020341_);
  and g_112383_(_020331_, _020341_, _020342_);
  or g_112384_(_020330_, _020342_, _020343_);
  not g_112385_(_020343_, _020344_);
  and g_112386_(_020325_, _020326_, _020345_);
  or g_112387_(_020324_, _020328_, _020346_);
  and g_112388_(_020314_, _020346_, _020347_);
  or g_112389_(_020313_, _020345_, _020348_);
  and g_112390_(_020343_, _020347_, _020350_);
  or g_112391_(_020344_, _020348_, _020351_);
  and g_112392_(out[387], out[388], _020352_);
  or g_112393_(out[389], _020352_, _020353_);
  or g_112394_(out[390], _020353_, _020354_);
  or g_112395_(out[391], _020354_, _020355_);
  or g_112396_(out[392], _020355_, _020356_);
  and g_112397_(out[393], _020356_, _020357_);
  or g_112398_(out[394], _020357_, _020358_);
  xor g_112399_(out[394], _020357_, _020359_);
  xor g_112400_(_004685_, _020357_, _020361_);
  and g_112401_(_020142_, _020302_, _020362_);
  or g_112402_(_020143_, _020301_, _020363_);
  and g_112403_(_020149_, _020301_, _020364_);
  or g_112404_(_020148_, _020302_, _020365_);
  and g_112405_(_020363_, _020365_, _020366_);
  or g_112406_(_020362_, _020364_, _020367_);
  and g_112407_(_020359_, _020366_, _020368_);
  or g_112408_(_020361_, _020367_, _020369_);
  and g_112409_(_020153_, _020155_, _020370_);
  or g_112410_(_020154_, _020156_, _020372_);
  xor g_112411_(out[395], _020358_, _020373_);
  xor g_112412_(_004663_, _020358_, _020374_);
  and g_112413_(_020370_, _020374_, _020375_);
  or g_112414_(_020372_, _020373_, _020376_);
  and g_112415_(_020369_, _020376_, _020377_);
  or g_112416_(_020368_, _020375_, _020378_);
  and g_112417_(_020372_, _020373_, _020379_);
  or g_112418_(_020370_, _020374_, _020380_);
  and g_112419_(_020361_, _020367_, _020381_);
  or g_112420_(_020359_, _020366_, _020383_);
  and g_112421_(_020380_, _020383_, _020384_);
  or g_112422_(_020379_, _020381_, _020385_);
  and g_112423_(_020377_, _020384_, _020386_);
  or g_112424_(_020378_, _020385_, _020387_);
  and g_112425_(_020168_, _020301_, _020388_);
  or g_112426_(_020169_, _020302_, _020389_);
  or g_112427_(_020170_, _020301_, _020390_);
  not g_112428_(_020390_, _020391_);
  or g_112429_(_020388_, _020391_, _020392_);
  and g_112430_(_020389_, _020390_, _020394_);
  xor g_112431_(out[393], _020356_, _020395_);
  xor g_112432_(_053830_, _020356_, _020396_);
  and g_112433_(_020394_, _020396_, _020397_);
  or g_112434_(_020392_, _020395_, _020398_);
  xor g_112435_(out[392], _020355_, _020399_);
  xor g_112436_(_053753_, _020355_, _020400_);
  or g_112437_(_020177_, _020301_, _020401_);
  not g_112438_(_020401_, _020402_);
  and g_112439_(_020185_, _020301_, _020403_);
  or g_112440_(_020183_, _020302_, _020405_);
  and g_112441_(_020401_, _020405_, _020406_);
  or g_112442_(_020402_, _020403_, _020407_);
  and g_112443_(_020399_, _020407_, _020408_);
  or g_112444_(_020400_, _020406_, _020409_);
  and g_112445_(_020398_, _020409_, _020410_);
  or g_112446_(_020397_, _020408_, _020411_);
  and g_112447_(_020392_, _020395_, _020412_);
  or g_112448_(_020394_, _020396_, _020413_);
  and g_112449_(_020400_, _020406_, _020414_);
  or g_112450_(_020399_, _020407_, _020416_);
  and g_112451_(_020413_, _020416_, _020417_);
  or g_112452_(_020412_, _020414_, _020418_);
  and g_112453_(_020410_, _020417_, _020419_);
  or g_112454_(_020411_, _020418_, _020420_);
  and g_112455_(_020386_, _020419_, _020421_);
  or g_112456_(_020387_, _020420_, _020422_);
  xor g_112457_(out[391], _020354_, _020423_);
  xor g_112458_(_053742_, _020354_, _020424_);
  or g_112459_(_020202_, _020301_, _020425_);
  not g_112460_(_020425_, _020427_);
  and g_112461_(_020210_, _020301_, _020428_);
  or g_112462_(_020209_, _020302_, _020429_);
  and g_112463_(_020425_, _020429_, _020430_);
  or g_112464_(_020427_, _020428_, _020431_);
  and g_112465_(_020423_, _020431_, _020432_);
  or g_112466_(_020424_, _020430_, _020433_);
  xor g_112467_(out[390], _020353_, _020434_);
  xor g_112468_(_053775_, _020353_, _020435_);
  and g_112469_(_020192_, _020302_, _020436_);
  or g_112470_(_020193_, _020301_, _020438_);
  and g_112471_(_020200_, _020301_, _020439_);
  or g_112472_(_020199_, _020302_, _020440_);
  and g_112473_(_020438_, _020440_, _020441_);
  or g_112474_(_020436_, _020439_, _020442_);
  and g_112475_(_020434_, _020441_, _020443_);
  or g_112476_(_020435_, _020442_, _020444_);
  and g_112477_(_020433_, _020444_, _020445_);
  or g_112478_(_020432_, _020443_, _020446_);
  and g_112479_(_020424_, _020430_, _020447_);
  or g_112480_(_020423_, _020431_, _020449_);
  and g_112481_(_020435_, _020442_, _020450_);
  or g_112482_(_020434_, _020441_, _020451_);
  and g_112483_(_020449_, _020451_, _020452_);
  or g_112484_(_020447_, _020450_, _020453_);
  and g_112485_(_020445_, _020452_, _020454_);
  or g_112486_(_020446_, _020453_, _020455_);
  xor g_112487_(out[387], out[388], _020456_);
  xor g_112488_(_053786_, out[388], _020457_);
  and g_112489_(_020234_, _020301_, _020458_);
  or g_112490_(_020235_, _020302_, _020460_);
  or g_112491_(_020229_, _020301_, _020461_);
  not g_112492_(_020461_, _020462_);
  or g_112493_(_020458_, _020462_, _020463_);
  and g_112494_(_020460_, _020461_, _020464_);
  and g_112495_(_020457_, _020464_, _020465_);
  or g_112496_(_020456_, _020463_, _020466_);
  xor g_112497_(out[389], _020352_, _020467_);
  xor g_112498_(_053764_, _020352_, _020468_);
  or g_112499_(_020219_, _020301_, _020469_);
  not g_112500_(_020469_, _020471_);
  and g_112501_(_020226_, _020301_, _020472_);
  or g_112502_(_020225_, _020302_, _020473_);
  and g_112503_(_020469_, _020473_, _020474_);
  or g_112504_(_020471_, _020472_, _020475_);
  and g_112505_(_020467_, _020475_, _020476_);
  or g_112506_(_020468_, _020474_, _020477_);
  and g_112507_(_020466_, _020477_, _020478_);
  or g_112508_(_020465_, _020476_, _020479_);
  and g_112509_(_020468_, _020474_, _020480_);
  or g_112510_(_020467_, _020475_, _020482_);
  and g_112511_(_020456_, _020463_, _020483_);
  or g_112512_(_020457_, _020464_, _020484_);
  and g_112513_(_020482_, _020484_, _020485_);
  or g_112514_(_020480_, _020483_, _020486_);
  and g_112515_(_020478_, _020485_, _020487_);
  or g_112516_(_020479_, _020486_, _020488_);
  and g_112517_(_020454_, _020487_, _020489_);
  or g_112518_(_020455_, _020488_, _020490_);
  and g_112519_(_020421_, _020489_, _020491_);
  or g_112520_(_020422_, _020490_, _020493_);
  and g_112521_(_020351_, _020491_, _020494_);
  or g_112522_(_020350_, _020493_, _020495_);
  and g_112523_(_020479_, _020482_, _020496_);
  or g_112524_(_020478_, _020480_, _020497_);
  and g_112525_(_020454_, _020496_, _020498_);
  or g_112526_(_020455_, _020497_, _020499_);
  and g_112527_(_020446_, _020449_, _020500_);
  or g_112528_(_020445_, _020447_, _020501_);
  and g_112529_(_020499_, _020501_, _020502_);
  or g_112530_(_020498_, _020500_, _020504_);
  and g_112531_(_020421_, _020504_, _020505_);
  or g_112532_(_020422_, _020502_, _020506_);
  and g_112533_(_020411_, _020413_, _020507_);
  or g_112534_(_020410_, _020412_, _020508_);
  and g_112535_(_020386_, _020507_, _020509_);
  or g_112536_(_020387_, _020508_, _020510_);
  and g_112537_(_020378_, _020380_, _020511_);
  or g_112538_(_020377_, _020379_, _020512_);
  and g_112539_(_020510_, _020512_, _020513_);
  or g_112540_(_020509_, _020511_, _020515_);
  or g_112541_(_020505_, _020515_, _020516_);
  and g_112542_(_020495_, _020513_, _020517_);
  and g_112543_(_020506_, _020517_, _020518_);
  or g_112544_(_020494_, _020516_, _020519_);
  and g_112545_(_004674_, _020336_, _020520_);
  or g_112546_(_020330_, _020520_, _020521_);
  or g_112547_(_020341_, _020521_, _020522_);
  or g_112548_(_020493_, _020522_, _020523_);
  not g_112549_(_020523_, _020524_);
  and g_112550_(_020519_, _020523_, _020526_);
  or g_112551_(_020518_, _020524_, _020527_);
  and g_112552_(_020306_, _020527_, _020528_);
  and g_112553_(_053819_, _020526_, _020529_);
  or g_112554_(_020528_, _020529_, _020530_);
  or g_112555_(_053786_, _020527_, _020531_);
  not g_112556_(_020531_, _020532_);
  and g_112557_(_020312_, _020527_, _020533_);
  not g_112558_(_020533_, _020534_);
  and g_112559_(_020531_, _020534_, _020535_);
  or g_112560_(_020532_, _020533_, _020537_);
  and g_112561_(out[403], _020535_, _020538_);
  or g_112562_(_053885_, _020537_, _020539_);
  and g_112563_(_020321_, _020527_, _020540_);
  not g_112564_(_020540_, _020541_);
  or g_112565_(out[386], _020527_, _020542_);
  not g_112566_(_020542_, _020543_);
  and g_112567_(_020541_, _020542_, _020544_);
  or g_112568_(_020540_, _020543_, _020545_);
  and g_112569_(out[402], _020545_, _020546_);
  or g_112570_(_020538_, _020546_, _020548_);
  and g_112571_(_053885_, _020537_, _020549_);
  or g_112572_(out[403], _020535_, _020550_);
  and g_112573_(_053907_, _020544_, _020551_);
  or g_112574_(out[402], _020545_, _020552_);
  or g_112575_(_020549_, _020551_, _020553_);
  or g_112576_(_020548_, _020553_, _020554_);
  or g_112577_(out[401], _020530_, _020555_);
  and g_112578_(_020337_, _020527_, _020556_);
  not g_112579_(_020556_, _020557_);
  or g_112580_(out[384], _020527_, _020559_);
  not g_112581_(_020559_, _020560_);
  and g_112582_(_020557_, _020559_, _020561_);
  or g_112583_(_020556_, _020560_, _020562_);
  and g_112584_(out[400], _020562_, _020563_);
  xor g_112585_(_053918_, _020530_, _020564_);
  or g_112586_(_020563_, _020564_, _020565_);
  and g_112587_(_020555_, _020565_, _020566_);
  or g_112588_(_020554_, _020566_, _020567_);
  not g_112589_(_020567_, _020568_);
  and g_112590_(_020539_, _020552_, _020570_);
  or g_112591_(_020538_, _020551_, _020571_);
  and g_112592_(_020550_, _020571_, _020572_);
  or g_112593_(_020549_, _020570_, _020573_);
  and g_112594_(_020567_, _020573_, _020574_);
  or g_112595_(_020568_, _020572_, _020575_);
  and g_112596_(out[403], out[404], _020576_);
  or g_112597_(out[405], _020576_, _020577_);
  or g_112598_(out[406], _020577_, _020578_);
  or g_112599_(out[407], _020578_, _020579_);
  or g_112600_(out[408], _020579_, _020581_);
  and g_112601_(out[409], _020581_, _020582_);
  or g_112602_(out[410], _020582_, _020583_);
  xor g_112603_(out[410], _020582_, _020584_);
  xor g_112604_(_004718_, _020582_, _020585_);
  and g_112605_(_020359_, _020526_, _020586_);
  or g_112606_(_020361_, _020527_, _020587_);
  and g_112607_(_020367_, _020527_, _020588_);
  or g_112608_(_020366_, _020526_, _020589_);
  and g_112609_(_020587_, _020589_, _020590_);
  or g_112610_(_020586_, _020588_, _020592_);
  and g_112611_(_020584_, _020590_, _020593_);
  or g_112612_(_020585_, _020592_, _020594_);
  and g_112613_(_020370_, _020373_, _020595_);
  or g_112614_(_020372_, _020374_, _020596_);
  xor g_112615_(out[411], _020583_, _020597_);
  xor g_112616_(_004696_, _020583_, _020598_);
  and g_112617_(_020595_, _020598_, _020599_);
  or g_112618_(_020596_, _020597_, _020600_);
  and g_112619_(_020594_, _020600_, _020601_);
  or g_112620_(_020593_, _020599_, _020603_);
  and g_112621_(_020585_, _020592_, _020604_);
  or g_112622_(_020584_, _020590_, _020605_);
  and g_112623_(_020596_, _020597_, _020606_);
  or g_112624_(_020595_, _020598_, _020607_);
  or g_112625_(_020396_, _020527_, _020608_);
  not g_112626_(_020608_, _020609_);
  and g_112627_(_020394_, _020527_, _020610_);
  not g_112628_(_020610_, _020611_);
  and g_112629_(_020608_, _020611_, _020612_);
  or g_112630_(_020609_, _020610_, _020614_);
  xor g_112631_(out[409], _020581_, _020615_);
  xor g_112632_(_053929_, _020581_, _020616_);
  and g_112633_(_020612_, _020615_, _020617_);
  or g_112634_(_020614_, _020616_, _020618_);
  xor g_112635_(out[408], _020579_, _020619_);
  xor g_112636_(_053852_, _020579_, _020620_);
  or g_112637_(_020399_, _020527_, _020621_);
  not g_112638_(_020621_, _020622_);
  and g_112639_(_020407_, _020527_, _020623_);
  not g_112640_(_020623_, _020625_);
  and g_112641_(_020621_, _020625_, _020626_);
  or g_112642_(_020622_, _020623_, _020627_);
  and g_112643_(_020619_, _020627_, _020628_);
  or g_112644_(_020620_, _020626_, _020629_);
  and g_112645_(_020614_, _020616_, _020630_);
  or g_112646_(_020612_, _020615_, _020631_);
  and g_112647_(_020629_, _020631_, _020632_);
  or g_112648_(_020628_, _020630_, _020633_);
  and g_112649_(_020620_, _020626_, _020634_);
  or g_112650_(_020619_, _020627_, _020636_);
  and g_112651_(_020605_, _020607_, _020637_);
  or g_112652_(_020604_, _020606_, _020638_);
  and g_112653_(_020601_, _020637_, _020639_);
  or g_112654_(_020603_, _020638_, _020640_);
  and g_112655_(_020618_, _020636_, _020641_);
  or g_112656_(_020617_, _020634_, _020642_);
  and g_112657_(_020632_, _020641_, _020643_);
  or g_112658_(_020633_, _020642_, _020644_);
  and g_112659_(_020639_, _020643_, _020645_);
  or g_112660_(_020640_, _020644_, _020647_);
  xor g_112661_(out[407], _020578_, _020648_);
  xor g_112662_(_053841_, _020578_, _020649_);
  or g_112663_(_020423_, _020527_, _020650_);
  not g_112664_(_020650_, _020651_);
  and g_112665_(_020431_, _020527_, _020652_);
  not g_112666_(_020652_, _020653_);
  and g_112667_(_020650_, _020653_, _020654_);
  or g_112668_(_020651_, _020652_, _020655_);
  and g_112669_(_020648_, _020655_, _020656_);
  or g_112670_(_020649_, _020654_, _020658_);
  xor g_112671_(out[406], _020577_, _020659_);
  xor g_112672_(_053874_, _020577_, _020660_);
  or g_112673_(_020435_, _020527_, _020661_);
  not g_112674_(_020661_, _020662_);
  and g_112675_(_020442_, _020527_, _020663_);
  not g_112676_(_020663_, _020664_);
  and g_112677_(_020661_, _020664_, _020665_);
  or g_112678_(_020662_, _020663_, _020666_);
  and g_112679_(_020659_, _020665_, _020667_);
  or g_112680_(_020660_, _020666_, _020669_);
  and g_112681_(_020658_, _020669_, _020670_);
  or g_112682_(_020656_, _020667_, _020671_);
  and g_112683_(_020660_, _020666_, _020672_);
  or g_112684_(_020659_, _020665_, _020673_);
  and g_112685_(_020649_, _020654_, _020674_);
  or g_112686_(_020648_, _020655_, _020675_);
  and g_112687_(_020673_, _020675_, _020676_);
  or g_112688_(_020672_, _020674_, _020677_);
  and g_112689_(_020670_, _020676_, _020678_);
  or g_112690_(_020671_, _020677_, _020680_);
  xor g_112691_(out[403], out[404], _020681_);
  xor g_112692_(_053885_, out[404], _020682_);
  or g_112693_(_020457_, _020527_, _020683_);
  not g_112694_(_020683_, _020684_);
  and g_112695_(_020464_, _020527_, _020685_);
  not g_112696_(_020685_, _020686_);
  and g_112697_(_020683_, _020686_, _020687_);
  or g_112698_(_020684_, _020685_, _020688_);
  and g_112699_(_020682_, _020688_, _020689_);
  or g_112700_(_020681_, _020687_, _020691_);
  xor g_112701_(out[405], _020576_, _020692_);
  xor g_112702_(_053863_, _020576_, _020693_);
  or g_112703_(_020467_, _020527_, _020694_);
  not g_112704_(_020694_, _020695_);
  and g_112705_(_020475_, _020527_, _020696_);
  not g_112706_(_020696_, _020697_);
  and g_112707_(_020694_, _020697_, _020698_);
  or g_112708_(_020695_, _020696_, _020699_);
  and g_112709_(_020692_, _020699_, _020700_);
  or g_112710_(_020693_, _020698_, _020702_);
  and g_112711_(_020691_, _020702_, _020703_);
  or g_112712_(_020689_, _020700_, _020704_);
  and g_112713_(_020693_, _020698_, _020705_);
  or g_112714_(_020692_, _020699_, _020706_);
  and g_112715_(_020681_, _020687_, _020707_);
  or g_112716_(_020682_, _020688_, _020708_);
  and g_112717_(_020706_, _020708_, _020709_);
  or g_112718_(_020705_, _020707_, _020710_);
  and g_112719_(_020703_, _020709_, _020711_);
  or g_112720_(_020704_, _020710_, _020713_);
  and g_112721_(_020678_, _020711_, _020714_);
  or g_112722_(_020680_, _020713_, _020715_);
  and g_112723_(_020645_, _020714_, _020716_);
  or g_112724_(_020647_, _020715_, _020717_);
  and g_112725_(_020575_, _020716_, _020718_);
  or g_112726_(_020574_, _020717_, _020719_);
  and g_112727_(_020704_, _020706_, _020720_);
  or g_112728_(_020703_, _020705_, _020721_);
  and g_112729_(_020678_, _020720_, _020722_);
  or g_112730_(_020680_, _020721_, _020724_);
  and g_112731_(_020671_, _020675_, _020725_);
  or g_112732_(_020670_, _020674_, _020726_);
  and g_112733_(_020724_, _020726_, _020727_);
  or g_112734_(_020722_, _020725_, _020728_);
  and g_112735_(_020645_, _020728_, _020729_);
  or g_112736_(_020647_, _020727_, _020730_);
  and g_112737_(_020603_, _020607_, _020731_);
  or g_112738_(_020601_, _020606_, _020732_);
  and g_112739_(_020633_, _020639_, _020733_);
  or g_112740_(_020632_, _020640_, _020735_);
  and g_112741_(_020618_, _020733_, _020736_);
  or g_112742_(_020617_, _020735_, _020737_);
  and g_112743_(_020732_, _020737_, _020738_);
  or g_112744_(_020731_, _020736_, _020739_);
  or g_112745_(_020729_, _020739_, _020740_);
  and g_112746_(_020719_, _020738_, _020741_);
  and g_112747_(_020730_, _020741_, _020742_);
  or g_112748_(_020718_, _020740_, _020743_);
  and g_112749_(_004707_, _020561_, _020744_);
  or g_112750_(out[400], _020562_, _020746_);
  or g_112751_(_020554_, _020565_, _020747_);
  not g_112752_(_020747_, _020748_);
  and g_112753_(_020716_, _020748_, _020749_);
  or g_112754_(_020717_, _020747_, _020750_);
  and g_112755_(_020746_, _020749_, _020751_);
  or g_112756_(_020744_, _020750_, _020752_);
  and g_112757_(_020743_, _020752_, _020753_);
  or g_112758_(_020742_, _020751_, _020754_);
  and g_112759_(_020530_, _020754_, _020755_);
  and g_112760_(_053918_, _020753_, _020757_);
  or g_112761_(_020755_, _020757_, _020758_);
  and g_112762_(_020545_, _020754_, _020759_);
  and g_112763_(_053907_, _020753_, _020760_);
  or g_112764_(_020759_, _020760_, _020761_);
  or g_112765_(out[418], _020761_, _020762_);
  and g_112766_(out[403], _020753_, _020763_);
  or g_112767_(_053885_, _020754_, _020764_);
  and g_112768_(_020537_, _020754_, _020765_);
  or g_112769_(_020535_, _020753_, _020766_);
  and g_112770_(_020764_, _020766_, _020768_);
  or g_112771_(_020763_, _020765_, _020769_);
  or g_112772_(_053984_, _020769_, _020770_);
  and g_112773_(_053984_, _020769_, _020771_);
  xor g_112774_(out[418], _020761_, _020772_);
  xor g_112775_(_054006_, _020761_, _020773_);
  xor g_112776_(out[419], _020768_, _020774_);
  xor g_112777_(_053984_, _020768_, _020775_);
  and g_112778_(_020772_, _020774_, _020776_);
  or g_112779_(_020773_, _020775_, _020777_);
  or g_112780_(out[417], _020758_, _020779_);
  and g_112781_(_020562_, _020754_, _020780_);
  and g_112782_(_004707_, _020753_, _020781_);
  or g_112783_(_020780_, _020781_, _020782_);
  and g_112784_(out[416], _020782_, _020783_);
  not g_112785_(_020783_, _020784_);
  xor g_112786_(out[417], _020758_, _020785_);
  xor g_112787_(_054017_, _020758_, _020786_);
  and g_112788_(_020784_, _020785_, _020787_);
  or g_112789_(_020783_, _020786_, _020788_);
  and g_112790_(_020779_, _020788_, _020790_);
  or g_112791_(_020777_, _020790_, _020791_);
  or g_112792_(_020762_, _020771_, _020792_);
  and g_112793_(_020770_, _020792_, _020793_);
  and g_112794_(_020791_, _020793_, _020794_);
  and g_112795_(_020595_, _020597_, _020795_);
  or g_112796_(_020596_, _020598_, _020796_);
  and g_112797_(out[419], out[420], _020797_);
  or g_112798_(out[421], _020797_, _020798_);
  or g_112799_(out[422], _020798_, _020799_);
  or g_112800_(out[423], _020799_, _020801_);
  or g_112801_(out[424], _020801_, _020802_);
  and g_112802_(out[425], _020802_, _020803_);
  or g_112803_(out[426], _020803_, _020804_);
  xor g_112804_(out[427], _020804_, _020805_);
  xor g_112805_(_004729_, _020804_, _020806_);
  or g_112806_(_020796_, _020805_, _020807_);
  and g_112807_(_020796_, _020805_, _020808_);
  xor g_112808_(_020796_, _020805_, _020809_);
  xor g_112809_(_020795_, _020805_, _020810_);
  xor g_112810_(out[426], _020803_, _020812_);
  not g_112811_(_020812_, _020813_);
  and g_112812_(_020584_, _020753_, _020814_);
  and g_112813_(_020592_, _020754_, _020815_);
  or g_112814_(_020814_, _020815_, _020816_);
  or g_112815_(_020813_, _020816_, _020817_);
  xor g_112816_(_054028_, _020802_, _020818_);
  and g_112817_(_020615_, _020753_, _020819_);
  and g_112818_(_020614_, _020754_, _020820_);
  or g_112819_(_020819_, _020820_, _020821_);
  or g_112820_(_020818_, _020821_, _020823_);
  xor g_112821_(out[424], _020801_, _020824_);
  and g_112822_(_020620_, _020753_, _020825_);
  and g_112823_(_020627_, _020754_, _020826_);
  or g_112824_(_020825_, _020826_, _020827_);
  and g_112825_(_020824_, _020827_, _020828_);
  not g_112826_(_020828_, _020829_);
  and g_112827_(_020818_, _020821_, _020830_);
  not g_112828_(_020830_, _020831_);
  and g_112829_(_020829_, _020831_, _020832_);
  or g_112830_(_020828_, _020830_, _020834_);
  or g_112831_(_020824_, _020827_, _020835_);
  xor g_112832_(_020813_, _020816_, _020836_);
  xor g_112833_(_020812_, _020816_, _020837_);
  and g_112834_(_020809_, _020836_, _020838_);
  or g_112835_(_020810_, _020837_, _020839_);
  and g_112836_(_020823_, _020835_, _020840_);
  not g_112837_(_020840_, _020841_);
  and g_112838_(_020832_, _020840_, _020842_);
  or g_112839_(_020834_, _020841_, _020843_);
  and g_112840_(_020838_, _020842_, _020845_);
  or g_112841_(_020839_, _020843_, _020846_);
  xor g_112842_(out[423], _020799_, _020847_);
  and g_112843_(_020649_, _020753_, _020848_);
  or g_112844_(_020648_, _020754_, _020849_);
  and g_112845_(_020655_, _020754_, _020850_);
  or g_112846_(_020654_, _020753_, _020851_);
  and g_112847_(_020849_, _020851_, _020852_);
  or g_112848_(_020848_, _020850_, _020853_);
  and g_112849_(_020847_, _020853_, _020854_);
  xor g_112850_(out[422], _020798_, _020856_);
  and g_112851_(_020659_, _020753_, _020857_);
  or g_112852_(_020660_, _020754_, _020858_);
  and g_112853_(_020666_, _020754_, _020859_);
  or g_112854_(_020665_, _020753_, _020860_);
  and g_112855_(_020858_, _020860_, _020861_);
  or g_112856_(_020857_, _020859_, _020862_);
  and g_112857_(_020856_, _020861_, _020863_);
  or g_112858_(_020854_, _020863_, _020864_);
  or g_112859_(_020847_, _020853_, _020865_);
  xor g_112860_(_020847_, _020853_, _020867_);
  xor g_112861_(_020847_, _020852_, _020868_);
  xor g_112862_(_020856_, _020861_, _020869_);
  xor g_112863_(_020856_, _020862_, _020870_);
  and g_112864_(_020867_, _020869_, _020871_);
  or g_112865_(_020868_, _020870_, _020872_);
  xor g_112866_(out[421], _020797_, _020873_);
  and g_112867_(_020693_, _020753_, _020874_);
  and g_112868_(_020699_, _020754_, _020875_);
  or g_112869_(_020874_, _020875_, _020876_);
  and g_112870_(_020873_, _020876_, _020878_);
  not g_112871_(_020878_, _020879_);
  xor g_112872_(_053984_, out[420], _020880_);
  and g_112873_(_020681_, _020753_, _020881_);
  and g_112874_(_020688_, _020754_, _020882_);
  or g_112875_(_020881_, _020882_, _020883_);
  and g_112876_(_020880_, _020883_, _020884_);
  not g_112877_(_020884_, _020885_);
  and g_112878_(_020879_, _020885_, _020886_);
  or g_112879_(_020878_, _020884_, _020887_);
  or g_112880_(_020873_, _020876_, _020889_);
  or g_112881_(_020880_, _020883_, _020890_);
  and g_112882_(_020889_, _020890_, _020891_);
  not g_112883_(_020891_, _020892_);
  and g_112884_(_020886_, _020891_, _020893_);
  or g_112885_(_020887_, _020892_, _020894_);
  and g_112886_(_020871_, _020893_, _020895_);
  or g_112887_(_020872_, _020894_, _020896_);
  and g_112888_(_020845_, _020895_, _020897_);
  and g_112889_(_020823_, _020834_, _020898_);
  not g_112890_(_020898_, _020900_);
  or g_112891_(_020839_, _020900_, _020901_);
  or g_112892_(_020808_, _020817_, _020902_);
  and g_112893_(_020807_, _020902_, _020903_);
  and g_112894_(_020901_, _020903_, _020904_);
  and g_112895_(_020864_, _020865_, _020905_);
  and g_112896_(_020887_, _020889_, _020906_);
  and g_112897_(_020871_, _020906_, _020907_);
  or g_112898_(_020905_, _020907_, _020908_);
  not g_112899_(_020908_, _020909_);
  or g_112900_(_020794_, _020896_, _020911_);
  and g_112901_(_020909_, _020911_, _020912_);
  or g_112902_(_020846_, _020912_, _020913_);
  and g_112903_(_020904_, _020913_, _020914_);
  or g_112904_(out[416], _020782_, _020915_);
  and g_112905_(_020776_, _020915_, _020916_);
  and g_112906_(_020787_, _020916_, _020917_);
  and g_112907_(_020897_, _020917_, _020918_);
  or g_112908_(_020914_, _020918_, _020919_);
  not g_112909_(_020919_, _020920_);
  and g_112910_(_020758_, _020919_, _020922_);
  and g_112911_(_054017_, _020920_, _020923_);
  or g_112912_(_020922_, _020923_, _020924_);
  and g_112913_(out[419], _020920_, _020925_);
  and g_112914_(_020769_, _020919_, _020926_);
  or g_112915_(_020925_, _020926_, _020927_);
  or g_112916_(_054083_, _020927_, _020928_);
  and g_112917_(_020761_, _020919_, _020929_);
  and g_112918_(_054006_, _020920_, _020930_);
  or g_112919_(_020929_, _020930_, _020931_);
  and g_112920_(_054083_, _020927_, _020933_);
  or g_112921_(out[434], _020931_, _020934_);
  xor g_112922_(_054083_, _020927_, _020935_);
  xor g_112923_(out[435], _020927_, _020936_);
  xor g_112924_(out[434], _020931_, _020937_);
  xor g_112925_(_054105_, _020931_, _020938_);
  and g_112926_(_020935_, _020937_, _020939_);
  or g_112927_(_020936_, _020938_, _020940_);
  or g_112928_(out[433], _020924_, _020941_);
  and g_112929_(_020782_, _020919_, _020942_);
  and g_112930_(_004740_, _020920_, _020944_);
  or g_112931_(_020942_, _020944_, _020945_);
  and g_112932_(out[432], _020945_, _020946_);
  not g_112933_(_020946_, _020947_);
  xor g_112934_(out[433], _020924_, _020948_);
  xor g_112935_(_054116_, _020924_, _020949_);
  and g_112936_(_020947_, _020948_, _020950_);
  or g_112937_(_020946_, _020949_, _020951_);
  and g_112938_(_020941_, _020951_, _020952_);
  or g_112939_(_020940_, _020952_, _020953_);
  and g_112940_(_020928_, _020934_, _020955_);
  or g_112941_(_020933_, _020955_, _020956_);
  and g_112942_(_020953_, _020956_, _020957_);
  and g_112943_(out[435], out[436], _020958_);
  or g_112944_(out[437], _020958_, _020959_);
  or g_112945_(out[438], _020959_, _020960_);
  or g_112946_(out[439], _020960_, _020961_);
  or g_112947_(out[440], _020961_, _020962_);
  and g_112948_(out[441], _020962_, _020963_);
  or g_112949_(out[442], _020963_, _020964_);
  xor g_112950_(out[442], _020963_, _020966_);
  not g_112951_(_020966_, _020967_);
  or g_112952_(_020813_, _020919_, _020968_);
  not g_112953_(_020968_, _020969_);
  and g_112954_(_020816_, _020919_, _020970_);
  not g_112955_(_020970_, _020971_);
  and g_112956_(_020968_, _020971_, _020972_);
  or g_112957_(_020969_, _020970_, _020973_);
  and g_112958_(_020966_, _020972_, _020974_);
  or g_112959_(_020967_, _020973_, _020975_);
  and g_112960_(_020795_, _020805_, _020977_);
  or g_112961_(_020796_, _020806_, _020978_);
  xor g_112962_(out[443], _020964_, _020979_);
  xor g_112963_(_004762_, _020964_, _020980_);
  and g_112964_(_020977_, _020980_, _020981_);
  or g_112965_(_020978_, _020979_, _020982_);
  and g_112966_(_020975_, _020982_, _020983_);
  or g_112967_(_020974_, _020981_, _020984_);
  and g_112968_(_020978_, _020979_, _020985_);
  and g_112969_(_020967_, _020973_, _020986_);
  or g_112970_(_020985_, _020986_, _020988_);
  not g_112971_(_020988_, _020989_);
  and g_112972_(_020983_, _020989_, _020990_);
  or g_112973_(_020984_, _020988_, _020991_);
  xor g_112974_(out[440], _020961_, _020992_);
  not g_112975_(_020992_, _020993_);
  or g_112976_(_020824_, _020919_, _020994_);
  and g_112977_(_020827_, _020919_, _020995_);
  not g_112978_(_020995_, _020996_);
  and g_112979_(_020994_, _020996_, _020997_);
  not g_112980_(_020997_, _020999_);
  or g_112981_(_020993_, _020997_, _021000_);
  xor g_112982_(out[441], _020962_, _021001_);
  xor g_112983_(_054127_, _020962_, _021002_);
  or g_112984_(_020818_, _020919_, _021003_);
  and g_112985_(_020821_, _020919_, _021004_);
  not g_112986_(_021004_, _021005_);
  and g_112987_(_021003_, _021005_, _021006_);
  or g_112988_(_021001_, _021006_, _021007_);
  and g_112989_(_021000_, _021007_, _021008_);
  not g_112990_(_021008_, _021010_);
  and g_112991_(_021001_, _021006_, _021011_);
  not g_112992_(_021011_, _021012_);
  and g_112993_(_020993_, _020997_, _021013_);
  or g_112994_(_020992_, _020999_, _021014_);
  and g_112995_(_021012_, _021014_, _021015_);
  or g_112996_(_021011_, _021013_, _021016_);
  and g_112997_(_021008_, _021015_, _021017_);
  or g_112998_(_021010_, _021016_, _021018_);
  and g_112999_(_020990_, _021017_, _021019_);
  or g_113000_(_020991_, _021018_, _021021_);
  xor g_113001_(out[437], _020958_, _021022_);
  xor g_113002_(_054061_, _020958_, _021023_);
  or g_113003_(_020873_, _020919_, _021024_);
  not g_113004_(_021024_, _021025_);
  and g_113005_(_020876_, _020919_, _021026_);
  not g_113006_(_021026_, _021027_);
  and g_113007_(_021024_, _021027_, _021028_);
  or g_113008_(_021025_, _021026_, _021029_);
  and g_113009_(_021023_, _021028_, _021030_);
  xor g_113010_(out[438], _020959_, _021032_);
  xor g_113011_(_054072_, _020959_, _021033_);
  and g_113012_(_020861_, _020919_, _021034_);
  or g_113013_(_020862_, _020920_, _021035_);
  or g_113014_(_020856_, _020919_, _021036_);
  not g_113015_(_021036_, _021037_);
  or g_113016_(_021034_, _021037_, _021038_);
  and g_113017_(_021035_, _021036_, _021039_);
  and g_113018_(_021033_, _021039_, _021040_);
  or g_113019_(_021030_, _021040_, _021041_);
  xor g_113020_(out[439], _020960_, _021043_);
  not g_113021_(_021043_, _021044_);
  or g_113022_(_020847_, _020919_, _021045_);
  not g_113023_(_021045_, _021046_);
  and g_113024_(_020853_, _020919_, _021047_);
  or g_113025_(_020852_, _020920_, _021048_);
  and g_113026_(_021045_, _021048_, _021049_);
  or g_113027_(_021046_, _021047_, _021050_);
  and g_113028_(_021044_, _021049_, _021051_);
  xor g_113029_(out[435], out[436], _021052_);
  xor g_113030_(_054083_, out[436], _021054_);
  or g_113031_(_020880_, _020919_, _021055_);
  not g_113032_(_021055_, _021056_);
  and g_113033_(_020883_, _020919_, _021057_);
  not g_113034_(_021057_, _021058_);
  and g_113035_(_021055_, _021058_, _021059_);
  or g_113036_(_021056_, _021057_, _021060_);
  and g_113037_(_021052_, _021059_, _021061_);
  or g_113038_(_021051_, _021061_, _021062_);
  or g_113039_(_021041_, _021062_, _021063_);
  not g_113040_(_021063_, _021065_);
  and g_113041_(_021043_, _021050_, _021066_);
  or g_113042_(_021044_, _021049_, _021067_);
  and g_113043_(_021032_, _021038_, _021068_);
  or g_113044_(_021033_, _021039_, _021069_);
  and g_113045_(_021067_, _021069_, _021070_);
  or g_113046_(_021066_, _021068_, _021071_);
  and g_113047_(_021054_, _021060_, _021072_);
  or g_113048_(_021052_, _021059_, _021073_);
  and g_113049_(_021022_, _021029_, _021074_);
  or g_113050_(_021023_, _021028_, _021076_);
  and g_113051_(_021073_, _021076_, _021077_);
  or g_113052_(_021072_, _021074_, _021078_);
  and g_113053_(_021070_, _021077_, _021079_);
  or g_113054_(_021071_, _021078_, _021080_);
  and g_113055_(_021065_, _021079_, _021081_);
  or g_113056_(_021063_, _021080_, _021082_);
  and g_113057_(_021019_, _021081_, _021083_);
  or g_113058_(_021021_, _021082_, _021084_);
  or g_113059_(_020957_, _021084_, _021085_);
  or g_113060_(_021041_, _021077_, _021087_);
  and g_113061_(_021070_, _021087_, _021088_);
  or g_113062_(_021051_, _021088_, _021089_);
  or g_113063_(_021021_, _021089_, _021090_);
  or g_113064_(_020983_, _020985_, _021091_);
  or g_113065_(_021008_, _021011_, _021092_);
  or g_113066_(_020991_, _021092_, _021093_);
  and g_113067_(_021091_, _021093_, _021094_);
  and g_113068_(_021090_, _021094_, _021095_);
  and g_113069_(_021085_, _021095_, _021096_);
  or g_113070_(out[432], _020945_, _021098_);
  and g_113071_(_020939_, _021098_, _021099_);
  and g_113072_(_020950_, _021099_, _021100_);
  and g_113073_(_021083_, _021100_, _021101_);
  or g_113074_(_021096_, _021101_, _021102_);
  not g_113075_(_021102_, _021103_);
  and g_113076_(_020924_, _021102_, _021104_);
  not g_113077_(_021104_, _021105_);
  or g_113078_(out[433], _021102_, _021106_);
  not g_113079_(_021106_, _021107_);
  and g_113080_(_021105_, _021106_, _021109_);
  or g_113081_(_021104_, _021107_, _021110_);
  and g_113082_(out[451], out[452], _021111_);
  or g_113083_(out[453], _021111_, _021112_);
  or g_113084_(out[454], _021112_, _021113_);
  xor g_113085_(_054171_, _021112_, _021114_);
  and g_113086_(_021032_, _021103_, _021115_);
  and g_113087_(_021039_, _021102_, _021116_);
  or g_113088_(_021115_, _021116_, _021117_);
  or g_113089_(_021114_, _021117_, _021118_);
  not g_113090_(_021118_, _021120_);
  or g_113091_(out[455], _021113_, _021121_);
  xor g_113092_(out[455], _021113_, _021122_);
  or g_113093_(_021043_, _021102_, _021123_);
  not g_113094_(_021123_, _021124_);
  and g_113095_(_021050_, _021102_, _021125_);
  or g_113096_(_021124_, _021125_, _021126_);
  and g_113097_(_021122_, _021126_, _021127_);
  or g_113098_(_021120_, _021127_, _021128_);
  not g_113099_(_021128_, _021129_);
  and g_113100_(out[435], _021103_, _021131_);
  and g_113101_(_020927_, _021102_, _021132_);
  or g_113102_(_021131_, _021132_, _021133_);
  not g_113103_(_021133_, _021134_);
  and g_113104_(out[451], _021134_, _021135_);
  or g_113105_(_054182_, _021133_, _021136_);
  and g_113106_(_020931_, _021102_, _021137_);
  not g_113107_(_021137_, _021138_);
  or g_113108_(out[434], _021102_, _021139_);
  not g_113109_(_021139_, _021140_);
  and g_113110_(_021138_, _021139_, _021142_);
  or g_113111_(_021137_, _021140_, _021143_);
  and g_113112_(out[450], _021143_, _021144_);
  not g_113113_(_021144_, _021145_);
  and g_113114_(_020945_, _021102_, _021146_);
  not g_113115_(_021146_, _021147_);
  or g_113116_(out[432], _021102_, _021148_);
  not g_113117_(_021148_, _021149_);
  and g_113118_(_021147_, _021148_, _021150_);
  or g_113119_(_021146_, _021149_, _021151_);
  and g_113120_(out[448], _021151_, _021153_);
  or g_113121_(_004806_, _021150_, _021154_);
  and g_113122_(out[449], _021110_, _021155_);
  or g_113123_(_054215_, _021109_, _021156_);
  and g_113124_(_021154_, _021156_, _021157_);
  or g_113125_(_021153_, _021155_, _021158_);
  and g_113126_(_054204_, _021142_, _021159_);
  or g_113127_(out[450], _021143_, _021160_);
  and g_113128_(_054215_, _021109_, _021161_);
  or g_113129_(out[449], _021110_, _021162_);
  and g_113130_(_021160_, _021162_, _021164_);
  or g_113131_(_021159_, _021161_, _021165_);
  and g_113132_(_021158_, _021164_, _021166_);
  or g_113133_(_021157_, _021165_, _021167_);
  and g_113134_(_021145_, _021167_, _021168_);
  or g_113135_(_021144_, _021166_, _021169_);
  and g_113136_(_021136_, _021169_, _021170_);
  or g_113137_(_021135_, _021168_, _021171_);
  xor g_113138_(out[451], out[452], _021172_);
  or g_113139_(_021054_, _021102_, _021173_);
  or g_113140_(_021059_, _021103_, _021175_);
  and g_113141_(_021173_, _021175_, _021176_);
  and g_113142_(_021172_, _021176_, _021177_);
  not g_113143_(_021177_, _021178_);
  or g_113144_(out[451], _021134_, _021179_);
  and g_113145_(_021178_, _021179_, _021180_);
  not g_113146_(_021180_, _021181_);
  and g_113147_(_021171_, _021180_, _021182_);
  or g_113148_(_021170_, _021181_, _021183_);
  xor g_113149_(out[453], _021111_, _021184_);
  not g_113150_(_021184_, _021186_);
  or g_113151_(_021022_, _021102_, _021187_);
  or g_113152_(_021028_, _021103_, _021188_);
  and g_113153_(_021187_, _021188_, _021189_);
  not g_113154_(_021189_, _021190_);
  or g_113155_(_021186_, _021189_, _021191_);
  or g_113156_(_021172_, _021176_, _021192_);
  and g_113157_(_021191_, _021192_, _021193_);
  not g_113158_(_021193_, _021194_);
  and g_113159_(_021183_, _021193_, _021195_);
  or g_113160_(_021182_, _021194_, _021197_);
  or g_113161_(_021184_, _021190_, _021198_);
  and g_113162_(_021114_, _021117_, _021199_);
  not g_113163_(_021199_, _021200_);
  and g_113164_(_021198_, _021200_, _021201_);
  not g_113165_(_021201_, _021202_);
  and g_113166_(_021197_, _021201_, _021203_);
  or g_113167_(_021195_, _021202_, _021204_);
  and g_113168_(_021129_, _021204_, _021205_);
  or g_113169_(_021128_, _021203_, _021206_);
  or g_113170_(out[456], _021121_, _021208_);
  xor g_113171_(out[456], _021121_, _021209_);
  not g_113172_(_021209_, _021210_);
  and g_113173_(_020992_, _021103_, _021211_);
  and g_113174_(_020997_, _021102_, _021212_);
  or g_113175_(_021211_, _021212_, _021213_);
  not g_113176_(_021213_, _021214_);
  or g_113177_(_021210_, _021213_, _021215_);
  and g_113178_(out[457], _021208_, _021216_);
  xor g_113179_(out[457], _021208_, _021217_);
  not g_113180_(_021217_, _021219_);
  or g_113181_(_021002_, _021102_, _021220_);
  or g_113182_(_021006_, _021103_, _021221_);
  and g_113183_(_021220_, _021221_, _021222_);
  not g_113184_(_021222_, _021223_);
  and g_113185_(_021217_, _021222_, _021224_);
  or g_113186_(_021217_, _021222_, _021225_);
  xor g_113187_(_021217_, _021222_, _021226_);
  and g_113188_(_021215_, _021226_, _021227_);
  not g_113189_(_021227_, _021228_);
  or g_113190_(out[458], _021216_, _021230_);
  xor g_113191_(_004817_, _021216_, _021231_);
  and g_113192_(_020966_, _021103_, _021232_);
  and g_113193_(_020973_, _021102_, _021233_);
  or g_113194_(_021232_, _021233_, _021234_);
  or g_113195_(_021231_, _021234_, _021235_);
  or g_113196_(_020978_, _020980_, _021236_);
  not g_113197_(_021236_, _021237_);
  xor g_113198_(out[459], _021230_, _021238_);
  or g_113199_(_021236_, _021238_, _021239_);
  and g_113200_(_021235_, _021239_, _021241_);
  not g_113201_(_021241_, _021242_);
  and g_113202_(_021236_, _021238_, _021243_);
  and g_113203_(_021231_, _021234_, _021244_);
  or g_113204_(_021243_, _021244_, _021245_);
  not g_113205_(_021245_, _021246_);
  and g_113206_(_021210_, _021213_, _021247_);
  or g_113207_(_021209_, _021214_, _021248_);
  or g_113208_(_021122_, _021126_, _021249_);
  not g_113209_(_021249_, _021250_);
  and g_113210_(_021248_, _021249_, _021252_);
  or g_113211_(_021247_, _021250_, _021253_);
  and g_113212_(_021246_, _021252_, _021254_);
  or g_113213_(_021245_, _021253_, _021255_);
  and g_113214_(_021241_, _021254_, _021256_);
  or g_113215_(_021242_, _021255_, _021257_);
  and g_113216_(_021227_, _021256_, _021258_);
  or g_113217_(_021228_, _021257_, _021259_);
  and g_113218_(_021206_, _021258_, _021260_);
  or g_113219_(_021205_, _021259_, _021261_);
  or g_113220_(_021241_, _021243_, _021263_);
  and g_113221_(_021215_, _021225_, _021264_);
  or g_113222_(_021224_, _021245_, _021265_);
  or g_113223_(_021264_, _021265_, _021266_);
  and g_113224_(_021263_, _021266_, _021267_);
  not g_113225_(_021267_, _021268_);
  and g_113226_(_021261_, _021267_, _021269_);
  or g_113227_(_021260_, _021268_, _021270_);
  and g_113228_(_021164_, _021180_, _021271_);
  and g_113229_(_021193_, _021201_, _021272_);
  and g_113230_(_021271_, _021272_, _021274_);
  not g_113231_(_021274_, _021275_);
  and g_113232_(_004806_, _021150_, _021276_);
  or g_113233_(out[448], _021151_, _021277_);
  and g_113234_(_021136_, _021145_, _021278_);
  or g_113235_(_021135_, _021144_, _021279_);
  and g_113236_(_021277_, _021278_, _021280_);
  or g_113237_(_021276_, _021279_, _021281_);
  or g_113238_(_021128_, _021158_, _021282_);
  not g_113239_(_021282_, _021283_);
  and g_113240_(_021280_, _021283_, _021285_);
  or g_113241_(_021281_, _021282_, _021286_);
  and g_113242_(_021274_, _021285_, _021287_);
  or g_113243_(_021275_, _021286_, _021288_);
  and g_113244_(_021258_, _021287_, _021289_);
  or g_113245_(_021259_, _021288_, _021290_);
  and g_113246_(_021270_, _021290_, _021291_);
  or g_113247_(_021269_, _021289_, _021292_);
  and g_113248_(_021110_, _021292_, _021293_);
  or g_113249_(_021109_, _021291_, _021294_);
  and g_113250_(_054215_, _021291_, _021296_);
  or g_113251_(out[449], _021292_, _021297_);
  and g_113252_(_021294_, _021297_, _021298_);
  or g_113253_(_021293_, _021296_, _021299_);
  and g_113254_(out[467], out[468], _021300_);
  or g_113255_(out[469], _021300_, _021301_);
  or g_113256_(out[470], _021301_, _021302_);
  or g_113257_(out[471], _021302_, _021303_);
  or g_113258_(out[472], _021303_, _021304_);
  and g_113259_(out[473], _021304_, _021305_);
  or g_113260_(out[474], _021305_, _021307_);
  xor g_113261_(out[474], _021305_, _021308_);
  or g_113262_(_021231_, _021292_, _021309_);
  and g_113263_(_021234_, _021292_, _021310_);
  not g_113264_(_021310_, _021311_);
  and g_113265_(_021309_, _021311_, _021312_);
  and g_113266_(_021308_, _021312_, _021313_);
  not g_113267_(_021313_, _021314_);
  and g_113268_(_021237_, _021238_, _021315_);
  not g_113269_(_021315_, _021316_);
  xor g_113270_(out[475], _021307_, _021318_);
  not g_113271_(_021318_, _021319_);
  and g_113272_(_021315_, _021319_, _021320_);
  or g_113273_(_021316_, _021318_, _021321_);
  and g_113274_(_021314_, _021321_, _021322_);
  or g_113275_(_021313_, _021320_, _021323_);
  or g_113276_(_021308_, _021312_, _021324_);
  not g_113277_(_021324_, _021325_);
  and g_113278_(_021316_, _021318_, _021326_);
  or g_113279_(_021315_, _021319_, _021327_);
  and g_113280_(_021324_, _021327_, _021329_);
  or g_113281_(_021325_, _021326_, _021330_);
  and g_113282_(_021322_, _021329_, _021331_);
  or g_113283_(_021323_, _021330_, _021332_);
  xor g_113284_(out[472], _021303_, _021333_);
  not g_113285_(_021333_, _021334_);
  or g_113286_(_021210_, _021292_, _021335_);
  not g_113287_(_021335_, _021336_);
  and g_113288_(_021213_, _021292_, _021337_);
  or g_113289_(_021336_, _021337_, _021338_);
  not g_113290_(_021338_, _021340_);
  and g_113291_(_021333_, _021340_, _021341_);
  or g_113292_(_021334_, _021338_, _021342_);
  xor g_113293_(out[473], _021304_, _021343_);
  xor g_113294_(_054325_, _021304_, _021344_);
  or g_113295_(_021219_, _021292_, _021345_);
  not g_113296_(_021345_, _021346_);
  and g_113297_(_021223_, _021292_, _021347_);
  not g_113298_(_021347_, _021348_);
  and g_113299_(_021345_, _021348_, _021349_);
  or g_113300_(_021346_, _021347_, _021351_);
  and g_113301_(_021344_, _021351_, _021352_);
  or g_113302_(_021343_, _021349_, _021353_);
  and g_113303_(_021342_, _021353_, _021354_);
  or g_113304_(_021341_, _021352_, _021355_);
  or g_113305_(_021333_, _021340_, _021356_);
  and g_113306_(_021343_, _021349_, _021357_);
  or g_113307_(_021344_, _021351_, _021358_);
  and g_113308_(_021356_, _021358_, _021359_);
  and g_113309_(_021354_, _021359_, _021360_);
  and g_113310_(_021331_, _021360_, _021362_);
  not g_113311_(_021362_, _021363_);
  xor g_113312_(out[471], _021302_, _021364_);
  xor g_113313_(_054237_, _021302_, _021365_);
  or g_113314_(_021122_, _021292_, _021366_);
  not g_113315_(_021366_, _021367_);
  and g_113316_(_021126_, _021292_, _021368_);
  not g_113317_(_021368_, _021369_);
  and g_113318_(_021366_, _021369_, _021370_);
  or g_113319_(_021367_, _021368_, _021371_);
  and g_113320_(_021364_, _021371_, _021373_);
  xor g_113321_(out[469], _021300_, _021374_);
  xor g_113322_(_054259_, _021300_, _021375_);
  or g_113323_(_021184_, _021292_, _021376_);
  and g_113324_(_021190_, _021292_, _021377_);
  not g_113325_(_021377_, _021378_);
  and g_113326_(_021376_, _021378_, _021379_);
  not g_113327_(_021379_, _021380_);
  and g_113328_(_021375_, _021379_, _021381_);
  or g_113329_(_021373_, _021381_, _021382_);
  not g_113330_(_021382_, _021384_);
  or g_113331_(_021364_, _021371_, _021385_);
  xor g_113332_(out[470], _021301_, _021386_);
  not g_113333_(_021386_, _021387_);
  or g_113334_(_021114_, _021292_, _021388_);
  and g_113335_(_021117_, _021292_, _021389_);
  not g_113336_(_021389_, _021390_);
  and g_113337_(_021388_, _021390_, _021391_);
  not g_113338_(_021391_, _021392_);
  and g_113339_(_021386_, _021391_, _021393_);
  xor g_113340_(_021386_, _021391_, _021395_);
  and g_113341_(_021385_, _021395_, _021396_);
  not g_113342_(_021396_, _021397_);
  and g_113343_(_021384_, _021396_, _021398_);
  or g_113344_(_021382_, _021397_, _021399_);
  xor g_113345_(out[467], out[468], _021400_);
  xor g_113346_(_054281_, out[468], _021401_);
  or g_113347_(_021172_, _021292_, _021402_);
  not g_113348_(_021402_, _021403_);
  and g_113349_(_021176_, _021292_, _021404_);
  not g_113350_(_021404_, _021406_);
  and g_113351_(_021402_, _021406_, _021407_);
  or g_113352_(_021403_, _021404_, _021408_);
  and g_113353_(_021400_, _021408_, _021409_);
  or g_113354_(_021401_, _021407_, _021410_);
  and g_113355_(_021401_, _021407_, _021411_);
  or g_113356_(_021400_, _021408_, _021412_);
  and g_113357_(_021374_, _021380_, _021413_);
  or g_113358_(_021375_, _021379_, _021414_);
  and g_113359_(_021412_, _021414_, _021415_);
  or g_113360_(_021411_, _021413_, _021417_);
  and g_113361_(_021410_, _021415_, _021418_);
  or g_113362_(_021409_, _021417_, _021419_);
  and g_113363_(_021398_, _021418_, _021420_);
  or g_113364_(_021399_, _021419_, _021421_);
  or g_113365_(_054182_, _021292_, _021422_);
  not g_113366_(_021422_, _021423_);
  and g_113367_(_021133_, _021292_, _021424_);
  not g_113368_(_021424_, _021425_);
  and g_113369_(_021422_, _021425_, _021426_);
  or g_113370_(_021423_, _021424_, _021428_);
  and g_113371_(out[467], _021426_, _021429_);
  or g_113372_(_054281_, _021428_, _021430_);
  and g_113373_(_021143_, _021292_, _021431_);
  not g_113374_(_021431_, _021432_);
  or g_113375_(out[450], _021292_, _021433_);
  not g_113376_(_021433_, _021434_);
  and g_113377_(_021432_, _021433_, _021435_);
  or g_113378_(_021431_, _021434_, _021436_);
  and g_113379_(out[466], _021436_, _021437_);
  or g_113380_(_054303_, _021435_, _021439_);
  and g_113381_(_021430_, _021439_, _021440_);
  or g_113382_(_021429_, _021437_, _021441_);
  and g_113383_(_054281_, _021428_, _021442_);
  or g_113384_(out[467], _021426_, _021443_);
  and g_113385_(_054303_, _021435_, _021444_);
  or g_113386_(out[466], _021436_, _021445_);
  and g_113387_(_021443_, _021445_, _021446_);
  or g_113388_(_021442_, _021444_, _021447_);
  and g_113389_(_021440_, _021446_, _021448_);
  or g_113390_(_021441_, _021447_, _021450_);
  and g_113391_(_054314_, _021298_, _021451_);
  or g_113392_(out[465], _021299_, _021452_);
  or g_113393_(_054314_, _021298_, _021453_);
  not g_113394_(_021453_, _021454_);
  and g_113395_(_021151_, _021292_, _021455_);
  or g_113396_(_021150_, _021291_, _021456_);
  and g_113397_(_004806_, _021291_, _021457_);
  or g_113398_(out[448], _021292_, _021458_);
  and g_113399_(_021456_, _021458_, _021459_);
  or g_113400_(_021455_, _021457_, _021461_);
  and g_113401_(out[464], _021461_, _021462_);
  or g_113402_(_004839_, _021459_, _021463_);
  and g_113403_(_021452_, _021463_, _021464_);
  or g_113404_(_021451_, _021462_, _021465_);
  and g_113405_(_021453_, _021464_, _021466_);
  or g_113406_(_021454_, _021465_, _021467_);
  and g_113407_(_021452_, _021467_, _021468_);
  or g_113408_(_021451_, _021466_, _021469_);
  and g_113409_(_021448_, _021469_, _021470_);
  or g_113410_(_021450_, _021468_, _021472_);
  and g_113411_(_021443_, _021444_, _021473_);
  or g_113412_(_021429_, _021473_, _021474_);
  not g_113413_(_021474_, _021475_);
  and g_113414_(_021472_, _021475_, _021476_);
  or g_113415_(_021470_, _021474_, _021477_);
  and g_113416_(_021420_, _021477_, _021478_);
  or g_113417_(_021421_, _021476_, _021479_);
  and g_113418_(_021398_, _021417_, _021480_);
  or g_113419_(_021399_, _021415_, _021481_);
  or g_113420_(_021373_, _021393_, _021483_);
  and g_113421_(_021385_, _021483_, _021484_);
  not g_113422_(_021484_, _021485_);
  and g_113423_(_021481_, _021485_, _021486_);
  or g_113424_(_021480_, _021484_, _021487_);
  and g_113425_(_021479_, _021486_, _021488_);
  or g_113426_(_021478_, _021487_, _021489_);
  and g_113427_(_021362_, _021489_, _021490_);
  or g_113428_(_021363_, _021488_, _021491_);
  and g_113429_(_021323_, _021327_, _021492_);
  or g_113430_(_021322_, _021326_, _021494_);
  and g_113431_(_021355_, _021358_, _021495_);
  or g_113432_(_021354_, _021357_, _021496_);
  and g_113433_(_021331_, _021495_, _021497_);
  or g_113434_(_021332_, _021496_, _021498_);
  and g_113435_(_021494_, _021498_, _021499_);
  or g_113436_(_021492_, _021497_, _021500_);
  and g_113437_(_021491_, _021499_, _021501_);
  or g_113438_(_021490_, _021500_, _021502_);
  and g_113439_(_004839_, _021459_, _021503_);
  or g_113440_(_021450_, _021503_, _021505_);
  not g_113441_(_021505_, _021506_);
  and g_113442_(_021466_, _021506_, _021507_);
  and g_113443_(_021362_, _021507_, _021508_);
  and g_113444_(_021420_, _021508_, _021509_);
  not g_113445_(_021509_, _021510_);
  and g_113446_(_021502_, _021510_, _021511_);
  or g_113447_(_021501_, _021509_, _021512_);
  or g_113448_(_021298_, _021511_, _021513_);
  not g_113449_(_021513_, _021514_);
  and g_113450_(_054314_, _021511_, _021516_);
  or g_113451_(out[465], _021512_, _021517_);
  and g_113452_(_021513_, _021517_, _021518_);
  or g_113453_(_021514_, _021516_, _021519_);
  and g_113454_(out[484], out[483], _021520_);
  or g_113455_(out[485], _021520_, _021521_);
  or g_113456_(out[486], _021521_, _021522_);
  or g_113457_(out[487], _021522_, _021523_);
  or g_113458_(out[488], _021523_, _021524_);
  and g_113459_(out[489], _021524_, _021525_);
  or g_113460_(out[490], _021525_, _021527_);
  xor g_113461_(out[491], _021527_, _021528_);
  xor g_113462_(_054358_, _021527_, _021529_);
  and g_113463_(out[500], out[499], _021530_);
  or g_113464_(out[501], _021530_, _021531_);
  or g_113465_(out[502], _021531_, _021532_);
  or g_113466_(out[503], _021532_, _021533_);
  or g_113467_(out[504], _021533_, _021534_);
  and g_113468_(out[505], _021534_, _021535_);
  or g_113469_(out[506], _021535_, _021536_);
  xor g_113470_(out[507], _021536_, _021538_);
  xor g_113471_(_054479_, _021536_, _021539_);
  and g_113472_(_021529_, _021538_, _021540_);
  or g_113473_(_021528_, _021539_, _021541_);
  xor g_113474_(out[489], _021524_, _021542_);
  xor g_113475_(_054457_, _021524_, _021543_);
  xor g_113476_(out[505], _021534_, _021544_);
  xor g_113477_(_054589_, _021534_, _021545_);
  and g_113478_(_021542_, _021545_, _021546_);
  or g_113479_(_021543_, _021544_, _021547_);
  xor g_113480_(out[504], _021533_, _021549_);
  xor g_113481_(_054578_, _021533_, _021550_);
  xor g_113482_(out[488], _021523_, _021551_);
  xor g_113483_(_054446_, _021523_, _021552_);
  and g_113484_(_021550_, _021551_, _021553_);
  or g_113485_(_021549_, _021552_, _021554_);
  xor g_113486_(out[487], _021522_, _021555_);
  xor g_113487_(_054369_, _021522_, _021556_);
  xor g_113488_(out[503], _021532_, _021557_);
  xor g_113489_(_054490_, _021532_, _021558_);
  and g_113490_(_021555_, _021558_, _021560_);
  or g_113491_(_021556_, _021557_, _021561_);
  xor g_113492_(out[484], out[483], _021562_);
  xor g_113493_(_054402_, out[483], _021563_);
  xor g_113494_(out[500], out[499], _021564_);
  xor g_113495_(_054523_, out[499], _021565_);
  and g_113496_(_021563_, _021564_, _021566_);
  or g_113497_(_021562_, _021565_, _021567_);
  and g_113498_(_054435_, out[499], _021568_);
  or g_113499_(out[483], _054567_, _021569_);
  and g_113500_(out[482], _054556_, _021571_);
  or g_113501_(_054424_, out[498], _021572_);
  and g_113502_(_016609_, _021572_, _021573_);
  or g_113503_(_016598_, _021571_, _021574_);
  and g_113504_(_016653_, _021573_, _021575_);
  or g_113505_(_016642_, _021574_, _021576_);
  and g_113506_(_054424_, out[498], _021577_);
  or g_113507_(out[482], _054556_, _021578_);
  and g_113508_(out[483], _054567_, _021579_);
  or g_113509_(_054435_, out[499], _021580_);
  and g_113510_(_021578_, _021580_, _021582_);
  or g_113511_(_021577_, _021579_, _021583_);
  and g_113512_(_021576_, _021582_, _021584_);
  or g_113513_(_021575_, _021583_, _021585_);
  and g_113514_(_021569_, _021585_, _021586_);
  or g_113515_(_021568_, _021584_, _021587_);
  and g_113516_(_021567_, _021587_, _021588_);
  or g_113517_(_021566_, _021586_, _021589_);
  and g_113518_(_016895_, _021588_, _021590_);
  or g_113519_(_016884_, _021589_, _021591_);
  and g_113520_(_021562_, _021565_, _021593_);
  or g_113521_(_021563_, _021564_, _021594_);
  xor g_113522_(out[485], _021520_, _021595_);
  xor g_113523_(_054391_, _021520_, _021596_);
  xor g_113524_(out[501], _021530_, _021597_);
  xor g_113525_(_054512_, _021530_, _021598_);
  and g_113526_(_021596_, _021597_, _021599_);
  or g_113527_(_021595_, _021598_, _021600_);
  and g_113528_(_021594_, _021600_, _021601_);
  or g_113529_(_021593_, _021599_, _021602_);
  and g_113530_(_021591_, _021601_, _021604_);
  or g_113531_(_021590_, _021602_, _021605_);
  and g_113532_(_021595_, _021598_, _021606_);
  or g_113533_(_021596_, _021597_, _021607_);
  xor g_113534_(out[486], _021521_, _021608_);
  xor g_113535_(_054380_, _021521_, _021609_);
  xor g_113536_(out[502], _021531_, _021610_);
  xor g_113537_(_054501_, _021531_, _021611_);
  and g_113538_(_021608_, _021611_, _021612_);
  or g_113539_(_021609_, _021610_, _021613_);
  and g_113540_(_021607_, _021613_, _021615_);
  or g_113541_(_021606_, _021612_, _021616_);
  and g_113542_(_021605_, _021615_, _021617_);
  or g_113543_(_021604_, _021616_, _021618_);
  and g_113544_(_021556_, _021557_, _021619_);
  or g_113545_(_021555_, _021558_, _021620_);
  and g_113546_(_021609_, _021610_, _021621_);
  or g_113547_(_021608_, _021611_, _021622_);
  and g_113548_(_021620_, _021622_, _021623_);
  or g_113549_(_021619_, _021621_, _021624_);
  and g_113550_(_021618_, _021623_, _021626_);
  or g_113551_(_021617_, _021624_, _021627_);
  and g_113552_(_021549_, _021552_, _021628_);
  or g_113553_(_021550_, _021551_, _021629_);
  and g_113554_(_021554_, _021561_, _021630_);
  or g_113555_(_021553_, _021560_, _021631_);
  and g_113556_(_021627_, _021630_, _021632_);
  or g_113557_(_021626_, _021631_, _021633_);
  and g_113558_(_021547_, _021629_, _021634_);
  or g_113559_(_021546_, _021628_, _021635_);
  and g_113560_(_021633_, _021634_, _021637_);
  or g_113561_(_021632_, _021635_, _021638_);
  xor g_113562_(out[490], _021525_, _021639_);
  xor g_113563_(_054468_, _021525_, _021640_);
  xor g_113564_(out[506], _021535_, _021641_);
  xor g_113565_(_054600_, _021535_, _021642_);
  and g_113566_(_021639_, _021642_, _021643_);
  or g_113567_(_021640_, _021641_, _021644_);
  and g_113568_(_021543_, _021544_, _021645_);
  or g_113569_(_021542_, _021545_, _021646_);
  and g_113570_(_021644_, _021646_, _021648_);
  or g_113571_(_021643_, _021645_, _021649_);
  and g_113572_(_021638_, _021648_, _021650_);
  or g_113573_(_021637_, _021649_, _021651_);
  and g_113574_(_021528_, _021539_, _021652_);
  or g_113575_(_021529_, _021538_, _021653_);
  and g_113576_(_021640_, _021641_, _021654_);
  or g_113577_(_021639_, _021642_, _021655_);
  and g_113578_(_021653_, _021655_, _021656_);
  or g_113579_(_021652_, _021654_, _021657_);
  and g_113580_(_021651_, _021656_, _021659_);
  or g_113581_(_021650_, _021657_, _021660_);
  and g_113582_(_021541_, _021660_, _021661_);
  or g_113583_(_021540_, _021659_, _021662_);
  or g_113584_(out[481], _021661_, _021663_);
  or g_113585_(out[497], _021662_, _021664_);
  and g_113586_(_021663_, _021664_, _021665_);
  not g_113587_(_021665_, _021666_);
  and g_113588_(out[516], out[515], _021667_);
  or g_113589_(out[517], _021667_, _021668_);
  or g_113590_(out[518], _021668_, _021670_);
  or g_113591_(out[519], _021670_, _021671_);
  xor g_113592_(out[519], _021670_, _021672_);
  xor g_113593_(_054622_, _021670_, _021673_);
  and g_113594_(_021556_, _021662_, _021674_);
  or g_113595_(_021555_, _021661_, _021675_);
  and g_113596_(_021558_, _021661_, _021676_);
  or g_113597_(_021557_, _021662_, _021677_);
  and g_113598_(_021675_, _021677_, _021678_);
  or g_113599_(_021674_, _021676_, _021679_);
  and g_113600_(_021672_, _021679_, _021681_);
  or g_113601_(_021673_, _021678_, _021682_);
  xor g_113602_(out[518], _021668_, _021683_);
  xor g_113603_(_054633_, _021668_, _021684_);
  and g_113604_(_021608_, _021662_, _021685_);
  or g_113605_(_021609_, _021661_, _021686_);
  and g_113606_(_021610_, _021661_, _021687_);
  or g_113607_(_021611_, _021662_, _021688_);
  and g_113608_(_021686_, _021688_, _021689_);
  or g_113609_(_021685_, _021687_, _021690_);
  and g_113610_(_021683_, _021689_, _021692_);
  or g_113611_(_021684_, _021690_, _021693_);
  and g_113612_(_021682_, _021693_, _021694_);
  or g_113613_(_021681_, _021692_, _021695_);
  and g_113614_(_021684_, _021690_, _021696_);
  or g_113615_(_021683_, _021689_, _021697_);
  and g_113616_(_021673_, _021678_, _021698_);
  or g_113617_(_021672_, _021679_, _021699_);
  xor g_113618_(out[517], _021667_, _021700_);
  xor g_113619_(_054644_, _021667_, _021701_);
  and g_113620_(_021596_, _021662_, _021703_);
  or g_113621_(_021595_, _021661_, _021704_);
  and g_113622_(_021598_, _021661_, _021705_);
  or g_113623_(_021597_, _021662_, _021706_);
  and g_113624_(_021704_, _021706_, _021707_);
  or g_113625_(_021703_, _021705_, _021708_);
  and g_113626_(_021701_, _021707_, _021709_);
  or g_113627_(_021700_, _021708_, _021710_);
  and g_113628_(_021699_, _021710_, _021711_);
  or g_113629_(_021698_, _021709_, _021712_);
  and g_113630_(_021697_, _021711_, _021714_);
  or g_113631_(_021696_, _021712_, _021715_);
  and g_113632_(_021694_, _021714_, _021716_);
  or g_113633_(_021695_, _021715_, _021717_);
  xor g_113634_(out[516], out[515], _021718_);
  xor g_113635_(_054655_, out[515], _021719_);
  and g_113636_(_021564_, _021661_, _021720_);
  or g_113637_(_021565_, _021662_, _021721_);
  and g_113638_(_021562_, _021662_, _021722_);
  or g_113639_(_021563_, _021661_, _021723_);
  and g_113640_(_021721_, _021723_, _021725_);
  or g_113641_(_021720_, _021722_, _021726_);
  and g_113642_(_021719_, _021726_, _021727_);
  or g_113643_(_021718_, _021725_, _021728_);
  and g_113644_(_021700_, _021708_, _021729_);
  or g_113645_(_021701_, _021707_, _021730_);
  and g_113646_(_021728_, _021730_, _021731_);
  or g_113647_(_021727_, _021729_, _021732_);
  and g_113648_(_021718_, _021725_, _021733_);
  or g_113649_(_021719_, _021726_, _021734_);
  and g_113650_(_021731_, _021734_, _021736_);
  or g_113651_(_021732_, _021733_, _021737_);
  and g_113652_(_021716_, _021736_, _021738_);
  or g_113653_(_021717_, _021737_, _021739_);
  and g_113654_(_021639_, _021662_, _021740_);
  or g_113655_(_021640_, _021661_, _021741_);
  and g_113656_(_021641_, _021661_, _021742_);
  or g_113657_(_021642_, _021662_, _021743_);
  and g_113658_(_021741_, _021743_, _021744_);
  or g_113659_(_021740_, _021742_, _021745_);
  or g_113660_(out[520], _021671_, _021747_);
  and g_113661_(out[521], _021747_, _021748_);
  or g_113662_(out[522], _021748_, _021749_);
  xor g_113663_(out[522], _021748_, _021750_);
  xor g_113664_(_054732_, _021748_, _021751_);
  and g_113665_(_021744_, _021750_, _021752_);
  or g_113666_(_021745_, _021751_, _021753_);
  and g_113667_(_021528_, _021538_, _021754_);
  or g_113668_(_021529_, _021539_, _021755_);
  xor g_113669_(out[523], _021749_, _021756_);
  xor g_113670_(_054611_, _021749_, _021758_);
  and g_113671_(_021754_, _021758_, _021759_);
  or g_113672_(_021755_, _021756_, _021760_);
  and g_113673_(_021753_, _021760_, _021761_);
  or g_113674_(_021752_, _021759_, _021762_);
  and g_113675_(_021745_, _021751_, _021763_);
  or g_113676_(_021744_, _021750_, _021764_);
  and g_113677_(_021755_, _021756_, _021765_);
  or g_113678_(_021754_, _021758_, _021766_);
  and g_113679_(_021764_, _021766_, _021767_);
  or g_113680_(_021763_, _021765_, _021769_);
  and g_113681_(_021761_, _021767_, _021770_);
  or g_113682_(_021762_, _021769_, _021771_);
  xor g_113683_(out[520], _021671_, _021772_);
  xor g_113684_(_054710_, _021671_, _021773_);
  and g_113685_(_021552_, _021662_, _021774_);
  or g_113686_(_021551_, _021661_, _021775_);
  and g_113687_(_021550_, _021661_, _021776_);
  or g_113688_(_021549_, _021662_, _021777_);
  and g_113689_(_021775_, _021777_, _021778_);
  or g_113690_(_021774_, _021776_, _021780_);
  and g_113691_(_021772_, _021780_, _021781_);
  or g_113692_(_021773_, _021778_, _021782_);
  xor g_113693_(out[521], _021747_, _021783_);
  xor g_113694_(_054721_, _021747_, _021784_);
  and g_113695_(_021542_, _021662_, _021785_);
  or g_113696_(_021543_, _021661_, _021786_);
  and g_113697_(_021544_, _021661_, _021787_);
  or g_113698_(_021545_, _021662_, _021788_);
  and g_113699_(_021786_, _021788_, _021789_);
  or g_113700_(_021785_, _021787_, _021791_);
  and g_113701_(_021784_, _021791_, _021792_);
  or g_113702_(_021783_, _021789_, _021793_);
  and g_113703_(_021782_, _021793_, _021794_);
  or g_113704_(_021781_, _021792_, _021795_);
  and g_113705_(_021773_, _021778_, _021796_);
  or g_113706_(_021772_, _021780_, _021797_);
  and g_113707_(_021783_, _021789_, _021798_);
  or g_113708_(_021784_, _021791_, _021799_);
  and g_113709_(_021797_, _021799_, _021800_);
  or g_113710_(_021796_, _021798_, _021802_);
  and g_113711_(_021794_, _021800_, _021803_);
  or g_113712_(_021795_, _021802_, _021804_);
  and g_113713_(_021770_, _021803_, _021805_);
  or g_113714_(_021771_, _021804_, _021806_);
  or g_113715_(_054567_, _021662_, _021807_);
  or g_113716_(_054435_, _021661_, _021808_);
  and g_113717_(_021807_, _021808_, _021809_);
  and g_113718_(out[515], _021809_, _021810_);
  or g_113719_(out[482], _021661_, _021811_);
  or g_113720_(out[498], _021662_, _021813_);
  and g_113721_(_021811_, _021813_, _021814_);
  or g_113722_(out[515], _021809_, _021815_);
  and g_113723_(_054688_, _021814_, _021816_);
  xor g_113724_(_054699_, _021809_, _021817_);
  xor g_113725_(out[514], _021814_, _021818_);
  or g_113726_(_021817_, _021818_, _021819_);
  not g_113727_(_021819_, _021820_);
  and g_113728_(_054347_, _021662_, _021821_);
  or g_113729_(out[480], _021661_, _021822_);
  and g_113730_(_054545_, _021661_, _021824_);
  or g_113731_(out[496], _021662_, _021825_);
  and g_113732_(_021822_, _021825_, _021826_);
  or g_113733_(_021821_, _021824_, _021827_);
  and g_113734_(out[512], _021827_, _021828_);
  or g_113735_(_054677_, _021826_, _021829_);
  and g_113736_(_054666_, _021665_, _021830_);
  or g_113737_(out[513], _021666_, _021831_);
  xor g_113738_(_054666_, _021665_, _021832_);
  xor g_113739_(out[513], _021665_, _021833_);
  and g_113740_(_021829_, _021832_, _021835_);
  or g_113741_(_021828_, _021833_, _021836_);
  and g_113742_(_054677_, _021826_, _021837_);
  or g_113743_(out[512], _021827_, _021838_);
  and g_113744_(_021835_, _021838_, _021839_);
  or g_113745_(_021836_, _021837_, _021840_);
  and g_113746_(_021820_, _021839_, _021841_);
  or g_113747_(_021819_, _021840_, _021842_);
  and g_113748_(_021805_, _021841_, _021843_);
  or g_113749_(_021806_, _021842_, _021844_);
  and g_113750_(_021738_, _021843_, _021846_);
  or g_113751_(_021739_, _021844_, _021847_);
  and g_113752_(_021831_, _021836_, _021848_);
  or g_113753_(_021830_, _021835_, _021849_);
  and g_113754_(_021820_, _021849_, _021850_);
  or g_113755_(_021819_, _021848_, _021851_);
  or g_113756_(_021810_, _021816_, _021852_);
  and g_113757_(_021815_, _021852_, _021853_);
  not g_113758_(_021853_, _021854_);
  and g_113759_(_021851_, _021854_, _021855_);
  or g_113760_(_021850_, _021853_, _021857_);
  and g_113761_(_021738_, _021857_, _021858_);
  or g_113762_(_021739_, _021855_, _021859_);
  and g_113763_(_021716_, _021732_, _021860_);
  or g_113764_(_021717_, _021731_, _021861_);
  and g_113765_(_021695_, _021699_, _021862_);
  or g_113766_(_021694_, _021698_, _021863_);
  and g_113767_(_021861_, _021863_, _021864_);
  or g_113768_(_021860_, _021862_, _021865_);
  and g_113769_(_021859_, _021864_, _021866_);
  or g_113770_(_021858_, _021865_, _021868_);
  and g_113771_(_021805_, _021868_, _021869_);
  or g_113772_(_021806_, _021866_, _021870_);
  and g_113773_(_021795_, _021799_, _021871_);
  or g_113774_(_021794_, _021798_, _021872_);
  and g_113775_(_021770_, _021871_, _021873_);
  or g_113776_(_021771_, _021872_, _021874_);
  and g_113777_(_021762_, _021766_, _021875_);
  or g_113778_(_021761_, _021765_, _021876_);
  and g_113779_(_021874_, _021876_, _021877_);
  or g_113780_(_021873_, _021875_, _021879_);
  and g_113781_(_021870_, _021877_, _021880_);
  or g_113782_(_021869_, _021879_, _021881_);
  and g_113783_(_021847_, _021881_, _021882_);
  or g_113784_(_021846_, _021880_, _021883_);
  or g_113785_(_021665_, _021882_, _021884_);
  or g_113786_(out[513], _021883_, _021885_);
  and g_113787_(_021884_, _021885_, _021886_);
  not g_113788_(_021886_, _021887_);
  and g_113789_(out[532], out[531], _021888_);
  or g_113790_(out[533], _021888_, _021890_);
  or g_113791_(out[534], _021890_, _021891_);
  or g_113792_(out[535], _021891_, _021892_);
  or g_113793_(out[536], _021892_, _021893_);
  and g_113794_(out[537], _021893_, _021894_);
  or g_113795_(out[538], _021894_, _021895_);
  xor g_113796_(out[538], _021894_, _021896_);
  xor g_113797_(_054864_, _021894_, _021897_);
  and g_113798_(_021750_, _021882_, _021898_);
  or g_113799_(_021751_, _021883_, _021899_);
  and g_113800_(_021745_, _021883_, _021901_);
  or g_113801_(_021744_, _021882_, _021902_);
  and g_113802_(_021899_, _021902_, _021903_);
  or g_113803_(_021898_, _021901_, _021904_);
  and g_113804_(_021896_, _021903_, _021905_);
  or g_113805_(_021897_, _021904_, _021906_);
  and g_113806_(_021754_, _021756_, _021907_);
  or g_113807_(_021755_, _021758_, _021908_);
  xor g_113808_(out[539], _021895_, _021909_);
  xor g_113809_(_054743_, _021895_, _021910_);
  and g_113810_(_021907_, _021910_, _021912_);
  or g_113811_(_021908_, _021909_, _021913_);
  and g_113812_(_021906_, _021913_, _021914_);
  or g_113813_(_021905_, _021912_, _021915_);
  and g_113814_(_021897_, _021904_, _021916_);
  or g_113815_(_021896_, _021903_, _021917_);
  and g_113816_(_021908_, _021909_, _021918_);
  or g_113817_(_021907_, _021910_, _021919_);
  xor g_113818_(out[537], _021893_, _021920_);
  xor g_113819_(_054853_, _021893_, _021921_);
  and g_113820_(_021783_, _021882_, _021923_);
  or g_113821_(_021784_, _021883_, _021924_);
  and g_113822_(_021791_, _021883_, _021925_);
  or g_113823_(_021789_, _021882_, _021926_);
  and g_113824_(_021924_, _021926_, _021927_);
  or g_113825_(_021923_, _021925_, _021928_);
  and g_113826_(_021920_, _021927_, _021929_);
  or g_113827_(_021921_, _021928_, _021930_);
  xor g_113828_(out[536], _021892_, _021931_);
  xor g_113829_(_054842_, _021892_, _021932_);
  and g_113830_(_021773_, _021882_, _021934_);
  or g_113831_(_021772_, _021883_, _021935_);
  and g_113832_(_021780_, _021883_, _021936_);
  or g_113833_(_021778_, _021882_, _021937_);
  and g_113834_(_021935_, _021937_, _021938_);
  or g_113835_(_021934_, _021936_, _021939_);
  and g_113836_(_021931_, _021939_, _021940_);
  or g_113837_(_021932_, _021938_, _021941_);
  and g_113838_(_021921_, _021928_, _021942_);
  or g_113839_(_021920_, _021927_, _021943_);
  and g_113840_(_021941_, _021943_, _021945_);
  or g_113841_(_021940_, _021942_, _021946_);
  and g_113842_(_021932_, _021938_, _021947_);
  or g_113843_(_021931_, _021939_, _021948_);
  and g_113844_(_021917_, _021919_, _021949_);
  or g_113845_(_021916_, _021918_, _021950_);
  and g_113846_(_021914_, _021949_, _021951_);
  or g_113847_(_021915_, _021950_, _021952_);
  and g_113848_(_021930_, _021948_, _021953_);
  or g_113849_(_021929_, _021947_, _021954_);
  and g_113850_(_021945_, _021953_, _021956_);
  or g_113851_(_021946_, _021954_, _021957_);
  and g_113852_(_021951_, _021956_, _021958_);
  or g_113853_(_021952_, _021957_, _021959_);
  xor g_113854_(out[534], _021890_, _021960_);
  xor g_113855_(_054765_, _021890_, _021961_);
  and g_113856_(_021683_, _021882_, _021962_);
  or g_113857_(_021684_, _021883_, _021963_);
  and g_113858_(_021690_, _021883_, _021964_);
  or g_113859_(_021689_, _021882_, _021965_);
  and g_113860_(_021963_, _021965_, _021967_);
  or g_113861_(_021962_, _021964_, _021968_);
  and g_113862_(_021960_, _021967_, _021969_);
  or g_113863_(_021961_, _021968_, _021970_);
  xor g_113864_(out[535], _021891_, _021971_);
  xor g_113865_(_054754_, _021891_, _021972_);
  and g_113866_(_021673_, _021882_, _021973_);
  or g_113867_(_021672_, _021883_, _021974_);
  and g_113868_(_021679_, _021883_, _021975_);
  or g_113869_(_021678_, _021882_, _021976_);
  and g_113870_(_021974_, _021976_, _021978_);
  or g_113871_(_021973_, _021975_, _021979_);
  and g_113872_(_021971_, _021979_, _021980_);
  or g_113873_(_021972_, _021978_, _021981_);
  and g_113874_(_021970_, _021981_, _021982_);
  or g_113875_(_021969_, _021980_, _021983_);
  and g_113876_(_021972_, _021978_, _021984_);
  or g_113877_(_021971_, _021979_, _021985_);
  and g_113878_(_021961_, _021968_, _021986_);
  or g_113879_(_021960_, _021967_, _021987_);
  and g_113880_(_021985_, _021987_, _021989_);
  or g_113881_(_021984_, _021986_, _021990_);
  and g_113882_(_021982_, _021989_, _021991_);
  or g_113883_(_021983_, _021990_, _021992_);
  xor g_113884_(out[533], _021888_, _021993_);
  xor g_113885_(_054776_, _021888_, _021994_);
  and g_113886_(_021701_, _021882_, _021995_);
  or g_113887_(_021700_, _021883_, _021996_);
  and g_113888_(_021708_, _021883_, _021997_);
  or g_113889_(_021707_, _021882_, _021998_);
  and g_113890_(_021996_, _021998_, _022000_);
  or g_113891_(_021995_, _021997_, _022001_);
  and g_113892_(_021993_, _022001_, _022002_);
  or g_113893_(_021994_, _022000_, _022003_);
  xor g_113894_(out[532], out[531], _022004_);
  xor g_113895_(_054787_, out[531], _022005_);
  and g_113896_(_021718_, _021882_, _022006_);
  or g_113897_(_021719_, _021883_, _022007_);
  and g_113898_(_021726_, _021883_, _022008_);
  or g_113899_(_021725_, _021882_, _022009_);
  and g_113900_(_022007_, _022009_, _022011_);
  or g_113901_(_022006_, _022008_, _022012_);
  and g_113902_(_022005_, _022012_, _022013_);
  or g_113903_(_022004_, _022011_, _022014_);
  and g_113904_(_022003_, _022014_, _022015_);
  or g_113905_(_022002_, _022013_, _022016_);
  and g_113906_(_022004_, _022011_, _022017_);
  or g_113907_(_022005_, _022012_, _022018_);
  and g_113908_(_021994_, _022000_, _022019_);
  or g_113909_(_021993_, _022001_, _022020_);
  and g_113910_(_022018_, _022020_, _022022_);
  or g_113911_(_022017_, _022019_, _022023_);
  and g_113912_(_022015_, _022022_, _022024_);
  or g_113913_(_022016_, _022023_, _022025_);
  and g_113914_(_021991_, _022024_, _022026_);
  or g_113915_(_021992_, _022025_, _022027_);
  or g_113916_(_054699_, _021883_, _022028_);
  or g_113917_(_021809_, _021882_, _022029_);
  and g_113918_(_022028_, _022029_, _022030_);
  and g_113919_(out[531], _022030_, _022031_);
  or g_113920_(_021814_, _021882_, _022033_);
  or g_113921_(out[514], _021883_, _022034_);
  and g_113922_(_022033_, _022034_, _022035_);
  or g_113923_(out[531], _022030_, _022036_);
  and g_113924_(_054820_, _022035_, _022037_);
  xor g_113925_(_054831_, _022030_, _022038_);
  xor g_113926_(out[530], _022035_, _022039_);
  or g_113927_(_022038_, _022039_, _022040_);
  not g_113928_(_022040_, _022041_);
  and g_113929_(_054798_, _021886_, _022042_);
  or g_113930_(out[529], _021887_, _022044_);
  and g_113931_(_021827_, _021883_, _022045_);
  or g_113932_(_021826_, _021882_, _022046_);
  and g_113933_(_054677_, _021882_, _022047_);
  or g_113934_(out[512], _021883_, _022048_);
  and g_113935_(_022046_, _022048_, _022049_);
  or g_113936_(_022045_, _022047_, _022050_);
  and g_113937_(out[528], _022050_, _022051_);
  or g_113938_(_054809_, _022049_, _022052_);
  xor g_113939_(_054798_, _021886_, _022053_);
  xor g_113940_(out[529], _021886_, _022055_);
  and g_113941_(_022052_, _022053_, _022056_);
  or g_113942_(_022051_, _022055_, _022057_);
  and g_113943_(_022044_, _022057_, _022058_);
  or g_113944_(_022042_, _022056_, _022059_);
  and g_113945_(_022041_, _022059_, _022060_);
  or g_113946_(_022040_, _022058_, _022061_);
  and g_113947_(_022036_, _022037_, _022062_);
  or g_113948_(_022031_, _022062_, _022063_);
  not g_113949_(_022063_, _022064_);
  and g_113950_(_022061_, _022064_, _022066_);
  or g_113951_(_022060_, _022063_, _022067_);
  and g_113952_(_022026_, _022067_, _022068_);
  or g_113953_(_022027_, _022066_, _022069_);
  and g_113954_(_021983_, _021985_, _022070_);
  or g_113955_(_021982_, _021984_, _022071_);
  and g_113956_(_022016_, _022020_, _022072_);
  or g_113957_(_022015_, _022019_, _022073_);
  and g_113958_(_021991_, _022072_, _022074_);
  or g_113959_(_021992_, _022073_, _022075_);
  and g_113960_(_022071_, _022075_, _022077_);
  or g_113961_(_022070_, _022074_, _022078_);
  and g_113962_(_022069_, _022077_, _022079_);
  or g_113963_(_022068_, _022078_, _022080_);
  and g_113964_(_021958_, _022080_, _022081_);
  or g_113965_(_021959_, _022079_, _022082_);
  and g_113966_(_021915_, _021919_, _022083_);
  or g_113967_(_021914_, _021918_, _022084_);
  and g_113968_(_021930_, _021946_, _022085_);
  or g_113969_(_021929_, _021945_, _022086_);
  and g_113970_(_021951_, _022085_, _022088_);
  or g_113971_(_021952_, _022086_, _022089_);
  and g_113972_(_022084_, _022089_, _022090_);
  or g_113973_(_022083_, _022088_, _022091_);
  and g_113974_(_022082_, _022090_, _022092_);
  or g_113975_(_022081_, _022091_, _022093_);
  and g_113976_(_054809_, _022049_, _022094_);
  or g_113977_(out[528], _022050_, _022095_);
  or g_113978_(_022040_, _022057_, _022096_);
  not g_113979_(_022096_, _022097_);
  and g_113980_(_022095_, _022097_, _022099_);
  or g_113981_(_022094_, _022096_, _022100_);
  and g_113982_(_022026_, _022099_, _022101_);
  or g_113983_(_022027_, _022100_, _022102_);
  and g_113984_(_021958_, _022101_, _022103_);
  or g_113985_(_021959_, _022102_, _022104_);
  and g_113986_(_022093_, _022104_, _022105_);
  or g_113987_(_022092_, _022103_, _022106_);
  or g_113988_(_021886_, _022105_, _022107_);
  or g_113989_(out[529], _022106_, _022108_);
  and g_113990_(_022107_, _022108_, _022110_);
  not g_113991_(_022110_, _022111_);
  and g_113992_(_021907_, _021909_, _022112_);
  or g_113993_(_021908_, _021910_, _022113_);
  and g_113994_(out[548], out[547], _022114_);
  or g_113995_(out[549], _022114_, _022115_);
  or g_113996_(out[550], _022115_, _022116_);
  or g_113997_(out[551], _022116_, _022117_);
  or g_113998_(out[552], _022117_, _022118_);
  and g_113999_(out[553], _022118_, _022119_);
  or g_114000_(out[554], _022119_, _022121_);
  xor g_114001_(out[555], _022121_, _022122_);
  xor g_114002_(_054875_, _022121_, _022123_);
  and g_114003_(_022112_, _022123_, _022124_);
  or g_114004_(_022113_, _022122_, _022125_);
  and g_114005_(_022113_, _022122_, _022126_);
  or g_114006_(_022112_, _022123_, _022127_);
  xor g_114007_(out[554], _022119_, _022128_);
  not g_114008_(_022128_, _022129_);
  and g_114009_(_021904_, _022106_, _022130_);
  or g_114010_(_021903_, _022105_, _022132_);
  and g_114011_(_021896_, _022105_, _022133_);
  or g_114012_(_021897_, _022106_, _022134_);
  and g_114013_(_022132_, _022134_, _022135_);
  or g_114014_(_022130_, _022133_, _022136_);
  and g_114015_(_022129_, _022136_, _022137_);
  or g_114016_(_022128_, _022135_, _022138_);
  and g_114017_(_022128_, _022135_, _022139_);
  or g_114018_(_022129_, _022136_, _022140_);
  xor g_114019_(out[553], _022118_, _022141_);
  xor g_114020_(_054985_, _022118_, _022143_);
  and g_114021_(_021928_, _022106_, _022144_);
  or g_114022_(_021927_, _022105_, _022145_);
  and g_114023_(_021920_, _022105_, _022146_);
  or g_114024_(_021921_, _022106_, _022147_);
  and g_114025_(_022145_, _022147_, _022148_);
  or g_114026_(_022144_, _022146_, _022149_);
  and g_114027_(_022141_, _022148_, _022150_);
  or g_114028_(_022143_, _022149_, _022151_);
  xor g_114029_(out[552], _022117_, _022152_);
  xor g_114030_(_054974_, _022117_, _022154_);
  and g_114031_(_021939_, _022106_, _022155_);
  or g_114032_(_021938_, _022105_, _022156_);
  and g_114033_(_021932_, _022105_, _022157_);
  or g_114034_(_021931_, _022106_, _022158_);
  and g_114035_(_022156_, _022158_, _022159_);
  or g_114036_(_022155_, _022157_, _022160_);
  and g_114037_(_022152_, _022160_, _022161_);
  or g_114038_(_022154_, _022159_, _022162_);
  and g_114039_(_022143_, _022149_, _022163_);
  or g_114040_(_022141_, _022148_, _022165_);
  and g_114041_(_022162_, _022165_, _022166_);
  or g_114042_(_022161_, _022163_, _022167_);
  and g_114043_(_022154_, _022159_, _022168_);
  or g_114044_(_022152_, _022160_, _022169_);
  and g_114045_(_022125_, _022138_, _022170_);
  or g_114046_(_022124_, _022137_, _022171_);
  and g_114047_(_022127_, _022140_, _022172_);
  or g_114048_(_022126_, _022139_, _022173_);
  and g_114049_(_022170_, _022172_, _022174_);
  or g_114050_(_022171_, _022173_, _022176_);
  and g_114051_(_022151_, _022169_, _022177_);
  or g_114052_(_022150_, _022168_, _022178_);
  and g_114053_(_022166_, _022177_, _022179_);
  or g_114054_(_022167_, _022178_, _022180_);
  and g_114055_(_022174_, _022179_, _022181_);
  or g_114056_(_022176_, _022180_, _022182_);
  xor g_114057_(out[550], _022115_, _022183_);
  xor g_114058_(_054897_, _022115_, _022184_);
  and g_114059_(_021968_, _022106_, _022185_);
  or g_114060_(_021967_, _022105_, _022187_);
  and g_114061_(_021960_, _022105_, _022188_);
  or g_114062_(_021961_, _022106_, _022189_);
  and g_114063_(_022187_, _022189_, _022190_);
  or g_114064_(_022185_, _022188_, _022191_);
  and g_114065_(_022183_, _022190_, _022192_);
  or g_114066_(_022184_, _022191_, _022193_);
  xor g_114067_(out[551], _022116_, _022194_);
  xor g_114068_(_054886_, _022116_, _022195_);
  and g_114069_(_021979_, _022106_, _022196_);
  or g_114070_(_021978_, _022105_, _022198_);
  and g_114071_(_021972_, _022105_, _022199_);
  or g_114072_(_021971_, _022106_, _022200_);
  and g_114073_(_022198_, _022200_, _022201_);
  or g_114074_(_022196_, _022199_, _022202_);
  and g_114075_(_022194_, _022202_, _022203_);
  or g_114076_(_022195_, _022201_, _022204_);
  and g_114077_(_022193_, _022204_, _022205_);
  or g_114078_(_022192_, _022203_, _022206_);
  and g_114079_(_022184_, _022191_, _022207_);
  or g_114080_(_022183_, _022190_, _022209_);
  and g_114081_(_022195_, _022201_, _022210_);
  or g_114082_(_022194_, _022202_, _022211_);
  xor g_114083_(out[549], _022114_, _022212_);
  xor g_114084_(_054908_, _022114_, _022213_);
  and g_114085_(_022001_, _022106_, _022214_);
  or g_114086_(_022000_, _022105_, _022215_);
  and g_114087_(_021994_, _022105_, _022216_);
  or g_114088_(_021993_, _022106_, _022217_);
  and g_114089_(_022215_, _022217_, _022218_);
  or g_114090_(_022214_, _022216_, _022220_);
  and g_114091_(_022213_, _022218_, _022221_);
  or g_114092_(_022212_, _022220_, _022222_);
  and g_114093_(_022211_, _022222_, _022223_);
  or g_114094_(_022210_, _022221_, _022224_);
  and g_114095_(_022209_, _022223_, _022225_);
  or g_114096_(_022207_, _022224_, _022226_);
  and g_114097_(_022205_, _022225_, _022227_);
  or g_114098_(_022206_, _022226_, _022228_);
  xor g_114099_(out[548], out[547], _022229_);
  xor g_114100_(_054919_, out[547], _022231_);
  and g_114101_(_022004_, _022105_, _022232_);
  or g_114102_(_022005_, _022106_, _022233_);
  and g_114103_(_022012_, _022106_, _022234_);
  or g_114104_(_022011_, _022105_, _022235_);
  and g_114105_(_022233_, _022235_, _022236_);
  or g_114106_(_022232_, _022234_, _022237_);
  and g_114107_(_022231_, _022237_, _022238_);
  or g_114108_(_022229_, _022236_, _022239_);
  and g_114109_(_022212_, _022220_, _022240_);
  or g_114110_(_022213_, _022218_, _022242_);
  and g_114111_(_022239_, _022242_, _022243_);
  or g_114112_(_022238_, _022240_, _022244_);
  and g_114113_(_022229_, _022236_, _022245_);
  or g_114114_(_022231_, _022237_, _022246_);
  and g_114115_(_022243_, _022246_, _022247_);
  or g_114116_(_022244_, _022245_, _022248_);
  and g_114117_(_022227_, _022247_, _022249_);
  or g_114118_(_022228_, _022248_, _022250_);
  or g_114119_(_054831_, _022106_, _022251_);
  or g_114120_(_022030_, _022105_, _022253_);
  and g_114121_(_022251_, _022253_, _022254_);
  and g_114122_(out[547], _022254_, _022255_);
  or g_114123_(_022035_, _022105_, _022256_);
  or g_114124_(out[530], _022106_, _022257_);
  and g_114125_(_022256_, _022257_, _022258_);
  or g_114126_(out[547], _022254_, _022259_);
  and g_114127_(_054952_, _022258_, _022260_);
  xor g_114128_(out[547], _022254_, _022261_);
  xor g_114129_(_054963_, _022254_, _022262_);
  xor g_114130_(_054952_, _022258_, _022264_);
  xor g_114131_(out[546], _022258_, _022265_);
  and g_114132_(_022261_, _022264_, _022266_);
  or g_114133_(_022262_, _022265_, _022267_);
  and g_114134_(_054930_, _022110_, _022268_);
  or g_114135_(out[545], _022111_, _022269_);
  and g_114136_(_022050_, _022106_, _022270_);
  or g_114137_(_022049_, _022105_, _022271_);
  and g_114138_(_054809_, _022105_, _022272_);
  or g_114139_(out[528], _022106_, _022273_);
  and g_114140_(_022271_, _022273_, _022275_);
  or g_114141_(_022270_, _022272_, _022276_);
  and g_114142_(out[544], _022276_, _022277_);
  or g_114143_(_054941_, _022275_, _022278_);
  xor g_114144_(_054930_, _022110_, _022279_);
  xor g_114145_(out[545], _022110_, _022280_);
  and g_114146_(_022278_, _022279_, _022281_);
  or g_114147_(_022277_, _022280_, _022282_);
  and g_114148_(_022269_, _022282_, _022283_);
  or g_114149_(_022268_, _022281_, _022284_);
  and g_114150_(_022266_, _022284_, _022286_);
  or g_114151_(_022267_, _022283_, _022287_);
  and g_114152_(_022259_, _022260_, _022288_);
  or g_114153_(_022255_, _022288_, _022289_);
  not g_114154_(_022289_, _022290_);
  and g_114155_(_022287_, _022290_, _022291_);
  or g_114156_(_022286_, _022289_, _022292_);
  and g_114157_(_022249_, _022292_, _022293_);
  or g_114158_(_022250_, _022291_, _022294_);
  and g_114159_(_022227_, _022244_, _022295_);
  or g_114160_(_022228_, _022243_, _022297_);
  and g_114161_(_022206_, _022211_, _022298_);
  or g_114162_(_022205_, _022210_, _022299_);
  and g_114163_(_022297_, _022299_, _022300_);
  or g_114164_(_022295_, _022298_, _022301_);
  and g_114165_(_022294_, _022300_, _022302_);
  or g_114166_(_022293_, _022301_, _022303_);
  and g_114167_(_022181_, _022303_, _022304_);
  or g_114168_(_022182_, _022302_, _022305_);
  and g_114169_(_022151_, _022167_, _022306_);
  or g_114170_(_022150_, _022166_, _022308_);
  and g_114171_(_022174_, _022306_, _022309_);
  or g_114172_(_022176_, _022308_, _022310_);
  and g_114173_(_022127_, _022139_, _022311_);
  or g_114174_(_022126_, _022140_, _022312_);
  and g_114175_(_022125_, _022312_, _022313_);
  or g_114176_(_022124_, _022311_, _022314_);
  and g_114177_(_022310_, _022313_, _022315_);
  or g_114178_(_022309_, _022314_, _022316_);
  and g_114179_(_022305_, _022315_, _022317_);
  or g_114180_(_022304_, _022316_, _022319_);
  and g_114181_(_054941_, _022275_, _022320_);
  or g_114182_(out[544], _022276_, _022321_);
  and g_114183_(_022266_, _022321_, _022322_);
  or g_114184_(_022267_, _022320_, _022323_);
  and g_114185_(_022281_, _022322_, _022324_);
  or g_114186_(_022282_, _022323_, _022325_);
  and g_114187_(_022181_, _022324_, _022326_);
  or g_114188_(_022182_, _022325_, _022327_);
  and g_114189_(_022249_, _022326_, _022328_);
  or g_114190_(_022250_, _022327_, _022330_);
  and g_114191_(_022319_, _022330_, _022331_);
  or g_114192_(_022317_, _022328_, _022332_);
  or g_114193_(_022110_, _022331_, _022333_);
  or g_114194_(out[545], _022332_, _022334_);
  and g_114195_(_022333_, _022334_, _022335_);
  not g_114196_(_022335_, _022336_);
  and g_114197_(_022128_, _022331_, _022337_);
  or g_114198_(_022129_, _022332_, _022338_);
  and g_114199_(_022136_, _022332_, _022339_);
  or g_114200_(_022135_, _022331_, _022341_);
  and g_114201_(_022338_, _022341_, _022342_);
  or g_114202_(_022337_, _022339_, _022343_);
  and g_114203_(out[564], out[563], _022344_);
  or g_114204_(out[565], _022344_, _022345_);
  or g_114205_(out[566], _022345_, _022346_);
  or g_114206_(out[567], _022346_, _022347_);
  or g_114207_(out[568], _022347_, _022348_);
  and g_114208_(out[569], _022348_, _022349_);
  or g_114209_(out[570], _022349_, _022350_);
  xor g_114210_(out[570], _022349_, _022352_);
  xor g_114211_(_055128_, _022349_, _022353_);
  and g_114212_(_022342_, _022352_, _022354_);
  or g_114213_(_022343_, _022353_, _022355_);
  and g_114214_(_022112_, _022122_, _022356_);
  or g_114215_(_022113_, _022123_, _022357_);
  xor g_114216_(out[571], _022350_, _022358_);
  xor g_114217_(_055007_, _022350_, _022359_);
  and g_114218_(_022356_, _022359_, _022360_);
  or g_114219_(_022357_, _022358_, _022361_);
  and g_114220_(_022355_, _022361_, _022363_);
  or g_114221_(_022354_, _022360_, _022364_);
  and g_114222_(_022343_, _022353_, _022365_);
  or g_114223_(_022342_, _022352_, _022366_);
  and g_114224_(_022357_, _022358_, _022367_);
  or g_114225_(_022356_, _022359_, _022368_);
  xor g_114226_(out[569], _022348_, _022369_);
  xor g_114227_(_055117_, _022348_, _022370_);
  and g_114228_(_022141_, _022331_, _022371_);
  or g_114229_(_022143_, _022332_, _022372_);
  and g_114230_(_022149_, _022332_, _022374_);
  or g_114231_(_022148_, _022331_, _022375_);
  and g_114232_(_022372_, _022375_, _022376_);
  or g_114233_(_022371_, _022374_, _022377_);
  and g_114234_(_022369_, _022376_, _022378_);
  or g_114235_(_022370_, _022377_, _022379_);
  and g_114236_(_022366_, _022368_, _022380_);
  or g_114237_(_022365_, _022367_, _022381_);
  and g_114238_(_022363_, _022380_, _022382_);
  or g_114239_(_022364_, _022381_, _022383_);
  and g_114240_(_022379_, _022382_, _022385_);
  or g_114241_(_022378_, _022383_, _022386_);
  and g_114242_(_022370_, _022377_, _022387_);
  or g_114243_(_022369_, _022376_, _022388_);
  xor g_114244_(out[568], _022347_, _022389_);
  xor g_114245_(_055106_, _022347_, _022390_);
  and g_114246_(_022154_, _022331_, _022391_);
  or g_114247_(_022152_, _022332_, _022392_);
  and g_114248_(_022160_, _022332_, _022393_);
  or g_114249_(_022159_, _022331_, _022394_);
  and g_114250_(_022392_, _022394_, _022396_);
  or g_114251_(_022391_, _022393_, _022397_);
  and g_114252_(_022389_, _022397_, _022398_);
  or g_114253_(_022390_, _022396_, _022399_);
  and g_114254_(_022388_, _022399_, _022400_);
  or g_114255_(_022387_, _022398_, _022401_);
  and g_114256_(_022390_, _022396_, _022402_);
  or g_114257_(_022389_, _022397_, _022403_);
  and g_114258_(_022400_, _022403_, _022404_);
  or g_114259_(_022401_, _022402_, _022405_);
  and g_114260_(_022385_, _022404_, _022407_);
  or g_114261_(_022386_, _022405_, _022408_);
  xor g_114262_(out[567], _022346_, _022409_);
  xor g_114263_(_055018_, _022346_, _022410_);
  and g_114264_(_022195_, _022331_, _022411_);
  or g_114265_(_022194_, _022332_, _022412_);
  and g_114266_(_022202_, _022332_, _022413_);
  or g_114267_(_022201_, _022331_, _022414_);
  and g_114268_(_022412_, _022414_, _022415_);
  or g_114269_(_022411_, _022413_, _022416_);
  and g_114270_(_022409_, _022416_, _022418_);
  or g_114271_(_022410_, _022415_, _022419_);
  xor g_114272_(out[566], _022345_, _022420_);
  xor g_114273_(_055029_, _022345_, _022421_);
  and g_114274_(_022183_, _022331_, _022422_);
  or g_114275_(_022184_, _022332_, _022423_);
  and g_114276_(_022191_, _022332_, _022424_);
  or g_114277_(_022190_, _022331_, _022425_);
  and g_114278_(_022423_, _022425_, _022426_);
  or g_114279_(_022422_, _022424_, _022427_);
  and g_114280_(_022420_, _022426_, _022429_);
  or g_114281_(_022421_, _022427_, _022430_);
  and g_114282_(_022419_, _022430_, _022431_);
  or g_114283_(_022418_, _022429_, _022432_);
  and g_114284_(_022410_, _022415_, _022433_);
  or g_114285_(_022409_, _022416_, _022434_);
  and g_114286_(_022421_, _022427_, _022435_);
  or g_114287_(_022420_, _022426_, _022436_);
  and g_114288_(_022434_, _022436_, _022437_);
  or g_114289_(_022433_, _022435_, _022438_);
  and g_114290_(_022431_, _022437_, _022440_);
  or g_114291_(_022432_, _022438_, _022441_);
  xor g_114292_(out[565], _022344_, _022442_);
  xor g_114293_(_055040_, _022344_, _022443_);
  and g_114294_(_022213_, _022331_, _022444_);
  or g_114295_(_022212_, _022332_, _022445_);
  and g_114296_(_022220_, _022332_, _022446_);
  or g_114297_(_022218_, _022331_, _022447_);
  and g_114298_(_022445_, _022447_, _022448_);
  or g_114299_(_022444_, _022446_, _022449_);
  and g_114300_(_022442_, _022449_, _022451_);
  or g_114301_(_022443_, _022448_, _022452_);
  xor g_114302_(out[564], out[563], _022453_);
  xor g_114303_(_055051_, out[563], _022454_);
  and g_114304_(_022229_, _022331_, _022455_);
  or g_114305_(_022231_, _022332_, _022456_);
  and g_114306_(_022237_, _022332_, _022457_);
  or g_114307_(_022236_, _022331_, _022458_);
  and g_114308_(_022456_, _022458_, _022459_);
  or g_114309_(_022455_, _022457_, _022460_);
  and g_114310_(_022454_, _022460_, _022462_);
  or g_114311_(_022453_, _022459_, _022463_);
  and g_114312_(_022452_, _022463_, _022464_);
  or g_114313_(_022451_, _022462_, _022465_);
  and g_114314_(_022453_, _022459_, _022466_);
  or g_114315_(_022454_, _022460_, _022467_);
  and g_114316_(_022443_, _022448_, _022468_);
  or g_114317_(_022442_, _022449_, _022469_);
  and g_114318_(_022467_, _022469_, _022470_);
  or g_114319_(_022466_, _022468_, _022471_);
  and g_114320_(_022464_, _022470_, _022473_);
  or g_114321_(_022465_, _022471_, _022474_);
  and g_114322_(_022440_, _022473_, _022475_);
  or g_114323_(_022441_, _022474_, _022476_);
  and g_114324_(_022407_, _022475_, _022477_);
  or g_114325_(_022408_, _022476_, _022478_);
  or g_114326_(_054963_, _022332_, _022479_);
  or g_114327_(_022254_, _022331_, _022480_);
  and g_114328_(_022479_, _022480_, _022481_);
  not g_114329_(_022481_, _022482_);
  and g_114330_(out[563], _022481_, _022484_);
  or g_114331_(_022258_, _022331_, _022485_);
  or g_114332_(out[546], _022332_, _022486_);
  and g_114333_(_022485_, _022486_, _022487_);
  or g_114334_(out[563], _022481_, _022488_);
  and g_114335_(_055084_, _022487_, _022489_);
  xor g_114336_(out[563], _022481_, _022490_);
  xor g_114337_(_055095_, _022481_, _022491_);
  xor g_114338_(_055084_, _022487_, _022492_);
  xor g_114339_(out[562], _022487_, _022493_);
  and g_114340_(_022490_, _022492_, _022495_);
  or g_114341_(_022491_, _022493_, _022496_);
  and g_114342_(_022276_, _022332_, _022497_);
  or g_114343_(_022275_, _022331_, _022498_);
  and g_114344_(_054941_, _022331_, _022499_);
  or g_114345_(out[544], _022332_, _022500_);
  and g_114346_(_022498_, _022500_, _022501_);
  or g_114347_(_022497_, _022499_, _022502_);
  and g_114348_(out[560], _022502_, _022503_);
  or g_114349_(_055073_, _022501_, _022504_);
  and g_114350_(_055062_, _022335_, _022506_);
  or g_114351_(out[561], _022336_, _022507_);
  xor g_114352_(_055062_, _022335_, _022508_);
  xor g_114353_(out[561], _022335_, _022509_);
  and g_114354_(_022504_, _022508_, _022510_);
  or g_114355_(_022503_, _022509_, _022511_);
  and g_114356_(_055073_, _022501_, _022512_);
  or g_114357_(out[560], _022502_, _022513_);
  and g_114358_(_022510_, _022513_, _022514_);
  or g_114359_(_022511_, _022512_, _022515_);
  and g_114360_(_022495_, _022514_, _022517_);
  or g_114361_(_022496_, _022515_, _022518_);
  and g_114362_(_022477_, _022517_, _022519_);
  or g_114363_(_022478_, _022518_, _022520_);
  and g_114364_(_022507_, _022511_, _022521_);
  or g_114365_(_022506_, _022510_, _022522_);
  and g_114366_(_022495_, _022522_, _022523_);
  or g_114367_(_022496_, _022521_, _022524_);
  and g_114368_(_022488_, _022489_, _022525_);
  or g_114369_(_022484_, _022525_, _022526_);
  not g_114370_(_022526_, _022528_);
  and g_114371_(_022524_, _022528_, _022529_);
  or g_114372_(_022523_, _022526_, _022530_);
  and g_114373_(_022477_, _022530_, _022531_);
  or g_114374_(_022478_, _022529_, _022532_);
  and g_114375_(_022432_, _022434_, _022533_);
  or g_114376_(_022431_, _022433_, _022534_);
  and g_114377_(_022465_, _022469_, _022535_);
  or g_114378_(_022464_, _022468_, _022536_);
  and g_114379_(_022440_, _022535_, _022537_);
  or g_114380_(_022441_, _022536_, _022539_);
  and g_114381_(_022534_, _022539_, _022540_);
  or g_114382_(_022533_, _022537_, _022541_);
  and g_114383_(_022407_, _022541_, _022542_);
  or g_114384_(_022408_, _022540_, _022543_);
  and g_114385_(_022385_, _022401_, _022544_);
  or g_114386_(_022386_, _022400_, _022545_);
  and g_114387_(_022364_, _022368_, _022546_);
  or g_114388_(_022363_, _022367_, _022547_);
  and g_114389_(_022545_, _022547_, _022548_);
  or g_114390_(_022544_, _022546_, _022550_);
  and g_114391_(_022543_, _022548_, _022551_);
  or g_114392_(_022542_, _022550_, _022552_);
  and g_114393_(_022532_, _022551_, _022553_);
  or g_114394_(_022531_, _022552_, _022554_);
  and g_114395_(_022520_, _022554_, _022555_);
  or g_114396_(_022519_, _022553_, _022556_);
  or g_114397_(_022335_, _022555_, _022557_);
  or g_114398_(out[561], _022556_, _022558_);
  and g_114399_(_022557_, _022558_, _022559_);
  not g_114400_(_022559_, _022561_);
  and g_114401_(_022356_, _022358_, _022562_);
  or g_114402_(_022357_, _022359_, _022563_);
  and g_114403_(out[580], out[579], _022564_);
  or g_114404_(out[581], _022564_, _022565_);
  or g_114405_(out[582], _022565_, _022566_);
  or g_114406_(out[583], _022566_, _022567_);
  or g_114407_(out[584], _022567_, _022568_);
  and g_114408_(out[585], _022568_, _022569_);
  or g_114409_(out[586], _022569_, _022570_);
  xor g_114410_(out[587], _022570_, _022572_);
  xor g_114411_(_055139_, _022570_, _022573_);
  and g_114412_(_022562_, _022573_, _022574_);
  or g_114413_(_022563_, _022572_, _022575_);
  and g_114414_(_022352_, _022555_, _022576_);
  or g_114415_(_022353_, _022556_, _022577_);
  and g_114416_(_022343_, _022556_, _022578_);
  or g_114417_(_022342_, _022555_, _022579_);
  and g_114418_(_022577_, _022579_, _022580_);
  or g_114419_(_022576_, _022578_, _022581_);
  xor g_114420_(out[586], _022569_, _022583_);
  xor g_114421_(_055260_, _022569_, _022584_);
  and g_114422_(_022580_, _022583_, _022585_);
  or g_114423_(_022581_, _022584_, _022586_);
  and g_114424_(_022575_, _022586_, _022587_);
  or g_114425_(_022574_, _022585_, _022588_);
  and g_114426_(_022581_, _022584_, _022589_);
  or g_114427_(_022580_, _022583_, _022590_);
  and g_114428_(_022563_, _022572_, _022591_);
  or g_114429_(_022562_, _022573_, _022592_);
  xor g_114430_(out[585], _022568_, _022594_);
  xor g_114431_(_055249_, _022568_, _022595_);
  and g_114432_(_022369_, _022555_, _022596_);
  or g_114433_(_022370_, _022556_, _022597_);
  and g_114434_(_022377_, _022556_, _022598_);
  or g_114435_(_022376_, _022555_, _022599_);
  and g_114436_(_022597_, _022599_, _022600_);
  or g_114437_(_022596_, _022598_, _022601_);
  and g_114438_(_022594_, _022600_, _022602_);
  or g_114439_(_022595_, _022601_, _022603_);
  xor g_114440_(out[584], _022567_, _022605_);
  xor g_114441_(_055238_, _022567_, _022606_);
  and g_114442_(_022390_, _022555_, _022607_);
  or g_114443_(_022389_, _022556_, _022608_);
  and g_114444_(_022397_, _022556_, _022609_);
  or g_114445_(_022396_, _022555_, _022610_);
  and g_114446_(_022608_, _022610_, _022611_);
  or g_114447_(_022607_, _022609_, _022612_);
  and g_114448_(_022605_, _022612_, _022613_);
  or g_114449_(_022606_, _022611_, _022614_);
  and g_114450_(_022595_, _022601_, _022616_);
  or g_114451_(_022594_, _022600_, _022617_);
  and g_114452_(_022614_, _022617_, _022618_);
  or g_114453_(_022613_, _022616_, _022619_);
  and g_114454_(_022606_, _022611_, _022620_);
  or g_114455_(_022605_, _022612_, _022621_);
  and g_114456_(_022590_, _022592_, _022622_);
  or g_114457_(_022589_, _022591_, _022623_);
  and g_114458_(_022587_, _022622_, _022624_);
  or g_114459_(_022588_, _022623_, _022625_);
  and g_114460_(_022603_, _022621_, _022627_);
  or g_114461_(_022602_, _022620_, _022628_);
  and g_114462_(_022618_, _022627_, _022629_);
  or g_114463_(_022619_, _022628_, _022630_);
  and g_114464_(_022624_, _022629_, _022631_);
  or g_114465_(_022625_, _022630_, _022632_);
  xor g_114466_(out[582], _022565_, _022633_);
  xor g_114467_(_055161_, _022565_, _022634_);
  and g_114468_(_022420_, _022555_, _022635_);
  or g_114469_(_022421_, _022556_, _022636_);
  and g_114470_(_022427_, _022556_, _022638_);
  or g_114471_(_022426_, _022555_, _022639_);
  and g_114472_(_022636_, _022639_, _022640_);
  or g_114473_(_022635_, _022638_, _022641_);
  and g_114474_(_022634_, _022641_, _022642_);
  or g_114475_(_022633_, _022640_, _022643_);
  xor g_114476_(out[581], _022564_, _022644_);
  xor g_114477_(_055172_, _022564_, _022645_);
  and g_114478_(_022443_, _022555_, _022646_);
  or g_114479_(_022442_, _022556_, _022647_);
  and g_114480_(_022449_, _022556_, _022649_);
  or g_114481_(_022448_, _022555_, _022650_);
  and g_114482_(_022647_, _022650_, _022651_);
  or g_114483_(_022646_, _022649_, _022652_);
  and g_114484_(_022645_, _022651_, _022653_);
  or g_114485_(_022644_, _022652_, _022654_);
  and g_114486_(_022643_, _022654_, _022655_);
  or g_114487_(_022642_, _022653_, _022656_);
  xor g_114488_(out[583], _022566_, _022657_);
  xor g_114489_(_055150_, _022566_, _022658_);
  and g_114490_(_022410_, _022555_, _022660_);
  or g_114491_(_022409_, _022556_, _022661_);
  and g_114492_(_022416_, _022556_, _022662_);
  or g_114493_(_022415_, _022555_, _022663_);
  and g_114494_(_022661_, _022663_, _022664_);
  or g_114495_(_022660_, _022662_, _022665_);
  and g_114496_(_022658_, _022664_, _022666_);
  or g_114497_(_022657_, _022665_, _022667_);
  xor g_114498_(out[580], out[579], _022668_);
  xor g_114499_(_055183_, out[579], _022669_);
  and g_114500_(_022453_, _022555_, _022671_);
  or g_114501_(_022454_, _022556_, _022672_);
  and g_114502_(_022460_, _022556_, _022673_);
  or g_114503_(_022459_, _022555_, _022674_);
  and g_114504_(_022672_, _022674_, _022675_);
  or g_114505_(_022671_, _022673_, _022676_);
  and g_114506_(_022668_, _022675_, _022677_);
  or g_114507_(_022669_, _022676_, _022678_);
  and g_114508_(_022667_, _022678_, _022679_);
  or g_114509_(_022666_, _022677_, _022680_);
  and g_114510_(_022655_, _022679_, _022682_);
  or g_114511_(_022656_, _022680_, _022683_);
  and g_114512_(_022633_, _022640_, _022684_);
  or g_114513_(_022634_, _022641_, _022685_);
  and g_114514_(_022657_, _022665_, _022686_);
  or g_114515_(_022658_, _022664_, _022687_);
  and g_114516_(_022685_, _022687_, _022688_);
  or g_114517_(_022684_, _022686_, _022689_);
  and g_114518_(_022644_, _022652_, _022690_);
  or g_114519_(_022645_, _022651_, _022691_);
  and g_114520_(_022669_, _022676_, _022693_);
  or g_114521_(_022668_, _022675_, _022694_);
  and g_114522_(_022691_, _022694_, _022695_);
  or g_114523_(_022690_, _022693_, _022696_);
  and g_114524_(_022688_, _022695_, _022697_);
  or g_114525_(_022689_, _022696_, _022698_);
  and g_114526_(_022682_, _022697_, _022699_);
  or g_114527_(_022683_, _022698_, _022700_);
  or g_114528_(_022487_, _022555_, _022701_);
  or g_114529_(out[562], _022556_, _022702_);
  and g_114530_(_022701_, _022702_, _022704_);
  not g_114531_(_022704_, _022705_);
  and g_114532_(_055216_, _022704_, _022706_);
  or g_114533_(out[578], _022705_, _022707_);
  and g_114534_(out[563], _022555_, _022708_);
  or g_114535_(_055095_, _022556_, _022709_);
  and g_114536_(_022482_, _022556_, _022710_);
  or g_114537_(_022481_, _022555_, _022711_);
  and g_114538_(_022709_, _022711_, _022712_);
  or g_114539_(_022708_, _022710_, _022713_);
  and g_114540_(out[579], _022712_, _022715_);
  or g_114541_(_055227_, _022713_, _022716_);
  and g_114542_(_055227_, _022713_, _022717_);
  or g_114543_(out[579], _022712_, _022718_);
  xor g_114544_(_055216_, _022704_, _022719_);
  xor g_114545_(out[578], _022704_, _022720_);
  and g_114546_(_022718_, _022719_, _022721_);
  or g_114547_(_022717_, _022720_, _022722_);
  and g_114548_(_022716_, _022721_, _022723_);
  or g_114549_(_022715_, _022722_, _022724_);
  and g_114550_(_055194_, _022559_, _022726_);
  or g_114551_(out[577], _022561_, _022727_);
  and g_114552_(_022502_, _022556_, _022728_);
  or g_114553_(_022501_, _022555_, _022729_);
  and g_114554_(_055073_, _022555_, _022730_);
  or g_114555_(out[560], _022556_, _022731_);
  and g_114556_(_022729_, _022731_, _022732_);
  or g_114557_(_022728_, _022730_, _022733_);
  and g_114558_(out[576], _022733_, _022734_);
  or g_114559_(_055205_, _022732_, _022735_);
  xor g_114560_(_055194_, _022559_, _022737_);
  xor g_114561_(out[577], _022559_, _022738_);
  and g_114562_(_022735_, _022737_, _022739_);
  or g_114563_(_022734_, _022738_, _022740_);
  and g_114564_(_022727_, _022740_, _022741_);
  or g_114565_(_022726_, _022739_, _022742_);
  and g_114566_(_022723_, _022742_, _022743_);
  or g_114567_(_022724_, _022741_, _022744_);
  and g_114568_(_022706_, _022718_, _022745_);
  or g_114569_(_022707_, _022717_, _022746_);
  and g_114570_(_022716_, _022746_, _022748_);
  or g_114571_(_022715_, _022745_, _022749_);
  and g_114572_(_022744_, _022748_, _022750_);
  or g_114573_(_022743_, _022749_, _022751_);
  and g_114574_(_022699_, _022751_, _022752_);
  or g_114575_(_022700_, _022750_, _022753_);
  and g_114576_(_022655_, _022696_, _022754_);
  or g_114577_(_022656_, _022695_, _022755_);
  and g_114578_(_022688_, _022755_, _022756_);
  or g_114579_(_022689_, _022754_, _022757_);
  and g_114580_(_022667_, _022757_, _022759_);
  or g_114581_(_022666_, _022756_, _022760_);
  and g_114582_(_022753_, _022760_, _022761_);
  or g_114583_(_022752_, _022759_, _022762_);
  and g_114584_(_022631_, _022762_, _022763_);
  or g_114585_(_022632_, _022761_, _022764_);
  and g_114586_(_022588_, _022592_, _022765_);
  or g_114587_(_022587_, _022591_, _022766_);
  and g_114588_(_022603_, _022619_, _022767_);
  or g_114589_(_022602_, _022618_, _022768_);
  and g_114590_(_022624_, _022767_, _022770_);
  or g_114591_(_022625_, _022768_, _022771_);
  and g_114592_(_022766_, _022771_, _022772_);
  or g_114593_(_022765_, _022770_, _022773_);
  and g_114594_(_022764_, _022772_, _022774_);
  or g_114595_(_022763_, _022773_, _022775_);
  and g_114596_(_055205_, _022732_, _022776_);
  or g_114597_(out[576], _022733_, _022777_);
  and g_114598_(_022739_, _022777_, _022778_);
  or g_114599_(_022740_, _022776_, _022779_);
  and g_114600_(_022723_, _022778_, _022781_);
  or g_114601_(_022724_, _022779_, _022782_);
  and g_114602_(_022631_, _022781_, _022783_);
  or g_114603_(_022632_, _022782_, _022784_);
  and g_114604_(_022699_, _022783_, _022785_);
  or g_114605_(_022700_, _022784_, _022786_);
  and g_114606_(_022775_, _022786_, _022787_);
  or g_114607_(_022774_, _022785_, _022788_);
  and g_114608_(_022561_, _022788_, _022789_);
  or g_114609_(_022559_, _022787_, _022790_);
  and g_114610_(_055194_, _022787_, _022792_);
  or g_114611_(out[577], _022788_, _022793_);
  and g_114612_(_022790_, _022793_, _022794_);
  or g_114613_(_022789_, _022792_, _022795_);
  and g_114614_(_022562_, _022572_, _022796_);
  or g_114615_(_022563_, _022573_, _022797_);
  and g_114616_(out[596], out[595], _022798_);
  or g_114617_(out[597], _022798_, _022799_);
  or g_114618_(out[598], _022799_, _022800_);
  or g_114619_(out[599], _022800_, _022801_);
  or g_114620_(out[600], _022801_, _022803_);
  and g_114621_(out[601], _022803_, _022804_);
  or g_114622_(out[602], _022804_, _022805_);
  xor g_114623_(out[603], _022805_, _022806_);
  xor g_114624_(_055271_, _022805_, _022807_);
  and g_114625_(_022796_, _022807_, _022808_);
  or g_114626_(_022797_, _022806_, _022809_);
  and g_114627_(_022581_, _022788_, _022810_);
  or g_114628_(_022580_, _022787_, _022811_);
  and g_114629_(_022583_, _022787_, _022812_);
  or g_114630_(_022584_, _022788_, _022814_);
  and g_114631_(_022811_, _022814_, _022815_);
  or g_114632_(_022810_, _022812_, _022816_);
  xor g_114633_(out[602], _022804_, _022817_);
  xor g_114634_(_055392_, _022804_, _022818_);
  and g_114635_(_022815_, _022817_, _022819_);
  or g_114636_(_022816_, _022818_, _022820_);
  and g_114637_(_022809_, _022820_, _022821_);
  or g_114638_(_022808_, _022819_, _022822_);
  xor g_114639_(out[601], _022803_, _022823_);
  xor g_114640_(_055381_, _022803_, _022825_);
  and g_114641_(_022601_, _022788_, _022826_);
  or g_114642_(_022600_, _022787_, _022827_);
  and g_114643_(_022594_, _022787_, _022828_);
  or g_114644_(_022595_, _022788_, _022829_);
  and g_114645_(_022827_, _022829_, _022830_);
  or g_114646_(_022826_, _022828_, _022831_);
  and g_114647_(_022823_, _022830_, _022832_);
  or g_114648_(_022825_, _022831_, _022833_);
  and g_114649_(_022797_, _022806_, _022834_);
  or g_114650_(_022796_, _022807_, _022836_);
  and g_114651_(_022816_, _022818_, _022837_);
  or g_114652_(_022815_, _022817_, _022838_);
  and g_114653_(_022836_, _022838_, _022839_);
  or g_114654_(_022834_, _022837_, _022840_);
  and g_114655_(_022833_, _022839_, _022841_);
  or g_114656_(_022832_, _022840_, _022842_);
  and g_114657_(_022821_, _022841_, _022843_);
  or g_114658_(_022822_, _022842_, _022844_);
  xor g_114659_(out[600], _022801_, _022845_);
  xor g_114660_(_055370_, _022801_, _022847_);
  and g_114661_(_022612_, _022788_, _022848_);
  or g_114662_(_022611_, _022787_, _022849_);
  and g_114663_(_022606_, _022787_, _022850_);
  or g_114664_(_022605_, _022788_, _022851_);
  and g_114665_(_022849_, _022851_, _022852_);
  or g_114666_(_022848_, _022850_, _022853_);
  and g_114667_(_022845_, _022853_, _022854_);
  or g_114668_(_022847_, _022852_, _022855_);
  and g_114669_(_022825_, _022831_, _022856_);
  or g_114670_(_022823_, _022830_, _022858_);
  and g_114671_(_022855_, _022858_, _022859_);
  or g_114672_(_022854_, _022856_, _022860_);
  or g_114673_(_022845_, _022853_, _022861_);
  and g_114674_(_022859_, _022861_, _022862_);
  and g_114675_(_022843_, _022862_, _022863_);
  not g_114676_(_022863_, _022864_);
  xor g_114677_(out[598], _022799_, _022865_);
  xor g_114678_(_055293_, _022799_, _022866_);
  and g_114679_(_022641_, _022788_, _022867_);
  or g_114680_(_022640_, _022787_, _022869_);
  and g_114681_(_022633_, _022787_, _022870_);
  or g_114682_(_022634_, _022788_, _022871_);
  and g_114683_(_022869_, _022871_, _022872_);
  or g_114684_(_022867_, _022870_, _022873_);
  and g_114685_(_022865_, _022872_, _022874_);
  or g_114686_(_022866_, _022873_, _022875_);
  xor g_114687_(out[599], _022800_, _022876_);
  xor g_114688_(_055282_, _022800_, _022877_);
  and g_114689_(_022665_, _022788_, _022878_);
  or g_114690_(_022664_, _022787_, _022880_);
  and g_114691_(_022658_, _022787_, _022881_);
  or g_114692_(_022657_, _022788_, _022882_);
  and g_114693_(_022880_, _022882_, _022883_);
  or g_114694_(_022878_, _022881_, _022884_);
  and g_114695_(_022876_, _022884_, _022885_);
  or g_114696_(_022877_, _022883_, _022886_);
  and g_114697_(_022875_, _022886_, _022887_);
  or g_114698_(_022874_, _022885_, _022888_);
  and g_114699_(_022877_, _022883_, _022889_);
  or g_114700_(_022876_, _022884_, _022891_);
  and g_114701_(_022866_, _022873_, _022892_);
  or g_114702_(_022865_, _022872_, _022893_);
  and g_114703_(_022891_, _022893_, _022894_);
  or g_114704_(_022889_, _022892_, _022895_);
  and g_114705_(_022887_, _022894_, _022896_);
  or g_114706_(_022888_, _022895_, _022897_);
  xor g_114707_(out[597], _022798_, _022898_);
  xor g_114708_(_055304_, _022798_, _022899_);
  and g_114709_(_022652_, _022788_, _022900_);
  or g_114710_(_022651_, _022787_, _022902_);
  and g_114711_(_022645_, _022787_, _022903_);
  or g_114712_(_022644_, _022788_, _022904_);
  and g_114713_(_022902_, _022904_, _022905_);
  or g_114714_(_022900_, _022903_, _022906_);
  and g_114715_(_022898_, _022906_, _022907_);
  or g_114716_(_022899_, _022905_, _022908_);
  xor g_114717_(out[596], out[595], _022909_);
  xor g_114718_(_055315_, out[595], _022910_);
  and g_114719_(_022668_, _022787_, _022911_);
  or g_114720_(_022669_, _022788_, _022913_);
  and g_114721_(_022676_, _022788_, _022914_);
  or g_114722_(_022675_, _022787_, _022915_);
  and g_114723_(_022913_, _022915_, _022916_);
  or g_114724_(_022911_, _022914_, _022917_);
  and g_114725_(_022910_, _022917_, _022918_);
  or g_114726_(_022909_, _022916_, _022919_);
  and g_114727_(_022908_, _022919_, _022920_);
  or g_114728_(_022907_, _022918_, _022921_);
  and g_114729_(_022899_, _022905_, _022922_);
  or g_114730_(_022898_, _022906_, _022924_);
  and g_114731_(_022909_, _022916_, _022925_);
  or g_114732_(_022910_, _022917_, _022926_);
  and g_114733_(_022924_, _022926_, _022927_);
  or g_114734_(_022922_, _022925_, _022928_);
  and g_114735_(_022920_, _022927_, _022929_);
  or g_114736_(_022921_, _022928_, _022930_);
  and g_114737_(_022896_, _022929_, _022931_);
  or g_114738_(_022897_, _022930_, _022932_);
  and g_114739_(out[579], _022787_, _022933_);
  not g_114740_(_022933_, _022935_);
  and g_114741_(_022713_, _022788_, _022936_);
  or g_114742_(_022712_, _022787_, _022937_);
  and g_114743_(_022935_, _022937_, _022938_);
  or g_114744_(_022933_, _022936_, _022939_);
  and g_114745_(out[595], _022938_, _022940_);
  or g_114746_(_055359_, _022939_, _022941_);
  or g_114747_(_022704_, _022787_, _022942_);
  or g_114748_(out[578], _022788_, _022943_);
  and g_114749_(_022942_, _022943_, _022944_);
  not g_114750_(_022944_, _022946_);
  and g_114751_(_055348_, _022944_, _022947_);
  or g_114752_(out[594], _022946_, _022948_);
  and g_114753_(_022941_, _022948_, _022949_);
  or g_114754_(_022940_, _022947_, _022950_);
  and g_114755_(_055359_, _022939_, _022951_);
  or g_114756_(out[595], _022938_, _022952_);
  and g_114757_(out[594], _022946_, _022953_);
  or g_114758_(_055348_, _022944_, _022954_);
  and g_114759_(_022952_, _022954_, _022955_);
  or g_114760_(_022951_, _022953_, _022957_);
  and g_114761_(_022949_, _022955_, _022958_);
  or g_114762_(_022950_, _022957_, _022959_);
  and g_114763_(_022733_, _022788_, _022960_);
  or g_114764_(_022732_, _022787_, _022961_);
  and g_114765_(_055205_, _022787_, _022962_);
  or g_114766_(out[576], _022788_, _022963_);
  and g_114767_(_022961_, _022963_, _022964_);
  or g_114768_(_022960_, _022962_, _022965_);
  and g_114769_(out[592], _022965_, _022966_);
  or g_114770_(_055337_, _022964_, _022968_);
  and g_114771_(out[593], _022795_, _022969_);
  or g_114772_(_055326_, _022794_, _022970_);
  and g_114773_(_022968_, _022970_, _022971_);
  or g_114774_(_022966_, _022969_, _022972_);
  and g_114775_(_055326_, _022794_, _022973_);
  not g_114776_(_022973_, _022974_);
  or g_114777_(out[592], _022965_, _022975_);
  and g_114778_(_022958_, _022975_, _022976_);
  and g_114779_(_022971_, _022976_, _022977_);
  and g_114780_(_022863_, _022931_, _022979_);
  and g_114781_(_022977_, _022979_, _022980_);
  not g_114782_(_022980_, _022981_);
  and g_114783_(_022974_, _022980_, _022982_);
  or g_114784_(_022973_, _022981_, _022983_);
  and g_114785_(_022972_, _022974_, _022984_);
  or g_114786_(_022971_, _022973_, _022985_);
  and g_114787_(_022958_, _022985_, _022986_);
  or g_114788_(_022959_, _022984_, _022987_);
  and g_114789_(_022947_, _022952_, _022988_);
  or g_114790_(_022948_, _022951_, _022990_);
  and g_114791_(_022941_, _022990_, _022991_);
  or g_114792_(_022940_, _022988_, _022992_);
  and g_114793_(_022987_, _022991_, _022993_);
  or g_114794_(_022986_, _022992_, _022994_);
  and g_114795_(_022931_, _022994_, _022995_);
  or g_114796_(_022932_, _022993_, _022996_);
  and g_114797_(_022888_, _022891_, _022997_);
  or g_114798_(_022887_, _022889_, _022998_);
  and g_114799_(_022921_, _022924_, _022999_);
  or g_114800_(_022920_, _022922_, _023001_);
  and g_114801_(_022896_, _022999_, _023002_);
  or g_114802_(_022897_, _023001_, _023003_);
  and g_114803_(_022998_, _023003_, _023004_);
  or g_114804_(_022997_, _023002_, _023005_);
  and g_114805_(_022996_, _023004_, _023006_);
  or g_114806_(_022995_, _023005_, _023007_);
  and g_114807_(_022863_, _023007_, _023008_);
  or g_114808_(_022864_, _023006_, _023009_);
  and g_114809_(_022843_, _022860_, _023010_);
  or g_114810_(_022844_, _022859_, _023012_);
  and g_114811_(_022822_, _022836_, _023013_);
  or g_114812_(_022821_, _022834_, _023014_);
  and g_114813_(_023012_, _023014_, _023015_);
  or g_114814_(_023010_, _023013_, _023016_);
  and g_114815_(_023009_, _023015_, _023017_);
  or g_114816_(_023008_, _023016_, _023018_);
  and g_114817_(_022983_, _023018_, _023019_);
  or g_114818_(_022982_, _023017_, _023020_);
  or g_114819_(_022794_, _023019_, _023021_);
  or g_114820_(out[593], _023020_, _023023_);
  and g_114821_(_023021_, _023023_, _023024_);
  not g_114822_(_023024_, _023025_);
  and g_114823_(_022817_, _023019_, _023026_);
  or g_114824_(_022818_, _023020_, _023027_);
  and g_114825_(_022816_, _023020_, _023028_);
  or g_114826_(_022815_, _023019_, _023029_);
  and g_114827_(_023027_, _023029_, _023030_);
  or g_114828_(_023026_, _023028_, _023031_);
  and g_114829_(out[612], out[611], _023032_);
  or g_114830_(out[613], _023032_, _023034_);
  or g_114831_(out[614], _023034_, _023035_);
  or g_114832_(out[615], _023035_, _023036_);
  or g_114833_(out[616], _023036_, _023037_);
  and g_114834_(out[617], _023037_, _023038_);
  or g_114835_(out[618], _023038_, _023039_);
  xor g_114836_(out[618], _023038_, _023040_);
  xor g_114837_(_055524_, _023038_, _023041_);
  and g_114838_(_023030_, _023040_, _023042_);
  or g_114839_(_023031_, _023041_, _023043_);
  and g_114840_(_022796_, _022806_, _023045_);
  or g_114841_(_022797_, _022807_, _023046_);
  xor g_114842_(out[619], _023039_, _023047_);
  xor g_114843_(_055403_, _023039_, _023048_);
  and g_114844_(_023045_, _023048_, _023049_);
  or g_114845_(_023046_, _023047_, _023050_);
  and g_114846_(_023043_, _023050_, _023051_);
  or g_114847_(_023042_, _023049_, _023052_);
  and g_114848_(_023031_, _023041_, _023053_);
  or g_114849_(_023030_, _023040_, _023054_);
  and g_114850_(_023046_, _023047_, _023056_);
  or g_114851_(_023045_, _023048_, _023057_);
  and g_114852_(_023054_, _023057_, _023058_);
  or g_114853_(_023053_, _023056_, _023059_);
  and g_114854_(_023051_, _023058_, _023060_);
  or g_114855_(_023052_, _023059_, _023061_);
  xor g_114856_(out[616], _023036_, _023062_);
  xor g_114857_(_055502_, _023036_, _023063_);
  and g_114858_(_022847_, _023019_, _023064_);
  or g_114859_(_022845_, _023020_, _023065_);
  and g_114860_(_022853_, _023020_, _023067_);
  or g_114861_(_022852_, _023019_, _023068_);
  and g_114862_(_023065_, _023068_, _023069_);
  or g_114863_(_023064_, _023067_, _023070_);
  and g_114864_(_023062_, _023070_, _023071_);
  or g_114865_(_023063_, _023069_, _023072_);
  xor g_114866_(out[617], _023037_, _023073_);
  xor g_114867_(_055513_, _023037_, _023074_);
  and g_114868_(_022823_, _023019_, _023075_);
  or g_114869_(_022825_, _023020_, _023076_);
  and g_114870_(_022831_, _023020_, _023078_);
  or g_114871_(_022830_, _023019_, _023079_);
  and g_114872_(_023076_, _023079_, _023080_);
  or g_114873_(_023075_, _023078_, _023081_);
  and g_114874_(_023074_, _023081_, _023082_);
  or g_114875_(_023073_, _023080_, _023083_);
  and g_114876_(_023072_, _023083_, _023084_);
  or g_114877_(_023071_, _023082_, _023085_);
  and g_114878_(_023073_, _023080_, _023086_);
  or g_114879_(_023074_, _023081_, _023087_);
  and g_114880_(_023063_, _023069_, _023089_);
  or g_114881_(_023062_, _023070_, _023090_);
  and g_114882_(_023087_, _023090_, _023091_);
  or g_114883_(_023086_, _023089_, _023092_);
  and g_114884_(_023084_, _023091_, _023093_);
  or g_114885_(_023085_, _023092_, _023094_);
  and g_114886_(_023060_, _023093_, _023095_);
  or g_114887_(_023061_, _023094_, _023096_);
  xor g_114888_(out[615], _023035_, _023097_);
  not g_114889_(_023097_, _023098_);
  and g_114890_(_022877_, _023019_, _023100_);
  or g_114891_(_022876_, _023020_, _023101_);
  and g_114892_(_022884_, _023020_, _023102_);
  or g_114893_(_022883_, _023019_, _023103_);
  and g_114894_(_023101_, _023103_, _023104_);
  or g_114895_(_023100_, _023102_, _023105_);
  and g_114896_(_023097_, _023105_, _023106_);
  or g_114897_(_023098_, _023104_, _023107_);
  xor g_114898_(out[614], _023034_, _023108_);
  xor g_114899_(_055425_, _023034_, _023109_);
  and g_114900_(_022865_, _023019_, _023111_);
  or g_114901_(_022866_, _023020_, _023112_);
  and g_114902_(_022873_, _023020_, _023113_);
  or g_114903_(_022872_, _023019_, _023114_);
  and g_114904_(_023112_, _023114_, _023115_);
  or g_114905_(_023111_, _023113_, _023116_);
  and g_114906_(_023108_, _023115_, _023117_);
  or g_114907_(_023109_, _023116_, _023118_);
  and g_114908_(_023107_, _023118_, _023119_);
  or g_114909_(_023106_, _023117_, _023120_);
  and g_114910_(_023109_, _023116_, _023122_);
  or g_114911_(_023108_, _023115_, _023123_);
  and g_114912_(_023098_, _023104_, _023124_);
  or g_114913_(_023097_, _023105_, _023125_);
  and g_114914_(_023123_, _023125_, _023126_);
  or g_114915_(_023122_, _023124_, _023127_);
  and g_114916_(_023119_, _023126_, _023128_);
  or g_114917_(_023120_, _023127_, _023129_);
  xor g_114918_(out[612], out[611], _023130_);
  xor g_114919_(_055447_, out[611], _023131_);
  and g_114920_(_022909_, _023019_, _023133_);
  or g_114921_(_022910_, _023020_, _023134_);
  and g_114922_(_022917_, _023020_, _023135_);
  or g_114923_(_022916_, _023019_, _023136_);
  and g_114924_(_023134_, _023136_, _023137_);
  or g_114925_(_023133_, _023135_, _023138_);
  and g_114926_(_023131_, _023138_, _023139_);
  or g_114927_(_023130_, _023137_, _023140_);
  xor g_114928_(out[613], _023032_, _023141_);
  xor g_114929_(_055436_, _023032_, _023142_);
  and g_114930_(_022899_, _023019_, _023144_);
  or g_114931_(_022898_, _023020_, _023145_);
  and g_114932_(_022906_, _023020_, _023146_);
  or g_114933_(_022905_, _023019_, _023147_);
  and g_114934_(_023145_, _023147_, _023148_);
  or g_114935_(_023144_, _023146_, _023149_);
  and g_114936_(_023141_, _023149_, _023150_);
  or g_114937_(_023142_, _023148_, _023151_);
  and g_114938_(_023140_, _023151_, _023152_);
  or g_114939_(_023139_, _023150_, _023153_);
  and g_114940_(_023142_, _023148_, _023155_);
  or g_114941_(_023141_, _023149_, _023156_);
  and g_114942_(_023130_, _023137_, _023157_);
  or g_114943_(_023131_, _023138_, _023158_);
  and g_114944_(_023156_, _023158_, _023159_);
  or g_114945_(_023155_, _023157_, _023160_);
  and g_114946_(_023152_, _023159_, _023161_);
  or g_114947_(_023153_, _023160_, _023162_);
  and g_114948_(_023128_, _023161_, _023163_);
  or g_114949_(_023129_, _023162_, _023164_);
  and g_114950_(_023095_, _023163_, _023166_);
  or g_114951_(_023096_, _023164_, _023167_);
  or g_114952_(_055359_, _023020_, _023168_);
  or g_114953_(_022938_, _023019_, _023169_);
  and g_114954_(_023168_, _023169_, _023170_);
  not g_114955_(_023170_, _023171_);
  and g_114956_(out[611], _023170_, _023172_);
  or g_114957_(_022944_, _023019_, _023173_);
  or g_114958_(out[594], _023020_, _023174_);
  and g_114959_(_023173_, _023174_, _023175_);
  and g_114960_(_055480_, _023175_, _023177_);
  or g_114961_(out[611], _023170_, _023178_);
  xor g_114962_(_055491_, _023170_, _023179_);
  xor g_114963_(out[610], _023175_, _023180_);
  or g_114964_(_023179_, _023180_, _023181_);
  not g_114965_(_023181_, _023182_);
  and g_114966_(_055458_, _023024_, _023183_);
  or g_114967_(out[609], _023025_, _023184_);
  and g_114968_(_022965_, _023020_, _023185_);
  or g_114969_(_022964_, _023019_, _023186_);
  and g_114970_(_055337_, _023019_, _023188_);
  or g_114971_(out[592], _023020_, _023189_);
  and g_114972_(_023186_, _023189_, _023190_);
  or g_114973_(_023185_, _023188_, _023191_);
  and g_114974_(out[608], _023191_, _023192_);
  or g_114975_(_055469_, _023190_, _023193_);
  xor g_114976_(_055458_, _023024_, _023194_);
  xor g_114977_(out[609], _023024_, _023195_);
  and g_114978_(_023193_, _023194_, _023196_);
  or g_114979_(_023192_, _023195_, _023197_);
  and g_114980_(_023184_, _023197_, _023199_);
  or g_114981_(_023183_, _023196_, _023200_);
  and g_114982_(_023182_, _023200_, _023201_);
  or g_114983_(_023181_, _023199_, _023202_);
  and g_114984_(_023177_, _023178_, _023203_);
  or g_114985_(_023172_, _023203_, _023204_);
  not g_114986_(_023204_, _023205_);
  and g_114987_(_023202_, _023205_, _023206_);
  or g_114988_(_023201_, _023204_, _023207_);
  and g_114989_(_023166_, _023207_, _023208_);
  or g_114990_(_023167_, _023206_, _023210_);
  and g_114991_(_023153_, _023156_, _023211_);
  or g_114992_(_023152_, _023155_, _023212_);
  and g_114993_(_023128_, _023211_, _023213_);
  or g_114994_(_023129_, _023212_, _023214_);
  or g_114995_(_023119_, _023124_, _023215_);
  not g_114996_(_023215_, _023216_);
  and g_114997_(_023214_, _023215_, _023217_);
  or g_114998_(_023213_, _023216_, _023218_);
  and g_114999_(_023095_, _023218_, _023219_);
  or g_115000_(_023096_, _023217_, _023221_);
  and g_115001_(_023052_, _023057_, _023222_);
  or g_115002_(_023051_, _023056_, _023223_);
  and g_115003_(_023085_, _023087_, _023224_);
  or g_115004_(_023084_, _023086_, _023225_);
  and g_115005_(_023060_, _023224_, _023226_);
  or g_115006_(_023061_, _023225_, _023227_);
  and g_115007_(_023223_, _023227_, _023228_);
  or g_115008_(_023222_, _023226_, _023229_);
  and g_115009_(_023210_, _023228_, _023230_);
  or g_115010_(_023208_, _023229_, _023232_);
  and g_115011_(_023221_, _023230_, _023233_);
  or g_115012_(_023219_, _023232_, _023234_);
  and g_115013_(_055469_, _023190_, _023235_);
  or g_115014_(_023181_, _023235_, _023236_);
  or g_115015_(_023197_, _023236_, _023237_);
  or g_115016_(_023167_, _023237_, _023238_);
  not g_115017_(_023238_, _023239_);
  and g_115018_(_023234_, _023238_, _023240_);
  or g_115019_(_023233_, _023239_, _023241_);
  or g_115020_(_023024_, _023240_, _023243_);
  or g_115021_(out[609], _023241_, _023244_);
  and g_115022_(_023243_, _023244_, _023245_);
  not g_115023_(_023245_, _023246_);
  and g_115024_(out[628], out[627], _023247_);
  or g_115025_(out[629], _023247_, _023248_);
  or g_115026_(out[630], _023248_, _023249_);
  xor g_115027_(out[630], _023248_, _023250_);
  xor g_115028_(_055557_, _023248_, _023251_);
  and g_115029_(_023108_, _023240_, _023252_);
  or g_115030_(_023109_, _023241_, _023254_);
  and g_115031_(_023116_, _023241_, _023255_);
  or g_115032_(_023115_, _023240_, _023256_);
  and g_115033_(_023254_, _023256_, _023257_);
  or g_115034_(_023252_, _023255_, _023258_);
  and g_115035_(_023250_, _023257_, _023259_);
  or g_115036_(_023251_, _023258_, _023260_);
  xor g_115037_(out[629], _023247_, _023261_);
  xor g_115038_(_055568_, _023247_, _023262_);
  or g_115039_(_023141_, _023241_, _023263_);
  not g_115040_(_023263_, _023265_);
  and g_115041_(_023149_, _023241_, _023266_);
  or g_115042_(_023148_, _023240_, _023267_);
  and g_115043_(_023263_, _023267_, _023268_);
  or g_115044_(_023265_, _023266_, _023269_);
  and g_115045_(_023262_, _023268_, _023270_);
  or g_115046_(_023261_, _023269_, _023271_);
  and g_115047_(_023260_, _023271_, _023272_);
  or g_115048_(_023259_, _023270_, _023273_);
  or g_115049_(out[631], _023249_, _023274_);
  xor g_115050_(out[631], _023249_, _023276_);
  xor g_115051_(_055546_, _023249_, _023277_);
  or g_115052_(_023097_, _023241_, _023278_);
  or g_115053_(_023104_, _023240_, _023279_);
  and g_115054_(_023278_, _023279_, _023280_);
  not g_115055_(_023280_, _023281_);
  or g_115056_(_023277_, _023280_, _023282_);
  and g_115057_(_023277_, _023280_, _023283_);
  xor g_115058_(_023277_, _023280_, _023284_);
  xor g_115059_(_023276_, _023280_, _023285_);
  and g_115060_(_023251_, _023258_, _023287_);
  or g_115061_(_023250_, _023257_, _023288_);
  and g_115062_(_023284_, _023288_, _023289_);
  or g_115063_(_023285_, _023287_, _023290_);
  and g_115064_(_023272_, _023289_, _023291_);
  or g_115065_(_023273_, _023290_, _023292_);
  xor g_115066_(out[628], out[627], _023293_);
  xor g_115067_(_055579_, out[627], _023294_);
  or g_115068_(_023131_, _023241_, _023295_);
  not g_115069_(_023295_, _023296_);
  and g_115070_(_023138_, _023241_, _023298_);
  not g_115071_(_023298_, _023299_);
  and g_115072_(_023295_, _023299_, _023300_);
  or g_115073_(_023296_, _023298_, _023301_);
  and g_115074_(_023294_, _023301_, _023302_);
  or g_115075_(_023293_, _023300_, _023303_);
  and g_115076_(_023261_, _023269_, _023304_);
  or g_115077_(_023262_, _023268_, _023305_);
  and g_115078_(_023303_, _023305_, _023306_);
  or g_115079_(_023302_, _023304_, _023307_);
  and g_115080_(_023293_, _023300_, _023309_);
  or g_115081_(_023294_, _023301_, _023310_);
  and g_115082_(_023306_, _023310_, _023311_);
  or g_115083_(_023307_, _023309_, _023312_);
  and g_115084_(_023291_, _023311_, _023313_);
  or g_115085_(_023292_, _023312_, _023314_);
  and g_115086_(_023045_, _023047_, _023315_);
  or g_115087_(_023046_, _023048_, _023316_);
  or g_115088_(out[632], _023274_, _023317_);
  and g_115089_(out[633], _023317_, _023318_);
  or g_115090_(out[634], _023318_, _023320_);
  xor g_115091_(out[635], _023320_, _023321_);
  xor g_115092_(_055535_, _023320_, _023322_);
  and g_115093_(_023315_, _023322_, _023323_);
  or g_115094_(_023316_, _023321_, _023324_);
  or g_115095_(_023041_, _023241_, _023325_);
  not g_115096_(_023325_, _023326_);
  and g_115097_(_023031_, _023241_, _023327_);
  not g_115098_(_023327_, _023328_);
  and g_115099_(_023325_, _023328_, _023329_);
  or g_115100_(_023326_, _023327_, _023331_);
  xor g_115101_(out[634], _023318_, _023332_);
  xor g_115102_(_055656_, _023318_, _023333_);
  and g_115103_(_023329_, _023332_, _023334_);
  or g_115104_(_023331_, _023333_, _023335_);
  and g_115105_(_023324_, _023335_, _023336_);
  or g_115106_(_023323_, _023334_, _023337_);
  and g_115107_(_023331_, _023333_, _023338_);
  or g_115108_(_023329_, _023332_, _023339_);
  and g_115109_(_023316_, _023321_, _023340_);
  or g_115110_(_023315_, _023322_, _023342_);
  and g_115111_(_023339_, _023342_, _023343_);
  or g_115112_(_023338_, _023340_, _023344_);
  and g_115113_(_023336_, _023343_, _023345_);
  or g_115114_(_023337_, _023344_, _023346_);
  xor g_115115_(out[632], _023274_, _023347_);
  xor g_115116_(_055634_, _023274_, _023348_);
  or g_115117_(_023062_, _023241_, _023349_);
  not g_115118_(_023349_, _023350_);
  and g_115119_(_023070_, _023241_, _023351_);
  not g_115120_(_023351_, _023353_);
  and g_115121_(_023349_, _023353_, _023354_);
  or g_115122_(_023350_, _023351_, _023355_);
  and g_115123_(_023347_, _023355_, _023356_);
  or g_115124_(_023348_, _023354_, _023357_);
  xor g_115125_(out[633], _023317_, _023358_);
  xor g_115126_(_055645_, _023317_, _023359_);
  or g_115127_(_023074_, _023241_, _023360_);
  not g_115128_(_023360_, _023361_);
  and g_115129_(_023081_, _023241_, _023362_);
  not g_115130_(_023362_, _023364_);
  and g_115131_(_023360_, _023364_, _023365_);
  or g_115132_(_023361_, _023362_, _023366_);
  and g_115133_(_023359_, _023366_, _023367_);
  or g_115134_(_023358_, _023365_, _023368_);
  and g_115135_(_023357_, _023368_, _023369_);
  or g_115136_(_023356_, _023367_, _023370_);
  and g_115137_(_023348_, _023354_, _023371_);
  or g_115138_(_023347_, _023355_, _023372_);
  and g_115139_(_023358_, _023365_, _023373_);
  or g_115140_(_023359_, _023366_, _023375_);
  and g_115141_(_023372_, _023375_, _023376_);
  or g_115142_(_023371_, _023373_, _023377_);
  and g_115143_(_023369_, _023376_, _023378_);
  or g_115144_(_023370_, _023377_, _023379_);
  and g_115145_(_023345_, _023378_, _023380_);
  or g_115146_(_023346_, _023379_, _023381_);
  or g_115147_(_023175_, _023240_, _023382_);
  or g_115148_(out[610], _023241_, _023383_);
  and g_115149_(_023382_, _023383_, _023384_);
  not g_115150_(_023384_, _023386_);
  and g_115151_(_055612_, _023384_, _023387_);
  or g_115152_(out[626], _023386_, _023388_);
  and g_115153_(out[611], _023240_, _023389_);
  or g_115154_(_055491_, _023241_, _023390_);
  and g_115155_(_023171_, _023241_, _023391_);
  or g_115156_(_023170_, _023240_, _023392_);
  and g_115157_(_023390_, _023392_, _023393_);
  or g_115158_(_023389_, _023391_, _023394_);
  and g_115159_(out[627], _023393_, _023395_);
  or g_115160_(_055623_, _023394_, _023397_);
  and g_115161_(_055623_, _023394_, _023398_);
  or g_115162_(out[627], _023393_, _023399_);
  xor g_115163_(_055612_, _023384_, _023400_);
  xor g_115164_(out[626], _023384_, _023401_);
  and g_115165_(_023399_, _023400_, _023402_);
  or g_115166_(_023398_, _023401_, _023403_);
  and g_115167_(_023397_, _023402_, _023404_);
  or g_115168_(_023395_, _023403_, _023405_);
  and g_115169_(_023191_, _023241_, _023406_);
  or g_115170_(_023190_, _023240_, _023408_);
  and g_115171_(_055469_, _023240_, _023409_);
  or g_115172_(out[608], _023241_, _023410_);
  and g_115173_(_023408_, _023410_, _023411_);
  or g_115174_(_023406_, _023409_, _023412_);
  and g_115175_(out[624], _023412_, _023413_);
  or g_115176_(_055601_, _023411_, _023414_);
  and g_115177_(_055590_, _023245_, _023415_);
  or g_115178_(out[625], _023246_, _023416_);
  xor g_115179_(_055590_, _023245_, _023417_);
  xor g_115180_(out[625], _023245_, _023419_);
  and g_115181_(_023414_, _023417_, _023420_);
  or g_115182_(_023413_, _023419_, _023421_);
  and g_115183_(_055601_, _023411_, _023422_);
  not g_115184_(_023422_, _023423_);
  and g_115185_(_023420_, _023423_, _023424_);
  and g_115186_(_023404_, _023424_, _023425_);
  and g_115187_(_023380_, _023425_, _023426_);
  and g_115188_(_023313_, _023426_, _023427_);
  not g_115189_(_023427_, _023428_);
  and g_115190_(_023416_, _023421_, _023430_);
  or g_115191_(_023415_, _023420_, _023431_);
  and g_115192_(_023404_, _023431_, _023432_);
  or g_115193_(_023405_, _023430_, _023433_);
  and g_115194_(_023387_, _023399_, _023434_);
  or g_115195_(_023388_, _023398_, _023435_);
  and g_115196_(_023397_, _023435_, _023436_);
  or g_115197_(_023395_, _023434_, _023437_);
  and g_115198_(_023433_, _023436_, _023438_);
  or g_115199_(_023432_, _023437_, _023439_);
  and g_115200_(_023313_, _023439_, _023441_);
  or g_115201_(_023314_, _023438_, _023442_);
  and g_115202_(_023291_, _023307_, _023443_);
  or g_115203_(_023292_, _023306_, _023444_);
  or g_115204_(_023260_, _023283_, _023445_);
  and g_115205_(_023282_, _023445_, _023446_);
  not g_115206_(_023446_, _023447_);
  and g_115207_(_023444_, _023446_, _023448_);
  or g_115208_(_023443_, _023447_, _023449_);
  and g_115209_(_023442_, _023448_, _023450_);
  or g_115210_(_023441_, _023449_, _023452_);
  and g_115211_(_023380_, _023452_, _023453_);
  or g_115212_(_023381_, _023450_, _023454_);
  and g_115213_(_023370_, _023375_, _023455_);
  or g_115214_(_023369_, _023373_, _023456_);
  and g_115215_(_023345_, _023455_, _023457_);
  or g_115216_(_023346_, _023456_, _023458_);
  and g_115217_(_023337_, _023342_, _023459_);
  or g_115218_(_023336_, _023340_, _023460_);
  and g_115219_(_023458_, _023460_, _023461_);
  or g_115220_(_023457_, _023459_, _023463_);
  and g_115221_(_023454_, _023461_, _023464_);
  or g_115222_(_023453_, _023463_, _023465_);
  and g_115223_(_023428_, _023465_, _023466_);
  or g_115224_(_023427_, _023464_, _023467_);
  or g_115225_(_023245_, _023466_, _023468_);
  or g_115226_(out[625], _023467_, _023469_);
  and g_115227_(_023468_, _023469_, _023470_);
  not g_115228_(_023470_, _023471_);
  and g_115229_(_023332_, _023466_, _023472_);
  not g_115230_(_023472_, _023474_);
  and g_115231_(_023331_, _023467_, _023475_);
  or g_115232_(_023329_, _023466_, _023476_);
  and g_115233_(_023474_, _023476_, _023477_);
  or g_115234_(_023472_, _023475_, _023478_);
  and g_115235_(out[644], out[643], _023479_);
  or g_115236_(out[645], _023479_, _023480_);
  or g_115237_(out[646], _023480_, _023481_);
  or g_115238_(out[647], _023481_, _023482_);
  or g_115239_(out[648], _023482_, _023483_);
  and g_115240_(out[649], _023483_, _023485_);
  or g_115241_(out[650], _023485_, _023486_);
  xor g_115242_(out[650], _023485_, _023487_);
  xor g_115243_(_055788_, _023485_, _023488_);
  and g_115244_(_023477_, _023487_, _023489_);
  or g_115245_(_023478_, _023488_, _023490_);
  and g_115246_(_023315_, _023321_, _023491_);
  or g_115247_(_023316_, _023322_, _023492_);
  xor g_115248_(out[651], _023486_, _023493_);
  xor g_115249_(_055667_, _023486_, _023494_);
  and g_115250_(_023491_, _023494_, _023496_);
  or g_115251_(_023492_, _023493_, _023497_);
  and g_115252_(_023490_, _023497_, _023498_);
  or g_115253_(_023489_, _023496_, _023499_);
  xor g_115254_(out[649], _023483_, _023500_);
  xor g_115255_(_055777_, _023483_, _023501_);
  and g_115256_(_023358_, _023466_, _023502_);
  not g_115257_(_023502_, _023503_);
  and g_115258_(_023366_, _023467_, _023504_);
  or g_115259_(_023365_, _023466_, _023505_);
  and g_115260_(_023503_, _023505_, _023507_);
  or g_115261_(_023502_, _023504_, _023508_);
  and g_115262_(_023500_, _023507_, _023509_);
  or g_115263_(_023501_, _023508_, _023510_);
  and g_115264_(_023492_, _023493_, _023511_);
  or g_115265_(_023491_, _023494_, _023512_);
  and g_115266_(_023478_, _023488_, _023513_);
  or g_115267_(_023477_, _023487_, _023514_);
  and g_115268_(_023512_, _023514_, _023515_);
  or g_115269_(_023511_, _023513_, _023516_);
  xor g_115270_(out[648], _023482_, _023518_);
  xor g_115271_(_055766_, _023482_, _023519_);
  and g_115272_(_023348_, _023466_, _023520_);
  or g_115273_(_023347_, _023467_, _023521_);
  and g_115274_(_023355_, _023467_, _023522_);
  or g_115275_(_023354_, _023466_, _023523_);
  and g_115276_(_023521_, _023523_, _023524_);
  or g_115277_(_023520_, _023522_, _023525_);
  and g_115278_(_023518_, _023525_, _023526_);
  or g_115279_(_023519_, _023524_, _023527_);
  and g_115280_(_023501_, _023508_, _023529_);
  or g_115281_(_023500_, _023507_, _023530_);
  and g_115282_(_023527_, _023530_, _023531_);
  or g_115283_(_023526_, _023529_, _023532_);
  and g_115284_(_023519_, _023524_, _023533_);
  or g_115285_(_023518_, _023525_, _023534_);
  and g_115286_(_023498_, _023515_, _023535_);
  or g_115287_(_023499_, _023516_, _023536_);
  and g_115288_(_023510_, _023534_, _023537_);
  or g_115289_(_023509_, _023533_, _023538_);
  and g_115290_(_023531_, _023537_, _023540_);
  or g_115291_(_023532_, _023538_, _023541_);
  and g_115292_(_023535_, _023540_, _023542_);
  or g_115293_(_023536_, _023541_, _023543_);
  xor g_115294_(out[647], _023481_, _023544_);
  not g_115295_(_023544_, _023545_);
  and g_115296_(_023277_, _023466_, _023546_);
  or g_115297_(_023276_, _023467_, _023547_);
  and g_115298_(_023281_, _023467_, _023548_);
  or g_115299_(_023280_, _023466_, _023549_);
  and g_115300_(_023547_, _023549_, _023551_);
  or g_115301_(_023546_, _023548_, _023552_);
  or g_115302_(_023545_, _023551_, _023553_);
  not g_115303_(_023553_, _023554_);
  xor g_115304_(out[646], _023480_, _023555_);
  xor g_115305_(_055689_, _023480_, _023556_);
  and g_115306_(_023250_, _023466_, _023557_);
  or g_115307_(_023251_, _023467_, _023558_);
  and g_115308_(_023258_, _023467_, _023559_);
  or g_115309_(_023257_, _023466_, _023560_);
  and g_115310_(_023558_, _023560_, _023562_);
  or g_115311_(_023557_, _023559_, _023563_);
  and g_115312_(_023555_, _023562_, _023564_);
  or g_115313_(_023556_, _023563_, _023565_);
  and g_115314_(_023553_, _023565_, _023566_);
  or g_115315_(_023554_, _023564_, _023567_);
  xor g_115316_(out[645], _023479_, _023568_);
  xor g_115317_(_055700_, _023479_, _023569_);
  and g_115318_(_023262_, _023466_, _023570_);
  or g_115319_(_023261_, _023467_, _023571_);
  and g_115320_(_023269_, _023467_, _023573_);
  not g_115321_(_023573_, _023574_);
  and g_115322_(_023571_, _023574_, _023575_);
  or g_115323_(_023570_, _023573_, _023576_);
  and g_115324_(_023569_, _023575_, _023577_);
  or g_115325_(_023568_, _023576_, _023578_);
  and g_115326_(_023545_, _023551_, _023579_);
  or g_115327_(_023544_, _023552_, _023580_);
  and g_115328_(_023556_, _023563_, _023581_);
  or g_115329_(_023555_, _023562_, _023582_);
  and g_115330_(_023580_, _023582_, _023584_);
  or g_115331_(_023579_, _023581_, _023585_);
  and g_115332_(_023578_, _023584_, _023586_);
  or g_115333_(_023577_, _023585_, _023587_);
  and g_115334_(_023566_, _023586_, _023588_);
  or g_115335_(_023567_, _023587_, _023589_);
  and g_115336_(_023568_, _023576_, _023590_);
  or g_115337_(_023569_, _023575_, _023591_);
  xor g_115338_(out[644], out[643], _023592_);
  xor g_115339_(_055711_, out[643], _023593_);
  and g_115340_(_023293_, _023466_, _023595_);
  not g_115341_(_023595_, _023596_);
  and g_115342_(_023301_, _023467_, _023597_);
  or g_115343_(_023300_, _023466_, _023598_);
  and g_115344_(_023596_, _023598_, _023599_);
  or g_115345_(_023595_, _023597_, _023600_);
  and g_115346_(_023593_, _023600_, _023601_);
  or g_115347_(_023592_, _023599_, _023602_);
  and g_115348_(_023591_, _023602_, _023603_);
  or g_115349_(_023590_, _023601_, _023604_);
  and g_115350_(_023592_, _023599_, _023606_);
  or g_115351_(_023593_, _023600_, _023607_);
  and g_115352_(_023603_, _023607_, _023608_);
  or g_115353_(_023604_, _023606_, _023609_);
  and g_115354_(_023588_, _023608_, _023610_);
  or g_115355_(_023589_, _023609_, _023611_);
  and g_115356_(out[627], _023466_, _023612_);
  not g_115357_(_023612_, _023613_);
  and g_115358_(_023394_, _023467_, _023614_);
  or g_115359_(_023393_, _023466_, _023615_);
  and g_115360_(_023613_, _023615_, _023617_);
  or g_115361_(_023612_, _023614_, _023618_);
  and g_115362_(out[643], _023617_, _023619_);
  or g_115363_(_055755_, _023618_, _023620_);
  or g_115364_(_023384_, _023466_, _023621_);
  not g_115365_(_023621_, _023622_);
  and g_115366_(_055612_, _023466_, _023623_);
  or g_115367_(out[626], _023467_, _023624_);
  and g_115368_(_023621_, _023624_, _023625_);
  or g_115369_(_023622_, _023623_, _023626_);
  and g_115370_(out[642], _023626_, _023628_);
  or g_115371_(_023619_, _023628_, _023629_);
  and g_115372_(_055755_, _023618_, _023630_);
  or g_115373_(out[643], _023617_, _023631_);
  and g_115374_(_055744_, _023625_, _023632_);
  or g_115375_(out[642], _023626_, _023633_);
  or g_115376_(_023630_, _023632_, _023634_);
  or g_115377_(_023629_, _023634_, _023635_);
  not g_115378_(_023635_, _023636_);
  and g_115379_(_055722_, _023470_, _023637_);
  or g_115380_(out[641], _023471_, _023639_);
  and g_115381_(_023412_, _023467_, _023640_);
  or g_115382_(_023411_, _023466_, _023641_);
  and g_115383_(_055601_, _023466_, _023642_);
  or g_115384_(out[624], _023467_, _023643_);
  and g_115385_(_023641_, _023643_, _023644_);
  or g_115386_(_023640_, _023642_, _023645_);
  and g_115387_(out[640], _023645_, _023646_);
  or g_115388_(_055733_, _023644_, _023647_);
  xor g_115389_(_055722_, _023470_, _023648_);
  xor g_115390_(out[641], _023470_, _023650_);
  and g_115391_(_023647_, _023648_, _023651_);
  or g_115392_(_023646_, _023650_, _023652_);
  and g_115393_(_023639_, _023652_, _023653_);
  or g_115394_(_023637_, _023651_, _023654_);
  and g_115395_(_023636_, _023654_, _023655_);
  or g_115396_(_023635_, _023653_, _023656_);
  and g_115397_(_023631_, _023632_, _023657_);
  or g_115398_(_023630_, _023633_, _023658_);
  and g_115399_(_023620_, _023658_, _023659_);
  or g_115400_(_023619_, _023657_, _023661_);
  and g_115401_(_023656_, _023659_, _023662_);
  or g_115402_(_023655_, _023661_, _023663_);
  and g_115403_(_023610_, _023663_, _023664_);
  or g_115404_(_023611_, _023662_, _023665_);
  and g_115405_(_023588_, _023604_, _023666_);
  or g_115406_(_023589_, _023603_, _023667_);
  or g_115407_(_023566_, _023579_, _023668_);
  not g_115408_(_023668_, _023669_);
  and g_115409_(_023667_, _023668_, _023670_);
  or g_115410_(_023666_, _023669_, _023672_);
  and g_115411_(_023665_, _023670_, _023673_);
  or g_115412_(_023664_, _023672_, _023674_);
  and g_115413_(_023542_, _023674_, _023675_);
  or g_115414_(_023543_, _023673_, _023676_);
  and g_115415_(_023510_, _023532_, _023677_);
  or g_115416_(_023509_, _023531_, _023678_);
  and g_115417_(_023535_, _023677_, _023679_);
  or g_115418_(_023536_, _023678_, _023680_);
  and g_115419_(_023499_, _023512_, _023681_);
  or g_115420_(_023498_, _023511_, _023683_);
  and g_115421_(_023680_, _023683_, _023684_);
  or g_115422_(_023679_, _023681_, _023685_);
  and g_115423_(_023676_, _023684_, _023686_);
  or g_115424_(_023675_, _023685_, _023687_);
  and g_115425_(_055733_, _023644_, _023688_);
  or g_115426_(_023635_, _023652_, _023689_);
  or g_115427_(_023688_, _023689_, _023690_);
  or g_115428_(_023543_, _023690_, _023691_);
  or g_115429_(_023611_, _023691_, _023692_);
  not g_115430_(_023692_, _023694_);
  and g_115431_(_023687_, _023692_, _023695_);
  or g_115432_(_023686_, _023694_, _023696_);
  and g_115433_(_023471_, _023696_, _023697_);
  or g_115434_(_023470_, _023695_, _023698_);
  and g_115435_(_055722_, _023695_, _023699_);
  or g_115436_(out[641], _023696_, _023700_);
  and g_115437_(_023698_, _023700_, _023701_);
  or g_115438_(_023697_, _023699_, _023702_);
  or g_115439_(_023488_, _023696_, _023703_);
  not g_115440_(_023703_, _023705_);
  and g_115441_(_023478_, _023696_, _023706_);
  not g_115442_(_023706_, _023707_);
  and g_115443_(_023703_, _023707_, _023708_);
  or g_115444_(_023705_, _023706_, _023709_);
  and g_115445_(out[660], out[659], _023710_);
  or g_115446_(out[661], _023710_, _023711_);
  or g_115447_(out[662], _023711_, _023712_);
  or g_115448_(out[663], _023712_, _023713_);
  or g_115449_(out[664], _023713_, _023714_);
  and g_115450_(out[665], _023714_, _023716_);
  or g_115451_(out[666], _023716_, _023717_);
  xor g_115452_(out[666], _023716_, _023718_);
  not g_115453_(_023718_, _023719_);
  and g_115454_(_023709_, _023719_, _023720_);
  or g_115455_(_023708_, _023718_, _023721_);
  and g_115456_(_023491_, _023493_, _023722_);
  or g_115457_(_023492_, _023494_, _023723_);
  xor g_115458_(out[667], _023717_, _023724_);
  xor g_115459_(_055799_, _023717_, _023725_);
  and g_115460_(_023722_, _023725_, _023727_);
  or g_115461_(_023723_, _023724_, _023728_);
  and g_115462_(_023723_, _023724_, _023729_);
  or g_115463_(_023722_, _023725_, _023730_);
  and g_115464_(_023708_, _023718_, _023731_);
  or g_115465_(_023709_, _023719_, _023732_);
  and g_115466_(_023721_, _023728_, _023733_);
  or g_115467_(_023720_, _023727_, _023734_);
  and g_115468_(_023730_, _023732_, _023735_);
  or g_115469_(_023729_, _023731_, _023736_);
  and g_115470_(_023733_, _023735_, _023738_);
  or g_115471_(_023734_, _023736_, _023739_);
  xor g_115472_(out[664], _023713_, _023740_);
  xor g_115473_(_055898_, _023713_, _023741_);
  or g_115474_(_023518_, _023696_, _023742_);
  not g_115475_(_023742_, _023743_);
  and g_115476_(_023525_, _023696_, _023744_);
  not g_115477_(_023744_, _023745_);
  and g_115478_(_023742_, _023745_, _023746_);
  or g_115479_(_023743_, _023744_, _023747_);
  and g_115480_(_023740_, _023747_, _023749_);
  or g_115481_(_023741_, _023746_, _023750_);
  xor g_115482_(out[665], _023714_, _023751_);
  xor g_115483_(_055909_, _023714_, _023752_);
  or g_115484_(_023501_, _023696_, _023753_);
  not g_115485_(_023753_, _023754_);
  and g_115486_(_023508_, _023696_, _023755_);
  not g_115487_(_023755_, _023756_);
  and g_115488_(_023753_, _023756_, _023757_);
  or g_115489_(_023754_, _023755_, _023758_);
  and g_115490_(_023752_, _023758_, _023760_);
  or g_115491_(_023751_, _023757_, _023761_);
  and g_115492_(_023750_, _023761_, _023762_);
  or g_115493_(_023749_, _023760_, _023763_);
  and g_115494_(_023741_, _023746_, _023764_);
  or g_115495_(_023740_, _023747_, _023765_);
  and g_115496_(_023751_, _023757_, _023766_);
  or g_115497_(_023752_, _023758_, _023767_);
  xor g_115498_(out[663], _023712_, _023768_);
  not g_115499_(_023768_, _023769_);
  or g_115500_(_023544_, _023696_, _023771_);
  or g_115501_(_023551_, _023695_, _023772_);
  and g_115502_(_023771_, _023772_, _023773_);
  not g_115503_(_023773_, _023774_);
  and g_115504_(_023769_, _023773_, _023775_);
  or g_115505_(_023768_, _023774_, _023776_);
  and g_115506_(_023767_, _023776_, _023777_);
  or g_115507_(_023766_, _023775_, _023778_);
  or g_115508_(_023764_, _023778_, _023779_);
  or g_115509_(_023763_, _023779_, _023780_);
  and g_115510_(_023762_, _023765_, _023782_);
  and g_115511_(_023738_, _023782_, _023783_);
  and g_115512_(_023777_, _023783_, _023784_);
  or g_115513_(_023739_, _023780_, _023785_);
  xor g_115514_(out[662], _023711_, _023786_);
  xor g_115515_(_055821_, _023711_, _023787_);
  or g_115516_(_023556_, _023696_, _023788_);
  not g_115517_(_023788_, _023789_);
  and g_115518_(_023563_, _023696_, _023790_);
  not g_115519_(_023790_, _023791_);
  and g_115520_(_023788_, _023791_, _023793_);
  or g_115521_(_023789_, _023790_, _023794_);
  or g_115522_(_023787_, _023794_, _023795_);
  or g_115523_(_023769_, _023773_, _023796_);
  and g_115524_(_023795_, _023796_, _023797_);
  not g_115525_(_023797_, _023798_);
  xor g_115526_(out[661], _023710_, _023799_);
  xor g_115527_(_055832_, _023710_, _023800_);
  or g_115528_(_023568_, _023696_, _023801_);
  not g_115529_(_023801_, _023802_);
  and g_115530_(_023576_, _023696_, _023804_);
  not g_115531_(_023804_, _023805_);
  and g_115532_(_023801_, _023805_, _023806_);
  or g_115533_(_023802_, _023804_, _023807_);
  or g_115534_(_023800_, _023806_, _023808_);
  xor g_115535_(out[660], out[659], _023809_);
  xor g_115536_(_055843_, out[659], _023810_);
  or g_115537_(_023593_, _023696_, _023811_);
  not g_115538_(_023811_, _023812_);
  and g_115539_(_023600_, _023696_, _023813_);
  not g_115540_(_023813_, _023815_);
  and g_115541_(_023811_, _023815_, _023816_);
  or g_115542_(_023812_, _023813_, _023817_);
  or g_115543_(_023809_, _023816_, _023818_);
  and g_115544_(_023808_, _023818_, _023819_);
  not g_115545_(_023819_, _023820_);
  or g_115546_(_055755_, _023696_, _023821_);
  not g_115547_(_023821_, _023822_);
  and g_115548_(_023618_, _023696_, _023823_);
  not g_115549_(_023823_, _023824_);
  and g_115550_(_023821_, _023824_, _023826_);
  or g_115551_(_023822_, _023823_, _023827_);
  and g_115552_(_055887_, _023827_, _023828_);
  or g_115553_(out[659], _023826_, _023829_);
  and g_115554_(_023809_, _023816_, _023830_);
  or g_115555_(_023810_, _023817_, _023831_);
  and g_115556_(_023829_, _023831_, _023832_);
  or g_115557_(_023828_, _023830_, _023833_);
  and g_115558_(out[659], _023826_, _023834_);
  not g_115559_(_023834_, _023835_);
  and g_115560_(_023626_, _023696_, _023837_);
  or g_115561_(_023625_, _023695_, _023838_);
  and g_115562_(_055744_, _023695_, _023839_);
  or g_115563_(out[642], _023696_, _023840_);
  and g_115564_(_023838_, _023840_, _023841_);
  or g_115565_(_023837_, _023839_, _023842_);
  and g_115566_(out[658], _023842_, _023843_);
  or g_115567_(_055876_, _023841_, _023844_);
  and g_115568_(_023645_, _023696_, _023845_);
  or g_115569_(_023644_, _023695_, _023846_);
  and g_115570_(_055733_, _023695_, _023848_);
  or g_115571_(out[640], _023696_, _023849_);
  and g_115572_(_023846_, _023849_, _023850_);
  or g_115573_(_023845_, _023848_, _023851_);
  and g_115574_(out[656], _023851_, _023852_);
  or g_115575_(_055865_, _023850_, _023853_);
  and g_115576_(out[657], _023702_, _023854_);
  or g_115577_(_055854_, _023701_, _023855_);
  and g_115578_(_023853_, _023855_, _023856_);
  or g_115579_(_023852_, _023854_, _023857_);
  and g_115580_(_055876_, _023841_, _023859_);
  or g_115581_(out[658], _023842_, _023860_);
  and g_115582_(_055854_, _023701_, _023861_);
  or g_115583_(out[657], _023702_, _023862_);
  and g_115584_(_023860_, _023862_, _023863_);
  or g_115585_(_023859_, _023861_, _023864_);
  and g_115586_(_023857_, _023863_, _023865_);
  or g_115587_(_023856_, _023864_, _023866_);
  and g_115588_(_023844_, _023866_, _023867_);
  or g_115589_(_023843_, _023865_, _023868_);
  and g_115590_(_023835_, _023868_, _023870_);
  or g_115591_(_023834_, _023867_, _023871_);
  and g_115592_(_023832_, _023871_, _023872_);
  or g_115593_(_023833_, _023870_, _023873_);
  and g_115594_(_023819_, _023873_, _023874_);
  or g_115595_(_023820_, _023872_, _023875_);
  or g_115596_(_023786_, _023793_, _023876_);
  or g_115597_(_023799_, _023807_, _023877_);
  and g_115598_(_023876_, _023877_, _023878_);
  not g_115599_(_023878_, _023879_);
  and g_115600_(_023875_, _023878_, _023881_);
  or g_115601_(_023874_, _023879_, _023882_);
  and g_115602_(_023797_, _023882_, _023883_);
  or g_115603_(_023798_, _023881_, _023884_);
  and g_115604_(_023784_, _023884_, _023885_);
  or g_115605_(_023785_, _023883_, _023886_);
  and g_115606_(_023763_, _023767_, _023887_);
  or g_115607_(_023762_, _023766_, _023888_);
  and g_115608_(_023738_, _023887_, _023889_);
  or g_115609_(_023739_, _023888_, _023890_);
  and g_115610_(_023730_, _023731_, _023892_);
  or g_115611_(_023729_, _023732_, _023893_);
  and g_115612_(_023728_, _023893_, _023894_);
  or g_115613_(_023727_, _023892_, _023895_);
  and g_115614_(_023890_, _023894_, _023896_);
  or g_115615_(_023889_, _023895_, _023897_);
  and g_115616_(_023886_, _023896_, _023898_);
  or g_115617_(_023885_, _023897_, _023899_);
  and g_115618_(_055865_, _023850_, _023900_);
  or g_115619_(out[656], _023851_, _023901_);
  and g_115620_(_023819_, _023878_, _023903_);
  and g_115621_(_023797_, _023856_, _023904_);
  and g_115622_(_023903_, _023904_, _023905_);
  not g_115623_(_023905_, _023906_);
  or g_115624_(_023834_, _023864_, _023907_);
  not g_115625_(_023907_, _023908_);
  and g_115626_(_023844_, _023901_, _023909_);
  or g_115627_(_023843_, _023900_, _023910_);
  and g_115628_(_023832_, _023909_, _023911_);
  or g_115629_(_023833_, _023910_, _023912_);
  and g_115630_(_023908_, _023911_, _023914_);
  or g_115631_(_023907_, _023912_, _023915_);
  and g_115632_(_023905_, _023914_, _023916_);
  or g_115633_(_023906_, _023915_, _023917_);
  and g_115634_(_023784_, _023916_, _023918_);
  or g_115635_(_023785_, _023917_, _023919_);
  and g_115636_(_023899_, _023919_, _023920_);
  or g_115637_(_023898_, _023918_, _023921_);
  or g_115638_(_023701_, _023920_, _023922_);
  or g_115639_(out[657], _023921_, _023923_);
  and g_115640_(_023922_, _023923_, _023925_);
  not g_115641_(_023925_, _023926_);
  and g_115642_(_023709_, _023921_, _023927_);
  or g_115643_(_023708_, _023920_, _023928_);
  and g_115644_(_023718_, _023920_, _023929_);
  or g_115645_(_023719_, _023921_, _023930_);
  and g_115646_(_023928_, _023930_, _023931_);
  or g_115647_(_023927_, _023929_, _023932_);
  and g_115648_(out[676], out[675], _023933_);
  or g_115649_(out[677], _023933_, _023934_);
  or g_115650_(out[678], _023934_, _023936_);
  or g_115651_(out[679], _023936_, _023937_);
  or g_115652_(out[680], _023937_, _023938_);
  and g_115653_(out[681], _023938_, _023939_);
  or g_115654_(out[682], _023939_, _023940_);
  xor g_115655_(out[682], _023939_, _023941_);
  xor g_115656_(_000087_, _023939_, _023942_);
  and g_115657_(_023931_, _023941_, _023943_);
  or g_115658_(_023932_, _023942_, _023944_);
  and g_115659_(_023722_, _023724_, _023945_);
  or g_115660_(_023723_, _023725_, _023947_);
  xor g_115661_(out[683], _023940_, _023948_);
  xor g_115662_(_055931_, _023940_, _023949_);
  and g_115663_(_023945_, _023949_, _023950_);
  or g_115664_(_023947_, _023948_, _023951_);
  and g_115665_(_023944_, _023951_, _023952_);
  or g_115666_(_023943_, _023950_, _023953_);
  and g_115667_(_023932_, _023942_, _023954_);
  or g_115668_(_023931_, _023941_, _023955_);
  and g_115669_(_023947_, _023948_, _023956_);
  or g_115670_(_023945_, _023949_, _023958_);
  and g_115671_(_023955_, _023958_, _023959_);
  or g_115672_(_023954_, _023956_, _023960_);
  and g_115673_(_023952_, _023959_, _023961_);
  or g_115674_(_023953_, _023960_, _023962_);
  xor g_115675_(out[681], _023938_, _023963_);
  xor g_115676_(_000076_, _023938_, _023964_);
  and g_115677_(_023758_, _023921_, _023965_);
  or g_115678_(_023757_, _023920_, _023966_);
  and g_115679_(_023751_, _023920_, _023967_);
  or g_115680_(_023752_, _023921_, _023969_);
  and g_115681_(_023966_, _023969_, _023970_);
  or g_115682_(_023965_, _023967_, _023971_);
  and g_115683_(_023964_, _023971_, _023972_);
  or g_115684_(_023963_, _023970_, _023973_);
  xor g_115685_(out[680], _023937_, _023974_);
  not g_115686_(_023974_, _023975_);
  and g_115687_(_023747_, _023921_, _023976_);
  or g_115688_(_023746_, _023920_, _023977_);
  and g_115689_(_023741_, _023920_, _023978_);
  or g_115690_(_023740_, _023921_, _023980_);
  and g_115691_(_023977_, _023980_, _023981_);
  or g_115692_(_023976_, _023978_, _023982_);
  and g_115693_(_023974_, _023982_, _023983_);
  or g_115694_(_023975_, _023981_, _023984_);
  and g_115695_(_023973_, _023984_, _023985_);
  or g_115696_(_023972_, _023983_, _023986_);
  and g_115697_(_023963_, _023970_, _023987_);
  or g_115698_(_023964_, _023971_, _023988_);
  and g_115699_(_023975_, _023981_, _023989_);
  or g_115700_(_023974_, _023982_, _023991_);
  and g_115701_(_023988_, _023991_, _023992_);
  or g_115702_(_023987_, _023989_, _023993_);
  and g_115703_(_023985_, _023992_, _023994_);
  or g_115704_(_023986_, _023993_, _023995_);
  and g_115705_(_023961_, _023994_, _023996_);
  or g_115706_(_023962_, _023995_, _023997_);
  xor g_115707_(out[679], _023936_, _023998_);
  xor g_115708_(_055942_, _023936_, _023999_);
  or g_115709_(_023773_, _023920_, _024000_);
  or g_115710_(_023768_, _023921_, _024002_);
  and g_115711_(_024000_, _024002_, _024003_);
  not g_115712_(_024003_, _024004_);
  and g_115713_(_023999_, _024003_, _024005_);
  or g_115714_(_023998_, _024004_, _024006_);
  and g_115715_(_023998_, _024004_, _024007_);
  or g_115716_(_023999_, _024003_, _024008_);
  and g_115717_(_024006_, _024008_, _024009_);
  or g_115718_(_024005_, _024007_, _024010_);
  xor g_115719_(out[678], _023934_, _024011_);
  not g_115720_(_024011_, _024013_);
  and g_115721_(_023794_, _023921_, _024014_);
  or g_115722_(_023793_, _023920_, _024015_);
  and g_115723_(_023786_, _023920_, _024016_);
  or g_115724_(_023787_, _023921_, _024017_);
  and g_115725_(_024015_, _024017_, _024018_);
  or g_115726_(_024014_, _024016_, _024019_);
  and g_115727_(_024011_, _024018_, _024020_);
  or g_115728_(_024013_, _024019_, _024021_);
  xor g_115729_(_024011_, _024018_, _024022_);
  xor g_115730_(_024013_, _024018_, _024024_);
  and g_115731_(_024009_, _024022_, _024025_);
  or g_115732_(_024010_, _024024_, _024026_);
  xor g_115733_(out[677], _023933_, _024027_);
  xor g_115734_(_055964_, _023933_, _024028_);
  and g_115735_(_023807_, _023921_, _024029_);
  or g_115736_(_023806_, _023920_, _024030_);
  and g_115737_(_023800_, _023920_, _024031_);
  or g_115738_(_023799_, _023921_, _024032_);
  and g_115739_(_024030_, _024032_, _024033_);
  or g_115740_(_024029_, _024031_, _024035_);
  and g_115741_(_024027_, _024035_, _024036_);
  or g_115742_(_024028_, _024033_, _024037_);
  xor g_115743_(out[676], out[675], _024038_);
  xor g_115744_(_000010_, out[675], _024039_);
  and g_115745_(_023809_, _023920_, _024040_);
  or g_115746_(_023810_, _023921_, _024041_);
  and g_115747_(_023817_, _023921_, _024042_);
  or g_115748_(_023816_, _023920_, _024043_);
  and g_115749_(_024041_, _024043_, _024044_);
  or g_115750_(_024040_, _024042_, _024046_);
  and g_115751_(_024039_, _024046_, _024047_);
  or g_115752_(_024038_, _024044_, _024048_);
  and g_115753_(_024037_, _024048_, _024049_);
  or g_115754_(_024036_, _024047_, _024050_);
  and g_115755_(_024038_, _024044_, _024051_);
  or g_115756_(_024039_, _024046_, _024052_);
  and g_115757_(_024028_, _024033_, _024053_);
  or g_115758_(_024027_, _024035_, _024054_);
  and g_115759_(_024052_, _024054_, _024055_);
  or g_115760_(_024051_, _024053_, _024057_);
  and g_115761_(_024049_, _024055_, _024058_);
  or g_115762_(_024050_, _024057_, _024059_);
  and g_115763_(_023996_, _024058_, _024060_);
  or g_115764_(_023997_, _024059_, _024061_);
  and g_115765_(_024025_, _024060_, _024062_);
  or g_115766_(_024026_, _024061_, _024063_);
  and g_115767_(out[659], _023920_, _024064_);
  not g_115768_(_024064_, _024065_);
  or g_115769_(_023826_, _023920_, _024066_);
  not g_115770_(_024066_, _024068_);
  and g_115771_(_024065_, _024066_, _024069_);
  or g_115772_(_024064_, _024068_, _024070_);
  or g_115773_(_000054_, _024070_, _024071_);
  not g_115774_(_024071_, _024072_);
  or g_115775_(_023841_, _023920_, _024073_);
  not g_115776_(_024073_, _024074_);
  and g_115777_(_055876_, _023920_, _024075_);
  not g_115778_(_024075_, _024076_);
  and g_115779_(_024073_, _024076_, _024077_);
  or g_115780_(_024074_, _024075_, _024079_);
  and g_115781_(out[674], _024079_, _024080_);
  or g_115782_(_000043_, _024077_, _024081_);
  and g_115783_(_024071_, _024081_, _024082_);
  or g_115784_(_024072_, _024080_, _024083_);
  and g_115785_(_000054_, _024070_, _024084_);
  or g_115786_(out[675], _024069_, _024085_);
  and g_115787_(_000043_, _024077_, _024086_);
  or g_115788_(out[674], _024079_, _024087_);
  and g_115789_(_024085_, _024087_, _024088_);
  or g_115790_(_024084_, _024086_, _024090_);
  and g_115791_(_024082_, _024088_, _024091_);
  or g_115792_(_024083_, _024090_, _024092_);
  and g_115793_(_023851_, _023921_, _024093_);
  or g_115794_(_023850_, _023920_, _024094_);
  and g_115795_(_055865_, _023920_, _024095_);
  or g_115796_(out[656], _023921_, _024096_);
  and g_115797_(_024094_, _024096_, _024097_);
  or g_115798_(_024093_, _024095_, _024098_);
  and g_115799_(out[672], _024098_, _024099_);
  or g_115800_(_000032_, _024097_, _024101_);
  and g_115801_(_000021_, _023925_, _024102_);
  or g_115802_(out[673], _023926_, _024103_);
  xor g_115803_(_000021_, _023925_, _024104_);
  xor g_115804_(out[673], _023925_, _024105_);
  and g_115805_(_024101_, _024104_, _024106_);
  or g_115806_(_024099_, _024105_, _024107_);
  or g_115807_(out[672], _024098_, _024108_);
  and g_115808_(_024106_, _024108_, _024109_);
  and g_115809_(_024091_, _024109_, _024110_);
  and g_115810_(_024062_, _024110_, _024112_);
  not g_115811_(_024112_, _024113_);
  and g_115812_(_024103_, _024107_, _024114_);
  or g_115813_(_024102_, _024106_, _024115_);
  and g_115814_(_024091_, _024115_, _024116_);
  or g_115815_(_024092_, _024114_, _024117_);
  and g_115816_(_024085_, _024086_, _024118_);
  or g_115817_(_024084_, _024087_, _024119_);
  and g_115818_(_024071_, _024119_, _024120_);
  or g_115819_(_024072_, _024118_, _024121_);
  and g_115820_(_024117_, _024120_, _024123_);
  or g_115821_(_024116_, _024121_, _024124_);
  and g_115822_(_024062_, _024124_, _024125_);
  or g_115823_(_024063_, _024123_, _024126_);
  and g_115824_(_024050_, _024054_, _024127_);
  or g_115825_(_024049_, _024053_, _024128_);
  and g_115826_(_024025_, _024127_, _024129_);
  or g_115827_(_024026_, _024128_, _024130_);
  and g_115828_(_024008_, _024021_, _024131_);
  or g_115829_(_024007_, _024020_, _024132_);
  and g_115830_(_024006_, _024132_, _024134_);
  or g_115831_(_024005_, _024131_, _024135_);
  and g_115832_(_024130_, _024135_, _024136_);
  or g_115833_(_024129_, _024134_, _024137_);
  and g_115834_(_023996_, _024137_, _024138_);
  or g_115835_(_023997_, _024136_, _024139_);
  and g_115836_(_023986_, _023988_, _024140_);
  or g_115837_(_023985_, _023987_, _024141_);
  and g_115838_(_023961_, _024140_, _024142_);
  or g_115839_(_023962_, _024141_, _024143_);
  and g_115840_(_023953_, _023958_, _024145_);
  or g_115841_(_023952_, _023956_, _024146_);
  and g_115842_(_024143_, _024146_, _024147_);
  or g_115843_(_024142_, _024145_, _024148_);
  and g_115844_(_024126_, _024147_, _024149_);
  or g_115845_(_024125_, _024148_, _024150_);
  and g_115846_(_024139_, _024149_, _024151_);
  or g_115847_(_024138_, _024150_, _024152_);
  and g_115848_(_024113_, _024152_, _024153_);
  or g_115849_(_024112_, _024151_, _024154_);
  or g_115850_(_023925_, _024153_, _024156_);
  or g_115851_(out[673], _024154_, _024157_);
  and g_115852_(_024156_, _024157_, _024158_);
  and g_115853_(_023945_, _023948_, _024159_);
  or g_115854_(_023947_, _023949_, _024160_);
  and g_115855_(out[692], out[691], _024161_);
  or g_115856_(out[693], _024161_, _024162_);
  or g_115857_(out[694], _024162_, _024163_);
  or g_115858_(out[695], _024163_, _024164_);
  or g_115859_(out[696], _024164_, _024165_);
  and g_115860_(out[697], _024165_, _024167_);
  or g_115861_(out[698], _024167_, _024168_);
  xor g_115862_(out[699], _024168_, _024169_);
  xor g_115863_(_000098_, _024168_, _024170_);
  or g_115864_(_024159_, _024170_, _024171_);
  and g_115865_(_023941_, _024153_, _024172_);
  or g_115866_(_023942_, _024154_, _024173_);
  and g_115867_(_023932_, _024154_, _024174_);
  or g_115868_(_023931_, _024153_, _024175_);
  and g_115869_(_024173_, _024175_, _024176_);
  or g_115870_(_024172_, _024174_, _024178_);
  xor g_115871_(out[698], _024167_, _024179_);
  xor g_115872_(_000219_, _024167_, _024180_);
  and g_115873_(_024176_, _024179_, _024181_);
  or g_115874_(_024178_, _024180_, _024182_);
  and g_115875_(_024159_, _024170_, _024183_);
  or g_115876_(_024160_, _024169_, _024184_);
  and g_115877_(_024182_, _024184_, _024185_);
  or g_115878_(_024181_, _024183_, _024186_);
  xor g_115879_(out[697], _024165_, _024187_);
  xor g_115880_(_000208_, _024165_, _024189_);
  or g_115881_(_023964_, _024154_, _024190_);
  not g_115882_(_024190_, _024191_);
  and g_115883_(_023971_, _024154_, _024192_);
  not g_115884_(_024192_, _024193_);
  and g_115885_(_024190_, _024193_, _024194_);
  or g_115886_(_024191_, _024192_, _024195_);
  and g_115887_(_024189_, _024195_, _024196_);
  or g_115888_(_024187_, _024194_, _024197_);
  xor g_115889_(out[696], _024164_, _024198_);
  xor g_115890_(_000197_, _024164_, _024200_);
  or g_115891_(_023974_, _024154_, _024201_);
  not g_115892_(_024201_, _024202_);
  and g_115893_(_023982_, _024154_, _024203_);
  not g_115894_(_024203_, _024204_);
  and g_115895_(_024201_, _024204_, _024205_);
  or g_115896_(_024202_, _024203_, _024206_);
  and g_115897_(_024198_, _024206_, _024207_);
  or g_115898_(_024200_, _024205_, _024208_);
  and g_115899_(_024197_, _024208_, _024209_);
  or g_115900_(_024196_, _024207_, _024211_);
  or g_115901_(_024176_, _024179_, _024212_);
  and g_115902_(_024187_, _024194_, _024213_);
  or g_115903_(_024189_, _024195_, _024214_);
  xor g_115904_(out[695], _024163_, _024215_);
  xor g_115905_(_000109_, _024163_, _024216_);
  and g_115906_(_023999_, _024153_, _024217_);
  or g_115907_(_023998_, _024154_, _024218_);
  and g_115908_(_024004_, _024154_, _024219_);
  or g_115909_(_024003_, _024153_, _024220_);
  and g_115910_(_024218_, _024220_, _024222_);
  or g_115911_(_024217_, _024219_, _024223_);
  and g_115912_(_024215_, _024223_, _024224_);
  or g_115913_(_024216_, _024222_, _024225_);
  xor g_115914_(out[694], _024162_, _024226_);
  xor g_115915_(_000120_, _024162_, _024227_);
  and g_115916_(_024011_, _024153_, _024228_);
  or g_115917_(_024013_, _024154_, _024229_);
  and g_115918_(_024019_, _024154_, _024230_);
  or g_115919_(_024018_, _024153_, _024231_);
  and g_115920_(_024229_, _024231_, _024233_);
  or g_115921_(_024228_, _024230_, _024234_);
  and g_115922_(_024226_, _024233_, _024235_);
  or g_115923_(_024227_, _024234_, _024236_);
  xor g_115924_(out[692], out[691], _024237_);
  xor g_115925_(_000142_, out[691], _024238_);
  or g_115926_(_024039_, _024154_, _024239_);
  not g_115927_(_024239_, _024240_);
  and g_115928_(_024046_, _024154_, _024241_);
  not g_115929_(_024241_, _024242_);
  and g_115930_(_024239_, _024242_, _024244_);
  or g_115931_(_024240_, _024241_, _024245_);
  and g_115932_(_024238_, _024245_, _024246_);
  or g_115933_(_024237_, _024244_, _024247_);
  xor g_115934_(out[693], _024161_, _024248_);
  xor g_115935_(_000131_, _024161_, _024249_);
  or g_115936_(_024027_, _024154_, _024250_);
  not g_115937_(_024250_, _024251_);
  and g_115938_(_024035_, _024154_, _024252_);
  not g_115939_(_024252_, _024253_);
  and g_115940_(_024250_, _024253_, _024255_);
  or g_115941_(_024251_, _024252_, _024256_);
  and g_115942_(_024248_, _024256_, _024257_);
  or g_115943_(_024249_, _024255_, _024258_);
  and g_115944_(_024247_, _024258_, _024259_);
  or g_115945_(_024246_, _024257_, _024260_);
  or g_115946_(_000054_, _024154_, _024261_);
  or g_115947_(_024069_, _024153_, _024262_);
  and g_115948_(_024261_, _024262_, _024263_);
  and g_115949_(out[691], _024263_, _024264_);
  or g_115950_(out[691], _024263_, _024266_);
  xor g_115951_(out[691], _024263_, _024267_);
  xor g_115952_(_000186_, _024263_, _024268_);
  or g_115953_(_024077_, _024153_, _024269_);
  or g_115954_(out[674], _024154_, _024270_);
  and g_115955_(_024269_, _024270_, _024271_);
  and g_115956_(_000175_, _024271_, _024272_);
  xor g_115957_(_000175_, _024271_, _024273_);
  xor g_115958_(out[690], _024271_, _024274_);
  and g_115959_(_024267_, _024273_, _024275_);
  or g_115960_(_024268_, _024274_, _024277_);
  and g_115961_(_000153_, _024158_, _024278_);
  and g_115962_(_024098_, _024154_, _024279_);
  not g_115963_(_024279_, _024280_);
  or g_115964_(out[672], _024154_, _024281_);
  not g_115965_(_024281_, _024282_);
  and g_115966_(_024280_, _024281_, _024283_);
  or g_115967_(_024279_, _024282_, _024284_);
  and g_115968_(out[688], _024284_, _024285_);
  or g_115969_(_000164_, _024283_, _024286_);
  or g_115970_(_000153_, _024158_, _024288_);
  and g_115971_(_024286_, _024288_, _024289_);
  xor g_115972_(out[689], _024158_, _024290_);
  or g_115973_(_024285_, _024290_, _024291_);
  or g_115974_(_024278_, _024289_, _024292_);
  and g_115975_(_024275_, _024292_, _024293_);
  and g_115976_(_024266_, _024272_, _024294_);
  or g_115977_(_024264_, _024294_, _024295_);
  or g_115978_(_024293_, _024295_, _024296_);
  and g_115979_(_024237_, _024244_, _024297_);
  or g_115980_(_024238_, _024245_, _024299_);
  and g_115981_(_024249_, _024255_, _024300_);
  or g_115982_(_024248_, _024256_, _024301_);
  and g_115983_(_024227_, _024234_, _024302_);
  or g_115984_(_024226_, _024233_, _024303_);
  and g_115985_(_024200_, _024205_, _024304_);
  or g_115986_(_024198_, _024206_, _024305_);
  and g_115987_(_024209_, _024305_, _024306_);
  or g_115988_(_024211_, _024304_, _024307_);
  and g_115989_(_024171_, _024212_, _024308_);
  not g_115990_(_024308_, _024310_);
  and g_115991_(_024185_, _024308_, _024311_);
  or g_115992_(_024186_, _024310_, _024312_);
  and g_115993_(_024214_, _024311_, _024313_);
  or g_115994_(_024213_, _024312_, _024314_);
  and g_115995_(_024306_, _024313_, _024315_);
  or g_115996_(_024307_, _024314_, _024316_);
  and g_115997_(_024216_, _024222_, _024317_);
  or g_115998_(_024215_, _024223_, _024318_);
  and g_115999_(_024235_, _024318_, _024319_);
  or g_116000_(_024236_, _024317_, _024321_);
  and g_116001_(_024236_, _024318_, _024322_);
  or g_116002_(_024235_, _024317_, _024323_);
  and g_116003_(_024225_, _024303_, _024324_);
  or g_116004_(_024224_, _024302_, _024325_);
  and g_116005_(_024322_, _024324_, _024326_);
  or g_116006_(_024323_, _024325_, _024327_);
  and g_116007_(_024260_, _024326_, _024328_);
  or g_116008_(_024259_, _024327_, _024329_);
  and g_116009_(_024301_, _024328_, _024330_);
  or g_116010_(_024300_, _024329_, _024332_);
  and g_116011_(_024321_, _024332_, _024333_);
  or g_116012_(_024319_, _024330_, _024334_);
  and g_116013_(_024225_, _024333_, _024335_);
  or g_116014_(_024224_, _024334_, _024336_);
  and g_116015_(_024315_, _024336_, _024337_);
  or g_116016_(_024316_, _024335_, _024338_);
  or g_116017_(_024209_, _024314_, _024339_);
  not g_116018_(_024339_, _024340_);
  and g_116019_(_024338_, _024339_, _024341_);
  or g_116020_(_024337_, _024340_, _024343_);
  and g_116021_(_024171_, _024186_, _024344_);
  and g_116022_(_024299_, _024301_, _024345_);
  or g_116023_(_024297_, _024300_, _024346_);
  and g_116024_(_024259_, _024326_, _024347_);
  or g_116025_(_024260_, _024327_, _024348_);
  and g_116026_(_024345_, _024347_, _024349_);
  or g_116027_(_024346_, _024348_, _024350_);
  and g_116028_(_024315_, _024349_, _024351_);
  or g_116029_(_024316_, _024350_, _024352_);
  and g_116030_(_024296_, _024351_, _024354_);
  or g_116031_(_024344_, _024354_, _024355_);
  not g_116032_(_024355_, _024356_);
  and g_116033_(_024341_, _024356_, _024357_);
  or g_116034_(_024343_, _024355_, _024358_);
  and g_116035_(_000164_, _024283_, _024359_);
  or g_116036_(out[688], _024284_, _024360_);
  or g_116037_(_024277_, _024291_, _024361_);
  or g_116038_(_024352_, _024361_, _024362_);
  not g_116039_(_024362_, _024363_);
  and g_116040_(_024360_, _024363_, _024365_);
  or g_116041_(_024359_, _024362_, _024366_);
  and g_116042_(_024358_, _024366_, _024367_);
  or g_116043_(_024357_, _024365_, _024368_);
  or g_116044_(_024158_, _024367_, _024369_);
  or g_116045_(out[689], _024368_, _024370_);
  and g_116046_(_024369_, _024370_, _024371_);
  and g_116047_(_024159_, _024169_, _024372_);
  or g_116048_(_024160_, _024170_, _024373_);
  and g_116049_(out[708], out[707], _024374_);
  or g_116050_(out[709], _024374_, _024376_);
  or g_116051_(out[710], _024376_, _024377_);
  or g_116052_(out[711], _024377_, _024378_);
  or g_116053_(out[712], _024378_, _024379_);
  and g_116054_(out[713], _024379_, _024380_);
  or g_116055_(out[714], _024380_, _024381_);
  xor g_116056_(out[715], _024381_, _024382_);
  xor g_116057_(_000230_, _024381_, _024383_);
  and g_116058_(_024372_, _024383_, _024384_);
  xor g_116059_(out[714], _024380_, _024385_);
  and g_116060_(_024179_, _024367_, _024387_);
  or g_116061_(_024180_, _024368_, _024388_);
  and g_116062_(_024178_, _024368_, _024389_);
  or g_116063_(_024176_, _024367_, _024390_);
  and g_116064_(_024388_, _024390_, _024391_);
  or g_116065_(_024387_, _024389_, _024392_);
  and g_116066_(_024385_, _024391_, _024393_);
  or g_116067_(_024384_, _024393_, _024394_);
  not g_116068_(_024394_, _024395_);
  or g_116069_(_024385_, _024391_, _024396_);
  or g_116070_(_024372_, _024383_, _024398_);
  xor g_116071_(out[713], _024379_, _024399_);
  not g_116072_(_024399_, _024400_);
  and g_116073_(_024187_, _024367_, _024401_);
  or g_116074_(_024189_, _024368_, _024402_);
  and g_116075_(_024195_, _024368_, _024403_);
  or g_116076_(_024194_, _024367_, _024404_);
  and g_116077_(_024402_, _024404_, _024405_);
  or g_116078_(_024401_, _024403_, _024406_);
  or g_116079_(_024400_, _024406_, _024407_);
  and g_116080_(_024398_, _024407_, _024409_);
  and g_116081_(_024396_, _024409_, _024410_);
  and g_116082_(_024395_, _024410_, _024411_);
  not g_116083_(_024411_, _024412_);
  and g_116084_(_024400_, _024406_, _024413_);
  xor g_116085_(out[712], _024378_, _024414_);
  not g_116086_(_024414_, _024415_);
  and g_116087_(_024200_, _024367_, _024416_);
  or g_116088_(_024198_, _024368_, _024417_);
  and g_116089_(_024206_, _024368_, _024418_);
  or g_116090_(_024205_, _024367_, _024420_);
  and g_116091_(_024417_, _024420_, _024421_);
  or g_116092_(_024416_, _024418_, _024422_);
  and g_116093_(_024414_, _024422_, _024423_);
  or g_116094_(_024413_, _024423_, _024424_);
  not g_116095_(_024424_, _024425_);
  and g_116096_(_024415_, _024421_, _024426_);
  or g_116097_(_024414_, _024422_, _024427_);
  and g_116098_(_024425_, _024427_, _024428_);
  or g_116099_(_024424_, _024426_, _024429_);
  and g_116100_(_024411_, _024428_, _024431_);
  or g_116101_(_024412_, _024429_, _024432_);
  xor g_116102_(out[710], _024376_, _024433_);
  and g_116103_(_024226_, _024367_, _024434_);
  or g_116104_(_024227_, _024368_, _024435_);
  and g_116105_(_024234_, _024368_, _024436_);
  or g_116106_(_024233_, _024367_, _024437_);
  and g_116107_(_024435_, _024437_, _024438_);
  or g_116108_(_024434_, _024436_, _024439_);
  and g_116109_(_024433_, _024438_, _024440_);
  xor g_116110_(out[711], _024377_, _024442_);
  and g_116111_(_024216_, _024367_, _024443_);
  or g_116112_(_024215_, _024368_, _024444_);
  and g_116113_(_024223_, _024368_, _024445_);
  or g_116114_(_024222_, _024367_, _024446_);
  and g_116115_(_024444_, _024446_, _024447_);
  or g_116116_(_024443_, _024445_, _024448_);
  and g_116117_(_024442_, _024448_, _024449_);
  or g_116118_(_024440_, _024449_, _024450_);
  or g_116119_(_024442_, _024448_, _024451_);
  not g_116120_(_024451_, _024453_);
  xor g_116121_(out[708], out[707], _024454_);
  not g_116122_(_024454_, _024455_);
  and g_116123_(_024237_, _024367_, _024456_);
  or g_116124_(_024238_, _024368_, _024457_);
  and g_116125_(_024245_, _024368_, _024458_);
  or g_116126_(_024244_, _024367_, _024459_);
  and g_116127_(_024457_, _024459_, _024460_);
  or g_116128_(_024456_, _024458_, _024461_);
  and g_116129_(_024454_, _024460_, _024462_);
  or g_116130_(_024453_, _024462_, _024464_);
  or g_116131_(_024450_, _024464_, _024465_);
  not g_116132_(_024465_, _024466_);
  and g_116133_(_024455_, _024461_, _024467_);
  xor g_116134_(out[709], _024374_, _024468_);
  and g_116135_(_024249_, _024367_, _024469_);
  or g_116136_(_024248_, _024368_, _024470_);
  and g_116137_(_024256_, _024368_, _024471_);
  or g_116138_(_024255_, _024367_, _024472_);
  and g_116139_(_024470_, _024472_, _024473_);
  or g_116140_(_024469_, _024471_, _024475_);
  and g_116141_(_024468_, _024475_, _024476_);
  or g_116142_(_024467_, _024476_, _024477_);
  not g_116143_(_024477_, _024478_);
  or g_116144_(_024433_, _024438_, _024479_);
  or g_116145_(_024468_, _024475_, _024480_);
  and g_116146_(_024479_, _024480_, _024481_);
  not g_116147_(_024481_, _024482_);
  and g_116148_(_024478_, _024481_, _024483_);
  or g_116149_(_024477_, _024482_, _024484_);
  and g_116150_(_024466_, _024483_, _024486_);
  or g_116151_(_024465_, _024484_, _024487_);
  or g_116152_(_024271_, _024367_, _024488_);
  or g_116153_(out[690], _024368_, _024489_);
  and g_116154_(_024488_, _024489_, _024490_);
  and g_116155_(_000307_, _024490_, _024491_);
  or g_116156_(_000186_, _024368_, _024492_);
  or g_116157_(_024263_, _024367_, _024493_);
  and g_116158_(_024492_, _024493_, _024494_);
  and g_116159_(out[707], _024494_, _024495_);
  or g_116160_(out[707], _024494_, _024497_);
  xor g_116161_(out[707], _024494_, _024498_);
  xor g_116162_(_000318_, _024494_, _024499_);
  xor g_116163_(_000307_, _024490_, _024500_);
  xor g_116164_(out[706], _024490_, _024501_);
  and g_116165_(_024498_, _024500_, _024502_);
  or g_116166_(_024499_, _024501_, _024503_);
  and g_116167_(_000285_, _024371_, _024504_);
  or g_116168_(_024283_, _024367_, _024505_);
  or g_116169_(out[688], _024368_, _024506_);
  and g_116170_(_024505_, _024506_, _024508_);
  not g_116171_(_024508_, _024509_);
  and g_116172_(out[704], _024509_, _024510_);
  or g_116173_(_000296_, _024508_, _024511_);
  xor g_116174_(_000285_, _024371_, _024512_);
  xor g_116175_(out[705], _024371_, _024513_);
  and g_116176_(_024511_, _024512_, _024514_);
  or g_116177_(_024510_, _024513_, _024515_);
  or g_116178_(_024504_, _024514_, _024516_);
  and g_116179_(_024502_, _024516_, _024517_);
  and g_116180_(_024491_, _024497_, _024519_);
  or g_116181_(_024495_, _024519_, _024520_);
  or g_116182_(_024517_, _024520_, _024521_);
  and g_116183_(_024486_, _024521_, _024522_);
  and g_116184_(_024477_, _024481_, _024523_);
  or g_116185_(_024450_, _024523_, _024524_);
  and g_116186_(_024451_, _024524_, _024525_);
  or g_116187_(_024522_, _024525_, _024526_);
  and g_116188_(_024431_, _024526_, _024527_);
  and g_116189_(_024394_, _024398_, _024528_);
  and g_116190_(_024411_, _024424_, _024530_);
  or g_116191_(_024528_, _024530_, _024531_);
  or g_116192_(_024527_, _024531_, _024532_);
  and g_116193_(_000296_, _024508_, _024533_);
  or g_116194_(_024503_, _024533_, _024534_);
  or g_116195_(_024515_, _024534_, _024535_);
  or g_116196_(_024487_, _024535_, _024536_);
  or g_116197_(_024432_, _024536_, _024537_);
  and g_116198_(_024532_, _024537_, _024538_);
  not g_116199_(_024538_, _024539_);
  or g_116200_(_024371_, _024538_, _024541_);
  not g_116201_(_024541_, _024542_);
  and g_116202_(_000285_, _024538_, _024543_);
  or g_116203_(out[705], _024539_, _024544_);
  and g_116204_(_024541_, _024544_, _024545_);
  or g_116205_(_024542_, _024543_, _024546_);
  and g_116206_(_024392_, _024539_, _024547_);
  or g_116207_(_024391_, _024538_, _024548_);
  and g_116208_(_024385_, _024538_, _024549_);
  not g_116209_(_024549_, _024550_);
  and g_116210_(_024548_, _024550_, _024552_);
  or g_116211_(_024547_, _024549_, _024553_);
  and g_116212_(out[724], out[723], _024554_);
  or g_116213_(out[725], _024554_, _024555_);
  or g_116214_(out[726], _024555_, _024556_);
  or g_116215_(out[727], _024556_, _024557_);
  or g_116216_(out[728], _024557_, _024558_);
  and g_116217_(out[729], _024558_, _024559_);
  or g_116218_(out[730], _024559_, _024560_);
  xor g_116219_(out[730], _024559_, _024561_);
  xor g_116220_(_000483_, _024559_, _024563_);
  and g_116221_(_024552_, _024561_, _024564_);
  or g_116222_(_024553_, _024563_, _024565_);
  and g_116223_(_024372_, _024382_, _024566_);
  or g_116224_(_024373_, _024383_, _024567_);
  xor g_116225_(out[731], _024560_, _024568_);
  xor g_116226_(_000362_, _024560_, _024569_);
  and g_116227_(_024566_, _024569_, _024570_);
  or g_116228_(_024567_, _024568_, _024571_);
  and g_116229_(_024565_, _024571_, _024572_);
  or g_116230_(_024564_, _024570_, _024574_);
  and g_116231_(_024567_, _024568_, _024575_);
  or g_116232_(_024566_, _024569_, _024576_);
  and g_116233_(_024553_, _024563_, _024577_);
  or g_116234_(_024552_, _024561_, _024578_);
  and g_116235_(_024576_, _024578_, _024579_);
  or g_116236_(_024575_, _024577_, _024580_);
  xor g_116237_(out[729], _024558_, _024581_);
  xor g_116238_(_000472_, _024558_, _024582_);
  and g_116239_(_024406_, _024539_, _024583_);
  or g_116240_(_024405_, _024538_, _024585_);
  and g_116241_(_024399_, _024538_, _024586_);
  not g_116242_(_024586_, _024587_);
  and g_116243_(_024585_, _024587_, _024588_);
  or g_116244_(_024583_, _024586_, _024589_);
  and g_116245_(_024581_, _024588_, _024590_);
  or g_116246_(_024582_, _024589_, _024591_);
  and g_116247_(_024572_, _024579_, _024592_);
  or g_116248_(_024574_, _024580_, _024593_);
  and g_116249_(_024591_, _024592_, _024594_);
  or g_116250_(_024590_, _024593_, _024596_);
  and g_116251_(_024582_, _024589_, _024597_);
  or g_116252_(_024581_, _024588_, _024598_);
  xor g_116253_(out[728], _024557_, _024599_);
  xor g_116254_(_000461_, _024557_, _024600_);
  and g_116255_(_024414_, _024538_, _024601_);
  not g_116256_(_024601_, _024602_);
  and g_116257_(_024421_, _024539_, _024603_);
  or g_116258_(_024422_, _024538_, _024604_);
  or g_116259_(_024601_, _024603_, _024605_);
  and g_116260_(_024602_, _024604_, _024607_);
  and g_116261_(_024599_, _024607_, _024608_);
  or g_116262_(_024600_, _024605_, _024609_);
  and g_116263_(_024598_, _024609_, _024610_);
  or g_116264_(_024597_, _024608_, _024611_);
  and g_116265_(_024600_, _024605_, _024612_);
  or g_116266_(_024599_, _024607_, _024613_);
  and g_116267_(_024610_, _024613_, _024614_);
  or g_116268_(_024611_, _024612_, _024615_);
  and g_116269_(_024594_, _024614_, _024616_);
  or g_116270_(_024596_, _024615_, _024618_);
  xor g_116271_(out[727], _024556_, _024619_);
  xor g_116272_(_000373_, _024556_, _024620_);
  and g_116273_(_024442_, _024538_, _024621_);
  not g_116274_(_024621_, _024622_);
  and g_116275_(_024447_, _024539_, _024623_);
  or g_116276_(_024448_, _024538_, _024624_);
  or g_116277_(_024621_, _024623_, _024625_);
  and g_116278_(_024622_, _024624_, _024626_);
  and g_116279_(_024619_, _024626_, _024627_);
  or g_116280_(_024620_, _024625_, _024629_);
  xor g_116281_(out[726], _024555_, _024630_);
  xor g_116282_(_000384_, _024555_, _024631_);
  and g_116283_(_024439_, _024539_, _024632_);
  or g_116284_(_024438_, _024538_, _024633_);
  and g_116285_(_024433_, _024538_, _024634_);
  not g_116286_(_024634_, _024635_);
  and g_116287_(_024633_, _024635_, _024636_);
  or g_116288_(_024632_, _024634_, _024637_);
  and g_116289_(_024630_, _024636_, _024638_);
  or g_116290_(_024631_, _024637_, _024640_);
  and g_116291_(_024629_, _024640_, _024641_);
  or g_116292_(_024627_, _024638_, _024642_);
  and g_116293_(_024631_, _024637_, _024643_);
  or g_116294_(_024630_, _024636_, _024644_);
  and g_116295_(_024620_, _024625_, _024645_);
  or g_116296_(_024619_, _024626_, _024646_);
  xor g_116297_(out[725], _024554_, _024647_);
  xor g_116298_(_000395_, _024554_, _024648_);
  and g_116299_(_024468_, _024538_, _024649_);
  not g_116300_(_024649_, _024651_);
  and g_116301_(_024473_, _024539_, _024652_);
  or g_116302_(_024475_, _024538_, _024653_);
  or g_116303_(_024649_, _024652_, _024654_);
  and g_116304_(_024651_, _024653_, _024655_);
  and g_116305_(_024648_, _024654_, _024656_);
  or g_116306_(_024647_, _024655_, _024657_);
  and g_116307_(_024646_, _024657_, _024658_);
  or g_116308_(_024645_, _024656_, _024659_);
  and g_116309_(_024644_, _024658_, _024660_);
  or g_116310_(_024643_, _024659_, _024662_);
  and g_116311_(_024641_, _024660_, _024663_);
  or g_116312_(_024642_, _024662_, _024664_);
  xor g_116313_(out[724], out[723], _024665_);
  xor g_116314_(_000406_, out[723], _024666_);
  and g_116315_(_024454_, _024538_, _024667_);
  not g_116316_(_024667_, _024668_);
  and g_116317_(_024461_, _024539_, _024669_);
  or g_116318_(_024460_, _024538_, _024670_);
  and g_116319_(_024668_, _024670_, _024671_);
  or g_116320_(_024667_, _024669_, _024673_);
  and g_116321_(_024665_, _024671_, _024674_);
  or g_116322_(_024666_, _024673_, _024675_);
  and g_116323_(_024647_, _024655_, _024676_);
  or g_116324_(_024648_, _024654_, _024677_);
  and g_116325_(_024666_, _024673_, _024678_);
  or g_116326_(_024665_, _024671_, _024679_);
  and g_116327_(_024677_, _024679_, _024680_);
  or g_116328_(_024676_, _024678_, _024681_);
  and g_116329_(_024675_, _024680_, _024682_);
  or g_116330_(_024674_, _024681_, _024684_);
  and g_116331_(_024663_, _024682_, _024685_);
  or g_116332_(_024664_, _024684_, _024686_);
  or g_116333_(_024490_, _024538_, _024687_);
  not g_116334_(_024687_, _024688_);
  and g_116335_(_000307_, _024538_, _024689_);
  or g_116336_(out[706], _024539_, _024690_);
  and g_116337_(_024687_, _024690_, _024691_);
  or g_116338_(_024688_, _024689_, _024692_);
  and g_116339_(_000439_, _024691_, _024693_);
  and g_116340_(out[707], _024538_, _024695_);
  not g_116341_(_024695_, _024696_);
  or g_116342_(_024494_, _024538_, _024697_);
  not g_116343_(_024697_, _024698_);
  and g_116344_(_024696_, _024697_, _024699_);
  or g_116345_(_024695_, _024698_, _024700_);
  and g_116346_(out[723], _024699_, _024701_);
  or g_116347_(out[723], _024699_, _024702_);
  xor g_116348_(out[723], _024699_, _024703_);
  xor g_116349_(_000450_, _024699_, _024704_);
  xor g_116350_(_000439_, _024691_, _024706_);
  xor g_116351_(out[722], _024691_, _024707_);
  and g_116352_(_024703_, _024706_, _024708_);
  or g_116353_(_024704_, _024707_, _024709_);
  and g_116354_(_000417_, _024545_, _024710_);
  or g_116355_(out[721], _024546_, _024711_);
  or g_116356_(_024508_, _024538_, _024712_);
  not g_116357_(_024712_, _024713_);
  and g_116358_(_000296_, _024538_, _024714_);
  or g_116359_(out[704], _024539_, _024715_);
  and g_116360_(_024712_, _024715_, _024717_);
  or g_116361_(_024713_, _024714_, _024718_);
  and g_116362_(out[720], _024718_, _024719_);
  or g_116363_(_000428_, _024717_, _024720_);
  xor g_116364_(_000417_, _024545_, _024721_);
  xor g_116365_(out[721], _024545_, _024722_);
  and g_116366_(_024720_, _024721_, _024723_);
  or g_116367_(_024719_, _024722_, _024724_);
  and g_116368_(_024711_, _024724_, _024725_);
  or g_116369_(_024710_, _024723_, _024726_);
  and g_116370_(_024708_, _024726_, _024728_);
  or g_116371_(_024709_, _024725_, _024729_);
  and g_116372_(_024693_, _024702_, _024730_);
  or g_116373_(_024701_, _024730_, _024731_);
  not g_116374_(_024731_, _024732_);
  and g_116375_(_024729_, _024732_, _024733_);
  or g_116376_(_024728_, _024731_, _024734_);
  and g_116377_(_024685_, _024734_, _024735_);
  or g_116378_(_024686_, _024733_, _024736_);
  and g_116379_(_024642_, _024646_, _024737_);
  or g_116380_(_024641_, _024645_, _024739_);
  and g_116381_(_024663_, _024681_, _024740_);
  or g_116382_(_024664_, _024680_, _024741_);
  and g_116383_(_024739_, _024741_, _024742_);
  or g_116384_(_024737_, _024740_, _024743_);
  and g_116385_(_024736_, _024742_, _024744_);
  or g_116386_(_024735_, _024743_, _024745_);
  and g_116387_(_024616_, _024745_, _024746_);
  or g_116388_(_024618_, _024744_, _024747_);
  and g_116389_(_024594_, _024611_, _024748_);
  or g_116390_(_024596_, _024610_, _024750_);
  and g_116391_(_024574_, _024576_, _024751_);
  or g_116392_(_024572_, _024575_, _024752_);
  and g_116393_(_024750_, _024752_, _024753_);
  or g_116394_(_024748_, _024751_, _024754_);
  and g_116395_(_024747_, _024753_, _024755_);
  or g_116396_(_024746_, _024754_, _024756_);
  and g_116397_(_000428_, _024717_, _024757_);
  or g_116398_(out[720], _024718_, _024758_);
  and g_116399_(_024708_, _024723_, _024759_);
  or g_116400_(_024709_, _024724_, _024761_);
  and g_116401_(_024758_, _024759_, _024762_);
  or g_116402_(_024757_, _024761_, _024763_);
  and g_116403_(_024616_, _024762_, _024764_);
  or g_116404_(_024618_, _024763_, _024765_);
  and g_116405_(_024685_, _024764_, _024766_);
  or g_116406_(_024686_, _024765_, _024767_);
  and g_116407_(_024756_, _024767_, _024768_);
  or g_116408_(_024755_, _024766_, _024769_);
  and g_116409_(_024546_, _024769_, _024770_);
  not g_116410_(_024770_, _024772_);
  or g_116411_(out[721], _024769_, _024773_);
  not g_116412_(_024773_, _024774_);
  and g_116413_(_024772_, _024773_, _024775_);
  or g_116414_(_024770_, _024774_, _024776_);
  and g_116415_(_024566_, _024568_, _024777_);
  or g_116416_(_024567_, _024569_, _024778_);
  and g_116417_(out[740], out[739], _024779_);
  or g_116418_(out[741], _024779_, _024780_);
  or g_116419_(out[742], _024780_, _024781_);
  or g_116420_(out[743], _024781_, _024783_);
  or g_116421_(out[744], _024783_, _024784_);
  and g_116422_(out[745], _024784_, _024785_);
  or g_116423_(out[746], _024785_, _024786_);
  xor g_116424_(out[747], _024786_, _024787_);
  xor g_116425_(_000494_, _024786_, _024788_);
  and g_116426_(_024778_, _024787_, _024789_);
  or g_116427_(_024777_, _024788_, _024790_);
  and g_116428_(_024553_, _024769_, _024791_);
  and g_116429_(_024561_, _024768_, _024792_);
  or g_116430_(_024791_, _024792_, _024794_);
  not g_116431_(_024794_, _024795_);
  xor g_116432_(out[746], _024785_, _024796_);
  xor g_116433_(_000615_, _024785_, _024797_);
  and g_116434_(_024795_, _024796_, _024798_);
  or g_116435_(_024794_, _024797_, _024799_);
  and g_116436_(_024777_, _024788_, _024800_);
  or g_116437_(_024778_, _024787_, _024801_);
  and g_116438_(_024799_, _024801_, _024802_);
  or g_116439_(_024798_, _024800_, _024803_);
  and g_116440_(_024790_, _024803_, _024805_);
  or g_116441_(_024789_, _024802_, _024806_);
  and g_116442_(_024794_, _024797_, _024807_);
  or g_116443_(_024795_, _024796_, _024808_);
  and g_116444_(_024790_, _024808_, _024809_);
  or g_116445_(_024789_, _024807_, _024810_);
  xor g_116446_(out[745], _024784_, _024811_);
  xor g_116447_(_000604_, _024784_, _024812_);
  and g_116448_(_024589_, _024769_, _024813_);
  and g_116449_(_024581_, _024768_, _024814_);
  or g_116450_(_024813_, _024814_, _024816_);
  not g_116451_(_024816_, _024817_);
  or g_116452_(_024812_, _024816_, _024818_);
  and g_116453_(_024802_, _024818_, _024819_);
  not g_116454_(_024819_, _024820_);
  and g_116455_(_024809_, _024819_, _024821_);
  or g_116456_(_024810_, _024820_, _024822_);
  xor g_116457_(out[744], _024783_, _024823_);
  not g_116458_(_024823_, _024824_);
  and g_116459_(_024607_, _024769_, _024825_);
  and g_116460_(_024600_, _024768_, _024827_);
  or g_116461_(_024825_, _024827_, _024828_);
  not g_116462_(_024828_, _024829_);
  and g_116463_(_024823_, _024828_, _024830_);
  not g_116464_(_024830_, _024831_);
  and g_116465_(_024812_, _024816_, _024832_);
  or g_116466_(_024811_, _024817_, _024833_);
  and g_116467_(_024831_, _024833_, _024834_);
  or g_116468_(_024830_, _024832_, _024835_);
  xor g_116469_(out[742], _024780_, _024836_);
  xor g_116470_(_000516_, _024780_, _024838_);
  and g_116471_(_024637_, _024769_, _024839_);
  or g_116472_(_024636_, _024768_, _024840_);
  and g_116473_(_024630_, _024768_, _024841_);
  or g_116474_(_024631_, _024769_, _024842_);
  and g_116475_(_024840_, _024842_, _024843_);
  or g_116476_(_024839_, _024841_, _024844_);
  and g_116477_(_024836_, _024843_, _024845_);
  or g_116478_(_024838_, _024844_, _024846_);
  xor g_116479_(out[743], _024781_, _024847_);
  xor g_116480_(_000505_, _024781_, _024849_);
  and g_116481_(_024626_, _024769_, _024850_);
  or g_116482_(_024625_, _024768_, _024851_);
  and g_116483_(_024620_, _024768_, _024852_);
  or g_116484_(_024619_, _024769_, _024853_);
  and g_116485_(_024851_, _024853_, _024854_);
  or g_116486_(_024850_, _024852_, _024855_);
  and g_116487_(_024847_, _024855_, _024856_);
  or g_116488_(_024849_, _024854_, _024857_);
  and g_116489_(_024846_, _024857_, _024858_);
  or g_116490_(_024845_, _024856_, _024860_);
  and g_116491_(_024849_, _024854_, _024861_);
  or g_116492_(_024847_, _024855_, _024862_);
  and g_116493_(_024838_, _024844_, _024863_);
  or g_116494_(_024836_, _024843_, _024864_);
  and g_116495_(_024862_, _024864_, _024865_);
  or g_116496_(_024861_, _024863_, _024866_);
  and g_116497_(_024858_, _024865_, _024867_);
  or g_116498_(_024860_, _024866_, _024868_);
  xor g_116499_(out[741], _024779_, _024869_);
  xor g_116500_(_000527_, _024779_, _024871_);
  and g_116501_(_024655_, _024769_, _024872_);
  not g_116502_(_024872_, _024873_);
  or g_116503_(_024647_, _024769_, _024874_);
  not g_116504_(_024874_, _024875_);
  and g_116505_(_024873_, _024874_, _024876_);
  or g_116506_(_024872_, _024875_, _024877_);
  and g_116507_(_024869_, _024877_, _024878_);
  or g_116508_(_024871_, _024876_, _024879_);
  xor g_116509_(out[740], out[739], _024880_);
  xor g_116510_(_000538_, out[739], _024882_);
  or g_116511_(_024666_, _024769_, _024883_);
  not g_116512_(_024883_, _024884_);
  and g_116513_(_024673_, _024769_, _024885_);
  not g_116514_(_024885_, _024886_);
  and g_116515_(_024883_, _024886_, _024887_);
  or g_116516_(_024884_, _024885_, _024888_);
  and g_116517_(_024882_, _024888_, _024889_);
  or g_116518_(_024880_, _024887_, _024890_);
  and g_116519_(_024879_, _024890_, _024891_);
  or g_116520_(_024878_, _024889_, _024893_);
  or g_116521_(_024869_, _024877_, _024894_);
  not g_116522_(_024894_, _024895_);
  or g_116523_(_024882_, _024888_, _024896_);
  not g_116524_(_024896_, _024897_);
  and g_116525_(_024894_, _024896_, _024898_);
  or g_116526_(_024893_, _024895_, _024899_);
  and g_116527_(_024891_, _024898_, _024900_);
  or g_116528_(_024868_, _024897_, _024901_);
  and g_116529_(_024867_, _024900_, _024902_);
  or g_116530_(_024899_, _024901_, _024904_);
  and g_116531_(_024692_, _024769_, _024905_);
  not g_116532_(_024905_, _024906_);
  or g_116533_(out[722], _024769_, _024907_);
  not g_116534_(_024907_, _024908_);
  and g_116535_(_024906_, _024907_, _024909_);
  or g_116536_(_024905_, _024908_, _024910_);
  and g_116537_(_000571_, _024909_, _024911_);
  or g_116538_(out[738], _024910_, _024912_);
  or g_116539_(_000450_, _024769_, _024913_);
  not g_116540_(_024913_, _024915_);
  and g_116541_(_024700_, _024769_, _024916_);
  not g_116542_(_024916_, _024917_);
  and g_116543_(_024913_, _024917_, _024918_);
  or g_116544_(_024915_, _024916_, _024919_);
  and g_116545_(out[739], _024918_, _024920_);
  or g_116546_(_000582_, _024919_, _024921_);
  and g_116547_(_000582_, _024919_, _024922_);
  or g_116548_(out[739], _024918_, _024923_);
  xor g_116549_(_000571_, _024909_, _024924_);
  xor g_116550_(out[738], _024909_, _024926_);
  and g_116551_(_024923_, _024924_, _024927_);
  or g_116552_(_024922_, _024926_, _024928_);
  and g_116553_(_024921_, _024927_, _024929_);
  or g_116554_(_024920_, _024928_, _024930_);
  and g_116555_(_000549_, _024775_, _024931_);
  or g_116556_(out[737], _024776_, _024932_);
  and g_116557_(_024718_, _024769_, _024933_);
  not g_116558_(_024933_, _024934_);
  or g_116559_(out[720], _024769_, _024935_);
  not g_116560_(_024935_, _024937_);
  and g_116561_(_024934_, _024935_, _024938_);
  or g_116562_(_024933_, _024937_, _024939_);
  and g_116563_(out[736], _024939_, _024940_);
  or g_116564_(_000560_, _024938_, _024941_);
  xor g_116565_(_000549_, _024775_, _024942_);
  xor g_116566_(out[737], _024775_, _024943_);
  and g_116567_(_024941_, _024942_, _024944_);
  or g_116568_(_024940_, _024943_, _024945_);
  and g_116569_(_024932_, _024945_, _024946_);
  or g_116570_(_024931_, _024944_, _024948_);
  and g_116571_(_024929_, _024948_, _024949_);
  or g_116572_(_024930_, _024946_, _024950_);
  and g_116573_(_024911_, _024923_, _024951_);
  or g_116574_(_024912_, _024922_, _024952_);
  and g_116575_(_024921_, _024952_, _024953_);
  or g_116576_(_024920_, _024951_, _024954_);
  and g_116577_(_024950_, _024953_, _024955_);
  or g_116578_(_024949_, _024954_, _024956_);
  and g_116579_(_024902_, _024956_, _024957_);
  or g_116580_(_024904_, _024955_, _024959_);
  and g_116581_(_024860_, _024862_, _024960_);
  or g_116582_(_024858_, _024861_, _024961_);
  and g_116583_(_024867_, _024893_, _024962_);
  or g_116584_(_024868_, _024891_, _024963_);
  and g_116585_(_024894_, _024962_, _024964_);
  or g_116586_(_024895_, _024963_, _024965_);
  and g_116587_(_024961_, _024965_, _024966_);
  or g_116588_(_024960_, _024964_, _024967_);
  and g_116589_(_024959_, _024966_, _024968_);
  or g_116590_(_024957_, _024967_, _024970_);
  and g_116591_(_024824_, _024829_, _024971_);
  or g_116592_(_024823_, _024828_, _024972_);
  and g_116593_(_024970_, _024972_, _024973_);
  or g_116594_(_024968_, _024971_, _024974_);
  and g_116595_(_024834_, _024974_, _024975_);
  or g_116596_(_024835_, _024973_, _024976_);
  and g_116597_(_024821_, _024976_, _024977_);
  or g_116598_(_024822_, _024975_, _024978_);
  and g_116599_(_024806_, _024978_, _024979_);
  or g_116600_(_024805_, _024977_, _024981_);
  or g_116601_(out[736], _024939_, _024982_);
  and g_116602_(_024972_, _024982_, _024983_);
  not g_116603_(_024983_, _024984_);
  and g_116604_(_024834_, _024983_, _024985_);
  or g_116605_(_024835_, _024984_, _024986_);
  and g_116606_(_024929_, _024985_, _024987_);
  or g_116607_(_024930_, _024986_, _024988_);
  and g_116608_(_024944_, _024987_, _024989_);
  or g_116609_(_024945_, _024988_, _024990_);
  and g_116610_(_024821_, _024902_, _024992_);
  or g_116611_(_024822_, _024904_, _024993_);
  and g_116612_(_024989_, _024992_, _024994_);
  or g_116613_(_024990_, _024993_, _024995_);
  and g_116614_(_024981_, _024995_, _024996_);
  or g_116615_(_024979_, _024994_, _024997_);
  and g_116616_(_024776_, _024997_, _024998_);
  and g_116617_(_000549_, _024996_, _024999_);
  or g_116618_(_024998_, _024999_, _025000_);
  and g_116619_(out[756], out[755], _025001_);
  or g_116620_(out[757], _025001_, _025003_);
  or g_116621_(out[758], _025003_, _025004_);
  or g_116622_(out[759], _025004_, _025005_);
  or g_116623_(out[760], _025005_, _025006_);
  and g_116624_(out[761], _025006_, _025007_);
  or g_116625_(out[762], _025007_, _025008_);
  xor g_116626_(out[762], _025007_, _025009_);
  xor g_116627_(_000747_, _025007_, _025010_);
  or g_116628_(_024797_, _024997_, _025011_);
  not g_116629_(_025011_, _025012_);
  and g_116630_(_024794_, _024997_, _025014_);
  not g_116631_(_025014_, _025015_);
  and g_116632_(_025011_, _025015_, _025016_);
  or g_116633_(_025012_, _025014_, _025017_);
  and g_116634_(_025009_, _025016_, _025018_);
  or g_116635_(_025010_, _025017_, _025019_);
  and g_116636_(_024777_, _024787_, _025020_);
  or g_116637_(_024778_, _024788_, _025021_);
  xor g_116638_(out[763], _025008_, _025022_);
  xor g_116639_(_000626_, _025008_, _025023_);
  and g_116640_(_025020_, _025023_, _025025_);
  or g_116641_(_025021_, _025022_, _025026_);
  and g_116642_(_025019_, _025026_, _025027_);
  or g_116643_(_025018_, _025025_, _025028_);
  and g_116644_(_025010_, _025017_, _025029_);
  or g_116645_(_025009_, _025016_, _025030_);
  and g_116646_(_025021_, _025022_, _025031_);
  or g_116647_(_025020_, _025023_, _025032_);
  xor g_116648_(_000736_, _025006_, _025033_);
  and g_116649_(_024811_, _024996_, _025034_);
  and g_116650_(_024816_, _024997_, _025036_);
  or g_116651_(_025034_, _025036_, _025037_);
  or g_116652_(_025033_, _025037_, _025038_);
  xor g_116653_(out[760], _025005_, _025039_);
  and g_116654_(_024828_, _024997_, _025040_);
  and g_116655_(_024824_, _024996_, _025041_);
  or g_116656_(_025040_, _025041_, _025042_);
  and g_116657_(_025039_, _025042_, _025043_);
  not g_116658_(_025043_, _025044_);
  and g_116659_(_025033_, _025037_, _025045_);
  not g_116660_(_025045_, _025047_);
  and g_116661_(_025044_, _025047_, _025048_);
  or g_116662_(_025043_, _025045_, _025049_);
  or g_116663_(_025039_, _025042_, _025050_);
  and g_116664_(_025030_, _025032_, _025051_);
  or g_116665_(_025029_, _025031_, _025052_);
  and g_116666_(_025027_, _025051_, _025053_);
  or g_116667_(_025028_, _025052_, _025054_);
  and g_116668_(_025038_, _025050_, _025055_);
  not g_116669_(_025055_, _025056_);
  and g_116670_(_025048_, _025055_, _025058_);
  or g_116671_(_025049_, _025056_, _025059_);
  and g_116672_(_025053_, _025058_, _025060_);
  or g_116673_(_025054_, _025059_, _025061_);
  xor g_116674_(out[759], _025004_, _025062_);
  not g_116675_(_025062_, _025063_);
  or g_116676_(_024847_, _024997_, _025064_);
  not g_116677_(_025064_, _025065_);
  and g_116678_(_024855_, _024997_, _025066_);
  or g_116679_(_024854_, _024996_, _025067_);
  and g_116680_(_025064_, _025067_, _025069_);
  or g_116681_(_025065_, _025066_, _025070_);
  and g_116682_(_025062_, _025070_, _025071_);
  not g_116683_(_025071_, _025072_);
  xor g_116684_(_000648_, _025003_, _025073_);
  and g_116685_(_024836_, _024996_, _025074_);
  and g_116686_(_024844_, _024997_, _025075_);
  or g_116687_(_025074_, _025075_, _025076_);
  or g_116688_(_025073_, _025076_, _025077_);
  not g_116689_(_025077_, _025078_);
  and g_116690_(_025072_, _025077_, _025080_);
  or g_116691_(_025071_, _025078_, _025081_);
  xor g_116692_(out[757], _025001_, _025082_);
  xor g_116693_(_000659_, _025001_, _025083_);
  or g_116694_(_024869_, _024997_, _025084_);
  not g_116695_(_025084_, _025085_);
  and g_116696_(_024877_, _024997_, _025086_);
  not g_116697_(_025086_, _025087_);
  and g_116698_(_025084_, _025087_, _025088_);
  or g_116699_(_025085_, _025086_, _025089_);
  and g_116700_(_025083_, _025088_, _025091_);
  or g_116701_(_025082_, _025089_, _025092_);
  and g_116702_(_025063_, _025069_, _025093_);
  or g_116703_(_025062_, _025070_, _025094_);
  and g_116704_(_025073_, _025076_, _025095_);
  not g_116705_(_025095_, _025096_);
  and g_116706_(_025094_, _025096_, _025097_);
  or g_116707_(_025093_, _025095_, _025098_);
  and g_116708_(_025092_, _025097_, _025099_);
  or g_116709_(_025091_, _025098_, _025100_);
  and g_116710_(_025080_, _025099_, _025102_);
  or g_116711_(_025081_, _025100_, _025103_);
  and g_116712_(_025082_, _025089_, _025104_);
  not g_116713_(_025104_, _025105_);
  xor g_116714_(_000670_, out[755], _025106_);
  and g_116715_(_024880_, _024996_, _025107_);
  and g_116716_(_024888_, _024997_, _025108_);
  or g_116717_(_025107_, _025108_, _025109_);
  and g_116718_(_025106_, _025109_, _025110_);
  not g_116719_(_025110_, _025111_);
  and g_116720_(_025105_, _025111_, _025113_);
  or g_116721_(_025104_, _025110_, _025114_);
  or g_116722_(_025106_, _025109_, _025115_);
  not g_116723_(_025115_, _025116_);
  and g_116724_(_025113_, _025115_, _025117_);
  or g_116725_(_025114_, _025116_, _025118_);
  and g_116726_(_025102_, _025117_, _025119_);
  or g_116727_(_025103_, _025118_, _025120_);
  and g_116728_(out[739], _024996_, _025121_);
  or g_116729_(_000582_, _024997_, _025122_);
  and g_116730_(_024919_, _024997_, _025124_);
  or g_116731_(_024918_, _024996_, _025125_);
  and g_116732_(_025122_, _025125_, _025126_);
  or g_116733_(_025121_, _025124_, _025127_);
  or g_116734_(_000714_, _025127_, _025128_);
  and g_116735_(_024910_, _024997_, _025129_);
  and g_116736_(_000571_, _024996_, _025130_);
  or g_116737_(_025129_, _025130_, _025131_);
  and g_116738_(_000714_, _025127_, _025132_);
  or g_116739_(out[754], _025131_, _025133_);
  xor g_116740_(out[755], _025126_, _025135_);
  xor g_116741_(_000714_, _025126_, _025136_);
  xor g_116742_(out[754], _025131_, _025137_);
  xor g_116743_(_000703_, _025131_, _025138_);
  and g_116744_(_025135_, _025137_, _025139_);
  or g_116745_(_025136_, _025138_, _025140_);
  or g_116746_(out[753], _025000_, _025141_);
  and g_116747_(_024939_, _024997_, _025142_);
  and g_116748_(_000560_, _024996_, _025143_);
  or g_116749_(_025142_, _025143_, _025144_);
  and g_116750_(out[752], _025144_, _025146_);
  not g_116751_(_025146_, _025147_);
  xor g_116752_(out[753], _025000_, _025148_);
  xor g_116753_(_000681_, _025000_, _025149_);
  and g_116754_(_025147_, _025148_, _025150_);
  or g_116755_(_025146_, _025149_, _025151_);
  and g_116756_(_025141_, _025151_, _025152_);
  or g_116757_(_025140_, _025152_, _025153_);
  or g_116758_(_025132_, _025133_, _025154_);
  and g_116759_(_025128_, _025154_, _025155_);
  and g_116760_(_025153_, _025155_, _025157_);
  or g_116761_(_025120_, _025157_, _025158_);
  or g_116762_(_025103_, _025113_, _025159_);
  and g_116763_(_025081_, _025094_, _025160_);
  not g_116764_(_025160_, _025161_);
  and g_116765_(_025159_, _025161_, _025162_);
  and g_116766_(_025158_, _025162_, _025163_);
  or g_116767_(_025061_, _025163_, _025164_);
  and g_116768_(_025038_, _025049_, _025165_);
  not g_116769_(_025165_, _025166_);
  or g_116770_(_025054_, _025166_, _025168_);
  or g_116771_(_025027_, _025031_, _025169_);
  and g_116772_(_025168_, _025169_, _025170_);
  and g_116773_(_025164_, _025170_, _025171_);
  or g_116774_(out[752], _025144_, _025172_);
  and g_116775_(_025139_, _025172_, _025173_);
  and g_116776_(_025150_, _025173_, _025174_);
  and g_116777_(_025060_, _025174_, _025175_);
  and g_116778_(_025119_, _025175_, _025176_);
  or g_116779_(_025171_, _025176_, _025177_);
  and g_116780_(_025000_, _025177_, _025179_);
  not g_116781_(_025179_, _025180_);
  or g_116782_(out[753], _025177_, _025181_);
  not g_116783_(_025181_, _025182_);
  and g_116784_(_025180_, _025181_, _025183_);
  or g_116785_(_025179_, _025182_, _025184_);
  and g_116786_(_025020_, _025022_, _025185_);
  or g_116787_(_025021_, _025023_, _025186_);
  and g_116788_(out[772], out[771], _025187_);
  or g_116789_(out[773], _025187_, _025188_);
  or g_116790_(out[774], _025188_, _025190_);
  or g_116791_(out[775], _025190_, _025191_);
  or g_116792_(out[776], _025191_, _025192_);
  and g_116793_(out[777], _025192_, _025193_);
  or g_116794_(out[778], _025193_, _025194_);
  xor g_116795_(out[779], _025194_, _025195_);
  xor g_116796_(_000758_, _025194_, _025196_);
  and g_116797_(_025185_, _025196_, _025197_);
  or g_116798_(_025185_, _025196_, _025198_);
  xor g_116799_(_025186_, _025195_, _025199_);
  or g_116800_(_025009_, _025177_, _025201_);
  not g_116801_(_025201_, _025202_);
  and g_116802_(_025016_, _025177_, _025203_);
  or g_116803_(_025202_, _025203_, _025204_);
  xor g_116804_(out[778], _025193_, _025205_);
  and g_116805_(_025204_, _025205_, _025206_);
  xor g_116806_(out[777], _025192_, _025207_);
  not g_116807_(_025207_, _025208_);
  or g_116808_(_025033_, _025177_, _025209_);
  not g_116809_(_025209_, _025210_);
  and g_116810_(_025037_, _025177_, _025212_);
  or g_116811_(_025210_, _025212_, _025213_);
  or g_116812_(_025208_, _025213_, _025214_);
  xor g_116813_(_025204_, _025205_, _025215_);
  and g_116814_(_025199_, _025215_, _025216_);
  and g_116815_(_025214_, _025216_, _025217_);
  and g_116816_(_025208_, _025213_, _025218_);
  xor g_116817_(out[776], _025191_, _025219_);
  or g_116818_(_025039_, _025177_, _025220_);
  not g_116819_(_025220_, _025221_);
  and g_116820_(_025042_, _025177_, _025223_);
  or g_116821_(_025221_, _025223_, _025224_);
  and g_116822_(_025219_, _025224_, _025225_);
  or g_116823_(_025218_, _025225_, _025226_);
  not g_116824_(_025226_, _025227_);
  or g_116825_(_025219_, _025224_, _025228_);
  and g_116826_(_025227_, _025228_, _025229_);
  and g_116827_(_025217_, _025229_, _025230_);
  xor g_116828_(out[775], _025190_, _025231_);
  not g_116829_(_025231_, _025232_);
  or g_116830_(_025062_, _025177_, _025234_);
  not g_116831_(_025234_, _025235_);
  and g_116832_(_025070_, _025177_, _025236_);
  not g_116833_(_025236_, _025237_);
  and g_116834_(_025234_, _025237_, _025238_);
  or g_116835_(_025235_, _025236_, _025239_);
  and g_116836_(_025231_, _025239_, _025240_);
  or g_116837_(_025232_, _025238_, _025241_);
  xor g_116838_(out[774], _025188_, _025242_);
  not g_116839_(_025242_, _025243_);
  or g_116840_(_025073_, _025177_, _025245_);
  not g_116841_(_025245_, _025246_);
  and g_116842_(_025076_, _025177_, _025247_);
  not g_116843_(_025247_, _025248_);
  and g_116844_(_025245_, _025248_, _025249_);
  or g_116845_(_025246_, _025247_, _025250_);
  and g_116846_(_025242_, _025249_, _025251_);
  or g_116847_(_025243_, _025250_, _025252_);
  and g_116848_(_025241_, _025252_, _025253_);
  or g_116849_(_025240_, _025251_, _025254_);
  or g_116850_(_025231_, _025239_, _025256_);
  or g_116851_(_025242_, _025249_, _025257_);
  and g_116852_(_025256_, _025257_, _025258_);
  and g_116853_(_025253_, _025258_, _025259_);
  xor g_116854_(out[772], out[771], _025260_);
  not g_116855_(_025260_, _025261_);
  or g_116856_(_025106_, _025177_, _025262_);
  not g_116857_(_025262_, _025263_);
  and g_116858_(_025109_, _025177_, _025264_);
  or g_116859_(_025263_, _025264_, _025265_);
  and g_116860_(_025261_, _025265_, _025267_);
  xor g_116861_(out[773], _025187_, _025268_);
  or g_116862_(_025082_, _025177_, _025269_);
  not g_116863_(_025269_, _025270_);
  and g_116864_(_025089_, _025177_, _025271_);
  or g_116865_(_025270_, _025271_, _025272_);
  and g_116866_(_025268_, _025272_, _025273_);
  or g_116867_(_025267_, _025273_, _025274_);
  not g_116868_(_025274_, _025275_);
  or g_116869_(_025268_, _025272_, _025276_);
  or g_116870_(_025261_, _025265_, _025278_);
  and g_116871_(_025276_, _025278_, _025279_);
  and g_116872_(_025275_, _025279_, _025280_);
  and g_116873_(_025259_, _025280_, _025281_);
  and g_116874_(_025230_, _025281_, _025282_);
  and g_116875_(_025126_, _025177_, _025283_);
  or g_116876_(out[755], _025177_, _025284_);
  not g_116877_(_025284_, _025285_);
  or g_116878_(_025283_, _025285_, _025286_);
  and g_116879_(out[771], _025286_, _025287_);
  and g_116880_(_025131_, _025177_, _025289_);
  not g_116881_(_025289_, _025290_);
  or g_116882_(out[754], _025177_, _025291_);
  and g_116883_(_025290_, _025291_, _025292_);
  or g_116884_(out[771], _025286_, _025293_);
  not g_116885_(_025293_, _025294_);
  and g_116886_(_000835_, _025292_, _025295_);
  or g_116887_(_025287_, _025294_, _025296_);
  xor g_116888_(out[770], _025292_, _025297_);
  or g_116889_(_025296_, _025297_, _025298_);
  or g_116890_(out[769], _025184_, _025300_);
  and g_116891_(_025144_, _025177_, _025301_);
  not g_116892_(_025301_, _025302_);
  or g_116893_(out[752], _025177_, _025303_);
  not g_116894_(_025303_, _025304_);
  and g_116895_(_025302_, _025303_, _025305_);
  or g_116896_(_025301_, _025304_, _025306_);
  and g_116897_(out[768], _025306_, _025307_);
  xor g_116898_(out[769], _025183_, _025308_);
  or g_116899_(_025307_, _025308_, _025309_);
  and g_116900_(_025300_, _025309_, _025311_);
  or g_116901_(_025298_, _025311_, _025312_);
  not g_116902_(_025312_, _025313_);
  and g_116903_(_025293_, _025295_, _025314_);
  or g_116904_(_025287_, _025314_, _025315_);
  or g_116905_(_025313_, _025315_, _025316_);
  and g_116906_(_025282_, _025316_, _025317_);
  and g_116907_(_025274_, _025276_, _025318_);
  and g_116908_(_025259_, _025318_, _025319_);
  and g_116909_(_025254_, _025256_, _025320_);
  or g_116910_(_025319_, _025320_, _025322_);
  and g_116911_(_025230_, _025322_, _025323_);
  and g_116912_(_025217_, _025226_, _025324_);
  and g_116913_(_025198_, _025206_, _025325_);
  or g_116914_(_025197_, _025325_, _025326_);
  or g_116915_(_025324_, _025326_, _025327_);
  or g_116916_(_025323_, _025327_, _025328_);
  or g_116917_(_025317_, _025328_, _025329_);
  or g_116918_(out[768], _025306_, _025330_);
  or g_116919_(_025298_, _025309_, _025331_);
  not g_116920_(_025331_, _025333_);
  and g_116921_(_025330_, _025333_, _025334_);
  and g_116922_(_025282_, _025334_, _025335_);
  not g_116923_(_025335_, _025336_);
  and g_116924_(_025329_, _025336_, _025337_);
  not g_116925_(_025337_, _025338_);
  and g_116926_(out[769], _025337_, _025339_);
  not g_116927_(_025339_, _025340_);
  and g_116928_(_025183_, _025338_, _025341_);
  or g_116929_(_025184_, _025337_, _025342_);
  or g_116930_(_025339_, _025341_, _025344_);
  and g_116931_(_025340_, _025342_, _025345_);
  and g_116932_(_025205_, _025337_, _025346_);
  not g_116933_(_025346_, _025347_);
  or g_116934_(_025204_, _025337_, _025348_);
  not g_116935_(_025348_, _025349_);
  and g_116936_(_025347_, _025348_, _025350_);
  or g_116937_(_025346_, _025349_, _025351_);
  and g_116938_(out[788], out[787], _025352_);
  or g_116939_(out[789], _025352_, _025353_);
  or g_116940_(out[790], _025353_, _025355_);
  or g_116941_(out[791], _025355_, _025356_);
  or g_116942_(out[792], _025356_, _025357_);
  and g_116943_(out[793], _025357_, _025358_);
  or g_116944_(out[794], _025358_, _025359_);
  xor g_116945_(out[794], _025358_, _025360_);
  xor g_116946_(_001011_, _025358_, _025361_);
  and g_116947_(_025350_, _025360_, _025362_);
  or g_116948_(_025351_, _025361_, _025363_);
  and g_116949_(_025185_, _025195_, _025364_);
  or g_116950_(_025186_, _025196_, _025366_);
  xor g_116951_(out[795], _025359_, _025367_);
  xor g_116952_(_000890_, _025359_, _025368_);
  and g_116953_(_025366_, _025367_, _025369_);
  or g_116954_(_025364_, _025368_, _025370_);
  and g_116955_(_025364_, _025368_, _025371_);
  or g_116956_(_025366_, _025367_, _025372_);
  and g_116957_(_025370_, _025372_, _025373_);
  or g_116958_(_025369_, _025371_, _025374_);
  and g_116959_(_025363_, _025373_, _025375_);
  or g_116960_(_025362_, _025374_, _025377_);
  or g_116961_(_025350_, _025360_, _025378_);
  xor g_116962_(_001000_, _025357_, _025379_);
  and g_116963_(_025207_, _025337_, _025380_);
  and g_116964_(_025213_, _025338_, _025381_);
  or g_116965_(_025380_, _025381_, _025382_);
  or g_116966_(_025379_, _025382_, _025383_);
  and g_116967_(_025378_, _025383_, _025384_);
  not g_116968_(_025384_, _025385_);
  and g_116969_(_025375_, _025384_, _025386_);
  or g_116970_(_025377_, _025385_, _025388_);
  xor g_116971_(out[792], _025356_, _025389_);
  not g_116972_(_025389_, _025390_);
  or g_116973_(_025224_, _025337_, _025391_);
  and g_116974_(_025219_, _025337_, _025392_);
  not g_116975_(_025392_, _025393_);
  and g_116976_(_025391_, _025393_, _025394_);
  not g_116977_(_025394_, _025395_);
  and g_116978_(_025389_, _025394_, _025396_);
  not g_116979_(_025396_, _025397_);
  and g_116980_(_025379_, _025382_, _025399_);
  not g_116981_(_025399_, _025400_);
  and g_116982_(_025397_, _025400_, _025401_);
  or g_116983_(_025396_, _025399_, _025402_);
  xor g_116984_(out[791], _025355_, _025403_);
  not g_116985_(_025403_, _025404_);
  and g_116986_(_025232_, _025337_, _025405_);
  and g_116987_(_025239_, _025338_, _025406_);
  or g_116988_(_025405_, _025406_, _025407_);
  not g_116989_(_025407_, _025408_);
  and g_116990_(_025403_, _025407_, _025410_);
  not g_116991_(_025410_, _025411_);
  xor g_116992_(_000912_, _025353_, _025412_);
  and g_116993_(_025242_, _025337_, _025413_);
  and g_116994_(_025250_, _025338_, _025414_);
  or g_116995_(_025413_, _025414_, _025415_);
  or g_116996_(_025412_, _025415_, _025416_);
  not g_116997_(_025416_, _025417_);
  and g_116998_(_025411_, _025416_, _025418_);
  or g_116999_(_025410_, _025417_, _025419_);
  xor g_117000_(out[789], _025352_, _025421_);
  or g_117001_(_025272_, _025337_, _025422_);
  and g_117002_(_025268_, _025337_, _025423_);
  not g_117003_(_025423_, _025424_);
  and g_117004_(_025422_, _025424_, _025425_);
  or g_117005_(_025421_, _025425_, _025426_);
  not g_117006_(_025426_, _025427_);
  and g_117007_(_025404_, _025408_, _025428_);
  or g_117008_(_025403_, _025407_, _025429_);
  and g_117009_(_025412_, _025415_, _025430_);
  not g_117010_(_025430_, _025432_);
  and g_117011_(_025429_, _025432_, _025433_);
  or g_117012_(_025428_, _025430_, _025434_);
  and g_117013_(_025426_, _025433_, _025435_);
  or g_117014_(_025427_, _025434_, _025436_);
  and g_117015_(_025418_, _025435_, _025437_);
  or g_117016_(_025419_, _025436_, _025438_);
  and g_117017_(_025421_, _025425_, _025439_);
  not g_117018_(_025439_, _025440_);
  xor g_117019_(_000934_, out[787], _025441_);
  and g_117020_(_025260_, _025337_, _025443_);
  and g_117021_(_025265_, _025338_, _025444_);
  or g_117022_(_025443_, _025444_, _025445_);
  and g_117023_(_025441_, _025445_, _025446_);
  not g_117024_(_025446_, _025447_);
  and g_117025_(_025440_, _025447_, _025448_);
  or g_117026_(_025439_, _025446_, _025449_);
  or g_117027_(_025441_, _025445_, _025450_);
  not g_117028_(_025450_, _025451_);
  and g_117029_(_025448_, _025450_, _025452_);
  or g_117030_(_025449_, _025451_, _025454_);
  and g_117031_(_025437_, _025452_, _025455_);
  or g_117032_(_025438_, _025454_, _025456_);
  or g_117033_(_025292_, _025337_, _025457_);
  not g_117034_(_025457_, _025458_);
  and g_117035_(_000835_, _025337_, _025459_);
  or g_117036_(_025458_, _025459_, _025460_);
  or g_117037_(out[786], _025460_, _025461_);
  not g_117038_(_025461_, _025462_);
  and g_117039_(out[771], _025337_, _025463_);
  not g_117040_(_025463_, _025465_);
  or g_117041_(_025286_, _025337_, _025466_);
  not g_117042_(_025466_, _025467_);
  and g_117043_(_025465_, _025466_, _025468_);
  or g_117044_(_025463_, _025467_, _025469_);
  and g_117045_(out[787], _025468_, _025470_);
  or g_117046_(_000978_, _025469_, _025471_);
  and g_117047_(_000978_, _025469_, _025472_);
  or g_117048_(out[787], _025468_, _025473_);
  xor g_117049_(out[786], _025460_, _025474_);
  xor g_117050_(_000967_, _025460_, _025476_);
  and g_117051_(_025473_, _025474_, _025477_);
  or g_117052_(_025472_, _025476_, _025478_);
  and g_117053_(_025471_, _025477_, _025479_);
  or g_117054_(_025470_, _025478_, _025480_);
  and g_117055_(out[768], _025337_, _025481_);
  not g_117056_(_025481_, _025482_);
  and g_117057_(_025305_, _025338_, _025483_);
  or g_117058_(_025306_, _025337_, _025484_);
  or g_117059_(_025481_, _025483_, _025485_);
  and g_117060_(_025482_, _025484_, _025487_);
  and g_117061_(out[784], _025487_, _025488_);
  or g_117062_(_000956_, _025485_, _025489_);
  and g_117063_(out[785], _025345_, _025490_);
  or g_117064_(_000945_, _025344_, _025491_);
  and g_117065_(_025489_, _025491_, _025492_);
  or g_117066_(_025488_, _025490_, _025493_);
  or g_117067_(out[785], _025345_, _025494_);
  not g_117068_(_025494_, _025495_);
  and g_117069_(_025493_, _025494_, _025496_);
  or g_117070_(_025492_, _025495_, _025498_);
  and g_117071_(_025479_, _025498_, _025499_);
  or g_117072_(_025480_, _025496_, _025500_);
  and g_117073_(_025462_, _025473_, _025501_);
  or g_117074_(_025461_, _025472_, _025502_);
  and g_117075_(_025471_, _025502_, _025503_);
  or g_117076_(_025470_, _025501_, _025504_);
  and g_117077_(_025500_, _025503_, _025505_);
  or g_117078_(_025499_, _025504_, _025506_);
  and g_117079_(_025455_, _025506_, _025507_);
  or g_117080_(_025456_, _025505_, _025509_);
  and g_117081_(_025437_, _025449_, _025510_);
  and g_117082_(_025419_, _025429_, _025511_);
  or g_117083_(_025510_, _025511_, _025512_);
  not g_117084_(_025512_, _025513_);
  and g_117085_(_025509_, _025513_, _025514_);
  or g_117086_(_025507_, _025512_, _025515_);
  and g_117087_(_025390_, _025395_, _025516_);
  or g_117088_(_025389_, _025394_, _025517_);
  and g_117089_(_025515_, _025517_, _025518_);
  or g_117090_(_025514_, _025516_, _025520_);
  and g_117091_(_025401_, _025517_, _025521_);
  and g_117092_(_025401_, _025520_, _025522_);
  or g_117093_(_025402_, _025518_, _025523_);
  and g_117094_(_025386_, _025523_, _025524_);
  or g_117095_(_025388_, _025522_, _025525_);
  and g_117096_(_025362_, _025370_, _025526_);
  or g_117097_(_025363_, _025369_, _025527_);
  or g_117098_(_025371_, _025526_, _025528_);
  and g_117099_(_025372_, _025527_, _025529_);
  and g_117100_(_025525_, _025529_, _025531_);
  or g_117101_(_025524_, _025528_, _025532_);
  or g_117102_(out[784], _025487_, _025533_);
  or g_117103_(_025480_, _025493_, _025534_);
  not g_117104_(_025534_, _025535_);
  and g_117105_(_025521_, _025533_, _025536_);
  not g_117106_(_025536_, _025537_);
  and g_117107_(_025535_, _025536_, _025538_);
  or g_117108_(_025534_, _025537_, _025539_);
  and g_117109_(_025455_, _025494_, _025540_);
  and g_117110_(_025386_, _025540_, _025542_);
  not g_117111_(_025542_, _025543_);
  and g_117112_(_025538_, _025542_, _025544_);
  or g_117113_(_025539_, _025543_, _025545_);
  and g_117114_(_025532_, _025545_, _025546_);
  or g_117115_(_025531_, _025544_, _025547_);
  and g_117116_(_025345_, _025547_, _025548_);
  and g_117117_(_000945_, _025546_, _025549_);
  or g_117118_(_025548_, _025549_, _025550_);
  and g_117119_(_025364_, _025367_, _025551_);
  or g_117120_(_025366_, _025368_, _025553_);
  and g_117121_(out[804], out[803], _025554_);
  or g_117122_(out[805], _025554_, _025555_);
  or g_117123_(out[806], _025555_, _025556_);
  or g_117124_(out[807], _025556_, _025557_);
  or g_117125_(out[808], _025557_, _025558_);
  and g_117126_(out[809], _025558_, _025559_);
  or g_117127_(out[810], _025559_, _025560_);
  xor g_117128_(out[811], _025560_, _025561_);
  xor g_117129_(_001022_, _025560_, _025562_);
  and g_117130_(_025551_, _025562_, _025564_);
  or g_117131_(_025553_, _025561_, _025565_);
  and g_117132_(_025360_, _025546_, _025566_);
  or g_117133_(_025361_, _025547_, _025567_);
  and g_117134_(_025351_, _025547_, _025568_);
  or g_117135_(_025350_, _025546_, _025569_);
  and g_117136_(_025567_, _025569_, _025570_);
  or g_117137_(_025566_, _025568_, _025571_);
  xor g_117138_(out[810], _025559_, _025572_);
  xor g_117139_(_001143_, _025559_, _025573_);
  and g_117140_(_025570_, _025572_, _025575_);
  or g_117141_(_025571_, _025573_, _025576_);
  and g_117142_(_025565_, _025576_, _025577_);
  or g_117143_(_025564_, _025575_, _025578_);
  and g_117144_(_025571_, _025573_, _025579_);
  or g_117145_(_025570_, _025572_, _025580_);
  and g_117146_(_025553_, _025561_, _025581_);
  or g_117147_(_025551_, _025562_, _025582_);
  xor g_117148_(out[809], _025558_, _025583_);
  or g_117149_(_025379_, _025547_, _025584_);
  and g_117150_(_025382_, _025547_, _025586_);
  not g_117151_(_025586_, _025587_);
  and g_117152_(_025584_, _025587_, _025588_);
  and g_117153_(_025583_, _025588_, _025589_);
  not g_117154_(_025589_, _025590_);
  and g_117155_(_025580_, _025582_, _025591_);
  or g_117156_(_025579_, _025581_, _025592_);
  and g_117157_(_025577_, _025591_, _025593_);
  or g_117158_(_025578_, _025592_, _025594_);
  and g_117159_(_025590_, _025593_, _025595_);
  or g_117160_(_025589_, _025594_, _025597_);
  or g_117161_(_025583_, _025588_, _025598_);
  not g_117162_(_025598_, _025599_);
  xor g_117163_(_001121_, _025557_, _025600_);
  or g_117164_(_025389_, _025547_, _025601_);
  or g_117165_(_025395_, _025546_, _025602_);
  and g_117166_(_025601_, _025602_, _025603_);
  or g_117167_(_025600_, _025603_, _025604_);
  not g_117168_(_025604_, _025605_);
  and g_117169_(_025598_, _025604_, _025606_);
  or g_117170_(_025599_, _025605_, _025608_);
  and g_117171_(_025600_, _025603_, _025609_);
  not g_117172_(_025609_, _025610_);
  and g_117173_(_025606_, _025610_, _025611_);
  or g_117174_(_025608_, _025609_, _025612_);
  and g_117175_(_025595_, _025611_, _025613_);
  or g_117176_(_025597_, _025612_, _025614_);
  xor g_117177_(out[806], _025555_, _025615_);
  or g_117178_(_025412_, _025547_, _025616_);
  and g_117179_(_025415_, _025547_, _025617_);
  not g_117180_(_025617_, _025619_);
  and g_117181_(_025616_, _025619_, _025620_);
  and g_117182_(_025615_, _025620_, _025621_);
  not g_117183_(_025621_, _025622_);
  xor g_117184_(out[807], _025556_, _025623_);
  xor g_117185_(_001033_, _025556_, _025624_);
  or g_117186_(_025403_, _025547_, _025625_);
  or g_117187_(_025408_, _025546_, _025626_);
  and g_117188_(_025625_, _025626_, _025627_);
  not g_117189_(_025627_, _025628_);
  or g_117190_(_025624_, _025627_, _025630_);
  not g_117191_(_025630_, _025631_);
  and g_117192_(_025622_, _025630_, _025632_);
  or g_117193_(_025621_, _025631_, _025633_);
  or g_117194_(_025615_, _025620_, _025634_);
  not g_117195_(_025634_, _025635_);
  and g_117196_(_025624_, _025627_, _025636_);
  or g_117197_(_025623_, _025628_, _025637_);
  and g_117198_(_025634_, _025637_, _025638_);
  or g_117199_(_025633_, _025636_, _025639_);
  and g_117200_(_025632_, _025638_, _025641_);
  or g_117201_(_025635_, _025639_, _025642_);
  xor g_117202_(_001055_, _025554_, _025643_);
  or g_117203_(_025421_, _025547_, _025644_);
  and g_117204_(_025425_, _025547_, _025645_);
  not g_117205_(_025645_, _025646_);
  and g_117206_(_025644_, _025646_, _025647_);
  or g_117207_(_025643_, _025647_, _025648_);
  not g_117208_(_025648_, _025649_);
  xor g_117209_(out[804], out[803], _025650_);
  or g_117210_(_025441_, _025547_, _025652_);
  and g_117211_(_025445_, _025547_, _025653_);
  not g_117212_(_025653_, _025654_);
  and g_117213_(_025652_, _025654_, _025655_);
  or g_117214_(_025650_, _025655_, _025656_);
  not g_117215_(_025656_, _025657_);
  and g_117216_(_025648_, _025656_, _025658_);
  or g_117217_(_025649_, _025657_, _025659_);
  and g_117218_(_025650_, _025655_, _025660_);
  and g_117219_(_025643_, _025647_, _025661_);
  or g_117220_(_025660_, _025661_, _025663_);
  not g_117221_(_025663_, _025664_);
  and g_117222_(_025658_, _025664_, _025665_);
  or g_117223_(_025659_, _025663_, _025666_);
  or g_117224_(_025642_, _025666_, _025667_);
  and g_117225_(_025613_, _025665_, _025668_);
  and g_117226_(_025641_, _025668_, _025669_);
  or g_117227_(_025614_, _025667_, _025670_);
  or g_117228_(_000978_, _025547_, _025671_);
  or g_117229_(_025468_, _025546_, _025672_);
  and g_117230_(_025671_, _025672_, _025674_);
  and g_117231_(out[803], _025674_, _025675_);
  and g_117232_(_025460_, _025547_, _025676_);
  not g_117233_(_025676_, _025677_);
  or g_117234_(out[786], _025547_, _025678_);
  not g_117235_(_025678_, _025679_);
  and g_117236_(_025677_, _025678_, _025680_);
  or g_117237_(_025676_, _025679_, _025681_);
  or g_117238_(out[803], _025674_, _025682_);
  and g_117239_(_001099_, _025680_, _025683_);
  xor g_117240_(out[803], _025674_, _025685_);
  xor g_117241_(_001110_, _025674_, _025686_);
  xor g_117242_(_001099_, _025680_, _025687_);
  xor g_117243_(out[802], _025680_, _025688_);
  and g_117244_(_025685_, _025687_, _025689_);
  or g_117245_(_025686_, _025688_, _025690_);
  and g_117246_(_025487_, _025547_, _025691_);
  and g_117247_(_000956_, _025546_, _025692_);
  or g_117248_(_025691_, _025692_, _025693_);
  and g_117249_(out[800], _025693_, _025694_);
  or g_117250_(out[801], _025550_, _025696_);
  xor g_117251_(_001077_, _025550_, _025697_);
  or g_117252_(_025694_, _025697_, _025698_);
  not g_117253_(_025698_, _025699_);
  or g_117254_(out[800], _025693_, _025700_);
  not g_117255_(_025700_, _025701_);
  or g_117256_(_025698_, _025701_, _025702_);
  and g_117257_(_025689_, _025699_, _025703_);
  and g_117258_(_025700_, _025703_, _025704_);
  or g_117259_(_025690_, _025702_, _025705_);
  and g_117260_(_025669_, _025704_, _025707_);
  or g_117261_(_025670_, _025705_, _025708_);
  and g_117262_(_025696_, _025698_, _025709_);
  not g_117263_(_025709_, _025710_);
  and g_117264_(_025689_, _025710_, _025711_);
  or g_117265_(_025690_, _025709_, _025712_);
  and g_117266_(_025682_, _025683_, _025713_);
  or g_117267_(_025675_, _025713_, _025714_);
  not g_117268_(_025714_, _025715_);
  and g_117269_(_025712_, _025715_, _025716_);
  or g_117270_(_025711_, _025714_, _025718_);
  and g_117271_(_025669_, _025718_, _025719_);
  or g_117272_(_025670_, _025716_, _025720_);
  or g_117273_(_025632_, _025636_, _025721_);
  or g_117274_(_025658_, _025661_, _025722_);
  or g_117275_(_025642_, _025722_, _025723_);
  and g_117276_(_025721_, _025723_, _025724_);
  or g_117277_(_025614_, _025724_, _025725_);
  not g_117278_(_025725_, _025726_);
  and g_117279_(_025578_, _025582_, _025727_);
  or g_117280_(_025577_, _025581_, _025729_);
  or g_117281_(_025597_, _025606_, _025730_);
  not g_117282_(_025730_, _025731_);
  and g_117283_(_025729_, _025730_, _025732_);
  and g_117284_(_025725_, _025732_, _025733_);
  or g_117285_(_025719_, _025731_, _025734_);
  or g_117286_(_025727_, _025734_, _025735_);
  and g_117287_(_025720_, _025733_, _025736_);
  or g_117288_(_025726_, _025735_, _025737_);
  and g_117289_(_025708_, _025737_, _025738_);
  or g_117290_(_025707_, _025736_, _025740_);
  and g_117291_(_025550_, _025740_, _025741_);
  and g_117292_(_001077_, _025738_, _025742_);
  or g_117293_(_025741_, _025742_, _025743_);
  and g_117294_(_025572_, _025738_, _025744_);
  or g_117295_(_025573_, _025740_, _025745_);
  and g_117296_(_025571_, _025740_, _025746_);
  or g_117297_(_025570_, _025738_, _025747_);
  and g_117298_(_025745_, _025747_, _025748_);
  or g_117299_(_025744_, _025746_, _025749_);
  and g_117300_(out[820], out[819], _025751_);
  or g_117301_(out[821], _025751_, _025752_);
  or g_117302_(out[822], _025752_, _025753_);
  or g_117303_(out[823], _025753_, _025754_);
  or g_117304_(out[824], _025754_, _025755_);
  and g_117305_(out[825], _025755_, _025756_);
  or g_117306_(out[826], _025756_, _025757_);
  xor g_117307_(out[826], _025756_, _025758_);
  xor g_117308_(_001275_, _025756_, _025759_);
  and g_117309_(_025748_, _025758_, _025760_);
  or g_117310_(_025749_, _025759_, _025762_);
  and g_117311_(_025551_, _025561_, _025763_);
  or g_117312_(_025553_, _025562_, _025764_);
  xor g_117313_(out[827], _025757_, _025765_);
  xor g_117314_(_001154_, _025757_, _025766_);
  and g_117315_(_025763_, _025766_, _025767_);
  or g_117316_(_025764_, _025765_, _025768_);
  and g_117317_(_025762_, _025768_, _025769_);
  or g_117318_(_025760_, _025767_, _025770_);
  and g_117319_(_025749_, _025759_, _025771_);
  or g_117320_(_025748_, _025758_, _025773_);
  and g_117321_(_025764_, _025765_, _025774_);
  or g_117322_(_025763_, _025766_, _025775_);
  xor g_117323_(out[825], _025755_, _025776_);
  xor g_117324_(_001264_, _025755_, _025777_);
  and g_117325_(_025583_, _025738_, _025778_);
  not g_117326_(_025778_, _025779_);
  or g_117327_(_025588_, _025738_, _025780_);
  not g_117328_(_025780_, _025781_);
  and g_117329_(_025779_, _025780_, _025782_);
  or g_117330_(_025778_, _025781_, _025784_);
  and g_117331_(_025776_, _025782_, _025785_);
  or g_117332_(_025777_, _025784_, _025786_);
  xor g_117333_(out[824], _025754_, _025787_);
  not g_117334_(_025787_, _025788_);
  and g_117335_(_025600_, _025738_, _025789_);
  not g_117336_(_025789_, _025790_);
  or g_117337_(_025603_, _025738_, _025791_);
  not g_117338_(_025791_, _025792_);
  and g_117339_(_025790_, _025791_, _025793_);
  or g_117340_(_025789_, _025792_, _025795_);
  and g_117341_(_025787_, _025795_, _025796_);
  or g_117342_(_025788_, _025793_, _025797_);
  and g_117343_(_025777_, _025784_, _025798_);
  or g_117344_(_025776_, _025782_, _025799_);
  and g_117345_(_025797_, _025799_, _025800_);
  or g_117346_(_025796_, _025798_, _025801_);
  and g_117347_(_025788_, _025793_, _025802_);
  or g_117348_(_025787_, _025795_, _025803_);
  and g_117349_(_025773_, _025775_, _025804_);
  or g_117350_(_025771_, _025774_, _025806_);
  and g_117351_(_025769_, _025804_, _025807_);
  or g_117352_(_025770_, _025806_, _025808_);
  and g_117353_(_025786_, _025803_, _025809_);
  or g_117354_(_025785_, _025802_, _025810_);
  and g_117355_(_025800_, _025809_, _025811_);
  or g_117356_(_025801_, _025810_, _025812_);
  and g_117357_(_025807_, _025811_, _025813_);
  or g_117358_(_025808_, _025812_, _025814_);
  xor g_117359_(out[823], _025753_, _025815_);
  xor g_117360_(_001165_, _025753_, _025817_);
  and g_117361_(_025624_, _025738_, _025818_);
  not g_117362_(_025818_, _025819_);
  or g_117363_(_025627_, _025738_, _025820_);
  not g_117364_(_025820_, _025821_);
  and g_117365_(_025819_, _025820_, _025822_);
  or g_117366_(_025818_, _025821_, _025823_);
  and g_117367_(_025815_, _025823_, _025824_);
  or g_117368_(_025817_, _025822_, _025825_);
  xor g_117369_(out[822], _025752_, _025826_);
  xor g_117370_(_001176_, _025752_, _025828_);
  and g_117371_(_025615_, _025738_, _025829_);
  not g_117372_(_025829_, _025830_);
  or g_117373_(_025620_, _025738_, _025831_);
  not g_117374_(_025831_, _025832_);
  and g_117375_(_025830_, _025831_, _025833_);
  or g_117376_(_025829_, _025832_, _025834_);
  and g_117377_(_025826_, _025833_, _025835_);
  or g_117378_(_025828_, _025834_, _025836_);
  and g_117379_(_025825_, _025836_, _025837_);
  or g_117380_(_025824_, _025835_, _025839_);
  and g_117381_(_025817_, _025822_, _025840_);
  or g_117382_(_025815_, _025823_, _025841_);
  and g_117383_(_025828_, _025834_, _025842_);
  or g_117384_(_025826_, _025833_, _025843_);
  and g_117385_(_025841_, _025843_, _025844_);
  or g_117386_(_025840_, _025842_, _025845_);
  and g_117387_(_025837_, _025844_, _025846_);
  or g_117388_(_025839_, _025845_, _025847_);
  xor g_117389_(_001198_, out[819], _025848_);
  and g_117390_(_025650_, _025738_, _025850_);
  or g_117391_(_025655_, _025738_, _025851_);
  not g_117392_(_025851_, _025852_);
  or g_117393_(_025850_, _025852_, _025853_);
  and g_117394_(_025848_, _025853_, _025854_);
  not g_117395_(_025854_, _025855_);
  xor g_117396_(out[821], _025751_, _025856_);
  and g_117397_(_025643_, _025738_, _025857_);
  or g_117398_(_025647_, _025738_, _025858_);
  not g_117399_(_025858_, _025859_);
  or g_117400_(_025857_, _025859_, _025861_);
  and g_117401_(_025856_, _025861_, _025862_);
  not g_117402_(_025862_, _025863_);
  and g_117403_(_025855_, _025863_, _025864_);
  or g_117404_(_025854_, _025862_, _025865_);
  or g_117405_(_025856_, _025861_, _025866_);
  or g_117406_(_025848_, _025853_, _025867_);
  and g_117407_(_025866_, _025867_, _025868_);
  not g_117408_(_025868_, _025869_);
  and g_117409_(_025864_, _025868_, _025870_);
  or g_117410_(_025865_, _025869_, _025872_);
  and g_117411_(_025813_, _025870_, _025873_);
  or g_117412_(_025814_, _025872_, _025874_);
  and g_117413_(_025846_, _025873_, _025875_);
  or g_117414_(_025847_, _025874_, _025876_);
  and g_117415_(_025681_, _025740_, _025877_);
  and g_117416_(_001099_, _025738_, _025878_);
  or g_117417_(_025877_, _025878_, _025879_);
  or g_117418_(out[818], _025879_, _025880_);
  not g_117419_(_025880_, _025881_);
  and g_117420_(out[803], _025738_, _025883_);
  not g_117421_(_025883_, _025884_);
  or g_117422_(_025674_, _025738_, _025885_);
  not g_117423_(_025885_, _025886_);
  and g_117424_(_025884_, _025885_, _025887_);
  or g_117425_(_025883_, _025886_, _025888_);
  and g_117426_(out[819], _025887_, _025889_);
  or g_117427_(_001242_, _025888_, _025890_);
  and g_117428_(_025880_, _025890_, _025891_);
  or g_117429_(_025881_, _025889_, _025892_);
  and g_117430_(_001242_, _025888_, _025894_);
  or g_117431_(out[819], _025887_, _025895_);
  xor g_117432_(out[818], _025879_, _025896_);
  and g_117433_(_025895_, _025896_, _025897_);
  and g_117434_(_025890_, _025897_, _025898_);
  not g_117435_(_025898_, _025899_);
  or g_117436_(out[817], _025743_, _025900_);
  and g_117437_(_025693_, _025740_, _025901_);
  and g_117438_(_001088_, _025738_, _025902_);
  or g_117439_(_025901_, _025902_, _025903_);
  and g_117440_(out[816], _025903_, _025905_);
  xor g_117441_(_001209_, _025743_, _025906_);
  or g_117442_(_025905_, _025906_, _025907_);
  not g_117443_(_025907_, _025908_);
  and g_117444_(_025900_, _025907_, _025909_);
  not g_117445_(_025909_, _025910_);
  and g_117446_(_025898_, _025910_, _025911_);
  or g_117447_(_025899_, _025909_, _025912_);
  and g_117448_(_025892_, _025895_, _025913_);
  or g_117449_(_025891_, _025894_, _025914_);
  and g_117450_(_025912_, _025914_, _025916_);
  or g_117451_(_025911_, _025913_, _025917_);
  and g_117452_(_025875_, _025917_, _025918_);
  or g_117453_(_025876_, _025916_, _025919_);
  and g_117454_(_025865_, _025866_, _025920_);
  not g_117455_(_025920_, _025921_);
  and g_117456_(_025846_, _025920_, _025922_);
  or g_117457_(_025847_, _025921_, _025923_);
  and g_117458_(_025839_, _025841_, _025924_);
  or g_117459_(_025837_, _025840_, _025925_);
  and g_117460_(_025923_, _025925_, _025927_);
  or g_117461_(_025922_, _025924_, _025928_);
  and g_117462_(_025813_, _025928_, _025929_);
  or g_117463_(_025814_, _025927_, _025930_);
  and g_117464_(_025786_, _025801_, _025931_);
  and g_117465_(_025807_, _025931_, _025932_);
  not g_117466_(_025932_, _025933_);
  and g_117467_(_025770_, _025775_, _025934_);
  or g_117468_(_025769_, _025774_, _025935_);
  and g_117469_(_025933_, _025935_, _025936_);
  or g_117470_(_025932_, _025934_, _025938_);
  or g_117471_(_025929_, _025938_, _025939_);
  and g_117472_(_025919_, _025936_, _025940_);
  and g_117473_(_025930_, _025940_, _025941_);
  or g_117474_(_025918_, _025939_, _025942_);
  or g_117475_(out[816], _025903_, _025943_);
  and g_117476_(_025898_, _025943_, _025944_);
  not g_117477_(_025944_, _025945_);
  and g_117478_(_025908_, _025944_, _025946_);
  or g_117479_(_025907_, _025945_, _025947_);
  and g_117480_(_025875_, _025946_, _025949_);
  or g_117481_(_025876_, _025947_, _025950_);
  and g_117482_(_025942_, _025950_, _025951_);
  or g_117483_(_025941_, _025949_, _025952_);
  and g_117484_(_025743_, _025952_, _025953_);
  and g_117485_(_001209_, _025951_, _025954_);
  or g_117486_(_025953_, _025954_, _025955_);
  and g_117487_(_025879_, _025952_, _025956_);
  and g_117488_(_001231_, _025951_, _025957_);
  or g_117489_(_025956_, _025957_, _025958_);
  or g_117490_(out[834], _025958_, _025960_);
  or g_117491_(_001242_, _025952_, _025961_);
  not g_117492_(_025961_, _025962_);
  and g_117493_(_025888_, _025952_, _025963_);
  or g_117494_(_025887_, _025951_, _025964_);
  and g_117495_(_025961_, _025964_, _025965_);
  or g_117496_(_025962_, _025963_, _025966_);
  or g_117497_(_001374_, _025966_, _025967_);
  and g_117498_(_025960_, _025967_, _025968_);
  and g_117499_(_001374_, _025966_, _025969_);
  xor g_117500_(out[834], _025958_, _025971_);
  xor g_117501_(out[835], _025965_, _025972_);
  and g_117502_(_025971_, _025972_, _025973_);
  not g_117503_(_025973_, _025974_);
  or g_117504_(out[833], _025955_, _025975_);
  and g_117505_(_025903_, _025952_, _025976_);
  and g_117506_(_001220_, _025951_, _025977_);
  or g_117507_(_025976_, _025977_, _025978_);
  and g_117508_(out[832], _025978_, _025979_);
  not g_117509_(_025979_, _025980_);
  xor g_117510_(out[833], _025955_, _025982_);
  xor g_117511_(_001341_, _025955_, _025983_);
  and g_117512_(_025980_, _025982_, _025984_);
  or g_117513_(_025979_, _025983_, _025985_);
  and g_117514_(_025975_, _025985_, _025986_);
  or g_117515_(_025974_, _025986_, _025987_);
  or g_117516_(_025968_, _025969_, _025988_);
  and g_117517_(_025987_, _025988_, _025989_);
  or g_117518_(_025759_, _025952_, _025990_);
  not g_117519_(_025990_, _025991_);
  and g_117520_(_025749_, _025952_, _025993_);
  or g_117521_(_025748_, _025951_, _025994_);
  and g_117522_(_025990_, _025994_, _025995_);
  or g_117523_(_025991_, _025993_, _025996_);
  and g_117524_(out[836], out[835], _025997_);
  or g_117525_(out[837], _025997_, _025998_);
  or g_117526_(out[838], _025998_, _025999_);
  or g_117527_(out[839], _025999_, _026000_);
  or g_117528_(out[840], _026000_, _026001_);
  and g_117529_(out[841], _026001_, _026002_);
  or g_117530_(out[842], _026002_, _026004_);
  xor g_117531_(out[842], _026002_, _026005_);
  xor g_117532_(_001407_, _026002_, _026006_);
  and g_117533_(_025995_, _026005_, _026007_);
  or g_117534_(_025996_, _026006_, _026008_);
  and g_117535_(_025763_, _025765_, _026009_);
  or g_117536_(_025764_, _025766_, _026010_);
  xor g_117537_(out[843], _026004_, _026011_);
  not g_117538_(_026011_, _026012_);
  or g_117539_(_026010_, _026011_, _026013_);
  not g_117540_(_026013_, _026015_);
  and g_117541_(_026008_, _026013_, _026016_);
  or g_117542_(_026007_, _026015_, _026017_);
  and g_117543_(_025996_, _026006_, _026018_);
  and g_117544_(_026010_, _026011_, _026019_);
  or g_117545_(_026017_, _026019_, _026020_);
  or g_117546_(_026018_, _026020_, _026021_);
  xor g_117547_(out[840], _026000_, _026022_);
  not g_117548_(_026022_, _026023_);
  or g_117549_(_025787_, _025952_, _026024_);
  not g_117550_(_026024_, _026026_);
  and g_117551_(_025795_, _025952_, _026027_);
  not g_117552_(_026027_, _026028_);
  and g_117553_(_026024_, _026028_, _026029_);
  or g_117554_(_026026_, _026027_, _026030_);
  and g_117555_(_026022_, _026030_, _026031_);
  or g_117556_(_026023_, _026029_, _026032_);
  xor g_117557_(out[841], _026001_, _026033_);
  not g_117558_(_026033_, _026034_);
  or g_117559_(_025777_, _025952_, _026035_);
  not g_117560_(_026035_, _026037_);
  and g_117561_(_025784_, _025952_, _026038_);
  not g_117562_(_026038_, _026039_);
  and g_117563_(_026035_, _026039_, _026040_);
  or g_117564_(_026037_, _026038_, _026041_);
  and g_117565_(_026034_, _026041_, _026042_);
  or g_117566_(_026033_, _026040_, _026043_);
  and g_117567_(_026032_, _026043_, _026044_);
  or g_117568_(_026031_, _026042_, _026045_);
  and g_117569_(_026033_, _026040_, _026046_);
  and g_117570_(_026023_, _026029_, _026048_);
  or g_117571_(_026046_, _026048_, _026049_);
  or g_117572_(_026045_, _026049_, _026050_);
  or g_117573_(_026021_, _026050_, _026051_);
  not g_117574_(_026051_, _026052_);
  xor g_117575_(out[839], _025999_, _026053_);
  not g_117576_(_026053_, _026054_);
  and g_117577_(_025817_, _025951_, _026055_);
  or g_117578_(_025815_, _025952_, _026056_);
  and g_117579_(_025823_, _025952_, _026057_);
  or g_117580_(_025822_, _025951_, _026059_);
  and g_117581_(_026056_, _026059_, _026060_);
  or g_117582_(_026055_, _026057_, _026061_);
  and g_117583_(_026053_, _026061_, _026062_);
  or g_117584_(_026054_, _026060_, _026063_);
  xor g_117585_(out[838], _025998_, _026064_);
  not g_117586_(_026064_, _026065_);
  and g_117587_(_025826_, _025951_, _026066_);
  or g_117588_(_025828_, _025952_, _026067_);
  and g_117589_(_025834_, _025952_, _026068_);
  or g_117590_(_025833_, _025951_, _026070_);
  and g_117591_(_026067_, _026070_, _026071_);
  or g_117592_(_026066_, _026068_, _026072_);
  and g_117593_(_026064_, _026071_, _026073_);
  or g_117594_(_026065_, _026072_, _026074_);
  and g_117595_(_026063_, _026074_, _026075_);
  or g_117596_(_026062_, _026073_, _026076_);
  and g_117597_(_026054_, _026060_, _026077_);
  and g_117598_(_026065_, _026072_, _026078_);
  or g_117599_(_026077_, _026078_, _026079_);
  or g_117600_(_026076_, _026079_, _026081_);
  not g_117601_(_026081_, _026082_);
  xor g_117602_(out[836], out[835], _026083_);
  not g_117603_(_026083_, _026084_);
  or g_117604_(_025848_, _025952_, _026085_);
  not g_117605_(_026085_, _026086_);
  and g_117606_(_025853_, _025952_, _026087_);
  not g_117607_(_026087_, _026088_);
  and g_117608_(_026085_, _026088_, _026089_);
  or g_117609_(_026086_, _026087_, _026090_);
  and g_117610_(_026084_, _026090_, _026092_);
  or g_117611_(_026083_, _026089_, _026093_);
  xor g_117612_(out[837], _025997_, _026094_);
  xor g_117613_(_001319_, _025997_, _026095_);
  or g_117614_(_025856_, _025952_, _026096_);
  not g_117615_(_026096_, _026097_);
  and g_117616_(_025861_, _025952_, _026098_);
  not g_117617_(_026098_, _026099_);
  and g_117618_(_026096_, _026099_, _026100_);
  or g_117619_(_026097_, _026098_, _026101_);
  and g_117620_(_026094_, _026101_, _026103_);
  or g_117621_(_026095_, _026100_, _026104_);
  and g_117622_(_026093_, _026104_, _026105_);
  or g_117623_(_026092_, _026103_, _026106_);
  and g_117624_(_026095_, _026100_, _026107_);
  and g_117625_(_026083_, _026089_, _026108_);
  or g_117626_(_026107_, _026108_, _026109_);
  not g_117627_(_026109_, _026110_);
  and g_117628_(_026105_, _026110_, _026111_);
  or g_117629_(_026106_, _026109_, _026112_);
  and g_117630_(_026082_, _026111_, _026114_);
  or g_117631_(_026081_, _026112_, _026115_);
  and g_117632_(_026052_, _026114_, _026116_);
  or g_117633_(_026051_, _026115_, _026117_);
  or g_117634_(_025989_, _026117_, _026118_);
  or g_117635_(_026081_, _026105_, _026119_);
  or g_117636_(_026107_, _026119_, _026120_);
  or g_117637_(_026075_, _026077_, _026121_);
  and g_117638_(_026120_, _026121_, _026122_);
  or g_117639_(_026051_, _026122_, _026123_);
  or g_117640_(_026044_, _026046_, _026125_);
  or g_117641_(_026021_, _026125_, _026126_);
  or g_117642_(_026016_, _026019_, _026127_);
  and g_117643_(_026126_, _026127_, _026128_);
  and g_117644_(_026118_, _026128_, _026129_);
  and g_117645_(_026123_, _026129_, _026130_);
  or g_117646_(out[832], _025978_, _026131_);
  and g_117647_(_025973_, _026131_, _026132_);
  and g_117648_(_025984_, _026132_, _026133_);
  and g_117649_(_026116_, _026133_, _026134_);
  or g_117650_(_026130_, _026134_, _026136_);
  not g_117651_(_026136_, _026137_);
  and g_117652_(_025955_, _026136_, _026138_);
  and g_117653_(_001341_, _026137_, _026139_);
  or g_117654_(_026138_, _026139_, _026140_);
  and g_117655_(_026005_, _026137_, _026141_);
  and g_117656_(_025996_, _026136_, _026142_);
  or g_117657_(_026141_, _026142_, _026143_);
  and g_117658_(out[852], out[851], _026144_);
  or g_117659_(out[853], _026144_, _026145_);
  or g_117660_(out[854], _026145_, _026147_);
  or g_117661_(out[855], _026147_, _026148_);
  or g_117662_(out[856], _026148_, _026149_);
  and g_117663_(out[857], _026149_, _026150_);
  or g_117664_(out[858], _026150_, _026151_);
  xor g_117665_(_001539_, _026150_, _026152_);
  or g_117666_(_026143_, _026152_, _026153_);
  not g_117667_(_026153_, _026154_);
  and g_117668_(_026009_, _026011_, _026155_);
  or g_117669_(_026010_, _026012_, _026156_);
  xor g_117670_(out[859], _026151_, _026158_);
  xor g_117671_(_001418_, _026151_, _026159_);
  and g_117672_(_026155_, _026159_, _026160_);
  or g_117673_(_026156_, _026158_, _026161_);
  and g_117674_(_026153_, _026161_, _026162_);
  or g_117675_(_026154_, _026160_, _026163_);
  and g_117676_(_026156_, _026158_, _026164_);
  or g_117677_(_026155_, _026159_, _026165_);
  and g_117678_(_026143_, _026152_, _026166_);
  or g_117679_(_026164_, _026166_, _026167_);
  not g_117680_(_026167_, _026169_);
  and g_117681_(_026162_, _026169_, _026170_);
  or g_117682_(_026163_, _026167_, _026171_);
  and g_117683_(_026023_, _026137_, _026172_);
  and g_117684_(_026030_, _026136_, _026173_);
  or g_117685_(_026172_, _026173_, _026174_);
  xor g_117686_(out[856], _026148_, _026175_);
  and g_117687_(_026174_, _026175_, _026176_);
  not g_117688_(_026176_, _026177_);
  xor g_117689_(_001528_, _026149_, _026178_);
  and g_117690_(_026033_, _026137_, _026180_);
  and g_117691_(_026041_, _026136_, _026181_);
  or g_117692_(_026180_, _026181_, _026182_);
  and g_117693_(_026178_, _026182_, _026183_);
  not g_117694_(_026183_, _026184_);
  and g_117695_(_026177_, _026184_, _026185_);
  or g_117696_(_026176_, _026183_, _026186_);
  or g_117697_(_026178_, _026182_, _026187_);
  or g_117698_(_026174_, _026175_, _026188_);
  and g_117699_(_026187_, _026188_, _026189_);
  not g_117700_(_026189_, _026191_);
  and g_117701_(_026185_, _026189_, _026192_);
  or g_117702_(_026186_, _026191_, _026193_);
  and g_117703_(_026170_, _026192_, _026194_);
  or g_117704_(_026171_, _026193_, _026195_);
  xor g_117705_(out[855], _026147_, _026196_);
  not g_117706_(_026196_, _026197_);
  and g_117707_(_026054_, _026137_, _026198_);
  and g_117708_(_026061_, _026136_, _026199_);
  or g_117709_(_026198_, _026199_, _026200_);
  not g_117710_(_026200_, _026202_);
  and g_117711_(_026196_, _026200_, _026203_);
  xor g_117712_(out[854], _026145_, _026204_);
  not g_117713_(_026204_, _026205_);
  and g_117714_(_026064_, _026137_, _026206_);
  or g_117715_(_026065_, _026136_, _026207_);
  and g_117716_(_026072_, _026136_, _026208_);
  or g_117717_(_026071_, _026137_, _026209_);
  and g_117718_(_026207_, _026209_, _026210_);
  or g_117719_(_026206_, _026208_, _026211_);
  and g_117720_(_026204_, _026210_, _026213_);
  or g_117721_(_026203_, _026213_, _026214_);
  and g_117722_(_026197_, _026202_, _026215_);
  or g_117723_(_026196_, _026200_, _026216_);
  and g_117724_(_026205_, _026211_, _026217_);
  or g_117725_(_026214_, _026217_, _026218_);
  xor g_117726_(_026196_, _026200_, _026219_);
  xor g_117727_(_026204_, _026210_, _026220_);
  and g_117728_(_026219_, _026220_, _026221_);
  or g_117729_(_026215_, _026218_, _026222_);
  xor g_117730_(out[853], _026144_, _026224_);
  and g_117731_(_026095_, _026137_, _026225_);
  and g_117732_(_026101_, _026136_, _026226_);
  or g_117733_(_026225_, _026226_, _026227_);
  and g_117734_(_026224_, _026227_, _026228_);
  not g_117735_(_026228_, _026229_);
  xor g_117736_(_001462_, out[851], _026230_);
  and g_117737_(_026083_, _026137_, _026231_);
  and g_117738_(_026090_, _026136_, _026232_);
  or g_117739_(_026231_, _026232_, _026233_);
  and g_117740_(_026230_, _026233_, _026235_);
  not g_117741_(_026235_, _026236_);
  and g_117742_(_026229_, _026236_, _026237_);
  or g_117743_(_026228_, _026235_, _026238_);
  or g_117744_(_026224_, _026227_, _026239_);
  or g_117745_(_026230_, _026233_, _026240_);
  and g_117746_(_026239_, _026240_, _026241_);
  not g_117747_(_026241_, _026242_);
  and g_117748_(_026237_, _026241_, _026243_);
  or g_117749_(_026238_, _026242_, _026244_);
  and g_117750_(_026221_, _026243_, _026246_);
  or g_117751_(_026222_, _026244_, _026247_);
  and g_117752_(_025965_, _026136_, _026248_);
  not g_117753_(_026248_, _026249_);
  or g_117754_(out[835], _026136_, _026250_);
  not g_117755_(_026250_, _026251_);
  or g_117756_(_026248_, _026251_, _026252_);
  and g_117757_(_026249_, _026250_, _026253_);
  and g_117758_(out[851], _026252_, _026254_);
  or g_117759_(_001506_, _026253_, _026255_);
  and g_117760_(_025958_, _026136_, _026257_);
  and g_117761_(_001363_, _026137_, _026258_);
  or g_117762_(_026257_, _026258_, _026259_);
  not g_117763_(_026259_, _026260_);
  or g_117764_(out[850], _026259_, _026261_);
  not g_117765_(_026261_, _026262_);
  and g_117766_(_026255_, _026261_, _026263_);
  or g_117767_(_026254_, _026262_, _026264_);
  and g_117768_(_001506_, _026253_, _026265_);
  or g_117769_(out[851], _026252_, _026266_);
  and g_117770_(out[850], _026259_, _026268_);
  or g_117771_(_001495_, _026260_, _026269_);
  and g_117772_(_026266_, _026269_, _026270_);
  or g_117773_(_026265_, _026268_, _026271_);
  and g_117774_(_026263_, _026270_, _026272_);
  or g_117775_(_026264_, _026271_, _026273_);
  or g_117776_(out[849], _026140_, _026274_);
  not g_117777_(_026274_, _026275_);
  and g_117778_(_025978_, _026136_, _026276_);
  not g_117779_(_026276_, _026277_);
  or g_117780_(out[832], _026136_, _026279_);
  not g_117781_(_026279_, _026280_);
  and g_117782_(_026277_, _026279_, _026281_);
  or g_117783_(_026276_, _026280_, _026282_);
  and g_117784_(out[848], _026282_, _026283_);
  or g_117785_(_001484_, _026281_, _026284_);
  xor g_117786_(out[849], _026140_, _026285_);
  xor g_117787_(_001473_, _026140_, _026286_);
  and g_117788_(_026284_, _026285_, _026287_);
  or g_117789_(_026283_, _026286_, _026288_);
  and g_117790_(_026274_, _026288_, _026290_);
  or g_117791_(_026275_, _026287_, _026291_);
  and g_117792_(_026272_, _026291_, _026292_);
  or g_117793_(_026273_, _026290_, _026293_);
  and g_117794_(_026262_, _026266_, _026294_);
  or g_117795_(_026261_, _026265_, _026295_);
  and g_117796_(_026255_, _026295_, _026296_);
  or g_117797_(_026254_, _026294_, _026297_);
  and g_117798_(_026293_, _026296_, _026298_);
  or g_117799_(_026292_, _026297_, _026299_);
  and g_117800_(_026246_, _026299_, _026301_);
  or g_117801_(_026247_, _026298_, _026302_);
  and g_117802_(_026214_, _026216_, _026303_);
  and g_117803_(_026238_, _026239_, _026304_);
  and g_117804_(_026221_, _026304_, _026305_);
  or g_117805_(_026303_, _026305_, _026306_);
  not g_117806_(_026306_, _026307_);
  and g_117807_(_026302_, _026307_, _026308_);
  or g_117808_(_026301_, _026306_, _026309_);
  and g_117809_(_026194_, _026309_, _026310_);
  or g_117810_(_026195_, _026308_, _026312_);
  and g_117811_(_026163_, _026165_, _026313_);
  or g_117812_(_026162_, _026164_, _026314_);
  and g_117813_(_026186_, _026187_, _026315_);
  not g_117814_(_026315_, _026316_);
  and g_117815_(_026170_, _026315_, _026317_);
  or g_117816_(_026171_, _026316_, _026318_);
  and g_117817_(_026314_, _026318_, _026319_);
  or g_117818_(_026313_, _026317_, _026320_);
  and g_117819_(_026312_, _026319_, _026321_);
  or g_117820_(_026310_, _026320_, _026323_);
  or g_117821_(out[848], _026282_, _026324_);
  not g_117822_(_026324_, _026325_);
  or g_117823_(_026273_, _026288_, _026326_);
  not g_117824_(_026326_, _026327_);
  and g_117825_(_026324_, _026327_, _026328_);
  or g_117826_(_026325_, _026326_, _026329_);
  and g_117827_(_026194_, _026246_, _026330_);
  or g_117828_(_026195_, _026247_, _026331_);
  and g_117829_(_026328_, _026330_, _026332_);
  or g_117830_(_026329_, _026331_, _026334_);
  and g_117831_(_026323_, _026334_, _026335_);
  or g_117832_(_026321_, _026332_, _026336_);
  and g_117833_(_026140_, _026336_, _026337_);
  and g_117834_(_001473_, _026335_, _026338_);
  or g_117835_(_026337_, _026338_, _026339_);
  and g_117836_(_026143_, _026336_, _026340_);
  not g_117837_(_026340_, _026341_);
  or g_117838_(_026152_, _026336_, _026342_);
  not g_117839_(_026342_, _026343_);
  and g_117840_(_026341_, _026342_, _026345_);
  or g_117841_(_026340_, _026343_, _026346_);
  and g_117842_(out[868], out[867], _026347_);
  or g_117843_(out[869], _026347_, _026348_);
  or g_117844_(out[870], _026348_, _026349_);
  or g_117845_(out[871], _026349_, _026350_);
  or g_117846_(out[872], _026350_, _026351_);
  and g_117847_(out[873], _026351_, _026352_);
  or g_117848_(out[874], _026352_, _026353_);
  xor g_117849_(out[874], _026352_, _026354_);
  not g_117850_(_026354_, _026356_);
  or g_117851_(_026346_, _026356_, _026357_);
  and g_117852_(_026155_, _026158_, _026358_);
  or g_117853_(_026156_, _026159_, _026359_);
  xor g_117854_(out[875], _026353_, _026360_);
  xor g_117855_(_001550_, _026353_, _026361_);
  or g_117856_(_026359_, _026360_, _026362_);
  and g_117857_(_026357_, _026362_, _026363_);
  or g_117858_(_026345_, _026354_, _026364_);
  and g_117859_(_026359_, _026360_, _026365_);
  xor g_117860_(out[873], _026351_, _026367_);
  and g_117861_(_026182_, _026336_, _026368_);
  not g_117862_(_026368_, _026369_);
  or g_117863_(_026178_, _026336_, _026370_);
  not g_117864_(_026370_, _026371_);
  and g_117865_(_026369_, _026370_, _026372_);
  or g_117866_(_026368_, _026371_, _026373_);
  and g_117867_(_026367_, _026372_, _026374_);
  not g_117868_(_026374_, _026375_);
  xor g_117869_(out[872], _026350_, _026376_);
  not g_117870_(_026376_, _026378_);
  and g_117871_(_026174_, _026336_, _026379_);
  not g_117872_(_026379_, _026380_);
  or g_117873_(_026175_, _026336_, _026381_);
  not g_117874_(_026381_, _026382_);
  and g_117875_(_026380_, _026381_, _026383_);
  or g_117876_(_026379_, _026382_, _026384_);
  or g_117877_(_026378_, _026383_, _026385_);
  or g_117878_(_026367_, _026372_, _026386_);
  and g_117879_(_026385_, _026386_, _026387_);
  not g_117880_(_026387_, _026389_);
  and g_117881_(_026378_, _026383_, _026390_);
  or g_117882_(_026376_, _026384_, _026391_);
  and g_117883_(_026363_, _026364_, _026392_);
  not g_117884_(_026392_, _026393_);
  or g_117885_(_026365_, _026393_, _026394_);
  not g_117886_(_026394_, _026395_);
  and g_117887_(_026375_, _026391_, _026396_);
  or g_117888_(_026374_, _026390_, _026397_);
  and g_117889_(_026387_, _026396_, _026398_);
  or g_117890_(_026389_, _026397_, _026400_);
  and g_117891_(_026395_, _026398_, _026401_);
  or g_117892_(_026394_, _026400_, _026402_);
  xor g_117893_(out[870], _026348_, _026403_);
  xor g_117894_(_001572_, _026348_, _026404_);
  and g_117895_(_026211_, _026336_, _026405_);
  or g_117896_(_026210_, _026335_, _026406_);
  or g_117897_(_026205_, _026336_, _026407_);
  not g_117898_(_026407_, _026408_);
  and g_117899_(_026406_, _026407_, _026409_);
  or g_117900_(_026405_, _026408_, _026411_);
  and g_117901_(_026403_, _026409_, _026412_);
  or g_117902_(_026404_, _026411_, _026413_);
  xor g_117903_(out[871], _026349_, _026414_);
  xor g_117904_(_001561_, _026349_, _026415_);
  and g_117905_(_026200_, _026336_, _026416_);
  not g_117906_(_026416_, _026417_);
  and g_117907_(_026197_, _026335_, _026418_);
  or g_117908_(_026196_, _026336_, _026419_);
  and g_117909_(_026417_, _026419_, _026420_);
  or g_117910_(_026416_, _026418_, _026422_);
  and g_117911_(_026414_, _026422_, _026423_);
  or g_117912_(_026415_, _026420_, _026424_);
  and g_117913_(_026413_, _026424_, _026425_);
  or g_117914_(_026412_, _026423_, _026426_);
  and g_117915_(_026404_, _026411_, _026427_);
  not g_117916_(_026427_, _026428_);
  and g_117917_(_026415_, _026420_, _026429_);
  not g_117918_(_026429_, _026430_);
  xor g_117919_(out[869], _026347_, _026431_);
  xor g_117920_(_001583_, _026347_, _026433_);
  and g_117921_(_026227_, _026336_, _026434_);
  not g_117922_(_026434_, _026435_);
  or g_117923_(_026224_, _026336_, _026436_);
  not g_117924_(_026436_, _026437_);
  and g_117925_(_026435_, _026436_, _026438_);
  or g_117926_(_026434_, _026437_, _026439_);
  and g_117927_(_026433_, _026438_, _026440_);
  not g_117928_(_026440_, _026441_);
  xor g_117929_(out[868], out[867], _026442_);
  not g_117930_(_026442_, _026444_);
  or g_117931_(_026230_, _026336_, _026445_);
  not g_117932_(_026445_, _026446_);
  and g_117933_(_026233_, _026336_, _026447_);
  not g_117934_(_026447_, _026448_);
  and g_117935_(_026445_, _026448_, _026449_);
  or g_117936_(_026446_, _026447_, _026450_);
  and g_117937_(_026442_, _026449_, _026451_);
  or g_117938_(_026444_, _026450_, _026452_);
  and g_117939_(_026444_, _026450_, _026453_);
  or g_117940_(_026442_, _026449_, _026455_);
  and g_117941_(_026431_, _026439_, _026456_);
  or g_117942_(_026433_, _026438_, _026457_);
  and g_117943_(_026455_, _026457_, _026458_);
  or g_117944_(_026453_, _026456_, _026459_);
  and g_117945_(_026441_, _026458_, _026460_);
  or g_117946_(_026440_, _026459_, _026461_);
  and g_117947_(_026425_, _026428_, _026462_);
  or g_117948_(_026426_, _026427_, _026463_);
  and g_117949_(_026430_, _026462_, _026464_);
  or g_117950_(_026429_, _026463_, _026466_);
  and g_117951_(_026452_, _026460_, _026467_);
  or g_117952_(_026451_, _026461_, _026468_);
  and g_117953_(_026464_, _026467_, _026469_);
  or g_117954_(_026466_, _026468_, _026470_);
  or g_117955_(_001506_, _026336_, _026471_);
  not g_117956_(_026471_, _026472_);
  and g_117957_(_026253_, _026336_, _026473_);
  or g_117958_(_026252_, _026335_, _026474_);
  and g_117959_(_026471_, _026474_, _026475_);
  or g_117960_(_026472_, _026473_, _026477_);
  or g_117961_(_001638_, _026477_, _026478_);
  and g_117962_(_026259_, _026336_, _026479_);
  and g_117963_(_001495_, _026335_, _026480_);
  or g_117964_(_026479_, _026480_, _026481_);
  and g_117965_(_001638_, _026477_, _026482_);
  or g_117966_(out[866], _026481_, _026483_);
  xor g_117967_(out[867], _026475_, _026484_);
  xor g_117968_(out[866], _026481_, _026485_);
  and g_117969_(_026484_, _026485_, _026486_);
  not g_117970_(_026486_, _026488_);
  or g_117971_(out[865], _026339_, _026489_);
  and g_117972_(_026282_, _026336_, _026490_);
  and g_117973_(_001484_, _026335_, _026491_);
  or g_117974_(_026490_, _026491_, _026492_);
  and g_117975_(out[864], _026492_, _026493_);
  not g_117976_(_026493_, _026494_);
  xor g_117977_(out[865], _026339_, _026495_);
  xor g_117978_(_001605_, _026339_, _026496_);
  and g_117979_(_026494_, _026495_, _026497_);
  or g_117980_(_026493_, _026496_, _026499_);
  and g_117981_(_026489_, _026499_, _026500_);
  or g_117982_(_026488_, _026500_, _026501_);
  or g_117983_(_026482_, _026483_, _026502_);
  and g_117984_(_026478_, _026502_, _026503_);
  and g_117985_(_026501_, _026503_, _026504_);
  or g_117986_(_026470_, _026504_, _026505_);
  or g_117987_(_026458_, _026466_, _026506_);
  or g_117988_(_026440_, _026506_, _026507_);
  or g_117989_(_026425_, _026429_, _026508_);
  and g_117990_(_026507_, _026508_, _026510_);
  and g_117991_(_026505_, _026510_, _026511_);
  or g_117992_(_026402_, _026511_, _026512_);
  or g_117993_(_026374_, _026387_, _026513_);
  or g_117994_(_026394_, _026513_, _026514_);
  or g_117995_(_026363_, _026365_, _026515_);
  and g_117996_(_026514_, _026515_, _026516_);
  and g_117997_(_026512_, _026516_, _026517_);
  or g_117998_(out[864], _026492_, _026518_);
  and g_117999_(_026486_, _026518_, _026519_);
  and g_118000_(_026497_, _026519_, _026521_);
  and g_118001_(_026401_, _026521_, _026522_);
  and g_118002_(_026469_, _026522_, _026523_);
  or g_118003_(_026517_, _026523_, _026524_);
  not g_118004_(_026524_, _026525_);
  and g_118005_(_026339_, _026524_, _026526_);
  not g_118006_(_026526_, _026527_);
  or g_118007_(out[865], _026524_, _026528_);
  not g_118008_(_026528_, _026529_);
  and g_118009_(_026527_, _026528_, _026530_);
  or g_118010_(_026526_, _026529_, _026532_);
  and g_118011_(_026358_, _026360_, _026533_);
  or g_118012_(_026359_, _026361_, _026534_);
  and g_118013_(out[884], out[883], _026535_);
  or g_118014_(out[885], _026535_, _026536_);
  or g_118015_(out[886], _026536_, _026537_);
  or g_118016_(out[887], _026537_, _026538_);
  or g_118017_(out[888], _026538_, _026539_);
  and g_118018_(out[889], _026539_, _026540_);
  or g_118019_(out[890], _026540_, _026541_);
  xor g_118020_(out[891], _026541_, _026543_);
  xor g_118021_(_001682_, _026541_, _026544_);
  and g_118022_(_026533_, _026544_, _026545_);
  or g_118023_(_026534_, _026543_, _026546_);
  and g_118024_(_026354_, _026525_, _026547_);
  or g_118025_(_026356_, _026524_, _026548_);
  and g_118026_(_026346_, _026524_, _026549_);
  or g_118027_(_026345_, _026525_, _026550_);
  and g_118028_(_026548_, _026550_, _026551_);
  or g_118029_(_026547_, _026549_, _026552_);
  xor g_118030_(out[890], _026540_, _026554_);
  xor g_118031_(_001803_, _026540_, _026555_);
  and g_118032_(_026551_, _026554_, _026556_);
  or g_118033_(_026552_, _026555_, _026557_);
  and g_118034_(_026546_, _026557_, _026558_);
  or g_118035_(_026545_, _026556_, _026559_);
  and g_118036_(_026534_, _026543_, _026560_);
  or g_118037_(_026533_, _026544_, _026561_);
  and g_118038_(_026552_, _026555_, _026562_);
  or g_118039_(_026551_, _026554_, _026563_);
  and g_118040_(_026561_, _026563_, _026565_);
  or g_118041_(_026560_, _026562_, _026566_);
  and g_118042_(_026558_, _026565_, _026567_);
  or g_118043_(_026559_, _026566_, _026568_);
  xor g_118044_(out[888], _026538_, _026569_);
  xor g_118045_(_001781_, _026538_, _026570_);
  or g_118046_(_026376_, _026524_, _026571_);
  not g_118047_(_026571_, _026572_);
  and g_118048_(_026384_, _026524_, _026573_);
  or g_118049_(_026383_, _026525_, _026574_);
  and g_118050_(_026571_, _026574_, _026576_);
  or g_118051_(_026572_, _026573_, _026577_);
  and g_118052_(_026569_, _026577_, _026578_);
  or g_118053_(_026570_, _026576_, _026579_);
  xor g_118054_(out[889], _026539_, _026580_);
  xor g_118055_(_001792_, _026539_, _026581_);
  and g_118056_(_026372_, _026524_, _026582_);
  or g_118057_(_026373_, _026525_, _026583_);
  or g_118058_(_026367_, _026524_, _026584_);
  not g_118059_(_026584_, _026585_);
  or g_118060_(_026582_, _026585_, _026587_);
  and g_118061_(_026583_, _026584_, _026588_);
  and g_118062_(_026581_, _026588_, _026589_);
  or g_118063_(_026580_, _026587_, _026590_);
  and g_118064_(_026579_, _026590_, _026591_);
  or g_118065_(_026578_, _026589_, _026592_);
  and g_118066_(_026580_, _026587_, _026593_);
  or g_118067_(_026581_, _026588_, _026594_);
  and g_118068_(_026570_, _026576_, _026595_);
  or g_118069_(_026569_, _026577_, _026596_);
  and g_118070_(_026594_, _026596_, _026598_);
  or g_118071_(_026593_, _026595_, _026599_);
  and g_118072_(_026591_, _026598_, _026600_);
  or g_118073_(_026592_, _026599_, _026601_);
  and g_118074_(_026567_, _026600_, _026602_);
  or g_118075_(_026568_, _026601_, _026603_);
  xor g_118076_(out[886], _026536_, _026604_);
  xor g_118077_(_001704_, _026536_, _026605_);
  or g_118078_(_026404_, _026524_, _026606_);
  not g_118079_(_026606_, _026607_);
  and g_118080_(_026411_, _026524_, _026609_);
  not g_118081_(_026609_, _026610_);
  and g_118082_(_026606_, _026610_, _026611_);
  or g_118083_(_026607_, _026609_, _026612_);
  and g_118084_(_026604_, _026611_, _026613_);
  or g_118085_(_026605_, _026612_, _026614_);
  xor g_118086_(out[887], _026537_, _026615_);
  xor g_118087_(_001693_, _026537_, _026616_);
  and g_118088_(_026420_, _026524_, _026617_);
  not g_118089_(_026617_, _026618_);
  and g_118090_(_026414_, _026525_, _026620_);
  or g_118091_(_026415_, _026524_, _026621_);
  or g_118092_(_026617_, _026620_, _026622_);
  and g_118093_(_026618_, _026621_, _026623_);
  and g_118094_(_026615_, _026623_, _026624_);
  or g_118095_(_026616_, _026622_, _026625_);
  and g_118096_(_026614_, _026625_, _026626_);
  or g_118097_(_026613_, _026624_, _026627_);
  and g_118098_(_026605_, _026612_, _026628_);
  or g_118099_(_026604_, _026611_, _026629_);
  and g_118100_(_026616_, _026622_, _026631_);
  or g_118101_(_026615_, _026623_, _026632_);
  xor g_118102_(out[885], _026535_, _026633_);
  xor g_118103_(_001715_, _026535_, _026634_);
  or g_118104_(_026431_, _026524_, _026635_);
  not g_118105_(_026635_, _026636_);
  and g_118106_(_026439_, _026524_, _026637_);
  or g_118107_(_026438_, _026525_, _026638_);
  and g_118108_(_026635_, _026638_, _026639_);
  or g_118109_(_026636_, _026637_, _026640_);
  and g_118110_(_026634_, _026639_, _026642_);
  or g_118111_(_026633_, _026640_, _026643_);
  xor g_118112_(out[884], out[883], _026644_);
  xor g_118113_(_001726_, out[883], _026645_);
  and g_118114_(_026442_, _026525_, _026646_);
  or g_118115_(_026444_, _026524_, _026647_);
  and g_118116_(_026450_, _026524_, _026648_);
  or g_118117_(_026449_, _026525_, _026649_);
  and g_118118_(_026647_, _026649_, _026650_);
  or g_118119_(_026646_, _026648_, _026651_);
  and g_118120_(_026644_, _026650_, _026653_);
  or g_118121_(_026645_, _026651_, _026654_);
  and g_118122_(_026645_, _026651_, _026655_);
  or g_118123_(_026644_, _026650_, _026656_);
  and g_118124_(_026633_, _026640_, _026657_);
  or g_118125_(_026634_, _026639_, _026658_);
  and g_118126_(_026656_, _026658_, _026659_);
  or g_118127_(_026655_, _026657_, _026660_);
  and g_118128_(_026643_, _026659_, _026661_);
  or g_118129_(_026642_, _026660_, _026662_);
  and g_118130_(_026626_, _026629_, _026664_);
  or g_118131_(_026627_, _026628_, _026665_);
  and g_118132_(_026632_, _026664_, _026666_);
  or g_118133_(_026631_, _026665_, _026667_);
  and g_118134_(_026654_, _026661_, _026668_);
  or g_118135_(_026653_, _026662_, _026669_);
  and g_118136_(_026666_, _026668_, _026670_);
  or g_118137_(_026667_, _026669_, _026671_);
  and g_118138_(_026481_, _026524_, _026672_);
  not g_118139_(_026672_, _026673_);
  or g_118140_(out[866], _026524_, _026675_);
  not g_118141_(_026675_, _026676_);
  and g_118142_(_026673_, _026675_, _026677_);
  or g_118143_(_026672_, _026676_, _026678_);
  and g_118144_(_001759_, _026677_, _026679_);
  or g_118145_(out[882], _026678_, _026680_);
  and g_118146_(_026475_, _026524_, _026681_);
  not g_118147_(_026681_, _026682_);
  or g_118148_(out[867], _026524_, _026683_);
  not g_118149_(_026683_, _026684_);
  or g_118150_(_026681_, _026684_, _026686_);
  and g_118151_(_026682_, _026683_, _026687_);
  and g_118152_(out[883], _026686_, _026688_);
  or g_118153_(_001770_, _026687_, _026689_);
  and g_118154_(_026680_, _026689_, _026690_);
  or g_118155_(_026679_, _026688_, _026691_);
  and g_118156_(_001770_, _026687_, _026692_);
  or g_118157_(out[883], _026686_, _026693_);
  and g_118158_(out[882], _026678_, _026694_);
  or g_118159_(_001759_, _026677_, _026695_);
  and g_118160_(_026693_, _026695_, _026697_);
  or g_118161_(_026692_, _026694_, _026698_);
  and g_118162_(_026690_, _026697_, _026699_);
  or g_118163_(_026691_, _026698_, _026700_);
  and g_118164_(_001737_, _026530_, _026701_);
  or g_118165_(out[881], _026532_, _026702_);
  and g_118166_(_026492_, _026524_, _026703_);
  not g_118167_(_026703_, _026704_);
  or g_118168_(out[864], _026524_, _026705_);
  not g_118169_(_026705_, _026706_);
  and g_118170_(_026704_, _026705_, _026708_);
  or g_118171_(_026703_, _026706_, _026709_);
  and g_118172_(out[880], _026709_, _026710_);
  or g_118173_(_001748_, _026708_, _026711_);
  xor g_118174_(_001737_, _026530_, _026712_);
  xor g_118175_(out[881], _026530_, _026713_);
  and g_118176_(_026711_, _026712_, _026714_);
  or g_118177_(_026710_, _026713_, _026715_);
  and g_118178_(_026702_, _026715_, _026716_);
  or g_118179_(_026701_, _026714_, _026717_);
  and g_118180_(_026699_, _026717_, _026719_);
  or g_118181_(_026700_, _026716_, _026720_);
  and g_118182_(_026679_, _026693_, _026721_);
  or g_118183_(_026680_, _026692_, _026722_);
  and g_118184_(_026689_, _026722_, _026723_);
  or g_118185_(_026688_, _026721_, _026724_);
  and g_118186_(_026720_, _026723_, _026725_);
  or g_118187_(_026719_, _026724_, _026726_);
  and g_118188_(_026670_, _026726_, _026727_);
  or g_118189_(_026671_, _026725_, _026728_);
  and g_118190_(_026660_, _026666_, _026730_);
  or g_118191_(_026659_, _026667_, _026731_);
  and g_118192_(_026643_, _026730_, _026732_);
  or g_118193_(_026642_, _026731_, _026733_);
  and g_118194_(_026627_, _026632_, _026734_);
  or g_118195_(_026626_, _026631_, _026735_);
  and g_118196_(_026733_, _026735_, _026736_);
  or g_118197_(_026732_, _026734_, _026737_);
  and g_118198_(_026728_, _026736_, _026738_);
  or g_118199_(_026727_, _026737_, _026739_);
  and g_118200_(_026602_, _026739_, _026741_);
  or g_118201_(_026603_, _026738_, _026742_);
  and g_118202_(_026592_, _026594_, _026743_);
  or g_118203_(_026591_, _026593_, _026744_);
  and g_118204_(_026567_, _026743_, _026745_);
  or g_118205_(_026568_, _026744_, _026746_);
  and g_118206_(_026559_, _026561_, _026747_);
  or g_118207_(_026558_, _026560_, _026748_);
  and g_118208_(_026746_, _026748_, _026749_);
  or g_118209_(_026745_, _026747_, _026750_);
  and g_118210_(_026742_, _026749_, _026752_);
  or g_118211_(_026741_, _026750_, _026753_);
  and g_118212_(_001748_, _026708_, _026754_);
  or g_118213_(out[880], _026709_, _026755_);
  and g_118214_(_026699_, _026714_, _026756_);
  or g_118215_(_026700_, _026715_, _026757_);
  and g_118216_(_026755_, _026756_, _026758_);
  or g_118217_(_026754_, _026757_, _026759_);
  and g_118218_(_026602_, _026758_, _026760_);
  or g_118219_(_026603_, _026759_, _026761_);
  and g_118220_(_026670_, _026760_, _026763_);
  or g_118221_(_026671_, _026761_, _026764_);
  and g_118222_(_026753_, _026764_, _026765_);
  or g_118223_(_026752_, _026763_, _026766_);
  and g_118224_(_026532_, _026766_, _026767_);
  and g_118225_(_001737_, _026765_, _026768_);
  or g_118226_(_026767_, _026768_, _026769_);
  or g_118227_(_026555_, _026766_, _026770_);
  not g_118228_(_026770_, _026771_);
  and g_118229_(_026552_, _026766_, _026772_);
  or g_118230_(_026551_, _026765_, _026774_);
  and g_118231_(_026770_, _026774_, _026775_);
  or g_118232_(_026771_, _026772_, _026776_);
  and g_118233_(out[900], out[899], _026777_);
  or g_118234_(out[901], _026777_, _026778_);
  or g_118235_(out[902], _026778_, _026779_);
  or g_118236_(out[903], _026779_, _026780_);
  or g_118237_(out[904], _026780_, _026781_);
  and g_118238_(out[905], _026781_, _026782_);
  or g_118239_(out[906], _026782_, _026783_);
  xor g_118240_(out[906], _026782_, _026785_);
  not g_118241_(_026785_, _026786_);
  and g_118242_(_026775_, _026785_, _026787_);
  or g_118243_(_026776_, _026786_, _026788_);
  and g_118244_(_026533_, _026543_, _026789_);
  or g_118245_(_026534_, _026544_, _026790_);
  xor g_118246_(out[907], _026783_, _026791_);
  xor g_118247_(_001814_, _026783_, _026792_);
  and g_118248_(_026789_, _026792_, _026793_);
  or g_118249_(_026790_, _026791_, _026794_);
  and g_118250_(_026788_, _026794_, _026796_);
  or g_118251_(_026787_, _026793_, _026797_);
  and g_118252_(_026776_, _026786_, _026798_);
  and g_118253_(_026790_, _026791_, _026799_);
  xor g_118254_(out[905], _026781_, _026800_);
  or g_118255_(_026581_, _026766_, _026801_);
  not g_118256_(_026801_, _026802_);
  and g_118257_(_026588_, _026766_, _026803_);
  not g_118258_(_026803_, _026804_);
  and g_118259_(_026801_, _026804_, _026805_);
  or g_118260_(_026802_, _026803_, _026807_);
  and g_118261_(_026800_, _026805_, _026808_);
  or g_118262_(_026797_, _026798_, _026809_);
  or g_118263_(_026799_, _026809_, _026810_);
  or g_118264_(_026808_, _026810_, _026811_);
  or g_118265_(_026800_, _026805_, _026812_);
  or g_118266_(_026569_, _026766_, _026813_);
  not g_118267_(_026813_, _026814_);
  and g_118268_(_026577_, _026766_, _026815_);
  not g_118269_(_026815_, _026816_);
  and g_118270_(_026813_, _026816_, _026818_);
  or g_118271_(_026814_, _026815_, _026819_);
  xor g_118272_(out[904], _026780_, _026820_);
  not g_118273_(_026820_, _026821_);
  or g_118274_(_026818_, _026821_, _026822_);
  and g_118275_(_026812_, _026822_, _026823_);
  or g_118276_(_026819_, _026820_, _026824_);
  and g_118277_(_026823_, _026824_, _026825_);
  not g_118278_(_026825_, _026826_);
  or g_118279_(_026811_, _026826_, _026827_);
  not g_118280_(_026827_, _026829_);
  xor g_118281_(_001847_, _026777_, _026830_);
  or g_118282_(_026633_, _026766_, _026831_);
  not g_118283_(_026831_, _026832_);
  and g_118284_(_026640_, _026766_, _026833_);
  not g_118285_(_026833_, _026834_);
  and g_118286_(_026831_, _026834_, _026835_);
  or g_118287_(_026832_, _026833_, _026836_);
  and g_118288_(_026830_, _026835_, _026837_);
  xor g_118289_(out[900], out[899], _026838_);
  or g_118290_(_026645_, _026766_, _026840_);
  or g_118291_(_026650_, _026765_, _026841_);
  and g_118292_(_026840_, _026841_, _026842_);
  and g_118293_(_026838_, _026842_, _026843_);
  or g_118294_(_026837_, _026843_, _026844_);
  xor g_118295_(out[902], _026778_, _026845_);
  not g_118296_(_026845_, _026846_);
  and g_118297_(_026604_, _026765_, _026847_);
  and g_118298_(_026612_, _026766_, _026848_);
  or g_118299_(_026847_, _026848_, _026849_);
  and g_118300_(_026846_, _026849_, _026851_);
  xor g_118301_(out[903], _026779_, _026852_);
  not g_118302_(_026852_, _026853_);
  or g_118303_(_026615_, _026766_, _026854_);
  or g_118304_(_026622_, _026765_, _026855_);
  and g_118305_(_026854_, _026855_, _026856_);
  and g_118306_(_026853_, _026856_, _026857_);
  or g_118307_(_026851_, _026857_, _026858_);
  or g_118308_(_026844_, _026858_, _026859_);
  not g_118309_(_026859_, _026860_);
  or g_118310_(_026846_, _026849_, _026862_);
  or g_118311_(_026853_, _026856_, _026863_);
  and g_118312_(_026862_, _026863_, _026864_);
  or g_118313_(_026830_, _026835_, _026865_);
  or g_118314_(_026838_, _026842_, _026866_);
  and g_118315_(_026865_, _026866_, _026867_);
  and g_118316_(_026864_, _026867_, _026868_);
  not g_118317_(_026868_, _026869_);
  and g_118318_(_026860_, _026868_, _026870_);
  or g_118319_(_026859_, _026869_, _026871_);
  and g_118320_(_026829_, _026870_, _026873_);
  or g_118321_(_026827_, _026871_, _026874_);
  and g_118322_(out[883], _026765_, _026875_);
  and g_118323_(_026687_, _026766_, _026876_);
  or g_118324_(_026875_, _026876_, _026877_);
  or g_118325_(_001902_, _026877_, _026878_);
  and g_118326_(_026678_, _026766_, _026879_);
  and g_118327_(_001759_, _026765_, _026880_);
  or g_118328_(_026879_, _026880_, _026881_);
  and g_118329_(_001902_, _026877_, _026882_);
  or g_118330_(out[898], _026881_, _026884_);
  xor g_118331_(_001902_, _026877_, _026885_);
  xor g_118332_(out[899], _026877_, _026886_);
  xor g_118333_(out[898], _026881_, _026887_);
  xor g_118334_(_001891_, _026881_, _026888_);
  and g_118335_(_026885_, _026887_, _026889_);
  or g_118336_(_026886_, _026888_, _026890_);
  or g_118337_(out[897], _026769_, _026891_);
  and g_118338_(_026709_, _026766_, _026892_);
  and g_118339_(_001748_, _026765_, _026893_);
  or g_118340_(_026892_, _026893_, _026895_);
  and g_118341_(out[896], _026895_, _026896_);
  not g_118342_(_026896_, _026897_);
  xor g_118343_(out[897], _026769_, _026898_);
  xor g_118344_(_001869_, _026769_, _026899_);
  and g_118345_(_026897_, _026898_, _026900_);
  or g_118346_(_026896_, _026899_, _026901_);
  and g_118347_(_026891_, _026901_, _026902_);
  or g_118348_(_026890_, _026902_, _026903_);
  or g_118349_(_026882_, _026884_, _026904_);
  and g_118350_(_026878_, _026904_, _026906_);
  and g_118351_(_026903_, _026906_, _026907_);
  or g_118352_(_026874_, _026907_, _026908_);
  or g_118353_(_026857_, _026864_, _026909_);
  or g_118354_(_026837_, _026858_, _026910_);
  or g_118355_(_026867_, _026910_, _026911_);
  and g_118356_(_026909_, _026911_, _026912_);
  or g_118357_(_026827_, _026912_, _026913_);
  or g_118358_(_026796_, _026799_, _026914_);
  or g_118359_(_026811_, _026823_, _026915_);
  and g_118360_(_026914_, _026915_, _026917_);
  and g_118361_(_026913_, _026917_, _026918_);
  and g_118362_(_026908_, _026918_, _026919_);
  or g_118363_(out[896], _026895_, _026920_);
  and g_118364_(_026889_, _026920_, _026921_);
  and g_118365_(_026900_, _026921_, _026922_);
  and g_118366_(_026873_, _026922_, _026923_);
  or g_118367_(_026919_, _026923_, _026924_);
  not g_118368_(_026924_, _026925_);
  and g_118369_(_026769_, _026924_, _026926_);
  and g_118370_(_001869_, _026925_, _026928_);
  or g_118371_(_026926_, _026928_, _026929_);
  and g_118372_(_026789_, _026791_, _026930_);
  or g_118373_(_026790_, _026792_, _026931_);
  and g_118374_(out[916], out[915], _026932_);
  or g_118375_(out[917], _026932_, _026933_);
  or g_118376_(out[918], _026933_, _026934_);
  or g_118377_(out[919], _026934_, _026935_);
  or g_118378_(out[920], _026935_, _026936_);
  and g_118379_(out[921], _026936_, _026937_);
  or g_118380_(out[922], _026937_, _026939_);
  xor g_118381_(out[923], _026939_, _026940_);
  xor g_118382_(_001946_, _026939_, _026941_);
  and g_118383_(_026930_, _026941_, _026942_);
  or g_118384_(_026931_, _026940_, _026943_);
  and g_118385_(_026776_, _026924_, _026944_);
  and g_118386_(_026785_, _026925_, _026945_);
  or g_118387_(_026944_, _026945_, _026946_);
  xor g_118388_(_002067_, _026937_, _026947_);
  or g_118389_(_026946_, _026947_, _026948_);
  not g_118390_(_026948_, _026950_);
  and g_118391_(_026943_, _026948_, _026951_);
  or g_118392_(_026942_, _026950_, _026952_);
  and g_118393_(_026946_, _026947_, _026953_);
  and g_118394_(_026931_, _026940_, _026954_);
  or g_118395_(_026953_, _026954_, _026955_);
  or g_118396_(_026952_, _026955_, _026956_);
  xor g_118397_(_002045_, _026935_, _026957_);
  or g_118398_(_026818_, _026925_, _026958_);
  or g_118399_(_026820_, _026924_, _026959_);
  and g_118400_(_026958_, _026959_, _026961_);
  or g_118401_(_026957_, _026961_, _026962_);
  not g_118402_(_026962_, _026963_);
  xor g_118403_(out[921], _026936_, _026964_);
  xor g_118404_(_002056_, _026936_, _026965_);
  and g_118405_(_026807_, _026924_, _026966_);
  and g_118406_(_026800_, _026925_, _026967_);
  or g_118407_(_026966_, _026967_, _026968_);
  not g_118408_(_026968_, _026969_);
  and g_118409_(_026965_, _026968_, _026970_);
  not g_118410_(_026970_, _026972_);
  and g_118411_(_026962_, _026972_, _026973_);
  or g_118412_(_026963_, _026970_, _026974_);
  and g_118413_(_026964_, _026969_, _026975_);
  or g_118414_(_026965_, _026968_, _026976_);
  and g_118415_(_026957_, _026961_, _026977_);
  and g_118416_(_026973_, _026976_, _026978_);
  or g_118417_(_026974_, _026975_, _026979_);
  or g_118418_(_026956_, _026977_, _026980_);
  not g_118419_(_026980_, _026981_);
  and g_118420_(_026978_, _026981_, _026983_);
  or g_118421_(_026979_, _026980_, _026984_);
  xor g_118422_(out[919], _026934_, _026985_);
  xor g_118423_(_001957_, _026934_, _026986_);
  or g_118424_(_026856_, _026925_, _026987_);
  not g_118425_(_026987_, _026988_);
  or g_118426_(_026852_, _026924_, _026989_);
  not g_118427_(_026989_, _026990_);
  and g_118428_(_026987_, _026989_, _026991_);
  or g_118429_(_026988_, _026990_, _026992_);
  and g_118430_(_026985_, _026992_, _026994_);
  or g_118431_(_026986_, _026991_, _026995_);
  xor g_118432_(out[918], _026933_, _026996_);
  xor g_118433_(_001968_, _026933_, _026997_);
  and g_118434_(_026849_, _026924_, _026998_);
  not g_118435_(_026998_, _026999_);
  and g_118436_(_026845_, _026925_, _027000_);
  or g_118437_(_026846_, _026924_, _027001_);
  and g_118438_(_026999_, _027001_, _027002_);
  or g_118439_(_026998_, _027000_, _027003_);
  and g_118440_(_026996_, _027002_, _027005_);
  or g_118441_(_026997_, _027003_, _027006_);
  and g_118442_(_026995_, _027006_, _027007_);
  or g_118443_(_026994_, _027005_, _027008_);
  and g_118444_(_026986_, _026991_, _027009_);
  or g_118445_(_027007_, _027009_, _027010_);
  and g_118446_(_026997_, _027003_, _027011_);
  or g_118447_(_027009_, _027011_, _027012_);
  or g_118448_(_027008_, _027012_, _027013_);
  xor g_118449_(_001979_, _026932_, _027014_);
  and g_118450_(_026836_, _026924_, _027016_);
  and g_118451_(_026830_, _026925_, _027017_);
  or g_118452_(_027016_, _027017_, _027018_);
  not g_118453_(_027018_, _027019_);
  or g_118454_(_027014_, _027019_, _027020_);
  and g_118455_(out[899], _026925_, _027021_);
  and g_118456_(_026877_, _026924_, _027022_);
  or g_118457_(_027021_, _027022_, _027023_);
  and g_118458_(_002034_, _027023_, _027024_);
  and g_118459_(_026881_, _026924_, _027025_);
  and g_118460_(_001891_, _026925_, _027027_);
  or g_118461_(_027025_, _027027_, _027028_);
  and g_118462_(out[914], _027028_, _027029_);
  or g_118463_(_027024_, _027029_, _027030_);
  or g_118464_(out[914], _027028_, _027031_);
  or g_118465_(out[913], _026929_, _027032_);
  and g_118466_(_027031_, _027032_, _027033_);
  or g_118467_(_002034_, _027023_, _027034_);
  xor g_118468_(out[916], out[915], _027035_);
  xor g_118469_(_001990_, out[915], _027036_);
  and g_118470_(_026842_, _026924_, _027038_);
  or g_118471_(_026838_, _026924_, _027039_);
  not g_118472_(_027039_, _027040_);
  or g_118473_(_027038_, _027040_, _027041_);
  or g_118474_(_027035_, _027041_, _027042_);
  and g_118475_(_027034_, _027042_, _027043_);
  and g_118476_(_026895_, _026924_, _027044_);
  and g_118477_(_001880_, _026925_, _027045_);
  or g_118478_(_027044_, _027045_, _027046_);
  and g_118479_(out[912], _027046_, _027047_);
  and g_118480_(out[913], _026929_, _027049_);
  or g_118481_(_027047_, _027049_, _027050_);
  or g_118482_(_027030_, _027050_, _027051_);
  and g_118483_(_027033_, _027050_, _027052_);
  or g_118484_(_027030_, _027052_, _027053_);
  and g_118485_(_027043_, _027053_, _027054_);
  and g_118486_(_027035_, _027041_, _027055_);
  and g_118487_(_027014_, _027019_, _027056_);
  or g_118488_(_027055_, _027056_, _027057_);
  not g_118489_(_027057_, _027058_);
  or g_118490_(_027054_, _027057_, _027060_);
  and g_118491_(_027020_, _027060_, _027061_);
  or g_118492_(_027013_, _027061_, _027062_);
  and g_118493_(_027010_, _027062_, _027063_);
  or g_118494_(_026984_, _027063_, _027064_);
  or g_118495_(_026973_, _026975_, _027065_);
  or g_118496_(_026956_, _027065_, _027066_);
  or g_118497_(_026951_, _026954_, _027067_);
  and g_118498_(_027066_, _027067_, _027068_);
  and g_118499_(_027064_, _027068_, _027069_);
  or g_118500_(out[912], _027046_, _027071_);
  and g_118501_(_027020_, _027071_, _027072_);
  and g_118502_(_027058_, _027072_, _027073_);
  and g_118503_(_027033_, _027043_, _027074_);
  and g_118504_(_027073_, _027074_, _027075_);
  or g_118505_(_027013_, _027051_, _027076_);
  not g_118506_(_027076_, _027077_);
  and g_118507_(_027075_, _027077_, _027078_);
  and g_118508_(_026983_, _027078_, _027079_);
  or g_118509_(_027069_, _027079_, _027080_);
  not g_118510_(_027080_, _027082_);
  and g_118511_(_026929_, _027080_, _027083_);
  and g_118512_(_002001_, _027082_, _027084_);
  or g_118513_(_027083_, _027084_, _027085_);
  and g_118514_(_026930_, _026940_, _027086_);
  not g_118515_(_027086_, _027087_);
  and g_118516_(out[932], out[931], _027088_);
  or g_118517_(out[933], _027088_, _027089_);
  or g_118518_(out[934], _027089_, _027090_);
  or g_118519_(out[935], _027090_, _027091_);
  or g_118520_(out[936], _027091_, _027093_);
  and g_118521_(out[937], _027093_, _027094_);
  or g_118522_(out[938], _027094_, _027095_);
  xor g_118523_(out[939], _027095_, _027096_);
  not g_118524_(_027096_, _027097_);
  and g_118525_(_027086_, _027097_, _027098_);
  or g_118526_(_027087_, _027096_, _027099_);
  or g_118527_(_026947_, _027080_, _027100_);
  not g_118528_(_027100_, _027101_);
  and g_118529_(_026946_, _027080_, _027102_);
  not g_118530_(_027102_, _027104_);
  and g_118531_(_027100_, _027104_, _027105_);
  or g_118532_(_027101_, _027102_, _027106_);
  xor g_118533_(out[938], _027094_, _027107_);
  xor g_118534_(_002177_, _027094_, _027108_);
  and g_118535_(_027105_, _027107_, _027109_);
  or g_118536_(_027106_, _027108_, _027110_);
  and g_118537_(_027099_, _027110_, _027111_);
  or g_118538_(_027098_, _027109_, _027112_);
  xor g_118539_(out[936], _027091_, _027113_);
  xor g_118540_(_002155_, _027091_, _027115_);
  or g_118541_(_026957_, _027080_, _027116_);
  not g_118542_(_027116_, _027117_);
  and g_118543_(_026961_, _027080_, _027118_);
  or g_118544_(_027117_, _027118_, _027119_);
  xor g_118545_(_002166_, _027093_, _027120_);
  or g_118546_(_026965_, _027080_, _027121_);
  not g_118547_(_027121_, _027122_);
  and g_118548_(_026968_, _027080_, _027123_);
  or g_118549_(_026969_, _027082_, _027124_);
  and g_118550_(_027121_, _027124_, _027126_);
  or g_118551_(_027122_, _027123_, _027127_);
  or g_118552_(_027120_, _027127_, _027128_);
  and g_118553_(_027087_, _027096_, _027129_);
  or g_118554_(_027086_, _027097_, _027130_);
  and g_118555_(_027106_, _027108_, _027131_);
  or g_118556_(_027105_, _027107_, _027132_);
  and g_118557_(_027130_, _027132_, _027133_);
  or g_118558_(_027129_, _027131_, _027134_);
  and g_118559_(_027120_, _027127_, _027135_);
  or g_118560_(_027115_, _027119_, _027137_);
  not g_118561_(_027137_, _027138_);
  or g_118562_(_027135_, _027138_, _027139_);
  xor g_118563_(_027120_, _027127_, _027140_);
  xor g_118564_(_027120_, _027126_, _027141_);
  and g_118565_(_027133_, _027140_, _027142_);
  or g_118566_(_027134_, _027141_, _027143_);
  xor g_118567_(_027115_, _027119_, _027144_);
  xor g_118568_(_027113_, _027119_, _027145_);
  and g_118569_(_027111_, _027144_, _027146_);
  or g_118570_(_027112_, _027145_, _027148_);
  and g_118571_(_027142_, _027146_, _027149_);
  or g_118572_(_027143_, _027148_, _027150_);
  xor g_118573_(out[934], _027089_, _027151_);
  not g_118574_(_027151_, _027152_);
  and g_118575_(_026996_, _027082_, _027153_);
  and g_118576_(_027003_, _027080_, _027154_);
  or g_118577_(_027153_, _027154_, _027155_);
  not g_118578_(_027155_, _027156_);
  and g_118579_(_027151_, _027156_, _027157_);
  xor g_118580_(out[935], _027090_, _027159_);
  and g_118581_(_026986_, _027082_, _027160_);
  and g_118582_(_026992_, _027080_, _027161_);
  or g_118583_(_027160_, _027161_, _027162_);
  not g_118584_(_027162_, _027163_);
  and g_118585_(_027159_, _027162_, _027164_);
  or g_118586_(_027157_, _027164_, _027165_);
  or g_118587_(_027159_, _027162_, _027166_);
  xor g_118588_(_027152_, _027155_, _027167_);
  xor g_118589_(_027151_, _027155_, _027168_);
  xor g_118590_(_027159_, _027162_, _027170_);
  xor g_118591_(_027159_, _027163_, _027171_);
  and g_118592_(_027167_, _027170_, _027172_);
  or g_118593_(_027168_, _027171_, _027173_);
  xor g_118594_(out[932], out[931], _027174_);
  or g_118595_(_027036_, _027080_, _027175_);
  or g_118596_(_027041_, _027082_, _027176_);
  and g_118597_(_027175_, _027176_, _027177_);
  or g_118598_(_027174_, _027177_, _027178_);
  not g_118599_(_027178_, _027179_);
  xor g_118600_(out[933], _027088_, _027181_);
  xor g_118601_(_002089_, _027088_, _027182_);
  and g_118602_(_027014_, _027082_, _027183_);
  and g_118603_(_027018_, _027080_, _027184_);
  or g_118604_(_027183_, _027184_, _027185_);
  not g_118605_(_027185_, _027186_);
  and g_118606_(_027181_, _027185_, _027187_);
  not g_118607_(_027187_, _027188_);
  and g_118608_(_027178_, _027188_, _027189_);
  or g_118609_(_027179_, _027187_, _027190_);
  and g_118610_(_027182_, _027186_, _027192_);
  or g_118611_(_027181_, _027185_, _027193_);
  and g_118612_(_027174_, _027177_, _027194_);
  not g_118613_(_027194_, _027195_);
  and g_118614_(_027193_, _027195_, _027196_);
  or g_118615_(_027192_, _027194_, _027197_);
  and g_118616_(_027189_, _027196_, _027198_);
  or g_118617_(_027190_, _027197_, _027199_);
  and g_118618_(_027172_, _027198_, _027200_);
  or g_118619_(_027173_, _027199_, _027201_);
  and g_118620_(out[915], _027082_, _027203_);
  and g_118621_(_027023_, _027080_, _027204_);
  or g_118622_(_027203_, _027204_, _027205_);
  or g_118623_(_002144_, _027205_, _027206_);
  and g_118624_(_002144_, _027205_, _027207_);
  xor g_118625_(_002144_, _027205_, _027208_);
  xor g_118626_(out[931], _027205_, _027209_);
  and g_118627_(_027028_, _027080_, _027210_);
  and g_118628_(_002023_, _027082_, _027211_);
  or g_118629_(_027210_, _027211_, _027212_);
  or g_118630_(out[930], _027212_, _027214_);
  xor g_118631_(out[930], _027212_, _027215_);
  xor g_118632_(_002133_, _027212_, _027216_);
  and g_118633_(_027208_, _027215_, _027217_);
  or g_118634_(_027209_, _027216_, _027218_);
  or g_118635_(out[929], _027085_, _027219_);
  xor g_118636_(out[929], _027085_, _027220_);
  xor g_118637_(_002111_, _027085_, _027221_);
  and g_118638_(_027046_, _027080_, _027222_);
  and g_118639_(_002012_, _027082_, _027223_);
  or g_118640_(_027222_, _027223_, _027225_);
  and g_118641_(out[928], _027225_, _027226_);
  not g_118642_(_027226_, _027227_);
  or g_118643_(_027221_, _027226_, _027228_);
  and g_118644_(_027217_, _027227_, _027229_);
  and g_118645_(_027220_, _027229_, _027230_);
  or g_118646_(_027218_, _027228_, _027231_);
  or g_118647_(_027218_, _027219_, _027232_);
  or g_118648_(_027207_, _027214_, _027233_);
  and g_118649_(_027206_, _027233_, _027234_);
  and g_118650_(_027232_, _027234_, _027236_);
  and g_118651_(_027231_, _027236_, _027237_);
  or g_118652_(_027201_, _027237_, _027238_);
  and g_118653_(_027165_, _027166_, _027239_);
  not g_118654_(_027239_, _027240_);
  or g_118655_(_027173_, _027189_, _027241_);
  or g_118656_(_027192_, _027241_, _027242_);
  and g_118657_(_027240_, _027242_, _027243_);
  and g_118658_(_027238_, _027243_, _027244_);
  or g_118659_(_027150_, _027244_, _027245_);
  and g_118660_(_027112_, _027130_, _027247_);
  and g_118661_(_027133_, _027139_, _027248_);
  and g_118662_(_027128_, _027248_, _027249_);
  or g_118663_(_027247_, _027249_, _027250_);
  not g_118664_(_027250_, _027251_);
  and g_118665_(_027245_, _027251_, _027252_);
  and g_118666_(_027200_, _027230_, _027253_);
  or g_118667_(out[928], _027225_, _027254_);
  and g_118668_(_027149_, _027254_, _027255_);
  and g_118669_(_027253_, _027255_, _027256_);
  or g_118670_(_027252_, _027256_, _027258_);
  not g_118671_(_027258_, _027259_);
  and g_118672_(_027085_, _027258_, _027260_);
  not g_118673_(_027260_, _027261_);
  or g_118674_(out[929], _027258_, _027262_);
  not g_118675_(_027262_, _027263_);
  and g_118676_(_027261_, _027262_, _027264_);
  or g_118677_(_027260_, _027263_, _027265_);
  or g_118678_(_002144_, _027258_, _027266_);
  not g_118679_(_027266_, _027267_);
  and g_118680_(_027205_, _027258_, _027269_);
  not g_118681_(_027269_, _027270_);
  and g_118682_(_027266_, _027270_, _027271_);
  or g_118683_(_027267_, _027269_, _027272_);
  and g_118684_(out[947], _027271_, _027273_);
  or g_118685_(_002254_, _027272_, _027274_);
  and g_118686_(_027212_, _027258_, _027275_);
  not g_118687_(_027275_, _027276_);
  or g_118688_(out[930], _027258_, _027277_);
  not g_118689_(_027277_, _027278_);
  and g_118690_(_027276_, _027277_, _027280_);
  or g_118691_(_027275_, _027278_, _027281_);
  and g_118692_(out[946], _027281_, _027282_);
  or g_118693_(_002243_, _027280_, _027283_);
  and g_118694_(_027274_, _027283_, _027284_);
  or g_118695_(_027273_, _027282_, _027285_);
  and g_118696_(_002254_, _027272_, _027286_);
  or g_118697_(out[947], _027271_, _027287_);
  and g_118698_(_002243_, _027280_, _027288_);
  or g_118699_(out[946], _027281_, _027289_);
  and g_118700_(_027287_, _027289_, _027291_);
  or g_118701_(_027286_, _027288_, _027292_);
  and g_118702_(_027284_, _027291_, _027293_);
  or g_118703_(_027285_, _027292_, _027294_);
  and g_118704_(_054336_, _027264_, _027295_);
  or g_118705_(out[945], _027265_, _027296_);
  and g_118706_(_027225_, _027258_, _027297_);
  not g_118707_(_027297_, _027298_);
  or g_118708_(out[928], _027258_, _027299_);
  and g_118709_(_027298_, _027299_, _027300_);
  not g_118710_(_027300_, _027302_);
  and g_118711_(out[944], _027302_, _027303_);
  or g_118712_(_002232_, _027300_, _027304_);
  xor g_118713_(_054336_, _027264_, _027305_);
  xor g_118714_(out[945], _027264_, _027306_);
  and g_118715_(_027304_, _027305_, _027307_);
  or g_118716_(_027303_, _027306_, _027308_);
  and g_118717_(_027296_, _027308_, _027309_);
  or g_118718_(_027295_, _027307_, _027310_);
  and g_118719_(_027293_, _027310_, _027311_);
  or g_118720_(_027294_, _027309_, _027313_);
  and g_118721_(_027287_, _027288_, _027314_);
  or g_118722_(_027286_, _027289_, _027315_);
  and g_118723_(_027274_, _027315_, _027316_);
  or g_118724_(_027273_, _027314_, _027317_);
  and g_118725_(_027313_, _027316_, _027318_);
  or g_118726_(_027311_, _027317_, _027319_);
  and g_118727_(_027086_, _027096_, _027320_);
  not g_118728_(_027320_, _027321_);
  and g_118729_(out[948], out[947], _027322_);
  or g_118730_(out[949], _027322_, _027324_);
  or g_118731_(out[950], _027324_, _027325_);
  or g_118732_(out[951], _027325_, _027326_);
  or g_118733_(out[952], _027326_, _027327_);
  and g_118734_(out[953], _027327_, _027328_);
  or g_118735_(out[954], _027328_, _027329_);
  xor g_118736_(out[955], _027329_, _027330_);
  not g_118737_(_027330_, _027331_);
  and g_118738_(_027321_, _027330_, _027332_);
  or g_118739_(_027320_, _027331_, _027333_);
  xor g_118740_(out[953], _027327_, _027335_);
  xor g_118741_(_002276_, _027327_, _027336_);
  or g_118742_(_027120_, _027258_, _027337_);
  not g_118743_(_027337_, _027338_);
  and g_118744_(_027127_, _027258_, _027339_);
  not g_118745_(_027339_, _027340_);
  and g_118746_(_027337_, _027340_, _027341_);
  or g_118747_(_027338_, _027339_, _027342_);
  and g_118748_(_027335_, _027341_, _027343_);
  or g_118749_(_027336_, _027342_, _027344_);
  xor g_118750_(out[954], _027328_, _027346_);
  xor g_118751_(_002287_, _027328_, _027347_);
  and g_118752_(_027107_, _027259_, _027348_);
  or g_118753_(_027108_, _027258_, _027349_);
  and g_118754_(_027106_, _027258_, _027350_);
  or g_118755_(_027105_, _027259_, _027351_);
  and g_118756_(_027349_, _027351_, _027352_);
  or g_118757_(_027348_, _027350_, _027353_);
  and g_118758_(_027347_, _027353_, _027354_);
  or g_118759_(_027346_, _027352_, _027355_);
  xor g_118760_(out[952], _027326_, _027357_);
  not g_118761_(_027357_, _027358_);
  and g_118762_(_027113_, _027259_, _027359_);
  and g_118763_(_027119_, _027258_, _027360_);
  or g_118764_(_027359_, _027360_, _027361_);
  not g_118765_(_027361_, _027362_);
  and g_118766_(_027358_, _027361_, _027363_);
  or g_118767_(_027357_, _027362_, _027364_);
  and g_118768_(_027320_, _027331_, _027365_);
  or g_118769_(_027321_, _027330_, _027366_);
  and g_118770_(_027346_, _027352_, _027368_);
  or g_118771_(_027347_, _027353_, _027369_);
  and g_118772_(_027366_, _027369_, _027370_);
  or g_118773_(_027365_, _027368_, _027371_);
  and g_118774_(_027336_, _027342_, _027372_);
  or g_118775_(_027335_, _027341_, _027373_);
  and g_118776_(_027357_, _027362_, _027374_);
  or g_118777_(_027358_, _027361_, _027375_);
  and g_118778_(_027373_, _027375_, _027376_);
  or g_118779_(_027372_, _027374_, _027377_);
  and g_118780_(_027344_, _027376_, _027379_);
  or g_118781_(_027343_, _027377_, _027380_);
  and g_118782_(_027333_, _027355_, _027381_);
  or g_118783_(_027332_, _027354_, _027382_);
  and g_118784_(_027370_, _027381_, _027383_);
  or g_118785_(_027371_, _027382_, _027384_);
  and g_118786_(_027364_, _027383_, _027385_);
  or g_118787_(_027363_, _027384_, _027386_);
  and g_118788_(_027379_, _027385_, _027387_);
  or g_118789_(_027380_, _027386_, _027388_);
  xor g_118790_(out[951], _027325_, _027390_);
  xor g_118791_(_002188_, _027325_, _027391_);
  or g_118792_(_027159_, _027258_, _027392_);
  not g_118793_(_027392_, _027393_);
  and g_118794_(_027162_, _027258_, _027394_);
  not g_118795_(_027394_, _027395_);
  and g_118796_(_027392_, _027395_, _027396_);
  or g_118797_(_027393_, _027394_, _027397_);
  and g_118798_(_027390_, _027397_, _027398_);
  or g_118799_(_027391_, _027396_, _027399_);
  xor g_118800_(out[950], _027324_, _027401_);
  xor g_118801_(_002199_, _027324_, _027402_);
  or g_118802_(_027152_, _027258_, _027403_);
  not g_118803_(_027403_, _027404_);
  and g_118804_(_027155_, _027258_, _027405_);
  not g_118805_(_027405_, _027406_);
  and g_118806_(_027403_, _027406_, _027407_);
  or g_118807_(_027404_, _027405_, _027408_);
  and g_118808_(_027401_, _027407_, _027409_);
  or g_118809_(_027402_, _027408_, _027410_);
  and g_118810_(_027399_, _027410_, _027412_);
  or g_118811_(_027398_, _027409_, _027413_);
  and g_118812_(_027391_, _027396_, _027414_);
  or g_118813_(_027390_, _027397_, _027415_);
  and g_118814_(_027402_, _027408_, _027416_);
  or g_118815_(_027401_, _027407_, _027417_);
  and g_118816_(_027415_, _027417_, _027418_);
  or g_118817_(_027414_, _027416_, _027419_);
  and g_118818_(_027412_, _027418_, _027420_);
  or g_118819_(_027413_, _027419_, _027421_);
  xor g_118820_(out[949], _027322_, _027423_);
  xor g_118821_(_002210_, _027322_, _027424_);
  or g_118822_(_027181_, _027258_, _027425_);
  or g_118823_(_027186_, _027259_, _027426_);
  and g_118824_(_027425_, _027426_, _027427_);
  not g_118825_(_027427_, _027428_);
  and g_118826_(_027423_, _027428_, _027429_);
  or g_118827_(_027424_, _027427_, _027430_);
  xor g_118828_(out[948], out[947], _027431_);
  xor g_118829_(_002221_, out[947], _027432_);
  or g_118830_(_027174_, _027258_, _027434_);
  not g_118831_(_027434_, _027435_);
  and g_118832_(_027177_, _027258_, _027436_);
  not g_118833_(_027436_, _027437_);
  and g_118834_(_027434_, _027437_, _027438_);
  or g_118835_(_027435_, _027436_, _027439_);
  and g_118836_(_027432_, _027438_, _027440_);
  or g_118837_(_027431_, _027439_, _027441_);
  and g_118838_(_027430_, _027441_, _027442_);
  or g_118839_(_027429_, _027440_, _027443_);
  and g_118840_(_027424_, _027427_, _027445_);
  or g_118841_(_027423_, _027428_, _027446_);
  and g_118842_(_027431_, _027439_, _027447_);
  or g_118843_(_027432_, _027438_, _027448_);
  and g_118844_(_027446_, _027448_, _027449_);
  or g_118845_(_027445_, _027447_, _027450_);
  and g_118846_(_027442_, _027449_, _027451_);
  or g_118847_(_027443_, _027450_, _027452_);
  and g_118848_(_027420_, _027451_, _027453_);
  or g_118849_(_027421_, _027452_, _027454_);
  and g_118850_(_027387_, _027453_, _027456_);
  or g_118851_(_027388_, _027454_, _027457_);
  and g_118852_(_027319_, _027456_, _027458_);
  or g_118853_(_027318_, _027457_, _027459_);
  and g_118854_(_027413_, _027415_, _027460_);
  or g_118855_(_027412_, _027414_, _027461_);
  or g_118856_(_027442_, _027445_, _027462_);
  or g_118857_(_027419_, _027462_, _027463_);
  and g_118858_(_027420_, _027443_, _027464_);
  and g_118859_(_027446_, _027464_, _027465_);
  and g_118860_(_027461_, _027463_, _027467_);
  or g_118861_(_027460_, _027465_, _027468_);
  and g_118862_(_027387_, _027468_, _027469_);
  or g_118863_(_027388_, _027467_, _027470_);
  and g_118864_(_027344_, _027355_, _027471_);
  or g_118865_(_027343_, _027354_, _027472_);
  and g_118866_(_027377_, _027471_, _027473_);
  or g_118867_(_027376_, _027472_, _027474_);
  and g_118868_(_027370_, _027474_, _027475_);
  or g_118869_(_027371_, _027473_, _027476_);
  and g_118870_(_027333_, _027476_, _027478_);
  or g_118871_(_027332_, _027475_, _027479_);
  and g_118872_(_027470_, _027479_, _027480_);
  or g_118873_(_027469_, _027478_, _027481_);
  and g_118874_(_027459_, _027480_, _027482_);
  or g_118875_(_027458_, _027481_, _027483_);
  and g_118876_(_002232_, _027300_, _027484_);
  or g_118877_(out[944], _027302_, _027485_);
  and g_118878_(_027293_, _027485_, _027486_);
  or g_118879_(_027294_, _027484_, _027487_);
  and g_118880_(_027307_, _027486_, _027489_);
  or g_118881_(_027308_, _027487_, _027490_);
  and g_118882_(_027456_, _027489_, _027491_);
  or g_118883_(_027457_, _027490_, _027492_);
  and g_118884_(_027483_, _027492_, _027493_);
  or g_118885_(_027482_, _027491_, _027494_);
  and g_118886_(_027265_, _027494_, _027495_);
  or g_118887_(_027264_, _027493_, _027496_);
  and g_118888_(_054336_, _027493_, _027497_);
  or g_118889_(out[945], _027494_, _027498_);
  and g_118890_(_027496_, _027498_, _027500_);
  or g_118891_(_027495_, _027497_, _027501_);
  and g_118892_(_021519_, _027500_, _027502_);
  and g_118893_(_021365_, _021511_, _027503_);
  not g_118894_(_027503_, _027504_);
  and g_118895_(_021371_, _021512_, _027505_);
  or g_118896_(_021370_, _021511_, _027506_);
  and g_118897_(_027504_, _027506_, _027507_);
  or g_118898_(_027503_, _027505_, _027508_);
  and g_118899_(_027390_, _027493_, _027509_);
  or g_118900_(_027391_, _027494_, _027511_);
  and g_118901_(_027396_, _027494_, _027512_);
  or g_118902_(_027397_, _027493_, _027513_);
  and g_118903_(_027511_, _027513_, _027514_);
  or g_118904_(_027509_, _027512_, _027515_);
  and g_118905_(_027507_, _027514_, _027516_);
  or g_118906_(_027502_, _027516_, _027517_);
  and g_118907_(_021308_, _021511_, _027518_);
  not g_118908_(_027518_, _027519_);
  or g_118909_(_021312_, _021511_, _027520_);
  not g_118910_(_027520_, _027522_);
  and g_118911_(_027519_, _027520_, _027523_);
  or g_118912_(_027518_, _027522_, _027524_);
  and g_118913_(_027346_, _027493_, _027525_);
  or g_118914_(_027347_, _027494_, _027526_);
  and g_118915_(_027353_, _027494_, _027527_);
  or g_118916_(_027352_, _027493_, _027528_);
  and g_118917_(_027526_, _027528_, _027529_);
  or g_118918_(_027525_, _027527_, _027530_);
  and g_118919_(_027524_, _027529_, _027531_);
  or g_118920_(_021435_, _021511_, _027533_);
  not g_118921_(_027533_, _027534_);
  and g_118922_(_054303_, _021511_, _027535_);
  or g_118923_(out[466], _021512_, _027536_);
  and g_118924_(_027533_, _027536_, _027537_);
  or g_118925_(_027534_, _027535_, _027538_);
  and g_118926_(_027281_, _027494_, _027539_);
  or g_118927_(_027280_, _027493_, _027540_);
  and g_118928_(_002243_, _027493_, _027541_);
  or g_118929_(out[946], _027494_, _027542_);
  and g_118930_(_027540_, _027542_, _027544_);
  or g_118931_(_027539_, _027541_, _027545_);
  and g_118932_(_027538_, _027544_, _027546_);
  or g_118933_(_027531_, _027546_, _027547_);
  or g_118934_(_027517_, _027547_, _027548_);
  or g_118935_(_021459_, _021511_, _027549_);
  or g_118936_(out[464], _021512_, _027550_);
  and g_118937_(_027549_, _027550_, _027551_);
  or g_118938_(_027300_, _027493_, _027552_);
  or g_118939_(out[944], _027494_, _027553_);
  and g_118940_(_027552_, _027553_, _027555_);
  xor g_118941_(_027551_, _027555_, _027556_);
  and g_118942_(_027523_, _027530_, _027557_);
  and g_118943_(_021315_, _021318_, _027558_);
  and g_118944_(_027320_, _027330_, _027559_);
  xor g_118945_(_027558_, _027559_, _027560_);
  or g_118946_(_027557_, _027560_, _027561_);
  or g_118947_(_027556_, _027561_, _027562_);
  or g_118948_(_027548_, _027562_, _027563_);
  and g_118949_(_021401_, _021511_, _027564_);
  or g_118950_(_021400_, _021512_, _027566_);
  and g_118951_(_021408_, _021512_, _027567_);
  or g_118952_(_021407_, _021511_, _027568_);
  and g_118953_(_027566_, _027568_, _027569_);
  or g_118954_(_027564_, _027567_, _027570_);
  and g_118955_(_027432_, _027493_, _027571_);
  or g_118956_(_027431_, _027494_, _027572_);
  and g_118957_(_027439_, _027494_, _027573_);
  or g_118958_(_027438_, _027493_, _027574_);
  and g_118959_(_027572_, _027574_, _027575_);
  or g_118960_(_027571_, _027573_, _027577_);
  and g_118961_(_027570_, _027575_, _027578_);
  and g_118962_(_021343_, _021511_, _027579_);
  or g_118963_(_021344_, _021512_, _027580_);
  and g_118964_(_021351_, _021512_, _027581_);
  or g_118965_(_021349_, _021511_, _027582_);
  and g_118966_(_027580_, _027582_, _027583_);
  or g_118967_(_027579_, _027581_, _027584_);
  and g_118968_(_027335_, _027493_, _027585_);
  or g_118969_(_027336_, _027494_, _027586_);
  and g_118970_(_027342_, _027494_, _027588_);
  or g_118971_(_027341_, _027493_, _027589_);
  and g_118972_(_027586_, _027589_, _027590_);
  or g_118973_(_027585_, _027588_, _027591_);
  and g_118974_(_027584_, _027590_, _027592_);
  or g_118975_(_027578_, _027592_, _027593_);
  or g_118976_(_021334_, _021512_, _027594_);
  or g_118977_(_021340_, _021511_, _027595_);
  and g_118978_(_027594_, _027595_, _027596_);
  or g_118979_(_027358_, _027494_, _027597_);
  or g_118980_(_027362_, _027493_, _027599_);
  and g_118981_(_027597_, _027599_, _027600_);
  xor g_118982_(_027596_, _027600_, _027601_);
  or g_118983_(_027593_, _027601_, _027602_);
  and g_118984_(_021386_, _021511_, _027603_);
  or g_118985_(_021387_, _021512_, _027604_);
  and g_118986_(_021392_, _021512_, _027605_);
  or g_118987_(_021391_, _021511_, _027606_);
  and g_118988_(_027604_, _027606_, _027607_);
  or g_118989_(_027603_, _027605_, _027608_);
  and g_118990_(_027407_, _027494_, _027610_);
  or g_118991_(_027408_, _027493_, _027611_);
  and g_118992_(_027402_, _027493_, _027612_);
  or g_118993_(_027401_, _027494_, _027613_);
  and g_118994_(_027611_, _027613_, _027614_);
  or g_118995_(_027610_, _027612_, _027615_);
  and g_118996_(_027608_, _027615_, _027616_);
  and g_118997_(_027508_, _027515_, _027617_);
  or g_118998_(_027616_, _027617_, _027618_);
  and g_118999_(_027537_, _027545_, _027619_);
  and g_119000_(_027569_, _027577_, _027621_);
  or g_119001_(_027619_, _027621_, _027622_);
  or g_119002_(_027618_, _027622_, _027623_);
  or g_119003_(_027602_, _027623_, _027624_);
  and g_119004_(out[467], _021511_, _027625_);
  or g_119005_(_054281_, _021512_, _027626_);
  or g_119006_(_021426_, _021511_, _027627_);
  not g_119007_(_027627_, _027628_);
  and g_119008_(_027626_, _027627_, _027629_);
  or g_119009_(_027625_, _027628_, _027630_);
  and g_119010_(out[947], _027493_, _027632_);
  or g_119011_(_002254_, _027494_, _027633_);
  and g_119012_(_027272_, _027494_, _027634_);
  or g_119013_(_027271_, _027493_, _027635_);
  and g_119014_(_027633_, _027635_, _027636_);
  or g_119015_(_027632_, _027634_, _027637_);
  and g_119016_(_027630_, _027636_, _027638_);
  and g_119017_(_027583_, _027591_, _027639_);
  and g_119018_(_027629_, _027637_, _027640_);
  or g_119019_(_027639_, _027640_, _027641_);
  or g_119020_(_027638_, _027641_, _027643_);
  and g_119021_(_021518_, _027501_, _027644_);
  and g_119022_(_027607_, _027614_, _027645_);
  or g_119023_(_027644_, _027645_, _027646_);
  or g_119024_(_021374_, _021512_, _027647_);
  or g_119025_(_021379_, _021511_, _027648_);
  and g_119026_(_027647_, _027648_, _027649_);
  or g_119027_(_027427_, _027493_, _027650_);
  or g_119028_(_027423_, _027494_, _027651_);
  and g_119029_(_027650_, _027651_, _027652_);
  xor g_119030_(_027649_, _027652_, _027654_);
  or g_119031_(_027646_, _027654_, _027655_);
  or g_119032_(_027643_, _027655_, _027656_);
  or g_119033_(_027624_, _027656_, _027657_);
  or g_119034_(_027563_, _027657_, _027658_);
  not g_119035_(_027658_, _027659_);
  or g_119036_(out[10], _003587_, _027660_);
  xor g_119037_(out[11], _027660_, _027661_);
  xor g_119038_(_002298_, _027660_, _027662_);
  or g_119039_(out[26], _003590_, _027663_);
  xor g_119040_(out[27], _027663_, _027665_);
  xor g_119041_(_002430_, _027663_, _027666_);
  and g_119042_(_027662_, _027665_, _027667_);
  or g_119043_(_027661_, _027666_, _027668_);
  xor g_119044_(out[10], _003587_, _027669_);
  xor g_119045_(_002419_, _003587_, _027670_);
  xor g_119046_(out[26], _003590_, _027671_);
  xor g_119047_(_002551_, _003590_, _027672_);
  and g_119048_(_027670_, _027671_, _027673_);
  or g_119049_(_027669_, _027672_, _027674_);
  and g_119050_(_027669_, _027672_, _027676_);
  or g_119051_(_027670_, _027671_, _027677_);
  and g_119052_(_003594_, _003699_, _027678_);
  or g_119053_(_003593_, _003698_, _027679_);
  and g_119054_(_027677_, _027679_, _027680_);
  or g_119055_(_027676_, _027678_, _027681_);
  and g_119056_(_027674_, _027681_, _027682_);
  or g_119057_(_027673_, _027680_, _027683_);
  and g_119058_(_027661_, _027666_, _027684_);
  or g_119059_(_027662_, _027665_, _027685_);
  and g_119060_(_027682_, _027685_, _027687_);
  or g_119061_(_027683_, _027684_, _027688_);
  and g_119062_(_027668_, _027688_, _027689_);
  or g_119063_(_027667_, _027687_, _027690_);
  and g_119064_(_003697_, _027690_, _027691_);
  or g_119065_(_003696_, _027689_, _027692_);
  and g_119066_(_003671_, _027692_, _027693_);
  or g_119067_(_003670_, _027691_, _027694_);
  or g_119068_(_003620_, _027693_, _027695_);
  or g_119069_(_003622_, _027694_, _027696_);
  and g_119070_(_027695_, _027696_, _027698_);
  not g_119071_(_027698_, _027699_);
  and g_119072_(_003652_, _027693_, _027700_);
  or g_119073_(_003650_, _027694_, _027701_);
  and g_119074_(_003649_, _027694_, _027702_);
  or g_119075_(_003648_, _027693_, _027703_);
  and g_119076_(_027701_, _027703_, _027704_);
  or g_119077_(_027700_, _027702_, _027705_);
  and g_119078_(_003854_, _027705_, _027706_);
  or g_119079_(_003855_, _027704_, _027707_);
  or g_119080_(_003616_, _027694_, _027709_);
  or g_119081_(_003614_, _027693_, _027710_);
  and g_119082_(_027709_, _027710_, _027711_);
  not g_119083_(_027711_, _027712_);
  and g_119084_(_003832_, _027711_, _027713_);
  or g_119085_(_003832_, _027711_, _027714_);
  and g_119086_(_003822_, _027698_, _027715_);
  xor g_119087_(_003832_, _027711_, _027716_);
  xor g_119088_(_003833_, _027711_, _027717_);
  xor g_119089_(_003822_, _027698_, _027718_);
  xor g_119090_(_003821_, _027698_, _027720_);
  and g_119091_(_027716_, _027718_, _027721_);
  or g_119092_(_027717_, _027720_, _027722_);
  and g_119093_(_027707_, _027721_, _027723_);
  or g_119094_(_027706_, _027722_, _027724_);
  and g_119095_(_003645_, _027693_, _027725_);
  or g_119096_(_003644_, _027694_, _027726_);
  and g_119097_(_003641_, _027694_, _027727_);
  or g_119098_(_003639_, _027693_, _027728_);
  and g_119099_(_027726_, _027728_, _027729_);
  or g_119100_(_027725_, _027727_, _027731_);
  and g_119101_(_003868_, _027729_, _027732_);
  or g_119102_(_003867_, _027731_, _027733_);
  and g_119103_(_003855_, _027704_, _027734_);
  or g_119104_(_003854_, _027705_, _027735_);
  and g_119105_(_027733_, _027735_, _027736_);
  or g_119106_(_027732_, _027734_, _027737_);
  and g_119107_(_003867_, _027731_, _027738_);
  or g_119108_(_003868_, _027729_, _027739_);
  and g_119109_(_027736_, _027739_, _027740_);
  or g_119110_(_027737_, _027738_, _027742_);
  and g_119111_(_027723_, _027740_, _027743_);
  or g_119112_(_027724_, _027742_, _027744_);
  or g_119113_(out[42], _003718_, _027745_);
  xor g_119114_(out[42], _003718_, _027746_);
  not g_119115_(_027746_, _027747_);
  and g_119116_(_027671_, _027693_, _027748_);
  or g_119117_(_027672_, _027694_, _027749_);
  and g_119118_(_027669_, _027694_, _027750_);
  or g_119119_(_027670_, _027693_, _027751_);
  and g_119120_(_027749_, _027751_, _027753_);
  or g_119121_(_027748_, _027750_, _027754_);
  and g_119122_(_027747_, _027754_, _027755_);
  or g_119123_(_027746_, _027753_, _027756_);
  xor g_119124_(out[43], _027745_, _027757_);
  xor g_119125_(_002562_, _027745_, _027758_);
  and g_119126_(_027666_, _027693_, _027759_);
  or g_119127_(_027665_, _027694_, _027760_);
  and g_119128_(_027662_, _027694_, _027761_);
  or g_119129_(_027661_, _027693_, _027762_);
  and g_119130_(_027760_, _027762_, _027764_);
  or g_119131_(_027759_, _027761_, _027765_);
  and g_119132_(_027757_, _027765_, _027766_);
  or g_119133_(_027758_, _027764_, _027767_);
  and g_119134_(_027756_, _027767_, _027768_);
  or g_119135_(_027755_, _027766_, _027769_);
  and g_119136_(_027746_, _027753_, _027770_);
  or g_119137_(_027747_, _027754_, _027771_);
  and g_119138_(_027758_, _027764_, _027772_);
  or g_119139_(_027757_, _027765_, _027773_);
  and g_119140_(_027771_, _027773_, _027775_);
  or g_119141_(_027770_, _027772_, _027776_);
  and g_119142_(_027768_, _027775_, _027777_);
  or g_119143_(_027769_, _027776_, _027778_);
  and g_119144_(_003601_, _027694_, _027779_);
  or g_119145_(_003600_, _027693_, _027780_);
  or g_119146_(_003602_, _027694_, _027781_);
  not g_119147_(_027781_, _027782_);
  and g_119148_(_027780_, _027781_, _027783_);
  or g_119149_(_027779_, _027782_, _027784_);
  and g_119150_(_003731_, _027783_, _027786_);
  or g_119151_(_003730_, _027784_, _027787_);
  and g_119152_(_003591_, _027693_, _027788_);
  or g_119153_(_003592_, _027694_, _027789_);
  and g_119154_(_003588_, _027694_, _027790_);
  or g_119155_(_003589_, _027693_, _027791_);
  and g_119156_(_027789_, _027791_, _027792_);
  or g_119157_(_027788_, _027790_, _027793_);
  and g_119158_(_003720_, _027793_, _027794_);
  or g_119159_(_003719_, _027792_, _027795_);
  and g_119160_(_027787_, _027795_, _027797_);
  or g_119161_(_027786_, _027794_, _027798_);
  and g_119162_(_003719_, _027792_, _027799_);
  or g_119163_(_003720_, _027793_, _027800_);
  and g_119164_(_003730_, _027784_, _027801_);
  or g_119165_(_003731_, _027783_, _027802_);
  and g_119166_(_027800_, _027802_, _027803_);
  or g_119167_(_027799_, _027801_, _027804_);
  and g_119168_(_027797_, _027803_, _027805_);
  or g_119169_(_027798_, _027804_, _027806_);
  and g_119170_(_027777_, _027805_, _027808_);
  or g_119171_(_027778_, _027806_, _027809_);
  or g_119172_(_002485_, _027694_, _027810_);
  or g_119173_(_002353_, _027693_, _027811_);
  and g_119174_(_027810_, _027811_, _027812_);
  and g_119175_(_002364_, _027694_, _027813_);
  or g_119176_(out[0], _027693_, _027814_);
  and g_119177_(_002496_, _027693_, _027815_);
  or g_119178_(out[16], _027694_, _027816_);
  and g_119179_(_027814_, _027816_, _027817_);
  or g_119180_(_027813_, _027815_, _027819_);
  and g_119181_(out[32], _027819_, _027820_);
  or g_119182_(_002628_, _027817_, _027821_);
  and g_119183_(out[33], _027812_, _027822_);
  not g_119184_(_027822_, _027823_);
  xor g_119185_(out[33], _027812_, _027824_);
  xor g_119186_(_002617_, _027812_, _027825_);
  and g_119187_(_027821_, _027824_, _027826_);
  or g_119188_(_027820_, _027825_, _027827_);
  and g_119189_(_005829_, _027693_, _027828_);
  and g_119190_(_005862_, _027694_, _027830_);
  or g_119191_(_027828_, _027830_, _027831_);
  not g_119192_(_027831_, _027832_);
  and g_119193_(_007842_, _027832_, _027833_);
  or g_119194_(_007853_, _027831_, _027834_);
  xor g_119195_(_007853_, _027831_, _027835_);
  xor g_119196_(_007842_, _027831_, _027836_);
  and g_119197_(_003674_, _027693_, _027837_);
  or g_119198_(_003675_, _027694_, _027838_);
  and g_119199_(_003672_, _027694_, _027839_);
  not g_119200_(_027839_, _027841_);
  and g_119201_(_027838_, _027841_, _027842_);
  or g_119202_(_027837_, _027839_, _027843_);
  and g_119203_(_003781_, _027843_, _027844_);
  or g_119204_(_003780_, _027842_, _027845_);
  and g_119205_(_003780_, _027842_, _027846_);
  or g_119206_(_003781_, _027843_, _027847_);
  or g_119207_(out[32], _027819_, _027848_);
  and g_119208_(_027835_, _027845_, _027849_);
  and g_119209_(_027847_, _027848_, _027850_);
  and g_119210_(_027826_, _027850_, _027852_);
  and g_119211_(_027849_, _027852_, _027853_);
  and g_119212_(_027743_, _027853_, _027854_);
  not g_119213_(_027854_, _027855_);
  and g_119214_(_027808_, _027854_, _027856_);
  or g_119215_(_027809_, _027855_, _027857_);
  and g_119216_(_027834_, _027847_, _027858_);
  or g_119217_(_027833_, _027846_, _027859_);
  and g_119218_(_027823_, _027827_, _027860_);
  or g_119219_(_027822_, _027826_, _027861_);
  and g_119220_(_027835_, _027861_, _027863_);
  or g_119221_(_027836_, _027860_, _027864_);
  and g_119222_(_027858_, _027864_, _027865_);
  or g_119223_(_027859_, _027863_, _027866_);
  and g_119224_(_027743_, _027845_, _027867_);
  or g_119225_(_027744_, _027844_, _027868_);
  and g_119226_(_027866_, _027867_, _027869_);
  or g_119227_(_027865_, _027868_, _027870_);
  and g_119228_(_027723_, _027737_, _027871_);
  and g_119229_(_027714_, _027715_, _027872_);
  or g_119230_(_027713_, _027872_, _027874_);
  or g_119231_(_027871_, _027874_, _027875_);
  not g_119232_(_027875_, _027876_);
  and g_119233_(_027870_, _027876_, _027877_);
  or g_119234_(_027869_, _027875_, _027878_);
  and g_119235_(_027808_, _027878_, _027879_);
  or g_119236_(_027809_, _027877_, _027880_);
  and g_119237_(_027798_, _027800_, _027881_);
  or g_119238_(_027778_, _027797_, _027882_);
  and g_119239_(_027777_, _027881_, _027883_);
  or g_119240_(_027799_, _027882_, _027885_);
  or g_119241_(_027766_, _027775_, _027886_);
  and g_119242_(_027767_, _027776_, _027887_);
  and g_119243_(_027885_, _027886_, _027888_);
  or g_119244_(_027883_, _027887_, _027889_);
  and g_119245_(_027880_, _027888_, _027890_);
  or g_119246_(_027879_, _027889_, _027891_);
  and g_119247_(_027857_, _027891_, _027892_);
  or g_119248_(_027856_, _027890_, _027893_);
  and g_119249_(_003781_, _027892_, _027894_);
  or g_119250_(_003780_, _027893_, _027896_);
  and g_119251_(_027842_, _027893_, _027897_);
  or g_119252_(_027843_, _027892_, _027898_);
  and g_119253_(_027896_, _027898_, _027899_);
  or g_119254_(_027894_, _027897_, _027900_);
  and g_119255_(_004060_, _027900_, _027901_);
  or g_119256_(_004061_, _027899_, _027902_);
  and g_119257_(_007842_, _027892_, _027903_);
  or g_119258_(_007853_, _027893_, _027904_);
  and g_119259_(_027831_, _027893_, _027905_);
  or g_119260_(_027832_, _027892_, _027907_);
  and g_119261_(_027904_, _027907_, _027908_);
  or g_119262_(_027903_, _027905_, _027909_);
  and g_119263_(_010834_, _027908_, _027910_);
  or g_119264_(_010845_, _027909_, _027911_);
  and g_119265_(_027902_, _027911_, _027912_);
  or g_119266_(_027901_, _027910_, _027913_);
  or g_119267_(_002617_, _027893_, _027914_);
  or g_119268_(_027812_, _027892_, _027915_);
  and g_119269_(_027914_, _027915_, _027916_);
  and g_119270_(out[49], _027916_, _027918_);
  not g_119271_(_027918_, _027919_);
  and g_119272_(_027819_, _027893_, _027920_);
  or g_119273_(_027817_, _027892_, _027921_);
  and g_119274_(_002628_, _027892_, _027922_);
  or g_119275_(out[32], _027893_, _027923_);
  and g_119276_(_027921_, _027923_, _027924_);
  or g_119277_(_027920_, _027922_, _027925_);
  and g_119278_(out[48], _027925_, _027926_);
  or g_119279_(_002760_, _027924_, _027927_);
  xor g_119280_(out[49], _027916_, _027929_);
  xor g_119281_(_002749_, _027916_, _027930_);
  and g_119282_(_027927_, _027929_, _027931_);
  or g_119283_(_027926_, _027930_, _027932_);
  and g_119284_(_027919_, _027932_, _027933_);
  or g_119285_(_027918_, _027931_, _027934_);
  and g_119286_(_010845_, _027909_, _027935_);
  or g_119287_(_010834_, _027908_, _027936_);
  and g_119288_(_027934_, _027936_, _027937_);
  or g_119289_(_027933_, _027935_, _027938_);
  and g_119290_(_027912_, _027938_, _027940_);
  or g_119291_(_027913_, _027937_, _027941_);
  and g_119292_(_027757_, _027764_, _027942_);
  or g_119293_(_027758_, _027765_, _027943_);
  or g_119294_(out[58], _003969_, _027944_);
  xor g_119295_(out[59], _027944_, _027945_);
  xor g_119296_(_002694_, _027944_, _027946_);
  and g_119297_(_027942_, _027946_, _027947_);
  or g_119298_(_027943_, _027945_, _027948_);
  xor g_119299_(out[58], _003969_, _027949_);
  xor g_119300_(_002815_, _003969_, _027951_);
  and g_119301_(_027754_, _027893_, _027952_);
  or g_119302_(_027753_, _027892_, _027953_);
  and g_119303_(_027746_, _027892_, _027954_);
  or g_119304_(_027747_, _027893_, _027955_);
  and g_119305_(_027953_, _027955_, _027956_);
  or g_119306_(_027952_, _027954_, _027957_);
  and g_119307_(_027949_, _027956_, _027958_);
  or g_119308_(_027951_, _027957_, _027959_);
  and g_119309_(_027948_, _027959_, _027960_);
  or g_119310_(_027947_, _027958_, _027962_);
  and g_119311_(_027951_, _027957_, _027963_);
  or g_119312_(_027949_, _027956_, _027964_);
  and g_119313_(_027943_, _027945_, _027965_);
  or g_119314_(_027942_, _027946_, _027966_);
  and g_119315_(_027964_, _027966_, _027967_);
  or g_119316_(_027963_, _027965_, _027968_);
  and g_119317_(_027960_, _027967_, _027969_);
  or g_119318_(_027962_, _027968_, _027970_);
  and g_119319_(_003730_, _027892_, _027971_);
  or g_119320_(_003731_, _027893_, _027973_);
  and g_119321_(_027783_, _027893_, _027974_);
  or g_119322_(_027784_, _027892_, _027975_);
  and g_119323_(_027973_, _027975_, _027976_);
  or g_119324_(_027971_, _027974_, _027977_);
  and g_119325_(_003976_, _027977_, _027978_);
  or g_119326_(_003975_, _027976_, _027979_);
  and g_119327_(_003719_, _027892_, _027980_);
  or g_119328_(_003720_, _027893_, _027981_);
  and g_119329_(_027793_, _027893_, _027982_);
  or g_119330_(_027792_, _027892_, _027984_);
  and g_119331_(_027981_, _027984_, _027985_);
  or g_119332_(_027980_, _027982_, _027986_);
  and g_119333_(_003972_, _027986_, _027987_);
  or g_119334_(_003971_, _027985_, _027988_);
  and g_119335_(_027979_, _027988_, _027989_);
  or g_119336_(_027978_, _027987_, _027990_);
  and g_119337_(_003971_, _027985_, _027991_);
  or g_119338_(_003972_, _027986_, _027992_);
  and g_119339_(_003975_, _027976_, _027993_);
  or g_119340_(_003976_, _027977_, _027995_);
  and g_119341_(_027992_, _027995_, _027996_);
  or g_119342_(_027991_, _027993_, _027997_);
  and g_119343_(_003833_, _027892_, _027998_);
  or g_119344_(_003832_, _027893_, _027999_);
  and g_119345_(_027711_, _027893_, _028000_);
  or g_119346_(_027712_, _027892_, _028001_);
  and g_119347_(_027999_, _028001_, _028002_);
  or g_119348_(_027998_, _028000_, _028003_);
  and g_119349_(_004009_, _028002_, _028004_);
  not g_119350_(_028004_, _028006_);
  and g_119351_(_003822_, _027892_, _028007_);
  or g_119352_(_003821_, _027893_, _028008_);
  and g_119353_(_027699_, _027893_, _028009_);
  or g_119354_(_027698_, _027892_, _028010_);
  and g_119355_(_028008_, _028010_, _028011_);
  or g_119356_(_028007_, _028009_, _028012_);
  and g_119357_(_004000_, _028011_, _028013_);
  or g_119358_(_003999_, _028012_, _028014_);
  and g_119359_(_004008_, _028003_, _028015_);
  or g_119360_(_004009_, _028002_, _028017_);
  and g_119361_(_003867_, _027892_, _028018_);
  or g_119362_(_003868_, _027893_, _028019_);
  and g_119363_(_027729_, _027893_, _028020_);
  or g_119364_(_027731_, _027892_, _028021_);
  and g_119365_(_028019_, _028021_, _028022_);
  or g_119366_(_028018_, _028020_, _028023_);
  and g_119367_(_004023_, _028023_, _028024_);
  or g_119368_(_004022_, _028022_, _028025_);
  and g_119369_(_003854_, _027892_, _028026_);
  or g_119370_(_003855_, _027893_, _028028_);
  and g_119371_(_027704_, _027893_, _028029_);
  or g_119372_(_027705_, _027892_, _028030_);
  and g_119373_(_028028_, _028030_, _028031_);
  or g_119374_(_028026_, _028029_, _028032_);
  and g_119375_(_004034_, _028032_, _028033_);
  or g_119376_(_004033_, _028031_, _028034_);
  and g_119377_(_028025_, _028034_, _028035_);
  or g_119378_(_028024_, _028033_, _028036_);
  and g_119379_(_004033_, _028031_, _028037_);
  or g_119380_(_004034_, _028032_, _028039_);
  and g_119381_(_004022_, _028022_, _028040_);
  or g_119382_(_004023_, _028023_, _028041_);
  and g_119383_(_027989_, _027996_, _028042_);
  or g_119384_(_027990_, _027997_, _028043_);
  and g_119385_(_027969_, _028042_, _028044_);
  or g_119386_(_027970_, _028043_, _028045_);
  xor g_119387_(_004000_, _028011_, _028046_);
  xor g_119388_(_003999_, _028011_, _028047_);
  and g_119389_(_028006_, _028046_, _028048_);
  or g_119390_(_028004_, _028047_, _028050_);
  and g_119391_(_028017_, _028048_, _028051_);
  or g_119392_(_028015_, _028050_, _028052_);
  and g_119393_(_028039_, _028051_, _028053_);
  or g_119394_(_028037_, _028052_, _028054_);
  and g_119395_(_028034_, _028041_, _028055_);
  or g_119396_(_028033_, _028040_, _028056_);
  and g_119397_(_028025_, _028055_, _028057_);
  or g_119398_(_028024_, _028056_, _028058_);
  and g_119399_(_028053_, _028057_, _028059_);
  or g_119400_(_028054_, _028058_, _028061_);
  and g_119401_(_028044_, _028059_, _028062_);
  or g_119402_(_028045_, _028061_, _028063_);
  and g_119403_(_004061_, _027899_, _028064_);
  or g_119404_(_004060_, _027900_, _028065_);
  and g_119405_(_027941_, _028062_, _028066_);
  or g_119406_(_027940_, _028063_, _028067_);
  and g_119407_(_028065_, _028066_, _028068_);
  or g_119408_(_028064_, _028067_, _028069_);
  and g_119409_(_028036_, _028039_, _028070_);
  or g_119410_(_028035_, _028037_, _028072_);
  and g_119411_(_028006_, _028013_, _028073_);
  or g_119412_(_028004_, _028014_, _028074_);
  and g_119413_(_028051_, _028070_, _028075_);
  or g_119414_(_028052_, _028072_, _028076_);
  and g_119415_(_028074_, _028076_, _028077_);
  or g_119416_(_028073_, _028075_, _028078_);
  and g_119417_(_028017_, _028077_, _028079_);
  or g_119418_(_028015_, _028078_, _028080_);
  and g_119419_(_028044_, _028080_, _028081_);
  or g_119420_(_028045_, _028079_, _028083_);
  and g_119421_(_027990_, _027992_, _028084_);
  or g_119422_(_027989_, _027991_, _028085_);
  and g_119423_(_027969_, _028084_, _028086_);
  or g_119424_(_027970_, _028085_, _028087_);
  and g_119425_(_027962_, _027966_, _028088_);
  or g_119426_(_027960_, _027965_, _028089_);
  and g_119427_(_028087_, _028089_, _028090_);
  or g_119428_(_028086_, _028088_, _028091_);
  and g_119429_(_028083_, _028090_, _028092_);
  or g_119430_(_028081_, _028091_, _028094_);
  and g_119431_(_028069_, _028092_, _028095_);
  or g_119432_(_028068_, _028094_, _028096_);
  and g_119433_(_002760_, _027924_, _028097_);
  not g_119434_(_028097_, _028098_);
  and g_119435_(_027936_, _028065_, _028099_);
  and g_119436_(_028098_, _028099_, _028100_);
  and g_119437_(_027912_, _028100_, _028101_);
  and g_119438_(_027931_, _028101_, _028102_);
  not g_119439_(_028102_, _028103_);
  and g_119440_(_028062_, _028102_, _028105_);
  or g_119441_(_028063_, _028103_, _028106_);
  and g_119442_(_028096_, _028106_, _028107_);
  or g_119443_(_028095_, _028105_, _028108_);
  or g_119444_(_004060_, _028108_, _028109_);
  or g_119445_(_027899_, _028107_, _028110_);
  and g_119446_(_028109_, _028110_, _028111_);
  or g_119447_(_004276_, _028111_, _028112_);
  and g_119448_(_027909_, _028108_, _028113_);
  and g_119449_(_010834_, _028107_, _028114_);
  or g_119450_(_028113_, _028114_, _028116_);
  and g_119451_(_004276_, _028111_, _028117_);
  or g_119452_(_026630_, _028116_, _028118_);
  xor g_119453_(_004276_, _028111_, _028119_);
  xor g_119454_(_004275_, _028111_, _028120_);
  xor g_119455_(_026630_, _028116_, _028121_);
  xor g_119456_(_026619_, _028116_, _028122_);
  and g_119457_(_028119_, _028121_, _028123_);
  or g_119458_(_028120_, _028122_, _028124_);
  or g_119459_(_002749_, _028108_, _028125_);
  or g_119460_(_027916_, _028107_, _028127_);
  and g_119461_(_028125_, _028127_, _028128_);
  and g_119462_(out[65], _028128_, _028129_);
  not g_119463_(_028129_, _028130_);
  or g_119464_(_028117_, _028118_, _028131_);
  and g_119465_(_028112_, _028131_, _028132_);
  not g_119466_(_028132_, _028133_);
  or g_119467_(_027924_, _028107_, _028134_);
  not g_119468_(_028134_, _028135_);
  and g_119469_(_002760_, _028107_, _028136_);
  not g_119470_(_028136_, _028138_);
  and g_119471_(_028134_, _028138_, _028139_);
  or g_119472_(_028135_, _028136_, _028140_);
  and g_119473_(out[64], _028140_, _028141_);
  or g_119474_(_002892_, _028139_, _028142_);
  xor g_119475_(out[65], _028128_, _028143_);
  xor g_119476_(_002881_, _028128_, _028144_);
  and g_119477_(_028142_, _028143_, _028145_);
  or g_119478_(_028141_, _028144_, _028146_);
  and g_119479_(_028130_, _028146_, _028147_);
  or g_119480_(_028129_, _028145_, _028149_);
  and g_119481_(_028123_, _028149_, _028150_);
  or g_119482_(_028124_, _028147_, _028151_);
  and g_119483_(_028132_, _028151_, _028152_);
  or g_119484_(_028133_, _028150_, _028153_);
  and g_119485_(_027942_, _027945_, _028154_);
  or g_119486_(_027943_, _027946_, _028155_);
  or g_119487_(out[74], _004183_, _028156_);
  xor g_119488_(out[75], _028156_, _028157_);
  xor g_119489_(_002826_, _028156_, _028158_);
  and g_119490_(_028154_, _028158_, _028160_);
  or g_119491_(_028155_, _028157_, _028161_);
  and g_119492_(_027957_, _028108_, _028162_);
  or g_119493_(_027956_, _028107_, _028163_);
  and g_119494_(_027949_, _028107_, _028164_);
  or g_119495_(_027951_, _028108_, _028165_);
  and g_119496_(_028163_, _028165_, _028166_);
  or g_119497_(_028162_, _028164_, _028167_);
  xor g_119498_(out[74], _004183_, _028168_);
  xor g_119499_(_002947_, _004183_, _028169_);
  and g_119500_(_028166_, _028168_, _028171_);
  or g_119501_(_028167_, _028169_, _028172_);
  and g_119502_(_028161_, _028172_, _028173_);
  or g_119503_(_028160_, _028171_, _028174_);
  and g_119504_(_028155_, _028157_, _028175_);
  or g_119505_(_028154_, _028158_, _028176_);
  and g_119506_(_028167_, _028169_, _028177_);
  or g_119507_(_028166_, _028168_, _028178_);
  and g_119508_(_028176_, _028178_, _028179_);
  or g_119509_(_028175_, _028177_, _028180_);
  and g_119510_(_028173_, _028179_, _028182_);
  or g_119511_(_028174_, _028180_, _028183_);
  and g_119512_(_003975_, _028107_, _028184_);
  or g_119513_(_003976_, _028108_, _028185_);
  and g_119514_(_027977_, _028108_, _028186_);
  or g_119515_(_027976_, _028107_, _028187_);
  and g_119516_(_028185_, _028187_, _028188_);
  or g_119517_(_028184_, _028186_, _028189_);
  and g_119518_(_004192_, _028189_, _028190_);
  or g_119519_(_004191_, _028188_, _028191_);
  and g_119520_(_003971_, _028107_, _028193_);
  or g_119521_(_003972_, _028108_, _028194_);
  and g_119522_(_027986_, _028108_, _028195_);
  or g_119523_(_027985_, _028107_, _028196_);
  and g_119524_(_028194_, _028196_, _028197_);
  or g_119525_(_028193_, _028195_, _028198_);
  and g_119526_(_004185_, _028198_, _028199_);
  or g_119527_(_004184_, _028197_, _028200_);
  and g_119528_(_028191_, _028200_, _028201_);
  or g_119529_(_028190_, _028199_, _028202_);
  and g_119530_(_004184_, _028197_, _028204_);
  or g_119531_(_004185_, _028198_, _028205_);
  and g_119532_(_004191_, _028188_, _028206_);
  or g_119533_(_004192_, _028189_, _028207_);
  and g_119534_(_028205_, _028207_, _028208_);
  or g_119535_(_028204_, _028206_, _028209_);
  and g_119536_(_028201_, _028208_, _028210_);
  or g_119537_(_028202_, _028209_, _028211_);
  and g_119538_(_028182_, _028210_, _028212_);
  or g_119539_(_028183_, _028211_, _028213_);
  or g_119540_(_003999_, _028108_, _028215_);
  or g_119541_(_028011_, _028107_, _028216_);
  and g_119542_(_028215_, _028216_, _028217_);
  not g_119543_(_028217_, _028218_);
  and g_119544_(_004222_, _028217_, _028219_);
  or g_119545_(_004221_, _028218_, _028220_);
  xor g_119546_(_004222_, _028217_, _028221_);
  xor g_119547_(_004221_, _028217_, _028222_);
  and g_119548_(_004009_, _028107_, _028223_);
  or g_119549_(_004008_, _028108_, _028224_);
  and g_119550_(_028003_, _028108_, _028226_);
  or g_119551_(_028002_, _028107_, _028227_);
  and g_119552_(_028224_, _028227_, _028228_);
  or g_119553_(_028223_, _028226_, _028229_);
  and g_119554_(_004215_, _028229_, _028230_);
  or g_119555_(_004216_, _028228_, _028231_);
  and g_119556_(_004033_, _028107_, _028232_);
  or g_119557_(_004034_, _028108_, _028233_);
  and g_119558_(_028032_, _028108_, _028234_);
  or g_119559_(_028031_, _028107_, _028235_);
  and g_119560_(_028233_, _028235_, _028237_);
  or g_119561_(_028232_, _028234_, _028238_);
  and g_119562_(_004249_, _028237_, _028239_);
  or g_119563_(_004250_, _028238_, _028240_);
  and g_119564_(_004022_, _028107_, _028241_);
  not g_119565_(_028241_, _028242_);
  or g_119566_(_028022_, _028107_, _028243_);
  not g_119567_(_028243_, _028244_);
  and g_119568_(_028242_, _028243_, _028245_);
  or g_119569_(_028241_, _028244_, _028246_);
  and g_119570_(_004239_, _028246_, _028248_);
  or g_119571_(_004238_, _028245_, _028249_);
  and g_119572_(_004250_, _028238_, _028250_);
  or g_119573_(_004249_, _028237_, _028251_);
  and g_119574_(_028249_, _028251_, _028252_);
  or g_119575_(_028248_, _028250_, _028253_);
  and g_119576_(_004216_, _028228_, _028254_);
  or g_119577_(_004215_, _028229_, _028255_);
  and g_119578_(_004238_, _028245_, _028256_);
  or g_119579_(_004239_, _028246_, _028257_);
  and g_119580_(_028252_, _028257_, _028259_);
  or g_119581_(_028253_, _028256_, _028260_);
  and g_119582_(_028231_, _028255_, _028261_);
  or g_119583_(_028230_, _028254_, _028262_);
  and g_119584_(_028221_, _028261_, _028263_);
  or g_119585_(_028222_, _028262_, _028264_);
  and g_119586_(_028240_, _028263_, _028265_);
  or g_119587_(_028239_, _028264_, _028266_);
  and g_119588_(_028259_, _028265_, _028267_);
  or g_119589_(_028260_, _028266_, _028268_);
  and g_119590_(_028212_, _028267_, _028270_);
  or g_119591_(_028213_, _028268_, _028271_);
  and g_119592_(_028174_, _028176_, _028272_);
  or g_119593_(_028173_, _028175_, _028273_);
  and g_119594_(_028202_, _028205_, _028274_);
  or g_119595_(_028201_, _028204_, _028275_);
  and g_119596_(_028182_, _028274_, _028276_);
  or g_119597_(_028183_, _028275_, _028277_);
  and g_119598_(_028273_, _028277_, _028278_);
  or g_119599_(_028272_, _028276_, _028279_);
  and g_119600_(_028153_, _028267_, _028281_);
  or g_119601_(_028152_, _028268_, _028282_);
  and g_119602_(_028253_, _028265_, _028283_);
  or g_119603_(_028252_, _028266_, _028284_);
  and g_119604_(_028219_, _028255_, _028285_);
  or g_119605_(_028220_, _028254_, _028286_);
  and g_119606_(_028231_, _028286_, _028287_);
  or g_119607_(_028230_, _028285_, _028288_);
  and g_119608_(_028284_, _028287_, _028289_);
  or g_119609_(_028283_, _028288_, _028290_);
  and g_119610_(_028282_, _028289_, _028292_);
  or g_119611_(_028281_, _028290_, _028293_);
  and g_119612_(_028212_, _028293_, _028294_);
  or g_119613_(_028213_, _028292_, _028295_);
  and g_119614_(_028278_, _028295_, _028296_);
  or g_119615_(_028279_, _028294_, _028297_);
  and g_119616_(_002892_, _028139_, _028298_);
  or g_119617_(out[64], _028140_, _028299_);
  and g_119618_(_028145_, _028299_, _028300_);
  or g_119619_(_028146_, _028298_, _028301_);
  and g_119620_(_028123_, _028300_, _028303_);
  or g_119621_(_028124_, _028301_, _028304_);
  and g_119622_(_028270_, _028303_, _028305_);
  or g_119623_(_028271_, _028304_, _028306_);
  and g_119624_(_028297_, _028306_, _028307_);
  or g_119625_(_028296_, _028305_, _028308_);
  or g_119626_(_004215_, _028308_, _028309_);
  or g_119627_(_028228_, _028307_, _028310_);
  and g_119628_(_028309_, _028310_, _028311_);
  or g_119629_(_004449_, _028311_, _028312_);
  and g_119630_(_004449_, _028311_, _028314_);
  xor g_119631_(_004448_, _028311_, _028315_);
  or g_119632_(_004250_, _028308_, _028316_);
  or g_119633_(_028237_, _028307_, _028317_);
  and g_119634_(_028316_, _028317_, _028318_);
  and g_119635_(_004473_, _028318_, _028319_);
  and g_119636_(_004222_, _028307_, _028320_);
  and g_119637_(_028218_, _028308_, _028321_);
  or g_119638_(_028320_, _028321_, _028322_);
  not g_119639_(_028322_, _028323_);
  or g_119640_(_004439_, _028322_, _028325_);
  xor g_119641_(_004440_, _028322_, _028326_);
  or g_119642_(_028315_, _028326_, _028327_);
  or g_119643_(_028319_, _028327_, _028328_);
  not g_119644_(_028328_, _028329_);
  and g_119645_(_028154_, _028157_, _028330_);
  or g_119646_(_028155_, _028158_, _028331_);
  or g_119647_(out[90], _004403_, _028332_);
  xor g_119648_(out[91], _028332_, _028333_);
  xor g_119649_(_002958_, _028332_, _028334_);
  and g_119650_(_028330_, _028334_, _028336_);
  or g_119651_(_028331_, _028333_, _028337_);
  and g_119652_(_028168_, _028307_, _028338_);
  or g_119653_(_028169_, _028308_, _028339_);
  and g_119654_(_028167_, _028308_, _028340_);
  or g_119655_(_028166_, _028307_, _028341_);
  and g_119656_(_028339_, _028341_, _028342_);
  or g_119657_(_028338_, _028340_, _028343_);
  xor g_119658_(out[90], _004403_, _028344_);
  xor g_119659_(_003079_, _004403_, _028345_);
  and g_119660_(_028342_, _028344_, _028347_);
  or g_119661_(_028343_, _028345_, _028348_);
  and g_119662_(_028337_, _028348_, _028349_);
  or g_119663_(_028336_, _028347_, _028350_);
  and g_119664_(_028343_, _028345_, _028351_);
  or g_119665_(_028342_, _028344_, _028352_);
  and g_119666_(_028331_, _028333_, _028353_);
  or g_119667_(_028330_, _028334_, _028354_);
  and g_119668_(_028352_, _028354_, _028355_);
  or g_119669_(_028351_, _028353_, _028356_);
  and g_119670_(_028349_, _028355_, _028358_);
  or g_119671_(_028350_, _028356_, _028359_);
  and g_119672_(_004191_, _028307_, _028360_);
  or g_119673_(_004192_, _028308_, _028361_);
  and g_119674_(_028189_, _028308_, _028362_);
  or g_119675_(_028188_, _028307_, _028363_);
  and g_119676_(_028361_, _028363_, _028364_);
  or g_119677_(_028360_, _028362_, _028365_);
  and g_119678_(_004409_, _028365_, _028366_);
  or g_119679_(_004408_, _028364_, _028367_);
  and g_119680_(_004184_, _028307_, _028369_);
  or g_119681_(_004185_, _028308_, _028370_);
  and g_119682_(_028198_, _028308_, _028371_);
  or g_119683_(_028197_, _028307_, _028372_);
  and g_119684_(_028370_, _028372_, _028373_);
  or g_119685_(_028369_, _028371_, _028374_);
  and g_119686_(_004405_, _028374_, _028375_);
  or g_119687_(_004404_, _028373_, _028376_);
  and g_119688_(_028367_, _028376_, _028377_);
  or g_119689_(_028366_, _028375_, _028378_);
  and g_119690_(_004404_, _028373_, _028380_);
  or g_119691_(_004405_, _028374_, _028381_);
  and g_119692_(_004408_, _028364_, _028382_);
  or g_119693_(_004409_, _028365_, _028383_);
  and g_119694_(_028381_, _028383_, _028384_);
  or g_119695_(_028380_, _028382_, _028385_);
  and g_119696_(_028377_, _028384_, _028386_);
  or g_119697_(_028378_, _028385_, _028387_);
  and g_119698_(_028358_, _028386_, _028388_);
  or g_119699_(_028359_, _028387_, _028389_);
  or g_119700_(_004239_, _028308_, _028391_);
  or g_119701_(_028245_, _028307_, _028392_);
  and g_119702_(_028391_, _028392_, _028393_);
  not g_119703_(_028393_, _028394_);
  and g_119704_(_004462_, _028393_, _028395_);
  not g_119705_(_028395_, _028396_);
  or g_119706_(_004462_, _028393_, _028397_);
  or g_119707_(_004473_, _028318_, _028398_);
  and g_119708_(_028397_, _028398_, _028399_);
  not g_119709_(_028399_, _028400_);
  and g_119710_(_028396_, _028399_, _028402_);
  or g_119711_(_028395_, _028400_, _028403_);
  and g_119712_(_028388_, _028402_, _028404_);
  or g_119713_(_028389_, _028403_, _028405_);
  and g_119714_(_028329_, _028404_, _028406_);
  or g_119715_(_028328_, _028405_, _028407_);
  or g_119716_(_004275_, _028308_, _028408_);
  or g_119717_(_028111_, _028307_, _028409_);
  and g_119718_(_028408_, _028409_, _028410_);
  not g_119719_(_028410_, _028411_);
  and g_119720_(_004501_, _028410_, _028413_);
  or g_119721_(_004500_, _028411_, _028414_);
  and g_119722_(_028116_, _028308_, _028415_);
  not g_119723_(_028415_, _028416_);
  or g_119724_(_026630_, _028308_, _028417_);
  not g_119725_(_028417_, _028418_);
  and g_119726_(_028416_, _028417_, _028419_);
  or g_119727_(_028415_, _028418_, _028420_);
  and g_119728_(_026586_, _028419_, _028421_);
  or g_119729_(_026597_, _028420_, _028422_);
  and g_119730_(_028414_, _028422_, _028424_);
  or g_119731_(_028413_, _028421_, _028425_);
  and g_119732_(_004500_, _028411_, _028426_);
  or g_119733_(_004501_, _028410_, _028427_);
  and g_119734_(_026597_, _028420_, _028428_);
  or g_119735_(_026586_, _028419_, _028429_);
  and g_119736_(_028427_, _028429_, _028430_);
  or g_119737_(_028426_, _028428_, _028431_);
  and g_119738_(_028424_, _028430_, _028432_);
  or g_119739_(_028425_, _028431_, _028433_);
  and g_119740_(_028406_, _028432_, _028435_);
  or g_119741_(_028407_, _028433_, _028436_);
  or g_119742_(_002881_, _028308_, _028437_);
  or g_119743_(_028128_, _028307_, _028438_);
  and g_119744_(_028437_, _028438_, _028439_);
  and g_119745_(out[81], _028439_, _028440_);
  not g_119746_(_028440_, _028441_);
  and g_119747_(_028435_, _028440_, _028442_);
  or g_119748_(_028436_, _028441_, _028443_);
  or g_119749_(_028328_, _028399_, _028444_);
  or g_119750_(_028314_, _028325_, _028446_);
  and g_119751_(_028312_, _028446_, _028447_);
  and g_119752_(_028444_, _028447_, _028448_);
  not g_119753_(_028448_, _028449_);
  and g_119754_(_028388_, _028449_, _028450_);
  or g_119755_(_028389_, _028448_, _028451_);
  and g_119756_(_028422_, _028427_, _028452_);
  or g_119757_(_028421_, _028426_, _028453_);
  and g_119758_(_028414_, _028453_, _028454_);
  or g_119759_(_028413_, _028452_, _028455_);
  and g_119760_(_028406_, _028454_, _028457_);
  or g_119761_(_028407_, _028455_, _028458_);
  and g_119762_(_028350_, _028354_, _028459_);
  or g_119763_(_028349_, _028353_, _028460_);
  and g_119764_(_028378_, _028381_, _028461_);
  or g_119765_(_028377_, _028380_, _028462_);
  and g_119766_(_028358_, _028461_, _028463_);
  or g_119767_(_028359_, _028462_, _028464_);
  and g_119768_(_028460_, _028464_, _028465_);
  or g_119769_(_028459_, _028463_, _028466_);
  and g_119770_(_028458_, _028465_, _028468_);
  or g_119771_(_028457_, _028466_, _028469_);
  and g_119772_(_028451_, _028468_, _028470_);
  or g_119773_(_028450_, _028469_, _028471_);
  and g_119774_(_028443_, _028470_, _028472_);
  or g_119775_(_028442_, _028471_, _028473_);
  and g_119776_(_028140_, _028308_, _028474_);
  not g_119777_(_028474_, _028475_);
  or g_119778_(out[64], _028308_, _028476_);
  not g_119779_(_028476_, _028477_);
  and g_119780_(_028475_, _028476_, _028479_);
  or g_119781_(_028474_, _028477_, _028480_);
  and g_119782_(out[80], _028480_, _028481_);
  or g_119783_(_003024_, _028479_, _028482_);
  xor g_119784_(out[81], _028439_, _028483_);
  xor g_119785_(_003013_, _028439_, _028484_);
  and g_119786_(_028482_, _028483_, _028485_);
  or g_119787_(_028481_, _028484_, _028486_);
  and g_119788_(_028435_, _028485_, _028487_);
  or g_119789_(_028436_, _028486_, _028488_);
  and g_119790_(_003024_, _028479_, _028490_);
  or g_119791_(out[80], _028480_, _028491_);
  and g_119792_(_028487_, _028490_, _028492_);
  or g_119793_(_028488_, _028491_, _028493_);
  and g_119794_(_028472_, _028493_, _028494_);
  or g_119795_(_028473_, _028492_, _028495_);
  or g_119796_(_004500_, _028494_, _028496_);
  or g_119797_(_028410_, _028495_, _028497_);
  and g_119798_(_028496_, _028497_, _028498_);
  not g_119799_(_028498_, _028499_);
  and g_119800_(_004599_, _028498_, _028501_);
  or g_119801_(_004599_, _028498_, _028502_);
  xor g_119802_(_004599_, _028498_, _028503_);
  xor g_119803_(_004598_, _028498_, _028504_);
  and g_119804_(_026586_, _028495_, _028505_);
  and g_119805_(_028420_, _028494_, _028506_);
  or g_119806_(_028505_, _028506_, _028507_);
  or g_119807_(_031217_, _028507_, _028508_);
  xor g_119808_(_031217_, _028507_, _028509_);
  xor g_119809_(_031206_, _028507_, _028510_);
  and g_119810_(_028503_, _028509_, _028512_);
  or g_119811_(_028504_, _028510_, _028513_);
  or g_119812_(_028439_, _028495_, _028514_);
  or g_119813_(_003013_, _028494_, _028515_);
  and g_119814_(_028514_, _028515_, _028516_);
  not g_119815_(_028516_, _028517_);
  and g_119816_(out[97], _028516_, _028518_);
  and g_119817_(out[80], _028473_, _028519_);
  or g_119818_(_003024_, _028472_, _028520_);
  and g_119819_(_028479_, _028494_, _028521_);
  not g_119820_(_028521_, _028523_);
  and g_119821_(_028520_, _028523_, _028524_);
  or g_119822_(_028519_, _028521_, _028525_);
  or g_119823_(_003156_, _028525_, _028526_);
  xor g_119824_(out[97], _028516_, _028527_);
  and g_119825_(_028526_, _028527_, _028528_);
  or g_119826_(_028518_, _028528_, _028529_);
  not g_119827_(_028529_, _028530_);
  and g_119828_(_028512_, _028529_, _028531_);
  or g_119829_(_028513_, _028530_, _028532_);
  and g_119830_(_028502_, _028508_, _028534_);
  or g_119831_(_028501_, _028534_, _028535_);
  not g_119832_(_028535_, _028536_);
  and g_119833_(_028532_, _028535_, _028537_);
  or g_119834_(_028531_, _028536_, _028538_);
  and g_119835_(_028330_, _028333_, _028539_);
  or g_119836_(_028331_, _028334_, _028540_);
  or g_119837_(out[106], _004650_, _028541_);
  xor g_119838_(out[107], _028541_, _028542_);
  xor g_119839_(_003090_, _028541_, _028543_);
  and g_119840_(_028539_, _028543_, _028545_);
  or g_119841_(_028540_, _028542_, _028546_);
  and g_119842_(_028344_, _028495_, _028547_);
  or g_119843_(_028345_, _028494_, _028548_);
  and g_119844_(_028343_, _028494_, _028549_);
  or g_119845_(_028342_, _028495_, _028550_);
  and g_119846_(_028548_, _028550_, _028551_);
  or g_119847_(_028547_, _028549_, _028552_);
  xor g_119848_(out[106], _004650_, _028553_);
  xor g_119849_(_003211_, _004650_, _028554_);
  and g_119850_(_028551_, _028553_, _028556_);
  or g_119851_(_028552_, _028554_, _028557_);
  and g_119852_(_028546_, _028557_, _028558_);
  or g_119853_(_028545_, _028556_, _028559_);
  and g_119854_(_028552_, _028554_, _028560_);
  or g_119855_(_028551_, _028553_, _028561_);
  and g_119856_(_028540_, _028542_, _028562_);
  or g_119857_(_028539_, _028543_, _028563_);
  and g_119858_(_028561_, _028563_, _028564_);
  or g_119859_(_028560_, _028562_, _028565_);
  and g_119860_(_028558_, _028564_, _028567_);
  or g_119861_(_028559_, _028565_, _028568_);
  and g_119862_(_028365_, _028494_, _028569_);
  not g_119863_(_028569_, _028570_);
  or g_119864_(_004409_, _028494_, _028571_);
  not g_119865_(_028571_, _028572_);
  and g_119866_(_028570_, _028571_, _028573_);
  or g_119867_(_028569_, _028572_, _028574_);
  and g_119868_(_004664_, _028574_, _028575_);
  or g_119869_(_004662_, _028573_, _028576_);
  or g_119870_(_004405_, _028494_, _028578_);
  not g_119871_(_028578_, _028579_);
  and g_119872_(_028374_, _028494_, _028580_);
  not g_119873_(_028580_, _028581_);
  and g_119874_(_028578_, _028581_, _028582_);
  or g_119875_(_028579_, _028580_, _028583_);
  and g_119876_(_004653_, _028583_, _028584_);
  or g_119877_(_004651_, _028582_, _028585_);
  and g_119878_(_028576_, _028585_, _028586_);
  or g_119879_(_028575_, _028584_, _028587_);
  and g_119880_(_004651_, _028582_, _028589_);
  or g_119881_(_004653_, _028583_, _028590_);
  and g_119882_(_004662_, _028573_, _028591_);
  or g_119883_(_004664_, _028574_, _028592_);
  and g_119884_(_028590_, _028592_, _028593_);
  or g_119885_(_028589_, _028591_, _028594_);
  and g_119886_(_028586_, _028593_, _028595_);
  or g_119887_(_028587_, _028594_, _028596_);
  and g_119888_(_028567_, _028595_, _028597_);
  or g_119889_(_028568_, _028596_, _028598_);
  or g_119890_(_028311_, _028495_, _028600_);
  or g_119891_(_004448_, _028494_, _028601_);
  and g_119892_(_028600_, _028601_, _028602_);
  not g_119893_(_028602_, _028603_);
  or g_119894_(_004692_, _028602_, _028604_);
  and g_119895_(_004692_, _028602_, _028605_);
  or g_119896_(_004691_, _028603_, _028606_);
  and g_119897_(_028604_, _028606_, _028607_);
  xor g_119898_(_004691_, _028602_, _028608_);
  or g_119899_(_028323_, _028495_, _028609_);
  or g_119900_(_004439_, _028494_, _028611_);
  and g_119901_(_028609_, _028611_, _028612_);
  not g_119902_(_028612_, _028613_);
  and g_119903_(_004702_, _028612_, _028614_);
  or g_119904_(_004701_, _028613_, _028615_);
  xor g_119905_(_004702_, _028612_, _028616_);
  xor g_119906_(_004701_, _028612_, _028617_);
  and g_119907_(_028607_, _028616_, _028618_);
  or g_119908_(_028608_, _028617_, _028619_);
  and g_119909_(_004474_, _028495_, _028620_);
  or g_119910_(_004473_, _028494_, _028622_);
  and g_119911_(_028318_, _028494_, _028623_);
  not g_119912_(_028623_, _028624_);
  or g_119913_(_028620_, _028623_, _028625_);
  and g_119914_(_028622_, _028624_, _028626_);
  or g_119915_(_004725_, _028625_, _028627_);
  or g_119916_(_004463_, _028494_, _028628_);
  not g_119917_(_028628_, _028629_);
  and g_119918_(_028394_, _028494_, _028630_);
  not g_119919_(_028630_, _028631_);
  and g_119920_(_028628_, _028631_, _028633_);
  or g_119921_(_028629_, _028630_, _028634_);
  or g_119922_(_004714_, _028633_, _028635_);
  and g_119923_(_028627_, _028635_, _028636_);
  and g_119924_(_004725_, _028625_, _028637_);
  or g_119925_(_004726_, _028626_, _028638_);
  or g_119926_(_004715_, _028634_, _028639_);
  and g_119927_(_028638_, _028639_, _028640_);
  xor g_119928_(_004715_, _028633_, _028641_);
  xor g_119929_(_004726_, _028625_, _028642_);
  and g_119930_(_028636_, _028640_, _028644_);
  or g_119931_(_028641_, _028642_, _028645_);
  and g_119932_(_028618_, _028644_, _028646_);
  or g_119933_(_028619_, _028645_, _028647_);
  and g_119934_(_028597_, _028646_, _028648_);
  or g_119935_(_028598_, _028647_, _028649_);
  and g_119936_(_028538_, _028648_, _028650_);
  or g_119937_(_028537_, _028649_, _028651_);
  or g_119938_(_028619_, _028637_, _028652_);
  or g_119939_(_028636_, _028652_, _028653_);
  and g_119940_(_028606_, _028614_, _028655_);
  or g_119941_(_028605_, _028615_, _028656_);
  and g_119942_(_028604_, _028653_, _028657_);
  not g_119943_(_028657_, _028658_);
  and g_119944_(_028656_, _028657_, _028659_);
  or g_119945_(_028655_, _028658_, _028660_);
  and g_119946_(_028597_, _028660_, _028661_);
  or g_119947_(_028598_, _028659_, _028662_);
  and g_119948_(_028559_, _028563_, _028663_);
  or g_119949_(_028558_, _028562_, _028664_);
  and g_119950_(_028567_, _028587_, _028666_);
  or g_119951_(_028568_, _028586_, _028667_);
  and g_119952_(_028590_, _028666_, _028668_);
  or g_119953_(_028589_, _028667_, _028669_);
  and g_119954_(_028651_, _028669_, _028670_);
  or g_119955_(_028650_, _028668_, _028671_);
  and g_119956_(_028662_, _028664_, _028672_);
  or g_119957_(_028663_, _028671_, _028673_);
  and g_119958_(_028670_, _028672_, _028674_);
  or g_119959_(_028661_, _028673_, _028675_);
  or g_119960_(out[96], _028524_, _028677_);
  and g_119961_(_028528_, _028677_, _028678_);
  not g_119962_(_028678_, _028679_);
  and g_119963_(_028512_, _028648_, _028680_);
  or g_119964_(_028513_, _028649_, _028681_);
  and g_119965_(_028678_, _028680_, _028682_);
  or g_119966_(_028679_, _028681_, _028683_);
  and g_119967_(_028675_, _028683_, _028684_);
  or g_119968_(_028674_, _028682_, _028685_);
  and g_119969_(_003156_, _028684_, _028686_);
  or g_119970_(out[96], _028685_, _028688_);
  and g_119971_(_028524_, _028685_, _028689_);
  or g_119972_(_028525_, _028684_, _028690_);
  and g_119973_(_028688_, _028690_, _028691_);
  or g_119974_(_028686_, _028689_, _028692_);
  and g_119975_(_028539_, _028542_, _028693_);
  or g_119976_(_028540_, _028543_, _028694_);
  or g_119977_(out[122], _004815_, _028695_);
  xor g_119978_(out[123], _028695_, _028696_);
  xor g_119979_(_003222_, _028695_, _028697_);
  and g_119980_(_028693_, _028697_, _028699_);
  or g_119981_(_028694_, _028696_, _028700_);
  and g_119982_(_028553_, _028684_, _028701_);
  and g_119983_(_028552_, _028685_, _028702_);
  or g_119984_(_028701_, _028702_, _028703_);
  xor g_119985_(_003343_, _004815_, _028704_);
  or g_119986_(_028703_, _028704_, _028705_);
  not g_119987_(_028705_, _028706_);
  and g_119988_(_028700_, _028705_, _028707_);
  or g_119989_(_028699_, _028706_, _028708_);
  and g_119990_(_028694_, _028696_, _028710_);
  or g_119991_(_028693_, _028697_, _028711_);
  and g_119992_(_028703_, _028704_, _028712_);
  or g_119993_(_028710_, _028712_, _028713_);
  not g_119994_(_028713_, _028714_);
  and g_119995_(_028707_, _028714_, _028715_);
  or g_119996_(_028708_, _028713_, _028716_);
  and g_119997_(_004651_, _028684_, _028717_);
  and g_119998_(_028583_, _028685_, _028718_);
  or g_119999_(_028717_, _028718_, _028719_);
  and g_120000_(_004818_, _028719_, _028721_);
  not g_120001_(_028721_, _028722_);
  and g_120002_(_004662_, _028684_, _028723_);
  and g_120003_(_028574_, _028685_, _028724_);
  or g_120004_(_028723_, _028724_, _028725_);
  and g_120005_(_004829_, _028725_, _028726_);
  not g_120006_(_028726_, _028727_);
  and g_120007_(_028722_, _028727_, _028728_);
  or g_120008_(_028721_, _028726_, _028729_);
  or g_120009_(_004818_, _028719_, _028730_);
  or g_120010_(_004829_, _028725_, _028732_);
  and g_120011_(_028730_, _028732_, _028733_);
  not g_120012_(_028733_, _028734_);
  and g_120013_(_028728_, _028733_, _028735_);
  or g_120014_(_028729_, _028734_, _028736_);
  and g_120015_(_028715_, _028735_, _028737_);
  or g_120016_(_028716_, _028736_, _028738_);
  and g_120017_(_004692_, _028684_, _028739_);
  or g_120018_(_004691_, _028685_, _028740_);
  and g_120019_(_028603_, _028685_, _028741_);
  or g_120020_(_028602_, _028684_, _028743_);
  and g_120021_(_028740_, _028743_, _028744_);
  or g_120022_(_028739_, _028741_, _028745_);
  or g_120023_(_004864_, _028744_, _028746_);
  and g_120024_(_004864_, _028744_, _028747_);
  xor g_120025_(_004864_, _028744_, _028748_);
  xor g_120026_(_004863_, _028744_, _028749_);
  and g_120027_(_004702_, _028684_, _028750_);
  and g_120028_(_028613_, _028685_, _028751_);
  or g_120029_(_028750_, _028751_, _028752_);
  or g_120030_(_004856_, _028752_, _028754_);
  and g_120031_(_004725_, _028684_, _028755_);
  and g_120032_(_028626_, _028685_, _028756_);
  or g_120033_(_028755_, _028756_, _028757_);
  or g_120034_(_004897_, _028757_, _028758_);
  not g_120035_(_028758_, _028759_);
  xor g_120036_(_004856_, _028752_, _028760_);
  xor g_120037_(_004857_, _028752_, _028761_);
  and g_120038_(_028748_, _028760_, _028762_);
  or g_120039_(_028749_, _028761_, _028763_);
  and g_120040_(_028758_, _028762_, _028765_);
  or g_120041_(_028759_, _028763_, _028766_);
  and g_120042_(_004714_, _028684_, _028767_);
  and g_120043_(_028634_, _028685_, _028768_);
  or g_120044_(_028767_, _028768_, _028769_);
  and g_120045_(_004886_, _028769_, _028770_);
  not g_120046_(_028770_, _028771_);
  and g_120047_(_004897_, _028757_, _028772_);
  not g_120048_(_028772_, _028773_);
  and g_120049_(_028771_, _028773_, _028774_);
  or g_120050_(_028770_, _028772_, _028776_);
  or g_120051_(_004886_, _028769_, _028777_);
  not g_120052_(_028777_, _028778_);
  and g_120053_(_028774_, _028777_, _028779_);
  or g_120054_(_028776_, _028778_, _028780_);
  and g_120055_(_028765_, _028779_, _028781_);
  or g_120056_(_028766_, _028780_, _028782_);
  and g_120057_(_004599_, _028684_, _028783_);
  and g_120058_(_028499_, _028685_, _028784_);
  or g_120059_(_028783_, _028784_, _028785_);
  or g_120060_(_004952_, _028785_, _028787_);
  and g_120061_(_004952_, _028785_, _028788_);
  xor g_120062_(_004952_, _028785_, _028789_);
  xor g_120063_(_004953_, _028785_, _028790_);
  and g_120064_(_028507_, _028685_, _028791_);
  and g_120065_(_031206_, _028684_, _028792_);
  or g_120066_(_028791_, _028792_, _028793_);
  not g_120067_(_028793_, _028794_);
  and g_120068_(_034121_, _028794_, _028795_);
  xor g_120069_(_034132_, _028793_, _028796_);
  xor g_120070_(_034121_, _028793_, _028798_);
  and g_120071_(_028789_, _028796_, _028799_);
  or g_120072_(_028790_, _028798_, _028800_);
  and g_120073_(out[97], _028684_, _028801_);
  or g_120074_(_003145_, _028685_, _028802_);
  and g_120075_(_028517_, _028685_, _028803_);
  or g_120076_(_028516_, _028684_, _028804_);
  and g_120077_(_028802_, _028804_, _028805_);
  or g_120078_(_028801_, _028803_, _028806_);
  and g_120079_(out[113], _028805_, _028807_);
  or g_120080_(_003277_, _028806_, _028809_);
  and g_120081_(out[112], _028692_, _028810_);
  or g_120082_(_003288_, _028691_, _028811_);
  xor g_120083_(out[113], _028805_, _028812_);
  xor g_120084_(_003277_, _028805_, _028813_);
  and g_120085_(_028811_, _028812_, _028814_);
  or g_120086_(_028810_, _028813_, _028815_);
  and g_120087_(_028809_, _028815_, _028816_);
  or g_120088_(_028807_, _028814_, _028817_);
  and g_120089_(_028799_, _028817_, _028818_);
  or g_120090_(_028800_, _028816_, _028820_);
  and g_120091_(_028787_, _028795_, _028821_);
  or g_120092_(_028788_, _028821_, _028822_);
  not g_120093_(_028822_, _028823_);
  and g_120094_(_028820_, _028823_, _028824_);
  or g_120095_(_028818_, _028822_, _028825_);
  and g_120096_(_028781_, _028825_, _028826_);
  or g_120097_(_028782_, _028824_, _028827_);
  and g_120098_(_028765_, _028776_, _028828_);
  or g_120099_(_028766_, _028774_, _028829_);
  or g_120100_(_028747_, _028754_, _028831_);
  and g_120101_(_028746_, _028831_, _028832_);
  not g_120102_(_028832_, _028833_);
  and g_120103_(_028829_, _028832_, _028834_);
  or g_120104_(_028828_, _028833_, _028835_);
  and g_120105_(_028827_, _028834_, _028836_);
  or g_120106_(_028826_, _028835_, _028837_);
  and g_120107_(_028737_, _028837_, _028838_);
  or g_120108_(_028738_, _028836_, _028839_);
  and g_120109_(_028708_, _028711_, _028840_);
  or g_120110_(_028707_, _028710_, _028842_);
  and g_120111_(_028729_, _028730_, _028843_);
  not g_120112_(_028843_, _028844_);
  and g_120113_(_028715_, _028843_, _028845_);
  or g_120114_(_028716_, _028844_, _028846_);
  and g_120115_(_028842_, _028846_, _028847_);
  or g_120116_(_028840_, _028845_, _028848_);
  and g_120117_(_028839_, _028847_, _028849_);
  or g_120118_(_028838_, _028848_, _028850_);
  or g_120119_(out[112], _028692_, _028851_);
  not g_120120_(_028851_, _028853_);
  or g_120121_(_028815_, _028853_, _028854_);
  or g_120122_(_028800_, _028854_, _028855_);
  or g_120123_(_028738_, _028855_, _028856_);
  not g_120124_(_028856_, _028857_);
  and g_120125_(_028781_, _028857_, _028858_);
  or g_120126_(_028782_, _028856_, _028859_);
  and g_120127_(_028850_, _028859_, _028860_);
  or g_120128_(_028849_, _028858_, _028861_);
  and g_120129_(_028692_, _028861_, _028862_);
  and g_120130_(_003288_, _028860_, _028864_);
  or g_120131_(_028862_, _028864_, _028865_);
  and g_120132_(_028693_, _028696_, _028866_);
  or g_120133_(_028694_, _028697_, _028867_);
  or g_120134_(out[138], _005042_, _028868_);
  xor g_120135_(out[139], _028868_, _028869_);
  xor g_120136_(_003354_, _028868_, _028870_);
  and g_120137_(_028866_, _028870_, _028871_);
  or g_120138_(_028867_, _028869_, _028872_);
  or g_120139_(_028704_, _028861_, _028873_);
  not g_120140_(_028873_, _028875_);
  and g_120141_(_028703_, _028861_, _028876_);
  or g_120142_(_028875_, _028876_, _028877_);
  xor g_120143_(_003475_, _005042_, _028878_);
  or g_120144_(_028877_, _028878_, _028879_);
  not g_120145_(_028879_, _028880_);
  and g_120146_(_028872_, _028879_, _028881_);
  or g_120147_(_028871_, _028880_, _028882_);
  and g_120148_(_028867_, _028869_, _028883_);
  or g_120149_(_028866_, _028870_, _028884_);
  and g_120150_(_028877_, _028878_, _028886_);
  or g_120151_(_028883_, _028886_, _028887_);
  not g_120152_(_028887_, _028888_);
  and g_120153_(_028881_, _028888_, _028889_);
  or g_120154_(_028882_, _028887_, _028890_);
  and g_120155_(_004827_, _028860_, _028891_);
  and g_120156_(_028725_, _028861_, _028892_);
  or g_120157_(_028891_, _028892_, _028893_);
  not g_120158_(_028893_, _028894_);
  and g_120159_(_005055_, _028893_, _028895_);
  or g_120160_(_005054_, _028894_, _028897_);
  and g_120161_(_004816_, _028860_, _028898_);
  and g_120162_(_028719_, _028861_, _028899_);
  or g_120163_(_028898_, _028899_, _028900_);
  not g_120164_(_028900_, _028901_);
  and g_120165_(_005044_, _028900_, _028902_);
  or g_120166_(_005043_, _028901_, _028903_);
  and g_120167_(_028897_, _028903_, _028904_);
  or g_120168_(_028895_, _028902_, _028905_);
  or g_120169_(_005044_, _028900_, _028906_);
  or g_120170_(_005055_, _028893_, _028908_);
  and g_120171_(_028906_, _028908_, _028909_);
  not g_120172_(_028909_, _028910_);
  and g_120173_(_028904_, _028909_, _028911_);
  or g_120174_(_028905_, _028910_, _028912_);
  and g_120175_(_028889_, _028911_, _028913_);
  or g_120176_(_028890_, _028912_, _028914_);
  and g_120177_(_004857_, _028860_, _028915_);
  and g_120178_(_028752_, _028861_, _028916_);
  or g_120179_(_028915_, _028916_, _028917_);
  or g_120180_(_005090_, _028917_, _028919_);
  not g_120181_(_028919_, _028920_);
  xor g_120182_(_005090_, _028917_, _028921_);
  xor g_120183_(_005091_, _028917_, _028922_);
  and g_120184_(_004896_, _028860_, _028923_);
  and g_120185_(_028757_, _028861_, _028924_);
  or g_120186_(_028923_, _028924_, _028925_);
  or g_120187_(_005119_, _028925_, _028926_);
  not g_120188_(_028926_, _028927_);
  and g_120189_(_004864_, _028860_, _028928_);
  and g_120190_(_028745_, _028861_, _028930_);
  or g_120191_(_028928_, _028930_, _028931_);
  or g_120192_(_005084_, _028931_, _028932_);
  and g_120193_(_005084_, _028931_, _028933_);
  xor g_120194_(_005084_, _028931_, _028934_);
  xor g_120195_(_005085_, _028931_, _028935_);
  and g_120196_(_028921_, _028934_, _028936_);
  or g_120197_(_028922_, _028935_, _028937_);
  and g_120198_(_028926_, _028936_, _028938_);
  or g_120199_(_028927_, _028937_, _028939_);
  and g_120200_(_004885_, _028860_, _028941_);
  and g_120201_(_028769_, _028861_, _028942_);
  or g_120202_(_028941_, _028942_, _028943_);
  or g_120203_(_005108_, _028943_, _028944_);
  and g_120204_(_005108_, _028943_, _028945_);
  not g_120205_(_028945_, _028946_);
  and g_120206_(_005119_, _028925_, _028947_);
  not g_120207_(_028947_, _028948_);
  and g_120208_(_028946_, _028948_, _028949_);
  or g_120209_(_028945_, _028947_, _028950_);
  and g_120210_(_028944_, _028949_, _028952_);
  and g_120211_(_028938_, _028952_, _028953_);
  and g_120212_(_028913_, _028953_, _028954_);
  or g_120213_(out[128], _028865_, _028955_);
  or g_120214_(_004952_, _028861_, _028956_);
  not g_120215_(_028956_, _028957_);
  and g_120216_(_028785_, _028861_, _028958_);
  not g_120217_(_028958_, _028959_);
  and g_120218_(_028956_, _028959_, _028960_);
  or g_120219_(_028957_, _028958_, _028961_);
  and g_120220_(_005145_, _028960_, _028963_);
  or g_120221_(_005144_, _028961_, _028964_);
  and g_120222_(_028793_, _028861_, _028965_);
  not g_120223_(_028965_, _028966_);
  or g_120224_(_034132_, _028861_, _028967_);
  not g_120225_(_028967_, _028968_);
  and g_120226_(_028966_, _028967_, _028969_);
  or g_120227_(_028965_, _028968_, _028970_);
  and g_120228_(_036200_, _028970_, _028971_);
  or g_120229_(_028963_, _028971_, _028972_);
  and g_120230_(_005144_, _028961_, _028974_);
  and g_120231_(_036189_, _028969_, _028975_);
  or g_120232_(_028974_, _028975_, _028976_);
  xor g_120233_(_005145_, _028960_, _028977_);
  xor g_120234_(_036189_, _028969_, _028978_);
  and g_120235_(_028977_, _028978_, _028979_);
  or g_120236_(_028972_, _028976_, _028980_);
  or g_120237_(_003277_, _028861_, _028981_);
  or g_120238_(_028805_, _028860_, _028982_);
  and g_120239_(_028981_, _028982_, _028983_);
  and g_120240_(out[129], _028983_, _028985_);
  xor g_120241_(out[129], _028983_, _028986_);
  xor g_120242_(_003409_, _028983_, _028987_);
  and g_120243_(out[128], _028865_, _028988_);
  not g_120244_(_028988_, _028989_);
  and g_120245_(_028986_, _028989_, _028990_);
  or g_120246_(_028987_, _028988_, _028991_);
  and g_120247_(_028979_, _028990_, _028992_);
  or g_120248_(_028980_, _028991_, _028993_);
  and g_120249_(_028954_, _028955_, _028994_);
  not g_120250_(_028994_, _028996_);
  and g_120251_(_028992_, _028994_, _028997_);
  or g_120252_(_028993_, _028996_, _028998_);
  and g_120253_(_028938_, _028950_, _028999_);
  or g_120254_(_028939_, _028949_, _029000_);
  and g_120255_(_028920_, _028932_, _029001_);
  or g_120256_(_028933_, _029001_, _029002_);
  not g_120257_(_029002_, _029003_);
  and g_120258_(_029000_, _029003_, _029004_);
  or g_120259_(_028999_, _029002_, _029005_);
  and g_120260_(_028913_, _029005_, _029007_);
  or g_120261_(_028914_, _029004_, _029008_);
  and g_120262_(_028979_, _028985_, _029009_);
  and g_120263_(_028964_, _028976_, _029010_);
  or g_120264_(_028992_, _029010_, _029011_);
  or g_120265_(_029009_, _029011_, _029012_);
  and g_120266_(_028954_, _029012_, _029013_);
  not g_120267_(_029013_, _029014_);
  and g_120268_(_028905_, _028906_, _029015_);
  not g_120269_(_029015_, _029016_);
  and g_120270_(_028889_, _029015_, _029018_);
  or g_120271_(_028890_, _029016_, _029019_);
  and g_120272_(_028882_, _028884_, _029020_);
  or g_120273_(_028881_, _028883_, _029021_);
  and g_120274_(_029008_, _029019_, _029022_);
  or g_120275_(_029007_, _029018_, _029023_);
  and g_120276_(_029014_, _029022_, _029024_);
  or g_120277_(_029013_, _029023_, _029025_);
  and g_120278_(_029021_, _029024_, _029026_);
  or g_120279_(_029020_, _029025_, _029027_);
  and g_120280_(_028998_, _029027_, _029029_);
  or g_120281_(_028997_, _029026_, _029030_);
  and g_120282_(_028865_, _029030_, _029031_);
  not g_120283_(_029031_, _029032_);
  or g_120284_(out[128], _029030_, _029033_);
  not g_120285_(_029033_, _029034_);
  and g_120286_(_029032_, _029033_, _029035_);
  or g_120287_(_029031_, _029034_, _029036_);
  and g_120288_(_005107_, _029029_, _029037_);
  and g_120289_(_028943_, _029030_, _029038_);
  or g_120290_(_029037_, _029038_, _029040_);
  not g_120291_(_029040_, _029041_);
  and g_120292_(_005309_, _029040_, _029042_);
  not g_120293_(_029042_, _029043_);
  and g_120294_(_005118_, _029029_, _029044_);
  and g_120295_(_028925_, _029030_, _029045_);
  or g_120296_(_029044_, _029045_, _029046_);
  and g_120297_(_005320_, _029046_, _029047_);
  not g_120298_(_029047_, _029048_);
  and g_120299_(_029043_, _029048_, _029049_);
  or g_120300_(_029042_, _029047_, _029051_);
  and g_120301_(_005308_, _029041_, _029052_);
  or g_120302_(_005309_, _029040_, _029053_);
  and g_120303_(_036189_, _029029_, _029054_);
  or g_120304_(_036200_, _029030_, _029055_);
  and g_120305_(_028970_, _029030_, _029056_);
  or g_120306_(_028969_, _029029_, _029057_);
  and g_120307_(_029055_, _029057_, _029058_);
  or g_120308_(_029054_, _029056_, _029059_);
  and g_120309_(_038466_, _029058_, _029060_);
  or g_120310_(_038477_, _029059_, _029062_);
  and g_120311_(_005145_, _029029_, _029063_);
  or g_120312_(_005144_, _029030_, _029064_);
  and g_120313_(_028961_, _029030_, _029065_);
  or g_120314_(_028960_, _029029_, _029066_);
  and g_120315_(_029064_, _029066_, _029067_);
  or g_120316_(_029063_, _029065_, _029068_);
  and g_120317_(_005375_, _029068_, _029069_);
  or g_120318_(_005376_, _029067_, _029070_);
  and g_120319_(_029062_, _029070_, _029071_);
  or g_120320_(_029060_, _029069_, _029073_);
  and g_120321_(_038477_, _029059_, _029074_);
  not g_120322_(_029074_, _029075_);
  or g_120323_(_005375_, _029068_, _029076_);
  not g_120324_(_029076_, _029077_);
  and g_120325_(_029071_, _029076_, _029078_);
  or g_120326_(_029073_, _029077_, _029079_);
  and g_120327_(_029075_, _029078_, _029080_);
  or g_120328_(_029074_, _029079_, _029081_);
  or g_120329_(_003409_, _029030_, _029082_);
  or g_120330_(_028983_, _029029_, _029084_);
  and g_120331_(_029082_, _029084_, _029085_);
  and g_120332_(out[145], _029085_, _029086_);
  not g_120333_(_029086_, _029087_);
  and g_120334_(out[144], _029036_, _029088_);
  or g_120335_(_003552_, _029035_, _029089_);
  xor g_120336_(out[145], _029085_, _029090_);
  xor g_120337_(_003541_, _029085_, _029091_);
  and g_120338_(_029089_, _029090_, _029092_);
  or g_120339_(_029088_, _029091_, _029093_);
  and g_120340_(_029087_, _029093_, _029095_);
  or g_120341_(_029086_, _029092_, _029096_);
  and g_120342_(_029080_, _029096_, _029097_);
  or g_120343_(_029081_, _029095_, _029098_);
  and g_120344_(_029073_, _029076_, _029099_);
  or g_120345_(_029071_, _029077_, _029100_);
  and g_120346_(_029098_, _029100_, _029101_);
  or g_120347_(_029097_, _029099_, _029102_);
  and g_120348_(_029053_, _029102_, _029103_);
  or g_120349_(_029052_, _029101_, _029104_);
  and g_120350_(_029049_, _029104_, _029106_);
  or g_120351_(_029051_, _029103_, _029107_);
  and g_120352_(_028866_, _028869_, _029108_);
  or g_120353_(_028867_, _028870_, _029109_);
  or g_120354_(out[154], _005244_, _029110_);
  xor g_120355_(out[155], _029110_, _029111_);
  xor g_120356_(_003486_, _029110_, _029112_);
  and g_120357_(_029108_, _029112_, _029113_);
  or g_120358_(_029109_, _029111_, _029114_);
  or g_120359_(_028878_, _029030_, _029115_);
  not g_120360_(_029115_, _029117_);
  and g_120361_(_028877_, _029030_, _029118_);
  or g_120362_(_029117_, _029118_, _029119_);
  xor g_120363_(_003607_, _005244_, _029120_);
  or g_120364_(_029119_, _029120_, _029121_);
  not g_120365_(_029121_, _029122_);
  and g_120366_(_029114_, _029121_, _029123_);
  or g_120367_(_029113_, _029122_, _029124_);
  and g_120368_(_029119_, _029120_, _029125_);
  and g_120369_(_029109_, _029111_, _029126_);
  or g_120370_(_029108_, _029112_, _029128_);
  or g_120371_(_029125_, _029126_, _029129_);
  not g_120372_(_029129_, _029130_);
  and g_120373_(_029123_, _029130_, _029131_);
  or g_120374_(_029124_, _029129_, _029132_);
  and g_120375_(_005054_, _029029_, _029133_);
  and g_120376_(_028893_, _029030_, _029134_);
  or g_120377_(_029133_, _029134_, _029135_);
  and g_120378_(_005258_, _029135_, _029136_);
  not g_120379_(_029136_, _029137_);
  and g_120380_(_005043_, _029029_, _029139_);
  and g_120381_(_028900_, _029030_, _029140_);
  or g_120382_(_029139_, _029140_, _029141_);
  and g_120383_(_005247_, _029141_, _029142_);
  not g_120384_(_029142_, _029143_);
  and g_120385_(_029137_, _029143_, _029144_);
  or g_120386_(_029136_, _029142_, _029145_);
  or g_120387_(_005247_, _029141_, _029146_);
  or g_120388_(_005258_, _029135_, _029147_);
  and g_120389_(_029146_, _029147_, _029148_);
  not g_120390_(_029148_, _029150_);
  and g_120391_(_029144_, _029148_, _029151_);
  or g_120392_(_029145_, _029150_, _029152_);
  and g_120393_(_029131_, _029151_, _029153_);
  or g_120394_(_029132_, _029152_, _029154_);
  or g_120395_(_005084_, _029030_, _029155_);
  not g_120396_(_029155_, _029156_);
  and g_120397_(_028931_, _029030_, _029157_);
  not g_120398_(_029157_, _029158_);
  and g_120399_(_029155_, _029158_, _029159_);
  or g_120400_(_029156_, _029157_, _029161_);
  and g_120401_(_005285_, _029161_, _029162_);
  or g_120402_(_005286_, _029159_, _029163_);
  or g_120403_(_005090_, _029030_, _029164_);
  not g_120404_(_029164_, _029165_);
  and g_120405_(_028917_, _029030_, _029166_);
  not g_120406_(_029166_, _029167_);
  and g_120407_(_029164_, _029167_, _029168_);
  or g_120408_(_029165_, _029166_, _029169_);
  and g_120409_(_005293_, _029168_, _029170_);
  or g_120410_(_005292_, _029169_, _029172_);
  and g_120411_(_029163_, _029172_, _029173_);
  or g_120412_(_029162_, _029170_, _029174_);
  or g_120413_(_005320_, _029046_, _029175_);
  not g_120414_(_029175_, _029176_);
  and g_120415_(_005286_, _029159_, _029177_);
  or g_120416_(_005285_, _029161_, _029178_);
  and g_120417_(_005292_, _029169_, _029179_);
  or g_120418_(_005293_, _029168_, _029180_);
  and g_120419_(_029178_, _029180_, _029181_);
  or g_120420_(_029177_, _029179_, _029183_);
  and g_120421_(_029175_, _029181_, _029184_);
  or g_120422_(_029176_, _029183_, _029185_);
  and g_120423_(_029173_, _029184_, _029186_);
  or g_120424_(_029174_, _029185_, _029187_);
  and g_120425_(_029153_, _029186_, _029188_);
  or g_120426_(_029154_, _029187_, _029189_);
  and g_120427_(_029107_, _029188_, _029190_);
  or g_120428_(_029106_, _029189_, _029191_);
  and g_120429_(_029170_, _029178_, _029192_);
  or g_120430_(_029172_, _029177_, _029194_);
  and g_120431_(_029163_, _029194_, _029195_);
  or g_120432_(_029162_, _029192_, _029196_);
  and g_120433_(_029153_, _029196_, _029197_);
  or g_120434_(_029154_, _029195_, _029198_);
  and g_120435_(_029145_, _029146_, _029199_);
  not g_120436_(_029199_, _029200_);
  and g_120437_(_029131_, _029199_, _029201_);
  or g_120438_(_029132_, _029200_, _029202_);
  and g_120439_(_029124_, _029128_, _029203_);
  or g_120440_(_029123_, _029126_, _029205_);
  and g_120441_(_029202_, _029205_, _029206_);
  or g_120442_(_029201_, _029203_, _029207_);
  and g_120443_(_029198_, _029206_, _029208_);
  or g_120444_(_029197_, _029207_, _029209_);
  and g_120445_(_029191_, _029208_, _029210_);
  or g_120446_(_029190_, _029209_, _029211_);
  or g_120447_(out[144], _029036_, _029212_);
  and g_120448_(_029053_, _029212_, _029213_);
  not g_120449_(_029213_, _029214_);
  and g_120450_(_029049_, _029213_, _029216_);
  or g_120451_(_029051_, _029214_, _029217_);
  and g_120452_(_029080_, _029216_, _029218_);
  or g_120453_(_029081_, _029217_, _029219_);
  and g_120454_(_029092_, _029218_, _029220_);
  or g_120455_(_029093_, _029219_, _029221_);
  and g_120456_(_029188_, _029220_, _029222_);
  or g_120457_(_029189_, _029221_, _029223_);
  and g_120458_(_029211_, _029223_, _029224_);
  or g_120459_(_029210_, _029222_, _029225_);
  and g_120460_(_029036_, _029225_, _029227_);
  and g_120461_(_003552_, _029224_, _029228_);
  or g_120462_(_029227_, _029228_, _029229_);
  and g_120463_(_005293_, _029224_, _029230_);
  and g_120464_(_029169_, _029225_, _029231_);
  or g_120465_(_029230_, _029231_, _029232_);
  and g_120466_(_029161_, _029225_, _029233_);
  or g_120467_(_029159_, _029224_, _029234_);
  or g_120468_(_005285_, _029225_, _029235_);
  not g_120469_(_029235_, _029236_);
  and g_120470_(_029234_, _029235_, _029238_);
  or g_120471_(_029233_, _029236_, _029239_);
  and g_120472_(_005494_, _029239_, _029240_);
  not g_120473_(_029240_, _029241_);
  or g_120474_(_005505_, _029232_, _029242_);
  and g_120475_(_005495_, _029238_, _029243_);
  and g_120476_(_005319_, _029224_, _029244_);
  and g_120477_(_029046_, _029225_, _029245_);
  or g_120478_(_029244_, _029245_, _029246_);
  or g_120479_(_005517_, _029246_, _029247_);
  not g_120480_(_029247_, _029249_);
  xor g_120481_(_005505_, _029232_, _029250_);
  xor g_120482_(_005506_, _029232_, _029251_);
  or g_120483_(_029243_, _029251_, _029252_);
  xor g_120484_(_005494_, _029239_, _029253_);
  and g_120485_(_029250_, _029253_, _029254_);
  or g_120486_(_029240_, _029252_, _029255_);
  or g_120487_(_029249_, _029255_, _029256_);
  and g_120488_(_029108_, _029111_, _029257_);
  or g_120489_(_029109_, _029112_, _029258_);
  or g_120490_(out[170], _005464_, _029260_);
  xor g_120491_(out[171], _029260_, _029261_);
  xor g_120492_(_003618_, _029260_, _029262_);
  and g_120493_(_029257_, _029262_, _029263_);
  or g_120494_(_029258_, _029261_, _029264_);
  or g_120495_(_029120_, _029225_, _029265_);
  not g_120496_(_029265_, _029266_);
  and g_120497_(_029119_, _029225_, _029267_);
  not g_120498_(_029267_, _029268_);
  and g_120499_(_029265_, _029268_, _029269_);
  or g_120500_(_029266_, _029267_, _029271_);
  xor g_120501_(out[170], _005464_, _029272_);
  xor g_120502_(_003739_, _005464_, _029273_);
  and g_120503_(_029269_, _029272_, _029274_);
  or g_120504_(_029271_, _029273_, _029275_);
  and g_120505_(_029264_, _029275_, _029276_);
  or g_120506_(_029263_, _029274_, _029277_);
  and g_120507_(_029271_, _029273_, _029278_);
  and g_120508_(_029258_, _029261_, _029279_);
  or g_120509_(_029278_, _029279_, _029280_);
  not g_120510_(_029280_, _029282_);
  and g_120511_(_029276_, _029282_, _029283_);
  or g_120512_(_029277_, _029280_, _029284_);
  and g_120513_(_005256_, _029224_, _029285_);
  and g_120514_(_029135_, _029225_, _029286_);
  or g_120515_(_029285_, _029286_, _029287_);
  not g_120516_(_029287_, _029288_);
  and g_120517_(_005482_, _029287_, _029289_);
  or g_120518_(_005481_, _029288_, _029290_);
  and g_120519_(_005245_, _029224_, _029291_);
  and g_120520_(_029141_, _029225_, _029293_);
  or g_120521_(_029291_, _029293_, _029294_);
  not g_120522_(_029294_, _029295_);
  and g_120523_(_005467_, _029294_, _029296_);
  or g_120524_(_005465_, _029295_, _029297_);
  and g_120525_(_029290_, _029297_, _029298_);
  or g_120526_(_029289_, _029296_, _029299_);
  or g_120527_(_005467_, _029294_, _029300_);
  or g_120528_(_005482_, _029287_, _029301_);
  and g_120529_(_029300_, _029301_, _029302_);
  not g_120530_(_029302_, _029304_);
  and g_120531_(_029298_, _029302_, _029305_);
  or g_120532_(_029299_, _029304_, _029306_);
  and g_120533_(_029283_, _029305_, _029307_);
  or g_120534_(_029284_, _029306_, _029308_);
  and g_120535_(_005308_, _029224_, _029309_);
  and g_120536_(_029040_, _029225_, _029310_);
  or g_120537_(_029309_, _029310_, _029311_);
  and g_120538_(_005530_, _029311_, _029312_);
  not g_120539_(_029312_, _029313_);
  and g_120540_(_005517_, _029246_, _029315_);
  not g_120541_(_029315_, _029316_);
  and g_120542_(_029313_, _029316_, _029317_);
  or g_120543_(_029312_, _029315_, _029318_);
  or g_120544_(_005530_, _029311_, _029319_);
  not g_120545_(_029319_, _029320_);
  or g_120546_(_029318_, _029320_, _029321_);
  or g_120547_(_029308_, _029321_, _029322_);
  and g_120548_(_029247_, _029319_, _029323_);
  and g_120549_(_029317_, _029323_, _029324_);
  and g_120550_(_029254_, _029324_, _029326_);
  and g_120551_(_029307_, _029326_, _029327_);
  or g_120552_(_029256_, _029322_, _029328_);
  or g_120553_(_005375_, _029225_, _029329_);
  not g_120554_(_029329_, _029330_);
  and g_120555_(_029068_, _029225_, _029331_);
  not g_120556_(_029331_, _029332_);
  and g_120557_(_029329_, _029332_, _029333_);
  or g_120558_(_029330_, _029331_, _029334_);
  or g_120559_(_005560_, _029333_, _029335_);
  and g_120560_(_005560_, _029333_, _029337_);
  xor g_120561_(_005560_, _029333_, _029338_);
  xor g_120562_(_005559_, _029333_, _029339_);
  and g_120563_(_029059_, _029225_, _029340_);
  and g_120564_(_038466_, _029224_, _029341_);
  or g_120565_(_029340_, _029341_, _029342_);
  or g_120566_(_040578_, _029342_, _029343_);
  xor g_120567_(_040578_, _029342_, _029344_);
  xor g_120568_(_040567_, _029342_, _029345_);
  and g_120569_(_029338_, _029344_, _029346_);
  or g_120570_(_029339_, _029345_, _029348_);
  or g_120571_(_003541_, _029225_, _029349_);
  or g_120572_(_029085_, _029224_, _029350_);
  and g_120573_(_029349_, _029350_, _029351_);
  and g_120574_(out[161], _029351_, _029352_);
  not g_120575_(_029352_, _029353_);
  and g_120576_(out[160], _029229_, _029354_);
  not g_120577_(_029354_, _029355_);
  xor g_120578_(out[161], _029351_, _029356_);
  xor g_120579_(_003673_, _029351_, _029357_);
  and g_120580_(_029355_, _029356_, _029359_);
  or g_120581_(_029354_, _029357_, _029360_);
  and g_120582_(_029353_, _029360_, _029361_);
  or g_120583_(_029348_, _029361_, _029362_);
  and g_120584_(_029335_, _029343_, _029363_);
  or g_120585_(_029337_, _029363_, _029364_);
  and g_120586_(_029362_, _029364_, _029365_);
  or g_120587_(_029328_, _029365_, _029366_);
  or g_120588_(_029256_, _029317_, _029367_);
  or g_120589_(_029242_, _029243_, _029368_);
  and g_120590_(_029241_, _029368_, _029370_);
  and g_120591_(_029367_, _029370_, _029371_);
  or g_120592_(_029308_, _029371_, _029372_);
  and g_120593_(_029299_, _029300_, _029373_);
  not g_120594_(_029373_, _029374_);
  or g_120595_(_029284_, _029374_, _029375_);
  or g_120596_(_029276_, _029279_, _029376_);
  and g_120597_(_029375_, _029376_, _029377_);
  and g_120598_(_029372_, _029377_, _029378_);
  and g_120599_(_029366_, _029378_, _029379_);
  or g_120600_(out[160], _029229_, _029381_);
  and g_120601_(_029346_, _029381_, _029382_);
  and g_120602_(_029359_, _029382_, _029383_);
  and g_120603_(_029327_, _029383_, _029384_);
  or g_120604_(_029379_, _029384_, _029385_);
  not g_120605_(_029385_, _029386_);
  and g_120606_(_029229_, _029385_, _029387_);
  and g_120607_(_003684_, _029386_, _029388_);
  or g_120608_(_029387_, _029388_, _029389_);
  and g_120609_(_029257_, _029261_, _029390_);
  or g_120610_(_029258_, _029262_, _029392_);
  or g_120611_(out[186], _005673_, _029393_);
  xor g_120612_(out[187], _029393_, _029394_);
  xor g_120613_(_003750_, _029393_, _029395_);
  and g_120614_(_029390_, _029395_, _029396_);
  or g_120615_(_029392_, _029394_, _029397_);
  or g_120616_(_029273_, _029385_, _029398_);
  not g_120617_(_029398_, _029399_);
  and g_120618_(_029271_, _029385_, _029400_);
  not g_120619_(_029400_, _029401_);
  and g_120620_(_029398_, _029401_, _029403_);
  or g_120621_(_029399_, _029400_, _029404_);
  xor g_120622_(out[186], _005673_, _029405_);
  xor g_120623_(_003871_, _005673_, _029406_);
  and g_120624_(_029403_, _029405_, _029407_);
  or g_120625_(_029404_, _029406_, _029408_);
  and g_120626_(_029397_, _029408_, _029409_);
  or g_120627_(_029396_, _029407_, _029410_);
  and g_120628_(_029404_, _029406_, _029411_);
  and g_120629_(_029392_, _029394_, _029412_);
  or g_120630_(_029411_, _029412_, _029414_);
  not g_120631_(_029414_, _029415_);
  and g_120632_(_029409_, _029415_, _029416_);
  or g_120633_(_029410_, _029414_, _029417_);
  and g_120634_(_005481_, _029386_, _029418_);
  and g_120635_(_029287_, _029385_, _029419_);
  or g_120636_(_029418_, _029419_, _029420_);
  and g_120637_(_005663_, _029420_, _029421_);
  not g_120638_(_029421_, _029422_);
  and g_120639_(_005465_, _029386_, _029423_);
  and g_120640_(_029294_, _029385_, _029425_);
  or g_120641_(_029423_, _029425_, _029426_);
  and g_120642_(_005676_, _029426_, _029427_);
  not g_120643_(_029427_, _029428_);
  and g_120644_(_029422_, _029428_, _029429_);
  or g_120645_(_029421_, _029427_, _029430_);
  or g_120646_(_005676_, _029426_, _029431_);
  or g_120647_(_005663_, _029420_, _029432_);
  and g_120648_(_029431_, _029432_, _029433_);
  not g_120649_(_029433_, _029434_);
  and g_120650_(_029429_, _029433_, _029436_);
  or g_120651_(_029430_, _029434_, _029437_);
  and g_120652_(_029416_, _029436_, _029438_);
  or g_120653_(_029417_, _029437_, _029439_);
  and g_120654_(_005506_, _029386_, _029440_);
  and g_120655_(_029232_, _029385_, _029441_);
  or g_120656_(_029440_, _029441_, _029442_);
  or g_120657_(_005714_, _029442_, _029443_);
  not g_120658_(_029443_, _029444_);
  xor g_120659_(_005714_, _029442_, _029445_);
  xor g_120660_(_005715_, _029442_, _029447_);
  and g_120661_(_005495_, _029386_, _029448_);
  and g_120662_(_029239_, _029385_, _029449_);
  or g_120663_(_029448_, _029449_, _029450_);
  and g_120664_(_005699_, _029450_, _029451_);
  or g_120665_(_005699_, _029450_, _029452_);
  xor g_120666_(_005699_, _029450_, _029453_);
  xor g_120667_(_005700_, _029450_, _029454_);
  and g_120668_(_029445_, _029453_, _029455_);
  or g_120669_(_029447_, _029454_, _029456_);
  and g_120670_(_005529_, _029386_, _029458_);
  and g_120671_(_029311_, _029385_, _029459_);
  or g_120672_(_029458_, _029459_, _029460_);
  and g_120673_(_005748_, _029460_, _029461_);
  not g_120674_(_029461_, _029462_);
  and g_120675_(_005516_, _029386_, _029463_);
  and g_120676_(_029246_, _029385_, _029464_);
  or g_120677_(_029463_, _029464_, _029465_);
  and g_120678_(_005726_, _029465_, _029466_);
  not g_120679_(_029466_, _029467_);
  and g_120680_(_029462_, _029467_, _029469_);
  or g_120681_(_029461_, _029466_, _029470_);
  or g_120682_(_005726_, _029465_, _029471_);
  or g_120683_(_005748_, _029460_, _029472_);
  and g_120684_(_029471_, _029472_, _029473_);
  not g_120685_(_029473_, _029474_);
  and g_120686_(_029469_, _029473_, _029475_);
  or g_120687_(_029470_, _029474_, _029476_);
  and g_120688_(_029455_, _029475_, _029477_);
  or g_120689_(_029456_, _029476_, _029478_);
  and g_120690_(_029438_, _029477_, _029480_);
  or g_120691_(_029439_, _029478_, _029481_);
  or g_120692_(_005559_, _029385_, _029482_);
  not g_120693_(_029482_, _029483_);
  and g_120694_(_029334_, _029385_, _029484_);
  or g_120695_(_029333_, _029386_, _029485_);
  and g_120696_(_029482_, _029485_, _029486_);
  or g_120697_(_029483_, _029484_, _029487_);
  or g_120698_(_005770_, _029486_, _029488_);
  and g_120699_(_029342_, _029385_, _029489_);
  and g_120700_(_040567_, _029386_, _029491_);
  or g_120701_(_029489_, _029491_, _029492_);
  or g_120702_(_042701_, _029492_, _029493_);
  and g_120703_(_005770_, _029486_, _029494_);
  xor g_120704_(_005770_, _029486_, _029495_);
  xor g_120705_(_005769_, _029486_, _029496_);
  xor g_120706_(_042701_, _029492_, _029497_);
  xor g_120707_(_042690_, _029492_, _029498_);
  and g_120708_(_029495_, _029497_, _029499_);
  or g_120709_(_029496_, _029498_, _029500_);
  or g_120710_(_003673_, _029385_, _029502_);
  or g_120711_(_029351_, _029386_, _029503_);
  and g_120712_(_029502_, _029503_, _029504_);
  and g_120713_(out[177], _029504_, _029505_);
  not g_120714_(_029505_, _029506_);
  and g_120715_(out[176], _029389_, _029507_);
  not g_120716_(_029507_, _029508_);
  xor g_120717_(out[177], _029504_, _029509_);
  xor g_120718_(_003805_, _029504_, _029510_);
  and g_120719_(_029508_, _029509_, _029511_);
  or g_120720_(_029507_, _029510_, _029513_);
  and g_120721_(_029506_, _029513_, _029514_);
  or g_120722_(_029500_, _029514_, _029515_);
  or g_120723_(_029493_, _029494_, _029516_);
  and g_120724_(_029488_, _029516_, _029517_);
  and g_120725_(_029515_, _029517_, _029518_);
  or g_120726_(_029481_, _029518_, _029519_);
  and g_120727_(_029455_, _029470_, _029520_);
  and g_120728_(_029471_, _029520_, _029521_);
  and g_120729_(_029444_, _029452_, _029522_);
  or g_120730_(_029451_, _029522_, _029524_);
  or g_120731_(_029521_, _029524_, _029525_);
  and g_120732_(_029438_, _029525_, _029526_);
  not g_120733_(_029526_, _029527_);
  or g_120734_(_029409_, _029412_, _029528_);
  and g_120735_(_029430_, _029431_, _029529_);
  not g_120736_(_029529_, _029530_);
  or g_120737_(_029417_, _029530_, _029531_);
  and g_120738_(_029528_, _029531_, _029532_);
  and g_120739_(_029519_, _029532_, _029533_);
  and g_120740_(_029527_, _029533_, _029535_);
  or g_120741_(out[176], _029389_, _029536_);
  and g_120742_(_029499_, _029536_, _029537_);
  and g_120743_(_029511_, _029537_, _029538_);
  and g_120744_(_029480_, _029538_, _029539_);
  or g_120745_(_029535_, _029539_, _029540_);
  not g_120746_(_029540_, _029541_);
  and g_120747_(_029389_, _029540_, _029542_);
  and g_120748_(_003816_, _029541_, _029543_);
  or g_120749_(_029542_, _029543_, _029544_);
  and g_120750_(_029390_, _029394_, _029546_);
  or g_120751_(_029392_, _029395_, _029547_);
  or g_120752_(out[202], _005898_, _029548_);
  xor g_120753_(out[203], _029548_, _029549_);
  xor g_120754_(_003882_, _029548_, _029550_);
  and g_120755_(_029546_, _029550_, _029551_);
  or g_120756_(_029547_, _029549_, _029552_);
  or g_120757_(_029406_, _029540_, _029553_);
  not g_120758_(_029553_, _029554_);
  and g_120759_(_029404_, _029540_, _029555_);
  not g_120760_(_029555_, _029557_);
  and g_120761_(_029553_, _029557_, _029558_);
  or g_120762_(_029554_, _029555_, _029559_);
  xor g_120763_(out[202], _005898_, _029560_);
  not g_120764_(_029560_, _029561_);
  and g_120765_(_029558_, _029560_, _029562_);
  or g_120766_(_029559_, _029561_, _029563_);
  and g_120767_(_029552_, _029563_, _029564_);
  or g_120768_(_029551_, _029562_, _029565_);
  and g_120769_(_029559_, _029561_, _029566_);
  and g_120770_(_029547_, _029549_, _029568_);
  or g_120771_(_029566_, _029568_, _029569_);
  or g_120772_(_029565_, _029569_, _029570_);
  or g_120773_(_005663_, _029540_, _029571_);
  not g_120774_(_029571_, _029572_);
  and g_120775_(_029420_, _029540_, _029573_);
  not g_120776_(_029573_, _029574_);
  and g_120777_(_029571_, _029574_, _029575_);
  or g_120778_(_029572_, _029573_, _029576_);
  or g_120779_(_005887_, _029575_, _029577_);
  or g_120780_(_005676_, _029540_, _029579_);
  not g_120781_(_029579_, _029580_);
  and g_120782_(_029426_, _029540_, _029581_);
  not g_120783_(_029581_, _029582_);
  and g_120784_(_029579_, _029582_, _029583_);
  or g_120785_(_029580_, _029581_, _029584_);
  or g_120786_(_005899_, _029583_, _029585_);
  and g_120787_(_029577_, _029585_, _029586_);
  not g_120788_(_029586_, _029587_);
  and g_120789_(_005899_, _029583_, _029588_);
  and g_120790_(_005887_, _029575_, _029590_);
  or g_120791_(_029588_, _029590_, _029591_);
  or g_120792_(_029587_, _029591_, _029592_);
  or g_120793_(_029570_, _029592_, _029593_);
  or g_120794_(_005714_, _029540_, _029594_);
  not g_120795_(_029594_, _029595_);
  and g_120796_(_029442_, _029540_, _029596_);
  not g_120797_(_029596_, _029597_);
  and g_120798_(_029594_, _029597_, _029598_);
  or g_120799_(_029595_, _029596_, _029599_);
  or g_120800_(_005934_, _029599_, _029601_);
  xor g_120801_(_005934_, _029598_, _029602_);
  or g_120802_(_005699_, _029540_, _029603_);
  not g_120803_(_029603_, _029604_);
  and g_120804_(_029450_, _029540_, _029605_);
  not g_120805_(_029605_, _029606_);
  and g_120806_(_029603_, _029606_, _029607_);
  or g_120807_(_029604_, _029605_, _029608_);
  or g_120808_(_005924_, _029607_, _029609_);
  and g_120809_(_005924_, _029607_, _029610_);
  xor g_120810_(_005923_, _029607_, _029612_);
  or g_120811_(_029602_, _029612_, _029613_);
  or g_120812_(_005748_, _029540_, _029614_);
  not g_120813_(_029614_, _029615_);
  and g_120814_(_029460_, _029540_, _029616_);
  not g_120815_(_029616_, _029617_);
  and g_120816_(_029614_, _029617_, _029618_);
  or g_120817_(_029615_, _029616_, _029619_);
  or g_120818_(_005954_, _029618_, _029620_);
  or g_120819_(_005726_, _029540_, _029621_);
  not g_120820_(_029621_, _029623_);
  and g_120821_(_029465_, _029540_, _029624_);
  not g_120822_(_029624_, _029625_);
  and g_120823_(_029621_, _029625_, _029626_);
  or g_120824_(_029623_, _029624_, _029627_);
  or g_120825_(_005965_, _029626_, _029628_);
  and g_120826_(_029620_, _029628_, _029629_);
  not g_120827_(_029629_, _029630_);
  and g_120828_(_005965_, _029626_, _029631_);
  and g_120829_(_005954_, _029618_, _029632_);
  or g_120830_(_029631_, _029632_, _029634_);
  or g_120831_(_029630_, _029634_, _029635_);
  or g_120832_(_029613_, _029635_, _029636_);
  or g_120833_(_029593_, _029636_, _029637_);
  or g_120834_(_005769_, _029540_, _029638_);
  not g_120835_(_029638_, _029639_);
  and g_120836_(_029487_, _029540_, _029640_);
  or g_120837_(_029486_, _029541_, _029641_);
  and g_120838_(_029638_, _029641_, _029642_);
  or g_120839_(_029639_, _029640_, _029643_);
  or g_120840_(_005986_, _029642_, _029645_);
  and g_120841_(_029492_, _029540_, _029646_);
  and g_120842_(_042690_, _029541_, _029647_);
  or g_120843_(_029646_, _029647_, _029648_);
  or g_120844_(_044538_, _029648_, _029649_);
  and g_120845_(_005986_, _029642_, _029650_);
  xor g_120846_(_005985_, _029642_, _029651_);
  xor g_120847_(_044527_, _029648_, _029652_);
  or g_120848_(_029651_, _029652_, _029653_);
  or g_120849_(_003805_, _029540_, _029654_);
  or g_120850_(_029504_, _029541_, _029656_);
  and g_120851_(_029654_, _029656_, _029657_);
  and g_120852_(out[193], _029657_, _029658_);
  not g_120853_(_029658_, _029659_);
  and g_120854_(out[192], _029544_, _029660_);
  xor g_120855_(_003937_, _029657_, _029661_);
  or g_120856_(_029660_, _029661_, _029662_);
  and g_120857_(_029659_, _029662_, _029663_);
  or g_120858_(_029653_, _029663_, _029664_);
  or g_120859_(_029649_, _029650_, _029665_);
  and g_120860_(_029645_, _029665_, _029667_);
  and g_120861_(_029664_, _029667_, _029668_);
  or g_120862_(_029637_, _029668_, _029669_);
  or g_120863_(_029613_, _029629_, _029670_);
  or g_120864_(_029631_, _029670_, _029671_);
  or g_120865_(_029601_, _029610_, _029672_);
  and g_120866_(_029609_, _029672_, _029673_);
  and g_120867_(_029671_, _029673_, _029674_);
  or g_120868_(_029593_, _029674_, _029675_);
  or g_120869_(_029564_, _029568_, _029676_);
  or g_120870_(_029586_, _029588_, _029678_);
  or g_120871_(_029570_, _029678_, _029679_);
  and g_120872_(_029676_, _029679_, _029680_);
  and g_120873_(_029675_, _029680_, _029681_);
  and g_120874_(_029669_, _029681_, _029682_);
  or g_120875_(out[192], _029544_, _029683_);
  or g_120876_(_029653_, _029662_, _029684_);
  or g_120877_(_029637_, _029684_, _029685_);
  not g_120878_(_029685_, _029686_);
  and g_120879_(_029683_, _029686_, _029687_);
  or g_120880_(_029682_, _029687_, _029689_);
  not g_120881_(_029689_, _029690_);
  and g_120882_(_029544_, _029689_, _029691_);
  not g_120883_(_029691_, _029692_);
  or g_120884_(out[192], _029689_, _029693_);
  not g_120885_(_029693_, _029694_);
  and g_120886_(_029692_, _029693_, _029695_);
  or g_120887_(_029691_, _029694_, _029696_);
  and g_120888_(_029560_, _029690_, _029697_);
  or g_120889_(_029561_, _029689_, _029698_);
  and g_120890_(_029559_, _029689_, _029700_);
  or g_120891_(_029558_, _029690_, _029701_);
  and g_120892_(_029698_, _029701_, _029702_);
  or g_120893_(_029697_, _029700_, _029703_);
  or g_120894_(out[218], _006110_, _029704_);
  xor g_120895_(out[218], _006110_, _029705_);
  not g_120896_(_029705_, _029706_);
  and g_120897_(_029702_, _029705_, _029707_);
  and g_120898_(_029546_, _029549_, _029708_);
  or g_120899_(_029547_, _029550_, _029709_);
  xor g_120900_(out[219], _029704_, _029711_);
  xor g_120901_(_003992_, _029704_, _029712_);
  and g_120902_(_029708_, _029712_, _029713_);
  or g_120903_(_029708_, _029712_, _029714_);
  xor g_120904_(_029709_, _029711_, _029715_);
  xor g_120905_(_029708_, _029711_, _029716_);
  xor g_120906_(_029702_, _029705_, _029717_);
  xor g_120907_(_029703_, _029705_, _029718_);
  and g_120908_(_029715_, _029717_, _029719_);
  or g_120909_(_029716_, _029718_, _029720_);
  and g_120910_(_005887_, _029690_, _029722_);
  and g_120911_(_029576_, _029689_, _029723_);
  or g_120912_(_029722_, _029723_, _029724_);
  and g_120913_(_006129_, _029724_, _029725_);
  not g_120914_(_029725_, _029726_);
  and g_120915_(_005899_, _029690_, _029727_);
  and g_120916_(_029584_, _029689_, _029728_);
  or g_120917_(_029727_, _029728_, _029729_);
  and g_120918_(_006112_, _029729_, _029730_);
  not g_120919_(_029730_, _029731_);
  and g_120920_(_029726_, _029731_, _029733_);
  or g_120921_(_029725_, _029730_, _029734_);
  or g_120922_(_006112_, _029729_, _029735_);
  and g_120923_(_029719_, _029734_, _029736_);
  and g_120924_(_029735_, _029736_, _029737_);
  and g_120925_(_029707_, _029714_, _029738_);
  or g_120926_(_029713_, _029738_, _029739_);
  or g_120927_(_029737_, _029739_, _029740_);
  or g_120928_(_006129_, _029724_, _029741_);
  and g_120929_(_029735_, _029741_, _029742_);
  not g_120930_(_029742_, _029744_);
  and g_120931_(_029733_, _029742_, _029745_);
  or g_120932_(_029734_, _029744_, _029746_);
  and g_120933_(_029719_, _029745_, _029747_);
  or g_120934_(_029720_, _029746_, _029748_);
  and g_120935_(_005924_, _029690_, _029749_);
  and g_120936_(_029608_, _029689_, _029750_);
  or g_120937_(_029749_, _029750_, _029751_);
  or g_120938_(_006146_, _029751_, _029752_);
  or g_120939_(_005934_, _029689_, _029753_);
  or g_120940_(_029598_, _029690_, _029755_);
  and g_120941_(_029753_, _029755_, _029756_);
  not g_120942_(_029756_, _029757_);
  and g_120943_(_006157_, _029756_, _029758_);
  and g_120944_(_006146_, _029751_, _029759_);
  or g_120945_(_029758_, _029759_, _029760_);
  and g_120946_(_029752_, _029760_, _029761_);
  and g_120947_(_029747_, _029761_, _029762_);
  or g_120948_(_029740_, _029762_, _029763_);
  not g_120949_(_029763_, _029764_);
  and g_120950_(_005965_, _029690_, _029766_);
  and g_120951_(_029627_, _029689_, _029767_);
  or g_120952_(_029766_, _029767_, _029768_);
  or g_120953_(_006180_, _029768_, _029769_);
  xor g_120954_(_006157_, _029756_, _029770_);
  xor g_120955_(_006146_, _029751_, _029771_);
  and g_120956_(_029770_, _029771_, _029772_);
  and g_120957_(_029769_, _029772_, _029773_);
  not g_120958_(_029773_, _029774_);
  and g_120959_(_029747_, _029773_, _029775_);
  or g_120960_(_029748_, _029774_, _029777_);
  and g_120961_(_005954_, _029690_, _029778_);
  and g_120962_(_029619_, _029689_, _029779_);
  or g_120963_(_029778_, _029779_, _029780_);
  and g_120964_(_006173_, _029780_, _029781_);
  and g_120965_(_006180_, _029768_, _029782_);
  or g_120966_(_029781_, _029782_, _029783_);
  not g_120967_(_029783_, _029784_);
  or g_120968_(_005985_, _029689_, _029785_);
  not g_120969_(_029785_, _029786_);
  and g_120970_(_029643_, _029689_, _029788_);
  or g_120971_(_029642_, _029690_, _029789_);
  and g_120972_(_029785_, _029789_, _029790_);
  or g_120973_(_029786_, _029788_, _029791_);
  or g_120974_(_006224_, _029791_, _029792_);
  or g_120975_(_006173_, _029780_, _029793_);
  and g_120976_(_029792_, _029793_, _029794_);
  not g_120977_(_029794_, _029795_);
  and g_120978_(_006224_, _029791_, _029796_);
  or g_120979_(_006226_, _029790_, _029797_);
  and g_120980_(_029648_, _029689_, _029799_);
  and g_120981_(_044527_, _029690_, _029800_);
  or g_120982_(_029799_, _029800_, _029801_);
  not g_120983_(_029801_, _029802_);
  and g_120984_(_046881_, _029802_, _029803_);
  or g_120985_(_046892_, _029801_, _029804_);
  and g_120986_(_029797_, _029804_, _029805_);
  or g_120987_(_029796_, _029803_, _029806_);
  and g_120988_(_046892_, _029801_, _029807_);
  or g_120989_(_046881_, _029802_, _029808_);
  and g_120990_(_029657_, _029689_, _029810_);
  not g_120991_(_029810_, _029811_);
  or g_120992_(out[193], _029689_, _029812_);
  not g_120993_(_029812_, _029813_);
  or g_120994_(_029810_, _029813_, _029814_);
  and g_120995_(_029811_, _029812_, _029815_);
  and g_120996_(out[209], _029814_, _029816_);
  or g_120997_(_004047_, _029815_, _029817_);
  or g_120998_(out[208], _029696_, _029818_);
  not g_120999_(_029818_, _029819_);
  and g_121000_(out[208], _029696_, _029821_);
  or g_121001_(_004058_, _029695_, _029822_);
  and g_121002_(_004047_, _029815_, _029823_);
  or g_121003_(out[209], _029814_, _029824_);
  and g_121004_(_029822_, _029824_, _029825_);
  or g_121005_(_029821_, _029823_, _029826_);
  and g_121006_(_029819_, _029825_, _029827_);
  or g_121007_(_029818_, _029826_, _029828_);
  and g_121008_(_029817_, _029828_, _029829_);
  or g_121009_(_029816_, _029827_, _029830_);
  and g_121010_(_029808_, _029830_, _029832_);
  or g_121011_(_029807_, _029829_, _029833_);
  and g_121012_(_029805_, _029833_, _029834_);
  or g_121013_(_029806_, _029832_, _029835_);
  and g_121014_(_029794_, _029835_, _029836_);
  or g_121015_(_029795_, _029834_, _029837_);
  and g_121016_(_029784_, _029837_, _029838_);
  or g_121017_(_029783_, _029836_, _029839_);
  and g_121018_(_029775_, _029839_, _029840_);
  or g_121019_(_029777_, _029838_, _029841_);
  and g_121020_(_029764_, _029841_, _029843_);
  or g_121021_(_029763_, _029840_, _029844_);
  and g_121022_(_029696_, _029843_, _029845_);
  and g_121023_(_004058_, _029844_, _029846_);
  or g_121024_(_029845_, _029846_, _029847_);
  and g_121025_(_029708_, _029711_, _029848_);
  or g_121026_(_029709_, _029712_, _029849_);
  or g_121027_(out[234], _006344_, _029850_);
  xor g_121028_(out[235], _029850_, _029851_);
  xor g_121029_(_004124_, _029850_, _029852_);
  and g_121030_(_029848_, _029852_, _029854_);
  or g_121031_(_029849_, _029851_, _029855_);
  or g_121032_(_029706_, _029843_, _029856_);
  not g_121033_(_029856_, _029857_);
  and g_121034_(_029703_, _029843_, _029858_);
  or g_121035_(_029702_, _029844_, _029859_);
  and g_121036_(_029856_, _029859_, _029860_);
  or g_121037_(_029857_, _029858_, _029861_);
  xor g_121038_(out[234], _006344_, _029862_);
  xor g_121039_(_004234_, _006344_, _029863_);
  and g_121040_(_029860_, _029862_, _029865_);
  or g_121041_(_029861_, _029863_, _029866_);
  and g_121042_(_029855_, _029866_, _029867_);
  or g_121043_(_029854_, _029865_, _029868_);
  and g_121044_(_029849_, _029851_, _029869_);
  and g_121045_(_029861_, _029863_, _029870_);
  or g_121046_(_029869_, _029870_, _029871_);
  not g_121047_(_029871_, _029872_);
  and g_121048_(_029867_, _029872_, _029873_);
  or g_121049_(_029868_, _029871_, _029874_);
  or g_121050_(_006129_, _029843_, _029876_);
  not g_121051_(_029876_, _029877_);
  and g_121052_(_029724_, _029843_, _029878_);
  not g_121053_(_029878_, _029879_);
  and g_121054_(_029876_, _029879_, _029880_);
  or g_121055_(_029877_, _029878_, _029881_);
  and g_121056_(_006369_, _029881_, _029882_);
  not g_121057_(_029882_, _029883_);
  or g_121058_(_006112_, _029843_, _029884_);
  not g_121059_(_029884_, _029885_);
  and g_121060_(_029729_, _029843_, _029887_);
  not g_121061_(_029887_, _029888_);
  and g_121062_(_029884_, _029888_, _029889_);
  or g_121063_(_029885_, _029887_, _029890_);
  and g_121064_(_006347_, _029890_, _029891_);
  not g_121065_(_029891_, _029892_);
  and g_121066_(_029883_, _029892_, _029893_);
  or g_121067_(_029882_, _029891_, _029894_);
  and g_121068_(_006367_, _029880_, _029895_);
  or g_121069_(_006369_, _029881_, _029896_);
  and g_121070_(_006345_, _029889_, _029898_);
  or g_121071_(_006347_, _029890_, _029899_);
  and g_121072_(_029896_, _029899_, _029900_);
  or g_121073_(_029895_, _029898_, _029901_);
  and g_121074_(_029893_, _029900_, _029902_);
  or g_121075_(_029894_, _029901_, _029903_);
  and g_121076_(_029873_, _029902_, _029904_);
  or g_121077_(_029874_, _029903_, _029905_);
  and g_121078_(_006147_, _029844_, _029906_);
  and g_121079_(_029751_, _029843_, _029907_);
  or g_121080_(_029906_, _029907_, _029909_);
  and g_121081_(_006389_, _029909_, _029910_);
  and g_121082_(_006157_, _029844_, _029911_);
  and g_121083_(_029757_, _029843_, _029912_);
  or g_121084_(_029911_, _029912_, _029913_);
  or g_121085_(_006405_, _029913_, _029914_);
  not g_121086_(_029914_, _029915_);
  or g_121087_(_006389_, _029909_, _029916_);
  xor g_121088_(_006405_, _029913_, _029917_);
  xor g_121089_(_006406_, _029913_, _029918_);
  xor g_121090_(_006389_, _029909_, _029920_);
  xor g_121091_(_006391_, _029909_, _029921_);
  and g_121092_(_029917_, _029920_, _029922_);
  or g_121093_(_029918_, _029921_, _029923_);
  or g_121094_(_006180_, _029843_, _029924_);
  not g_121095_(_029924_, _029925_);
  and g_121096_(_029768_, _029843_, _029926_);
  not g_121097_(_029926_, _029927_);
  and g_121098_(_029924_, _029927_, _029928_);
  or g_121099_(_029925_, _029926_, _029929_);
  or g_121100_(_006433_, _029928_, _029931_);
  or g_121101_(_006173_, _029843_, _029932_);
  not g_121102_(_029932_, _029933_);
  and g_121103_(_029780_, _029843_, _029934_);
  not g_121104_(_029934_, _029935_);
  and g_121105_(_029932_, _029935_, _029936_);
  or g_121106_(_029933_, _029934_, _029937_);
  or g_121107_(_006422_, _029936_, _029938_);
  and g_121108_(_029931_, _029938_, _029939_);
  or g_121109_(_006435_, _029929_, _029940_);
  not g_121110_(_029940_, _029942_);
  or g_121111_(_006424_, _029937_, _029943_);
  and g_121112_(_029940_, _029943_, _029944_);
  xor g_121113_(_006435_, _029928_, _029945_);
  xor g_121114_(_006424_, _029936_, _029946_);
  and g_121115_(_029939_, _029944_, _029947_);
  or g_121116_(_029945_, _029946_, _029948_);
  and g_121117_(_029922_, _029947_, _029949_);
  or g_121118_(_029923_, _029948_, _029950_);
  and g_121119_(_029904_, _029949_, _029951_);
  or g_121120_(_029905_, _029950_, _029953_);
  and g_121121_(_006226_, _029844_, _029954_);
  and g_121122_(_029791_, _029843_, _029955_);
  or g_121123_(_029954_, _029955_, _029956_);
  and g_121124_(_006292_, _029956_, _029957_);
  or g_121125_(_046892_, _029843_, _029958_);
  not g_121126_(_029958_, _029959_);
  and g_121127_(_029801_, _029843_, _029960_);
  not g_121128_(_029960_, _029961_);
  and g_121129_(_029958_, _029961_, _029962_);
  or g_121130_(_029959_, _029960_, _029964_);
  or g_121131_(_006292_, _029956_, _029965_);
  and g_121132_(_047816_, _029962_, _029966_);
  xor g_121133_(_006292_, _029956_, _029967_);
  xor g_121134_(_006293_, _029956_, _029968_);
  xor g_121135_(_047816_, _029962_, _029969_);
  xor g_121136_(_047827_, _029962_, _029970_);
  and g_121137_(_029967_, _029969_, _029971_);
  or g_121138_(_029968_, _029970_, _029972_);
  or g_121139_(_029814_, _029844_, _029973_);
  or g_121140_(_004047_, _029843_, _029975_);
  and g_121141_(_029973_, _029975_, _029976_);
  and g_121142_(out[225], _029976_, _029977_);
  not g_121143_(_029977_, _029978_);
  and g_121144_(out[224], _029847_, _029979_);
  not g_121145_(_029979_, _029980_);
  xor g_121146_(out[225], _029976_, _029981_);
  xor g_121147_(_004179_, _029976_, _029982_);
  and g_121148_(_029980_, _029981_, _029983_);
  or g_121149_(_029979_, _029982_, _029984_);
  and g_121150_(_029978_, _029984_, _029986_);
  or g_121151_(_029972_, _029986_, _029987_);
  and g_121152_(_029965_, _029966_, _029988_);
  or g_121153_(_029957_, _029988_, _029989_);
  not g_121154_(_029989_, _029990_);
  and g_121155_(_029987_, _029990_, _029991_);
  or g_121156_(_029953_, _029991_, _029992_);
  or g_121157_(_029939_, _029942_, _029993_);
  or g_121158_(_029923_, _029993_, _029994_);
  and g_121159_(_029915_, _029916_, _029995_);
  or g_121160_(_029910_, _029995_, _029997_);
  not g_121161_(_029997_, _029998_);
  and g_121162_(_029994_, _029998_, _029999_);
  or g_121163_(_029905_, _029999_, _030000_);
  or g_121164_(_029867_, _029869_, _030001_);
  or g_121165_(_029874_, _029893_, _030002_);
  or g_121166_(_029898_, _030002_, _030003_);
  and g_121167_(_030001_, _030003_, _030004_);
  and g_121168_(_029992_, _030004_, _030005_);
  and g_121169_(_030000_, _030005_, _030006_);
  or g_121170_(out[224], _029847_, _030008_);
  and g_121171_(_029971_, _030008_, _030009_);
  and g_121172_(_029983_, _030009_, _030010_);
  and g_121173_(_029951_, _030010_, _030011_);
  or g_121174_(_030006_, _030011_, _030012_);
  and g_121175_(_029847_, _030012_, _030013_);
  not g_121176_(_030013_, _030014_);
  or g_121177_(out[224], _030012_, _030015_);
  not g_121178_(_030015_, _030016_);
  and g_121179_(_030014_, _030015_, _030017_);
  or g_121180_(_030013_, _030016_, _030019_);
  and g_121181_(_029848_, _029851_, _030020_);
  or g_121182_(_029849_, _029852_, _030021_);
  or g_121183_(out[250], _006519_, _030022_);
  xor g_121184_(out[251], _030022_, _030023_);
  xor g_121185_(_004245_, _030022_, _030024_);
  and g_121186_(_030020_, _030024_, _030025_);
  or g_121187_(_030021_, _030023_, _030026_);
  or g_121188_(_029863_, _030012_, _030027_);
  not g_121189_(_030027_, _030028_);
  and g_121190_(_029861_, _030012_, _030030_);
  or g_121191_(_030028_, _030030_, _030031_);
  xor g_121192_(_004355_, _006519_, _030032_);
  or g_121193_(_030031_, _030032_, _030033_);
  not g_121194_(_030033_, _030034_);
  and g_121195_(_030026_, _030033_, _030035_);
  or g_121196_(_030025_, _030034_, _030036_);
  and g_121197_(_030021_, _030023_, _030037_);
  or g_121198_(_030020_, _030024_, _030038_);
  and g_121199_(_030036_, _030038_, _030039_);
  or g_121200_(_030035_, _030037_, _030041_);
  or g_121201_(_006369_, _030012_, _030042_);
  not g_121202_(_030042_, _030043_);
  and g_121203_(_029881_, _030012_, _030044_);
  or g_121204_(_030043_, _030044_, _030045_);
  not g_121205_(_030045_, _030046_);
  and g_121206_(_006530_, _030045_, _030047_);
  or g_121207_(_006529_, _030046_, _030048_);
  or g_121208_(_006347_, _030012_, _030049_);
  not g_121209_(_030049_, _030050_);
  and g_121210_(_029890_, _030012_, _030052_);
  or g_121211_(_030050_, _030052_, _030053_);
  not g_121212_(_030053_, _030054_);
  and g_121213_(_006521_, _030053_, _030055_);
  or g_121214_(_006520_, _030054_, _030056_);
  and g_121215_(_030048_, _030056_, _030057_);
  or g_121216_(_030047_, _030055_, _030058_);
  or g_121217_(_006389_, _030012_, _030059_);
  not g_121218_(_030059_, _030060_);
  and g_121219_(_029909_, _030012_, _030061_);
  not g_121220_(_030061_, _030063_);
  and g_121221_(_030059_, _030063_, _030064_);
  or g_121222_(_030060_, _030061_, _030065_);
  and g_121223_(_006546_, _030065_, _030066_);
  or g_121224_(_006547_, _030064_, _030067_);
  and g_121225_(_006547_, _030064_, _030068_);
  or g_121226_(_006546_, _030065_, _030069_);
  or g_121227_(_006405_, _030012_, _030070_);
  not g_121228_(_030070_, _030071_);
  and g_121229_(_029913_, _030012_, _030072_);
  not g_121230_(_030072_, _030074_);
  and g_121231_(_030070_, _030074_, _030075_);
  or g_121232_(_030071_, _030072_, _030076_);
  and g_121233_(_006554_, _030075_, _030077_);
  or g_121234_(_006553_, _030076_, _030078_);
  and g_121235_(_030069_, _030077_, _030079_);
  or g_121236_(_030068_, _030078_, _030080_);
  and g_121237_(_030067_, _030080_, _030081_);
  or g_121238_(_030066_, _030079_, _030082_);
  and g_121239_(_030067_, _030069_, _030083_);
  or g_121240_(_030066_, _030068_, _030085_);
  or g_121241_(_006435_, _030012_, _030086_);
  not g_121242_(_030086_, _030087_);
  and g_121243_(_029929_, _030012_, _030088_);
  or g_121244_(_030087_, _030088_, _030089_);
  not g_121245_(_030089_, _030090_);
  and g_121246_(_006569_, _030090_, _030091_);
  or g_121247_(_006570_, _030089_, _030092_);
  xor g_121248_(_006554_, _030075_, _030093_);
  xor g_121249_(_006553_, _030075_, _030094_);
  and g_121250_(_030083_, _030093_, _030096_);
  or g_121251_(_030085_, _030094_, _030097_);
  and g_121252_(_030092_, _030096_, _030098_);
  or g_121253_(_030091_, _030097_, _030099_);
  or g_121254_(_006424_, _030012_, _030100_);
  not g_121255_(_030100_, _030101_);
  and g_121256_(_029937_, _030012_, _030102_);
  or g_121257_(_030101_, _030102_, _030103_);
  not g_121258_(_030103_, _030104_);
  and g_121259_(_006584_, _030103_, _030105_);
  or g_121260_(_006583_, _030104_, _030107_);
  and g_121261_(_006570_, _030089_, _030108_);
  or g_121262_(_006569_, _030090_, _030109_);
  and g_121263_(_030107_, _030109_, _030110_);
  or g_121264_(_030105_, _030108_, _030111_);
  or g_121265_(_047827_, _030012_, _030112_);
  not g_121266_(_030112_, _030113_);
  and g_121267_(_029964_, _030012_, _030114_);
  or g_121268_(_030113_, _030114_, _030115_);
  not g_121269_(_030115_, _030116_);
  or g_121270_(_006292_, _030012_, _030118_);
  not g_121271_(_030118_, _030119_);
  and g_121272_(_029956_, _030012_, _030120_);
  not g_121273_(_030120_, _030121_);
  and g_121274_(_030118_, _030121_, _030122_);
  or g_121275_(_030119_, _030120_, _030123_);
  and g_121276_(_006600_, _030123_, _030124_);
  not g_121277_(_030124_, _030125_);
  and g_121278_(_050478_, _030116_, _030126_);
  or g_121279_(_050489_, _030115_, _030127_);
  and g_121280_(_006601_, _030122_, _030129_);
  or g_121281_(_006600_, _030123_, _030130_);
  xor g_121282_(_050489_, _030115_, _030131_);
  xor g_121283_(_050478_, _030115_, _030132_);
  and g_121284_(_030130_, _030131_, _030133_);
  or g_121285_(_030129_, _030132_, _030134_);
  and g_121286_(_030125_, _030133_, _030135_);
  or g_121287_(_030124_, _030134_, _030136_);
  and g_121288_(_029976_, _030012_, _030137_);
  or g_121289_(out[225], _030012_, _030138_);
  not g_121290_(_030138_, _030140_);
  or g_121291_(_030137_, _030140_, _030141_);
  and g_121292_(out[241], _030141_, _030142_);
  not g_121293_(_030142_, _030143_);
  and g_121294_(out[240], _030019_, _030144_);
  or g_121295_(_004300_, _030017_, _030145_);
  xor g_121296_(out[241], _030141_, _030146_);
  xor g_121297_(_053038_, _030141_, _030147_);
  and g_121298_(_030145_, _030146_, _030148_);
  or g_121299_(_030144_, _030147_, _030149_);
  and g_121300_(_030143_, _030149_, _030151_);
  or g_121301_(_030142_, _030148_, _030152_);
  and g_121302_(_030135_, _030152_, _030153_);
  or g_121303_(_030136_, _030151_, _030154_);
  and g_121304_(_030126_, _030130_, _030155_);
  or g_121305_(_030127_, _030129_, _030156_);
  and g_121306_(_030125_, _030156_, _030157_);
  or g_121307_(_030124_, _030155_, _030158_);
  and g_121308_(_030154_, _030157_, _030159_);
  or g_121309_(_030153_, _030158_, _030160_);
  and g_121310_(_006583_, _030104_, _030162_);
  or g_121311_(_006584_, _030103_, _030163_);
  and g_121312_(_030110_, _030163_, _030164_);
  or g_121313_(_030111_, _030162_, _030165_);
  and g_121314_(_030098_, _030164_, _030166_);
  or g_121315_(_030099_, _030165_, _030167_);
  and g_121316_(_030160_, _030166_, _030168_);
  or g_121317_(_030159_, _030167_, _030169_);
  and g_121318_(_030098_, _030111_, _030170_);
  or g_121319_(_030099_, _030110_, _030171_);
  and g_121320_(_030081_, _030171_, _030173_);
  or g_121321_(_030082_, _030170_, _030174_);
  and g_121322_(_030169_, _030173_, _030175_);
  or g_121323_(_030168_, _030174_, _030176_);
  and g_121324_(_006529_, _030046_, _030177_);
  or g_121325_(_006530_, _030045_, _030178_);
  and g_121326_(_030031_, _030032_, _030179_);
  or g_121327_(_030037_, _030179_, _030180_);
  not g_121328_(_030180_, _030181_);
  and g_121329_(_030035_, _030181_, _030182_);
  or g_121330_(_030036_, _030180_, _030184_);
  and g_121331_(_006520_, _030054_, _030185_);
  or g_121332_(_006521_, _030053_, _030186_);
  and g_121333_(_030058_, _030186_, _030187_);
  or g_121334_(_030057_, _030185_, _030188_);
  and g_121335_(_030182_, _030187_, _030189_);
  or g_121336_(_030184_, _030188_, _030190_);
  and g_121337_(_030178_, _030186_, _030191_);
  or g_121338_(_030177_, _030185_, _030192_);
  and g_121339_(_030057_, _030191_, _030193_);
  or g_121340_(_030058_, _030192_, _030195_);
  and g_121341_(_030182_, _030193_, _030196_);
  or g_121342_(_030184_, _030195_, _030197_);
  and g_121343_(_030176_, _030196_, _030198_);
  or g_121344_(_030175_, _030197_, _030199_);
  and g_121345_(_030041_, _030190_, _030200_);
  or g_121346_(_030039_, _030189_, _030201_);
  and g_121347_(_030199_, _030200_, _030202_);
  or g_121348_(_030198_, _030201_, _030203_);
  or g_121349_(out[240], _030019_, _030204_);
  not g_121350_(_030204_, _030206_);
  or g_121351_(_030149_, _030206_, _030207_);
  not g_121352_(_030207_, _030208_);
  and g_121353_(_030135_, _030208_, _030209_);
  or g_121354_(_030136_, _030207_, _030210_);
  and g_121355_(_030196_, _030209_, _030211_);
  or g_121356_(_030197_, _030210_, _030212_);
  and g_121357_(_030166_, _030211_, _030213_);
  or g_121358_(_030167_, _030212_, _030214_);
  and g_121359_(_030203_, _030214_, _030215_);
  or g_121360_(_030202_, _030213_, _030217_);
  and g_121361_(_030019_, _030217_, _030218_);
  and g_121362_(_004300_, _030215_, _030219_);
  or g_121363_(_030218_, _030219_, _030220_);
  and g_121364_(_030020_, _030023_, _030221_);
  or g_121365_(_030021_, _030024_, _030222_);
  or g_121366_(out[266], _006780_, _030223_);
  xor g_121367_(out[267], _030223_, _030224_);
  xor g_121368_(_004366_, _030223_, _030225_);
  and g_121369_(_030221_, _030225_, _030226_);
  or g_121370_(_030222_, _030224_, _030228_);
  and g_121371_(_030031_, _030217_, _030229_);
  not g_121372_(_030229_, _030230_);
  or g_121373_(_030032_, _030217_, _030231_);
  not g_121374_(_030231_, _030232_);
  and g_121375_(_030230_, _030231_, _030233_);
  or g_121376_(_030229_, _030232_, _030234_);
  xor g_121377_(out[266], _006780_, _030235_);
  xor g_121378_(_004421_, _006780_, _030236_);
  and g_121379_(_030233_, _030235_, _030237_);
  or g_121380_(_030234_, _030236_, _030239_);
  and g_121381_(_030228_, _030239_, _030240_);
  or g_121382_(_030226_, _030237_, _030241_);
  and g_121383_(_030234_, _030236_, _030242_);
  and g_121384_(_030222_, _030224_, _030243_);
  or g_121385_(_030242_, _030243_, _030244_);
  not g_121386_(_030244_, _030245_);
  and g_121387_(_030240_, _030245_, _030246_);
  or g_121388_(_030241_, _030244_, _030247_);
  and g_121389_(_006529_, _030215_, _030248_);
  and g_121390_(_030045_, _030217_, _030250_);
  or g_121391_(_030248_, _030250_, _030251_);
  not g_121392_(_030251_, _030252_);
  and g_121393_(_006771_, _030251_, _030253_);
  or g_121394_(_006770_, _030252_, _030254_);
  and g_121395_(_006520_, _030215_, _030255_);
  and g_121396_(_030053_, _030217_, _030256_);
  or g_121397_(_030255_, _030256_, _030257_);
  not g_121398_(_030257_, _030258_);
  and g_121399_(_006782_, _030257_, _030259_);
  or g_121400_(_006781_, _030258_, _030261_);
  and g_121401_(_030254_, _030261_, _030262_);
  or g_121402_(_030253_, _030259_, _030263_);
  or g_121403_(_006782_, _030257_, _030264_);
  or g_121404_(_006771_, _030251_, _030265_);
  and g_121405_(_030264_, _030265_, _030266_);
  not g_121406_(_030266_, _030267_);
  and g_121407_(_030262_, _030266_, _030268_);
  or g_121408_(_030263_, _030267_, _030269_);
  and g_121409_(_030246_, _030268_, _030270_);
  or g_121410_(_030247_, _030269_, _030272_);
  and g_121411_(_030076_, _030217_, _030273_);
  and g_121412_(_006554_, _030215_, _030274_);
  or g_121413_(_030273_, _030274_, _030275_);
  or g_121414_(_006803_, _030275_, _030276_);
  not g_121415_(_030276_, _030277_);
  and g_121416_(_006547_, _030215_, _030278_);
  or g_121417_(_006546_, _030217_, _030279_);
  and g_121418_(_030065_, _030217_, _030280_);
  or g_121419_(_030064_, _030215_, _030281_);
  and g_121420_(_030279_, _030281_, _030283_);
  or g_121421_(_030278_, _030280_, _030284_);
  and g_121422_(_006812_, _030284_, _030285_);
  or g_121423_(_006813_, _030283_, _030286_);
  and g_121424_(_030276_, _030286_, _030287_);
  or g_121425_(_030277_, _030285_, _030288_);
  and g_121426_(_006803_, _030275_, _030289_);
  or g_121427_(_006570_, _030217_, _030290_);
  not g_121428_(_030290_, _030291_);
  and g_121429_(_030089_, _030217_, _030292_);
  not g_121430_(_030292_, _030294_);
  and g_121431_(_030290_, _030294_, _030295_);
  or g_121432_(_030291_, _030292_, _030296_);
  and g_121433_(_006832_, _030295_, _030297_);
  or g_121434_(_006833_, _030296_, _030298_);
  or g_121435_(_030289_, _030297_, _030299_);
  or g_121436_(_030288_, _030299_, _030300_);
  or g_121437_(_006584_, _030217_, _030301_);
  not g_121438_(_030301_, _030302_);
  and g_121439_(_030103_, _030217_, _030303_);
  not g_121440_(_030303_, _030305_);
  and g_121441_(_030301_, _030305_, _030306_);
  or g_121442_(_030302_, _030303_, _030307_);
  and g_121443_(_006825_, _030307_, _030308_);
  or g_121444_(_006824_, _030306_, _030309_);
  and g_121445_(_006833_, _030296_, _030310_);
  or g_121446_(_006832_, _030295_, _030311_);
  and g_121447_(_030309_, _030311_, _030312_);
  or g_121448_(_030308_, _030310_, _030313_);
  and g_121449_(_006813_, _030283_, _030314_);
  or g_121450_(_006812_, _030284_, _030316_);
  or g_121451_(_006825_, _030307_, _030317_);
  xor g_121452_(_006803_, _030275_, _030318_);
  and g_121453_(_030286_, _030316_, _030319_);
  and g_121454_(_030318_, _030319_, _030320_);
  and g_121455_(_030312_, _030317_, _030321_);
  and g_121456_(_030298_, _030320_, _030322_);
  and g_121457_(_030270_, _030322_, _030323_);
  and g_121458_(_030321_, _030323_, _030324_);
  or g_121459_(out[256], _030220_, _030325_);
  and g_121460_(_030123_, _030217_, _030327_);
  and g_121461_(_006601_, _030215_, _030328_);
  or g_121462_(_030327_, _030328_, _030329_);
  or g_121463_(_006716_, _030329_, _030330_);
  and g_121464_(_030115_, _030217_, _030331_);
  and g_121465_(_050478_, _030215_, _030332_);
  or g_121466_(_030331_, _030332_, _030333_);
  and g_121467_(_006716_, _030329_, _030334_);
  or g_121468_(_051427_, _030333_, _030335_);
  not g_121469_(_030335_, _030336_);
  or g_121470_(_030334_, _030336_, _030338_);
  xor g_121471_(_006716_, _030329_, _030339_);
  xor g_121472_(_051427_, _030333_, _030340_);
  and g_121473_(_030339_, _030340_, _030341_);
  or g_121474_(_053038_, _030217_, _030342_);
  or g_121475_(_030141_, _030215_, _030343_);
  and g_121476_(_030342_, _030343_, _030344_);
  and g_121477_(out[256], _030220_, _030345_);
  not g_121478_(_030345_, _030346_);
  and g_121479_(out[257], _030344_, _030347_);
  xor g_121480_(out[257], _030344_, _030349_);
  and g_121481_(_030346_, _030349_, _030350_);
  and g_121482_(_030341_, _030350_, _030351_);
  and g_121483_(_030325_, _030351_, _030352_);
  and g_121484_(_030324_, _030352_, _030353_);
  not g_121485_(_030353_, _030354_);
  and g_121486_(_030330_, _030338_, _030355_);
  or g_121487_(_030347_, _030350_, _030356_);
  and g_121488_(_030341_, _030356_, _030357_);
  or g_121489_(_030355_, _030357_, _030358_);
  and g_121490_(_030324_, _030358_, _030360_);
  not g_121491_(_030360_, _030361_);
  or g_121492_(_030240_, _030243_, _030362_);
  not g_121493_(_030362_, _030363_);
  and g_121494_(_030263_, _030264_, _030364_);
  not g_121495_(_030364_, _030365_);
  and g_121496_(_030246_, _030364_, _030366_);
  or g_121497_(_030247_, _030365_, _030367_);
  and g_121498_(_030362_, _030367_, _030368_);
  or g_121499_(_030363_, _030366_, _030369_);
  or g_121500_(_030300_, _030312_, _030371_);
  and g_121501_(_030287_, _030371_, _030372_);
  or g_121502_(_030272_, _030314_, _030373_);
  and g_121503_(_030313_, _030322_, _030374_);
  and g_121504_(_030277_, _030316_, _030375_);
  or g_121505_(_030374_, _030375_, _030376_);
  or g_121506_(_030285_, _030376_, _030377_);
  and g_121507_(_030270_, _030377_, _030378_);
  or g_121508_(_030372_, _030373_, _030379_);
  and g_121509_(_030368_, _030379_, _030380_);
  or g_121510_(_030369_, _030378_, _030382_);
  and g_121511_(_030361_, _030380_, _030383_);
  or g_121512_(_030360_, _030382_, _030384_);
  and g_121513_(_030354_, _030384_, _030385_);
  or g_121514_(_030353_, _030383_, _030386_);
  and g_121515_(_030220_, _030386_, _030387_);
  and g_121516_(_004388_, _030385_, _030388_);
  or g_121517_(_030387_, _030388_, _030389_);
  or g_121518_(out[272], _030389_, _030390_);
  not g_121519_(_030390_, _030391_);
  or g_121520_(_053027_, _030386_, _030393_);
  or g_121521_(_030344_, _030385_, _030394_);
  and g_121522_(_030393_, _030394_, _030395_);
  and g_121523_(out[272], _030389_, _030396_);
  not g_121524_(_030396_, _030397_);
  and g_121525_(out[273], _030395_, _030398_);
  not g_121526_(_030398_, _030399_);
  xor g_121527_(out[273], _030395_, _030400_);
  xor g_121528_(_053126_, _030395_, _030401_);
  and g_121529_(_030397_, _030400_, _030402_);
  or g_121530_(_030396_, _030401_, _030404_);
  and g_121531_(_030221_, _030224_, _030405_);
  or g_121532_(_030222_, _030225_, _030406_);
  or g_121533_(out[282], _006904_, _030407_);
  xor g_121534_(out[283], _030407_, _030408_);
  not g_121535_(_030408_, _030409_);
  or g_121536_(_030406_, _030408_, _030410_);
  and g_121537_(_030235_, _030385_, _030411_);
  and g_121538_(_030234_, _030386_, _030412_);
  or g_121539_(_030411_, _030412_, _030413_);
  not g_121540_(_030413_, _030415_);
  xor g_121541_(out[282], _006904_, _030416_);
  not g_121542_(_030416_, _030417_);
  or g_121543_(_030413_, _030417_, _030418_);
  and g_121544_(_030410_, _030418_, _030419_);
  and g_121545_(_030406_, _030408_, _030420_);
  or g_121546_(_030405_, _030409_, _030421_);
  or g_121547_(_030415_, _030416_, _030422_);
  and g_121548_(_030421_, _030422_, _030423_);
  xor g_121549_(_030405_, _030408_, _030424_);
  xor g_121550_(_030413_, _030416_, _030426_);
  and g_121551_(_030419_, _030423_, _030427_);
  or g_121552_(_030424_, _030426_, _030428_);
  or g_121553_(_006771_, _030386_, _030429_);
  not g_121554_(_030429_, _030430_);
  and g_121555_(_030251_, _030386_, _030431_);
  not g_121556_(_030431_, _030432_);
  and g_121557_(_030429_, _030432_, _030433_);
  or g_121558_(_030430_, _030431_, _030434_);
  and g_121559_(_006922_, _030434_, _030435_);
  or g_121560_(_006921_, _030433_, _030437_);
  or g_121561_(_006782_, _030386_, _030438_);
  not g_121562_(_030438_, _030439_);
  and g_121563_(_030257_, _030386_, _030440_);
  not g_121564_(_030440_, _030441_);
  and g_121565_(_030438_, _030441_, _030442_);
  or g_121566_(_030439_, _030440_, _030443_);
  and g_121567_(_006906_, _030443_, _030444_);
  or g_121568_(_006905_, _030442_, _030445_);
  and g_121569_(_030437_, _030445_, _030446_);
  or g_121570_(_030435_, _030444_, _030448_);
  and g_121571_(_006905_, _030442_, _030449_);
  or g_121572_(_006906_, _030443_, _030450_);
  and g_121573_(_006921_, _030433_, _030451_);
  or g_121574_(_006922_, _030434_, _030452_);
  and g_121575_(_030450_, _030452_, _030453_);
  or g_121576_(_030449_, _030451_, _030454_);
  and g_121577_(_030446_, _030453_, _030455_);
  or g_121578_(_030448_, _030454_, _030456_);
  and g_121579_(_030427_, _030455_, _030457_);
  or g_121580_(_030428_, _030456_, _030459_);
  and g_121581_(_030275_, _030386_, _030460_);
  and g_121582_(_006804_, _030385_, _030461_);
  or g_121583_(_030460_, _030461_, _030462_);
  or g_121584_(_006949_, _030462_, _030463_);
  or g_121585_(_006812_, _030386_, _030464_);
  not g_121586_(_030464_, _030465_);
  and g_121587_(_030284_, _030386_, _030466_);
  not g_121588_(_030466_, _030467_);
  and g_121589_(_030464_, _030467_, _030468_);
  or g_121590_(_030465_, _030466_, _030470_);
  and g_121591_(_006944_, _030468_, _030471_);
  or g_121592_(_006944_, _030468_, _030472_);
  xor g_121593_(_006949_, _030462_, _030473_);
  xor g_121594_(_006950_, _030462_, _030474_);
  xor g_121595_(_006944_, _030468_, _030475_);
  xor g_121596_(_006943_, _030468_, _030476_);
  and g_121597_(_030473_, _030475_, _030477_);
  or g_121598_(_030474_, _030476_, _030478_);
  and g_121599_(_006832_, _030385_, _030479_);
  or g_121600_(_006833_, _030386_, _030481_);
  and g_121601_(_030296_, _030386_, _030482_);
  or g_121602_(_030295_, _030385_, _030483_);
  and g_121603_(_030481_, _030483_, _030484_);
  or g_121604_(_030479_, _030482_, _030485_);
  and g_121605_(_006978_, _030485_, _030486_);
  or g_121606_(_006977_, _030484_, _030487_);
  and g_121607_(_006824_, _030385_, _030488_);
  or g_121608_(_006825_, _030386_, _030489_);
  and g_121609_(_030307_, _030386_, _030490_);
  or g_121610_(_030306_, _030385_, _030492_);
  and g_121611_(_030489_, _030492_, _030493_);
  or g_121612_(_030488_, _030490_, _030494_);
  and g_121613_(_006968_, _030494_, _030495_);
  or g_121614_(_006967_, _030493_, _030496_);
  and g_121615_(_030487_, _030496_, _030497_);
  or g_121616_(_030486_, _030495_, _030498_);
  or g_121617_(_006968_, _030494_, _030499_);
  or g_121618_(_006978_, _030485_, _030500_);
  and g_121619_(_030499_, _030500_, _030501_);
  not g_121620_(_030501_, _030503_);
  and g_121621_(_030497_, _030501_, _030504_);
  or g_121622_(_030498_, _030503_, _030505_);
  and g_121623_(_030477_, _030504_, _030506_);
  or g_121624_(_030478_, _030505_, _030507_);
  and g_121625_(_030457_, _030506_, _030508_);
  or g_121626_(_030459_, _030507_, _030509_);
  and g_121627_(_006717_, _030385_, _030510_);
  and g_121628_(_030329_, _030386_, _030511_);
  or g_121629_(_030510_, _030511_, _030512_);
  not g_121630_(_030512_, _030514_);
  and g_121631_(_006996_, _030512_, _030515_);
  or g_121632_(_006997_, _030514_, _030516_);
  and g_121633_(_030333_, _030386_, _030517_);
  and g_121634_(_051426_, _030385_, _030518_);
  or g_121635_(_030517_, _030518_, _030519_);
  or g_121636_(_051642_, _030519_, _030520_);
  not g_121637_(_030520_, _030521_);
  or g_121638_(_030515_, _030521_, _030522_);
  and g_121639_(_006997_, _030514_, _030523_);
  or g_121640_(_006996_, _030512_, _030525_);
  and g_121641_(_051642_, _030519_, _030526_);
  or g_121642_(_030523_, _030526_, _030527_);
  or g_121643_(_030522_, _030527_, _030528_);
  and g_121644_(_030516_, _030525_, _030529_);
  xor g_121645_(_051642_, _030519_, _030530_);
  and g_121646_(_030508_, _030530_, _030531_);
  and g_121647_(_030529_, _030531_, _030532_);
  or g_121648_(_030509_, _030528_, _030533_);
  and g_121649_(_030402_, _030532_, _030534_);
  or g_121650_(_030404_, _030533_, _030536_);
  and g_121651_(_030390_, _030534_, _030537_);
  or g_121652_(_030391_, _030536_, _030538_);
  and g_121653_(_030498_, _030500_, _030539_);
  not g_121654_(_030539_, _030540_);
  and g_121655_(_030477_, _030539_, _030541_);
  or g_121656_(_030478_, _030540_, _030542_);
  or g_121657_(_030463_, _030471_, _030543_);
  and g_121658_(_030472_, _030543_, _030544_);
  not g_121659_(_030544_, _030545_);
  and g_121660_(_030542_, _030544_, _030547_);
  or g_121661_(_030541_, _030545_, _030548_);
  and g_121662_(_030457_, _030548_, _030549_);
  or g_121663_(_030459_, _030547_, _030550_);
  and g_121664_(_030521_, _030525_, _030551_);
  or g_121665_(_030520_, _030523_, _030552_);
  and g_121666_(_030516_, _030552_, _030553_);
  or g_121667_(_030515_, _030551_, _030554_);
  and g_121668_(_030508_, _030554_, _030555_);
  or g_121669_(_030509_, _030553_, _030556_);
  and g_121670_(_030448_, _030450_, _030558_);
  or g_121671_(_030428_, _030446_, _030559_);
  and g_121672_(_030427_, _030558_, _030560_);
  or g_121673_(_030449_, _030559_, _030561_);
  or g_121674_(_030419_, _030420_, _030562_);
  not g_121675_(_030562_, _030563_);
  and g_121676_(_030561_, _030562_, _030564_);
  or g_121677_(_030560_, _030563_, _030565_);
  and g_121678_(_030556_, _030564_, _030566_);
  or g_121679_(_030555_, _030565_, _030567_);
  and g_121680_(_030550_, _030566_, _030569_);
  or g_121681_(_030549_, _030567_, _030570_);
  and g_121682_(_030399_, _030404_, _030571_);
  or g_121683_(_030398_, _030402_, _030572_);
  or g_121684_(_030533_, _030571_, _030573_);
  and g_121685_(_030532_, _030572_, _030574_);
  and g_121686_(_030569_, _030573_, _030575_);
  or g_121687_(_030570_, _030574_, _030576_);
  and g_121688_(_030538_, _030576_, _030577_);
  or g_121689_(_030537_, _030575_, _030578_);
  and g_121690_(_030389_, _030578_, _030580_);
  and g_121691_(_004443_, _030577_, _030581_);
  or g_121692_(_030580_, _030581_, _030582_);
  and g_121693_(_030405_, _030408_, _030583_);
  or g_121694_(_030406_, _030409_, _030584_);
  or g_121695_(out[298], _007082_, _030585_);
  xor g_121696_(out[299], _030585_, _030586_);
  xor g_121697_(_004465_, _030585_, _030587_);
  and g_121698_(_030583_, _030587_, _030588_);
  or g_121699_(_030584_, _030586_, _030589_);
  and g_121700_(_030413_, _030578_, _030591_);
  not g_121701_(_030591_, _030592_);
  or g_121702_(_030417_, _030578_, _030593_);
  not g_121703_(_030593_, _030594_);
  and g_121704_(_030592_, _030593_, _030595_);
  or g_121705_(_030591_, _030594_, _030596_);
  xor g_121706_(out[298], _007082_, _030597_);
  xor g_121707_(_004487_, _007082_, _030598_);
  and g_121708_(_030595_, _030597_, _030599_);
  or g_121709_(_030596_, _030598_, _030600_);
  and g_121710_(_030589_, _030600_, _030602_);
  or g_121711_(_030588_, _030599_, _030603_);
  and g_121712_(_030596_, _030598_, _030604_);
  or g_121713_(_030595_, _030597_, _030605_);
  and g_121714_(_030584_, _030586_, _030606_);
  or g_121715_(_030583_, _030587_, _030607_);
  and g_121716_(_006905_, _030577_, _030608_);
  and g_121717_(_030443_, _030578_, _030609_);
  or g_121718_(_030608_, _030609_, _030610_);
  or g_121719_(_007085_, _030610_, _030611_);
  and g_121720_(_030434_, _030578_, _030613_);
  and g_121721_(_006921_, _030577_, _030614_);
  or g_121722_(_030613_, _030614_, _030615_);
  and g_121723_(_007100_, _030615_, _030616_);
  not g_121724_(_030616_, _030617_);
  and g_121725_(_007085_, _030610_, _030618_);
  not g_121726_(_030618_, _030619_);
  and g_121727_(_030617_, _030619_, _030620_);
  or g_121728_(_030616_, _030618_, _030621_);
  or g_121729_(_007100_, _030615_, _030622_);
  and g_121730_(_030605_, _030607_, _030624_);
  or g_121731_(_030604_, _030606_, _030625_);
  and g_121732_(_030602_, _030624_, _030626_);
  or g_121733_(_030603_, _030625_, _030627_);
  and g_121734_(_030611_, _030622_, _030628_);
  not g_121735_(_030628_, _030629_);
  and g_121736_(_030620_, _030628_, _030630_);
  or g_121737_(_030621_, _030629_, _030631_);
  and g_121738_(_030626_, _030630_, _030632_);
  or g_121739_(_030627_, _030631_, _030633_);
  and g_121740_(_030462_, _030578_, _030635_);
  and g_121741_(_006950_, _030577_, _030636_);
  or g_121742_(_030635_, _030636_, _030637_);
  or g_121743_(_007129_, _030637_, _030638_);
  not g_121744_(_030638_, _030639_);
  xor g_121745_(_007129_, _030637_, _030640_);
  xor g_121746_(_007130_, _030637_, _030641_);
  and g_121747_(_030470_, _030578_, _030642_);
  or g_121748_(_030468_, _030577_, _030643_);
  and g_121749_(_006944_, _030577_, _030644_);
  or g_121750_(_006943_, _030578_, _030646_);
  and g_121751_(_030643_, _030646_, _030647_);
  or g_121752_(_030642_, _030644_, _030648_);
  and g_121753_(_007121_, _030648_, _030649_);
  or g_121754_(_007122_, _030647_, _030650_);
  and g_121755_(_007122_, _030647_, _030651_);
  or g_121756_(_007121_, _030648_, _030652_);
  and g_121757_(_030650_, _030652_, _030653_);
  or g_121758_(_030649_, _030651_, _030654_);
  and g_121759_(_030640_, _030653_, _030655_);
  or g_121760_(_030641_, _030654_, _030657_);
  or g_121761_(_006968_, _030578_, _030658_);
  not g_121762_(_030658_, _030659_);
  and g_121763_(_030494_, _030578_, _030660_);
  not g_121764_(_030660_, _030661_);
  and g_121765_(_030658_, _030661_, _030662_);
  or g_121766_(_030659_, _030660_, _030663_);
  and g_121767_(_007146_, _030663_, _030664_);
  or g_121768_(_007145_, _030662_, _030665_);
  and g_121769_(_030485_, _030578_, _030666_);
  not g_121770_(_030666_, _030668_);
  or g_121771_(_006978_, _030578_, _030669_);
  not g_121772_(_030669_, _030670_);
  and g_121773_(_030668_, _030669_, _030671_);
  or g_121774_(_030666_, _030670_, _030672_);
  and g_121775_(_007154_, _030672_, _030673_);
  or g_121776_(_007153_, _030671_, _030674_);
  and g_121777_(_030665_, _030674_, _030675_);
  or g_121778_(_030664_, _030673_, _030676_);
  or g_121779_(_007154_, _030672_, _030677_);
  not g_121780_(_030677_, _030679_);
  or g_121781_(_007146_, _030663_, _030680_);
  and g_121782_(_030677_, _030680_, _030681_);
  not g_121783_(_030681_, _030682_);
  and g_121784_(_030675_, _030681_, _030683_);
  or g_121785_(_030676_, _030682_, _030684_);
  and g_121786_(_030655_, _030683_, _030685_);
  or g_121787_(_030657_, _030684_, _030686_);
  and g_121788_(_030632_, _030685_, _030687_);
  or g_121789_(_030633_, _030686_, _030688_);
  and g_121790_(_030512_, _030578_, _030690_);
  not g_121791_(_030690_, _030691_);
  or g_121792_(_006996_, _030578_, _030692_);
  not g_121793_(_030692_, _030693_);
  and g_121794_(_030691_, _030692_, _030694_);
  or g_121795_(_030690_, _030693_, _030695_);
  and g_121796_(_007174_, _030695_, _030696_);
  or g_121797_(_007175_, _030694_, _030697_);
  and g_121798_(_007175_, _030694_, _030698_);
  or g_121799_(_007174_, _030695_, _030699_);
  and g_121800_(_030697_, _030699_, _030701_);
  or g_121801_(_030696_, _030698_, _030702_);
  and g_121802_(_030519_, _030578_, _030703_);
  and g_121803_(_051641_, _030577_, _030704_);
  or g_121804_(_030703_, _030704_, _030705_);
  not g_121805_(_030705_, _030706_);
  and g_121806_(_051816_, _030706_, _030707_);
  or g_121807_(_051817_, _030705_, _030708_);
  xor g_121808_(_051817_, _030705_, _030709_);
  xor g_121809_(_051816_, _030705_, _030710_);
  and g_121810_(_030701_, _030709_, _030712_);
  or g_121811_(_030702_, _030710_, _030713_);
  or g_121812_(_030395_, _030577_, _030714_);
  or g_121813_(_053126_, _030578_, _030715_);
  and g_121814_(_030714_, _030715_, _030716_);
  and g_121815_(out[289], _030716_, _030717_);
  not g_121816_(_030717_, _030718_);
  and g_121817_(out[288], _030582_, _030719_);
  not g_121818_(_030719_, _030720_);
  xor g_121819_(out[289], _030716_, _030721_);
  xor g_121820_(_053225_, _030716_, _030723_);
  and g_121821_(_030720_, _030721_, _030724_);
  or g_121822_(_030719_, _030723_, _030725_);
  and g_121823_(_030718_, _030725_, _030726_);
  or g_121824_(_030717_, _030724_, _030727_);
  and g_121825_(_030712_, _030727_, _030728_);
  or g_121826_(_030713_, _030726_, _030729_);
  and g_121827_(_030697_, _030708_, _030730_);
  or g_121828_(_030696_, _030707_, _030731_);
  and g_121829_(_030699_, _030731_, _030732_);
  or g_121830_(_030698_, _030730_, _030734_);
  and g_121831_(_030729_, _030734_, _030735_);
  or g_121832_(_030728_, _030732_, _030736_);
  and g_121833_(_030687_, _030736_, _030737_);
  or g_121834_(_030688_, _030735_, _030738_);
  and g_121835_(_030655_, _030676_, _030739_);
  or g_121836_(_030657_, _030675_, _030740_);
  and g_121837_(_030677_, _030739_, _030741_);
  or g_121838_(_030679_, _030740_, _030742_);
  and g_121839_(_030639_, _030652_, _030743_);
  or g_121840_(_030638_, _030651_, _030745_);
  and g_121841_(_030650_, _030745_, _030746_);
  or g_121842_(_030649_, _030743_, _030747_);
  and g_121843_(_030742_, _030746_, _030748_);
  or g_121844_(_030741_, _030747_, _030749_);
  and g_121845_(_030632_, _030749_, _030750_);
  or g_121846_(_030633_, _030748_, _030751_);
  and g_121847_(_030611_, _030621_, _030752_);
  not g_121848_(_030752_, _030753_);
  and g_121849_(_030626_, _030752_, _030754_);
  or g_121850_(_030627_, _030753_, _030756_);
  and g_121851_(_030603_, _030607_, _030757_);
  or g_121852_(_030602_, _030606_, _030758_);
  and g_121853_(_030756_, _030758_, _030759_);
  or g_121854_(_030754_, _030757_, _030760_);
  and g_121855_(_030751_, _030759_, _030761_);
  or g_121856_(_030750_, _030760_, _030762_);
  and g_121857_(_030738_, _030761_, _030763_);
  or g_121858_(_030737_, _030762_, _030764_);
  or g_121859_(out[288], _030582_, _030765_);
  not g_121860_(_030765_, _030767_);
  and g_121861_(_030712_, _030765_, _030768_);
  or g_121862_(_030713_, _030767_, _030769_);
  and g_121863_(_030724_, _030768_, _030770_);
  or g_121864_(_030725_, _030769_, _030771_);
  and g_121865_(_030687_, _030770_, _030772_);
  or g_121866_(_030688_, _030771_, _030773_);
  and g_121867_(_030764_, _030773_, _030774_);
  or g_121868_(_030763_, _030772_, _030775_);
  and g_121869_(_030582_, _030775_, _030776_);
  and g_121870_(_004476_, _030774_, _030778_);
  or g_121871_(_030776_, _030778_, _030779_);
  and g_121872_(_030583_, _030586_, _030780_);
  or g_121873_(_030584_, _030587_, _030781_);
  or g_121874_(out[314], _007252_, _030782_);
  xor g_121875_(out[315], _030782_, _030783_);
  xor g_121876_(_004498_, _030782_, _030784_);
  and g_121877_(_030780_, _030784_, _030785_);
  or g_121878_(_030781_, _030783_, _030786_);
  or g_121879_(_030598_, _030775_, _030787_);
  not g_121880_(_030787_, _030789_);
  and g_121881_(_030596_, _030775_, _030790_);
  or g_121882_(_030595_, _030774_, _030791_);
  and g_121883_(_030787_, _030791_, _030792_);
  or g_121884_(_030789_, _030790_, _030793_);
  xor g_121885_(out[314], _007252_, _030794_);
  xor g_121886_(_004520_, _007252_, _030795_);
  and g_121887_(_030792_, _030794_, _030796_);
  or g_121888_(_030793_, _030795_, _030797_);
  and g_121889_(_030786_, _030797_, _030798_);
  or g_121890_(_030785_, _030796_, _030800_);
  and g_121891_(_030781_, _030783_, _030801_);
  and g_121892_(_030793_, _030795_, _030802_);
  or g_121893_(_030800_, _030802_, _030803_);
  or g_121894_(_030801_, _030803_, _030804_);
  or g_121895_(_007100_, _030775_, _030805_);
  not g_121896_(_030805_, _030806_);
  and g_121897_(_030615_, _030775_, _030807_);
  not g_121898_(_030807_, _030808_);
  and g_121899_(_030805_, _030808_, _030809_);
  or g_121900_(_030806_, _030807_, _030811_);
  and g_121901_(_007264_, _030811_, _030812_);
  or g_121902_(_007263_, _030809_, _030813_);
  or g_121903_(_007085_, _030775_, _030814_);
  not g_121904_(_030814_, _030815_);
  and g_121905_(_030610_, _030775_, _030816_);
  not g_121906_(_030816_, _030817_);
  and g_121907_(_030814_, _030817_, _030818_);
  or g_121908_(_030815_, _030816_, _030819_);
  and g_121909_(_007254_, _030819_, _030820_);
  or g_121910_(_007253_, _030818_, _030822_);
  and g_121911_(_030813_, _030822_, _030823_);
  or g_121912_(_030812_, _030820_, _030824_);
  and g_121913_(_007263_, _030809_, _030825_);
  and g_121914_(_007253_, _030818_, _030826_);
  or g_121915_(_030825_, _030826_, _030827_);
  or g_121916_(_030824_, _030827_, _030828_);
  or g_121917_(_030804_, _030828_, _030829_);
  or g_121918_(_007154_, _030775_, _030830_);
  not g_121919_(_030830_, _030831_);
  and g_121920_(_030672_, _030775_, _030833_);
  not g_121921_(_030833_, _030834_);
  and g_121922_(_030830_, _030834_, _030835_);
  or g_121923_(_030831_, _030833_, _030836_);
  or g_121924_(_007302_, _030835_, _030837_);
  or g_121925_(_007146_, _030775_, _030838_);
  not g_121926_(_030838_, _030839_);
  and g_121927_(_030663_, _030775_, _030840_);
  not g_121928_(_030840_, _030841_);
  and g_121929_(_030838_, _030841_, _030842_);
  or g_121930_(_030839_, _030840_, _030844_);
  or g_121931_(_007317_, _030842_, _030845_);
  and g_121932_(_030837_, _030845_, _030846_);
  not g_121933_(_030846_, _030847_);
  and g_121934_(_007122_, _030774_, _030848_);
  or g_121935_(_007121_, _030775_, _030849_);
  and g_121936_(_030648_, _030775_, _030850_);
  or g_121937_(_030647_, _030774_, _030851_);
  and g_121938_(_030849_, _030851_, _030852_);
  or g_121939_(_030848_, _030850_, _030853_);
  or g_121940_(_007284_, _030852_, _030855_);
  and g_121941_(_007284_, _030852_, _030856_);
  xor g_121942_(_007283_, _030852_, _030857_);
  and g_121943_(_007130_, _030774_, _030858_);
  and g_121944_(_030637_, _030775_, _030859_);
  or g_121945_(_030858_, _030859_, _030860_);
  or g_121946_(_007293_, _030860_, _030861_);
  and g_121947_(_007302_, _030835_, _030862_);
  xor g_121948_(_007294_, _030860_, _030863_);
  or g_121949_(_030857_, _030863_, _030864_);
  or g_121950_(_030862_, _030864_, _030866_);
  or g_121951_(_030846_, _030866_, _030867_);
  or g_121952_(_030856_, _030861_, _030868_);
  and g_121953_(_030855_, _030868_, _030869_);
  and g_121954_(_030867_, _030869_, _030870_);
  or g_121955_(_030829_, _030870_, _030871_);
  and g_121956_(_007317_, _030842_, _030872_);
  or g_121957_(_030866_, _030872_, _030873_);
  or g_121958_(_030829_, _030873_, _030874_);
  not g_121959_(_030874_, _030875_);
  and g_121960_(_030846_, _030875_, _030877_);
  or g_121961_(_030847_, _030874_, _030878_);
  or g_121962_(_007174_, _030775_, _030879_);
  not g_121963_(_030879_, _030880_);
  and g_121964_(_030695_, _030775_, _030881_);
  not g_121965_(_030881_, _030882_);
  and g_121966_(_030879_, _030882_, _030883_);
  or g_121967_(_030880_, _030881_, _030884_);
  or g_121968_(_007343_, _030883_, _030885_);
  and g_121969_(_030705_, _030775_, _030886_);
  and g_121970_(_051816_, _030774_, _030888_);
  or g_121971_(_030886_, _030888_, _030889_);
  or g_121972_(_051958_, _030889_, _030890_);
  and g_121973_(_007343_, _030883_, _030891_);
  xor g_121974_(_007343_, _030883_, _030892_);
  xor g_121975_(_007342_, _030883_, _030893_);
  xor g_121976_(_051958_, _030889_, _030894_);
  xor g_121977_(_051957_, _030889_, _030895_);
  and g_121978_(_030892_, _030894_, _030896_);
  or g_121979_(_030893_, _030895_, _030897_);
  or g_121980_(_053225_, _030775_, _030899_);
  or g_121981_(_030716_, _030774_, _030900_);
  and g_121982_(_030899_, _030900_, _030901_);
  and g_121983_(out[305], _030901_, _030902_);
  not g_121984_(_030902_, _030903_);
  and g_121985_(out[304], _030779_, _030904_);
  not g_121986_(_030904_, _030905_);
  xor g_121987_(out[305], _030901_, _030906_);
  xor g_121988_(_053324_, _030901_, _030907_);
  and g_121989_(_030905_, _030906_, _030908_);
  or g_121990_(_030904_, _030907_, _030910_);
  and g_121991_(_030903_, _030910_, _030911_);
  or g_121992_(_030897_, _030911_, _030912_);
  or g_121993_(_030890_, _030891_, _030913_);
  and g_121994_(_030885_, _030913_, _030914_);
  and g_121995_(_030912_, _030914_, _030915_);
  or g_121996_(_030878_, _030915_, _030916_);
  or g_121997_(_030798_, _030801_, _030917_);
  or g_121998_(_030823_, _030826_, _030918_);
  or g_121999_(_030804_, _030918_, _030919_);
  and g_122000_(_030917_, _030919_, _030921_);
  and g_122001_(_030916_, _030921_, _030922_);
  and g_122002_(_030871_, _030922_, _030923_);
  or g_122003_(out[304], _030779_, _030924_);
  and g_122004_(_030896_, _030924_, _030925_);
  and g_122005_(_030908_, _030925_, _030926_);
  and g_122006_(_030877_, _030926_, _030927_);
  or g_122007_(_030923_, _030927_, _030928_);
  not g_122008_(_030928_, _030929_);
  and g_122009_(_030779_, _030928_, _030930_);
  not g_122010_(_030930_, _030932_);
  or g_122011_(out[304], _030928_, _030933_);
  not g_122012_(_030933_, _030934_);
  and g_122013_(_030932_, _030933_, _030935_);
  or g_122014_(_030930_, _030934_, _030936_);
  and g_122015_(_030780_, _030783_, _030937_);
  or g_122016_(_030781_, _030784_, _030938_);
  or g_122017_(out[330], _007418_, _030939_);
  xor g_122018_(out[331], _030939_, _030940_);
  xor g_122019_(_004531_, _030939_, _030941_);
  and g_122020_(_030937_, _030941_, _030943_);
  or g_122021_(_030938_, _030940_, _030944_);
  and g_122022_(_030794_, _030929_, _030945_);
  or g_122023_(_030795_, _030928_, _030946_);
  and g_122024_(_030793_, _030928_, _030947_);
  not g_122025_(_030947_, _030948_);
  and g_122026_(_030946_, _030948_, _030949_);
  or g_122027_(_030945_, _030947_, _030950_);
  xor g_122028_(out[330], _007418_, _030951_);
  xor g_122029_(_004553_, _007418_, _030952_);
  and g_122030_(_030949_, _030951_, _030954_);
  or g_122031_(_030950_, _030952_, _030955_);
  and g_122032_(_030944_, _030955_, _030956_);
  or g_122033_(_030943_, _030954_, _030957_);
  and g_122034_(_030950_, _030952_, _030958_);
  and g_122035_(_030938_, _030940_, _030959_);
  or g_122036_(_030958_, _030959_, _030960_);
  not g_122037_(_030960_, _030961_);
  and g_122038_(_030956_, _030961_, _030962_);
  or g_122039_(_030957_, _030960_, _030963_);
  and g_122040_(_007263_, _030929_, _030965_);
  and g_122041_(_030811_, _030928_, _030966_);
  or g_122042_(_030965_, _030966_, _030967_);
  not g_122043_(_030967_, _030968_);
  and g_122044_(_007429_, _030967_, _030969_);
  or g_122045_(_007428_, _030968_, _030970_);
  and g_122046_(_007253_, _030929_, _030971_);
  and g_122047_(_030819_, _030928_, _030972_);
  or g_122048_(_030971_, _030972_, _030973_);
  and g_122049_(_007420_, _030973_, _030974_);
  not g_122050_(_030974_, _030976_);
  and g_122051_(_030970_, _030976_, _030977_);
  or g_122052_(_030969_, _030974_, _030978_);
  or g_122053_(_007420_, _030973_, _030979_);
  or g_122054_(_007429_, _030967_, _030980_);
  and g_122055_(_030979_, _030980_, _030981_);
  not g_122056_(_030981_, _030982_);
  and g_122057_(_030977_, _030981_, _030983_);
  or g_122058_(_030978_, _030982_, _030984_);
  and g_122059_(_030962_, _030983_, _030985_);
  or g_122060_(_030963_, _030984_, _030987_);
  and g_122061_(_007294_, _030929_, _030988_);
  and g_122062_(_030860_, _030928_, _030989_);
  or g_122063_(_030988_, _030989_, _030990_);
  or g_122064_(_007514_, _030990_, _030991_);
  not g_122065_(_030991_, _030992_);
  xor g_122066_(_007514_, _030990_, _030993_);
  or g_122067_(_007283_, _030928_, _030994_);
  not g_122068_(_030994_, _030995_);
  and g_122069_(_030853_, _030928_, _030996_);
  or g_122070_(_030852_, _030929_, _030998_);
  and g_122071_(_030994_, _030998_, _030999_);
  or g_122072_(_030995_, _030996_, _031000_);
  and g_122073_(_007503_, _031000_, _031001_);
  or g_122074_(_007504_, _030999_, _031002_);
  or g_122075_(_007503_, _031000_, _031003_);
  and g_122076_(_030993_, _031003_, _031004_);
  not g_122077_(_031004_, _031005_);
  and g_122078_(_031002_, _031004_, _031006_);
  or g_122079_(_031001_, _031005_, _031007_);
  and g_122080_(_007302_, _030929_, _031009_);
  and g_122081_(_030836_, _030928_, _031010_);
  or g_122082_(_031009_, _031010_, _031011_);
  and g_122083_(_007526_, _031011_, _031012_);
  and g_122084_(_007317_, _030929_, _031013_);
  and g_122085_(_030844_, _030928_, _031014_);
  or g_122086_(_031013_, _031014_, _031015_);
  and g_122087_(_007546_, _031015_, _031016_);
  or g_122088_(_031012_, _031016_, _031017_);
  or g_122089_(_007526_, _031011_, _031018_);
  xor g_122090_(_007546_, _031015_, _031020_);
  xor g_122091_(_007544_, _031015_, _031021_);
  xor g_122092_(_007526_, _031011_, _031022_);
  xor g_122093_(_007525_, _031011_, _031023_);
  and g_122094_(_031020_, _031022_, _031024_);
  or g_122095_(_031021_, _031023_, _031025_);
  and g_122096_(_031006_, _031024_, _031026_);
  or g_122097_(_031007_, _031025_, _031027_);
  and g_122098_(_030985_, _031026_, _031028_);
  or g_122099_(_030987_, _031027_, _031029_);
  and g_122100_(_007343_, _030929_, _031031_);
  and g_122101_(_030884_, _030928_, _031032_);
  or g_122102_(_031031_, _031032_, _031033_);
  and g_122103_(_007462_, _031033_, _031034_);
  or g_122104_(_007462_, _031033_, _031035_);
  xor g_122105_(_007462_, _031033_, _031036_);
  xor g_122106_(_007463_, _031033_, _031037_);
  and g_122107_(_030889_, _030928_, _031038_);
  and g_122108_(_051957_, _030929_, _031039_);
  or g_122109_(_031038_, _031039_, _031040_);
  or g_122110_(_052168_, _031040_, _031042_);
  not g_122111_(_031042_, _031043_);
  xor g_122112_(_052168_, _031040_, _031044_);
  xor g_122113_(_052167_, _031040_, _031045_);
  and g_122114_(_031036_, _031044_, _031046_);
  or g_122115_(_031037_, _031045_, _031047_);
  and g_122116_(_030901_, _030928_, _031048_);
  not g_122117_(_031048_, _031049_);
  or g_122118_(out[305], _030928_, _031050_);
  not g_122119_(_031050_, _031051_);
  or g_122120_(_031048_, _031051_, _031053_);
  and g_122121_(_031049_, _031050_, _031054_);
  and g_122122_(out[321], _031053_, _031055_);
  or g_122123_(_053423_, _031054_, _031056_);
  and g_122124_(out[320], _030936_, _031057_);
  or g_122125_(_004542_, _030935_, _031058_);
  xor g_122126_(out[321], _031053_, _031059_);
  xor g_122127_(_053423_, _031053_, _031060_);
  and g_122128_(_031058_, _031059_, _031061_);
  or g_122129_(_031057_, _031060_, _031062_);
  and g_122130_(_031056_, _031062_, _031064_);
  or g_122131_(_031055_, _031061_, _031065_);
  and g_122132_(_031046_, _031065_, _031066_);
  or g_122133_(_031047_, _031064_, _031067_);
  or g_122134_(_031034_, _031043_, _031068_);
  and g_122135_(_031035_, _031068_, _031069_);
  not g_122136_(_031069_, _031070_);
  and g_122137_(_031067_, _031070_, _031071_);
  or g_122138_(_031066_, _031069_, _031072_);
  and g_122139_(_031028_, _031072_, _031073_);
  or g_122140_(_031029_, _031071_, _031075_);
  and g_122141_(_031017_, _031018_, _031076_);
  and g_122142_(_031006_, _031076_, _031077_);
  or g_122143_(_030992_, _031001_, _031078_);
  and g_122144_(_031003_, _031078_, _031079_);
  or g_122145_(_031077_, _031079_, _031080_);
  and g_122146_(_030985_, _031080_, _031081_);
  not g_122147_(_031081_, _031082_);
  or g_122148_(_030956_, _030959_, _031083_);
  not g_122149_(_031083_, _031084_);
  and g_122150_(_030978_, _030979_, _031086_);
  and g_122151_(_030962_, _031086_, _031087_);
  not g_122152_(_031087_, _031088_);
  or g_122153_(_031084_, _031087_, _031089_);
  or g_122154_(_031081_, _031089_, _031090_);
  and g_122155_(_031075_, _031088_, _031091_);
  and g_122156_(_031082_, _031083_, _031092_);
  and g_122157_(_031091_, _031092_, _031093_);
  or g_122158_(_031073_, _031090_, _031094_);
  or g_122159_(out[320], _030936_, _031095_);
  and g_122160_(_031046_, _031095_, _031097_);
  not g_122161_(_031097_, _031098_);
  and g_122162_(_031061_, _031097_, _031099_);
  or g_122163_(_031062_, _031098_, _031100_);
  and g_122164_(_031028_, _031099_, _031101_);
  or g_122165_(_031029_, _031100_, _031102_);
  and g_122166_(_031094_, _031102_, _031103_);
  or g_122167_(_031093_, _031101_, _031104_);
  and g_122168_(_030936_, _031104_, _031105_);
  and g_122169_(_004542_, _031103_, _031106_);
  or g_122170_(_031105_, _031106_, _031108_);
  or g_122171_(out[346], _007673_, _031109_);
  xor g_122172_(out[346], _007673_, _031110_);
  or g_122173_(_030952_, _031104_, _031111_);
  not g_122174_(_031111_, _031112_);
  and g_122175_(_030950_, _031104_, _031113_);
  not g_122176_(_031113_, _031114_);
  and g_122177_(_031111_, _031114_, _031115_);
  or g_122178_(_031112_, _031113_, _031116_);
  and g_122179_(_030937_, _030940_, _031117_);
  or g_122180_(_030938_, _030941_, _031119_);
  xor g_122181_(out[347], _031109_, _031120_);
  xor g_122182_(_004564_, _031109_, _031121_);
  or g_122183_(_031117_, _031121_, _031122_);
  and g_122184_(_031117_, _031121_, _031123_);
  xor g_122185_(_031119_, _031120_, _031124_);
  xor g_122186_(_031117_, _031120_, _031125_);
  and g_122187_(_031110_, _031115_, _031126_);
  xor g_122188_(_031110_, _031115_, _031127_);
  xor g_122189_(_031110_, _031116_, _031128_);
  and g_122190_(_031124_, _031127_, _031130_);
  or g_122191_(_031125_, _031128_, _031131_);
  and g_122192_(_007419_, _031103_, _031132_);
  and g_122193_(_030973_, _031104_, _031133_);
  or g_122194_(_031132_, _031133_, _031134_);
  not g_122195_(_031134_, _031135_);
  and g_122196_(_007675_, _031134_, _031136_);
  or g_122197_(_007674_, _031135_, _031137_);
  and g_122198_(_007428_, _031103_, _031138_);
  and g_122199_(_030967_, _031104_, _031139_);
  or g_122200_(_031138_, _031139_, _031141_);
  not g_122201_(_031141_, _031142_);
  and g_122202_(_007682_, _031141_, _031143_);
  or g_122203_(_007681_, _031142_, _031144_);
  and g_122204_(_031137_, _031144_, _031145_);
  or g_122205_(_031136_, _031143_, _031146_);
  and g_122206_(_007674_, _031135_, _031147_);
  or g_122207_(_007675_, _031134_, _031148_);
  and g_122208_(_007681_, _031142_, _031149_);
  or g_122209_(_007682_, _031141_, _031150_);
  and g_122210_(_031148_, _031150_, _031152_);
  or g_122211_(_031147_, _031149_, _031153_);
  and g_122212_(_031145_, _031152_, _031154_);
  or g_122213_(_031146_, _031153_, _031155_);
  and g_122214_(_031130_, _031154_, _031156_);
  or g_122215_(_031131_, _031155_, _031157_);
  and g_122216_(_052167_, _031103_, _031158_);
  and g_122217_(_031040_, _031104_, _031159_);
  or g_122218_(_031158_, _031159_, _031160_);
  or g_122219_(_052355_, _031160_, _031161_);
  and g_122220_(_007463_, _031103_, _031163_);
  and g_122221_(_031033_, _031104_, _031164_);
  or g_122222_(_031163_, _031164_, _031165_);
  not g_122223_(_031165_, _031166_);
  and g_122224_(_007616_, _031165_, _031167_);
  or g_122225_(_007617_, _031166_, _031168_);
  and g_122226_(_031161_, _031168_, _031169_);
  or g_122227_(_053423_, _031104_, _031170_);
  or g_122228_(_031053_, _031103_, _031171_);
  and g_122229_(_031170_, _031171_, _031172_);
  and g_122230_(out[337], _031172_, _031174_);
  not g_122231_(_031174_, _031175_);
  and g_122232_(out[336], _031108_, _031176_);
  xor g_122233_(_053522_, _031172_, _031177_);
  or g_122234_(_031176_, _031177_, _031178_);
  and g_122235_(_031175_, _031178_, _031179_);
  xor g_122236_(_052354_, _031160_, _031180_);
  or g_122237_(_031167_, _031180_, _031181_);
  or g_122238_(_031179_, _031181_, _031182_);
  and g_122239_(_031169_, _031182_, _031183_);
  and g_122240_(_007504_, _031103_, _031185_);
  or g_122241_(_007503_, _031104_, _031186_);
  and g_122242_(_031000_, _031104_, _031187_);
  or g_122243_(_030999_, _031103_, _031188_);
  and g_122244_(_031186_, _031188_, _031189_);
  or g_122245_(_031185_, _031187_, _031190_);
  and g_122246_(_007702_, _031190_, _031191_);
  or g_122247_(_007514_, _031104_, _031192_);
  and g_122248_(_030990_, _031104_, _031193_);
  not g_122249_(_031193_, _031194_);
  and g_122250_(_031192_, _031194_, _031196_);
  and g_122251_(_007713_, _031196_, _031197_);
  or g_122252_(_007702_, _031190_, _031198_);
  and g_122253_(_007525_, _031103_, _031199_);
  and g_122254_(_031011_, _031104_, _031200_);
  or g_122255_(_031199_, _031200_, _031201_);
  or g_122256_(_007737_, _031201_, _031202_);
  not g_122257_(_031202_, _031203_);
  xor g_122258_(_007703_, _031189_, _031204_);
  xor g_122259_(_007702_, _031189_, _031205_);
  xor g_122260_(_007713_, _031196_, _031207_);
  xor g_122261_(_007712_, _031196_, _031208_);
  and g_122262_(_031204_, _031207_, _031209_);
  or g_122263_(_031205_, _031208_, _031210_);
  and g_122264_(_031202_, _031209_, _031211_);
  or g_122265_(_031203_, _031210_, _031212_);
  and g_122266_(_007544_, _031103_, _031213_);
  and g_122267_(_031015_, _031104_, _031214_);
  or g_122268_(_031213_, _031214_, _031215_);
  and g_122269_(_007726_, _031215_, _031216_);
  and g_122270_(_007737_, _031201_, _031218_);
  or g_122271_(_031216_, _031218_, _031219_);
  or g_122272_(_007726_, _031215_, _031220_);
  not g_122273_(_031220_, _031221_);
  or g_122274_(_031219_, _031221_, _031222_);
  or g_122275_(_031212_, _031222_, _031223_);
  and g_122276_(_007617_, _031166_, _031224_);
  or g_122277_(_007616_, _031165_, _031225_);
  or g_122278_(_031223_, _031224_, _031226_);
  or g_122279_(_031183_, _031226_, _031227_);
  and g_122280_(_031211_, _031219_, _031229_);
  and g_122281_(_031197_, _031198_, _031230_);
  or g_122282_(_031191_, _031230_, _031231_);
  or g_122283_(_031229_, _031231_, _031232_);
  not g_122284_(_031232_, _031233_);
  and g_122285_(_031227_, _031233_, _031234_);
  or g_122286_(_031157_, _031234_, _031235_);
  and g_122287_(_031146_, _031148_, _031236_);
  and g_122288_(_031130_, _031236_, _031237_);
  or g_122289_(_031123_, _031126_, _031238_);
  and g_122290_(_031122_, _031238_, _031240_);
  or g_122291_(_031237_, _031240_, _031241_);
  not g_122292_(_031241_, _031242_);
  and g_122293_(_031235_, _031242_, _031243_);
  or g_122294_(out[336], _031108_, _031244_);
  and g_122295_(_031225_, _031244_, _031245_);
  not g_122296_(_031245_, _031246_);
  or g_122297_(_031178_, _031246_, _031247_);
  or g_122298_(_031181_, _031247_, _031248_);
  or g_122299_(_031223_, _031248_, _031249_);
  not g_122300_(_031249_, _031251_);
  and g_122301_(_031156_, _031251_, _031252_);
  or g_122302_(_031243_, _031252_, _031253_);
  not g_122303_(_031253_, _031254_);
  and g_122304_(_031108_, _031253_, _031255_);
  and g_122305_(_004575_, _031254_, _031256_);
  or g_122306_(_031255_, _031256_, _031257_);
  and g_122307_(_031117_, _031120_, _031258_);
  or g_122308_(_031119_, _031121_, _031259_);
  or g_122309_(out[362], _007799_, _031260_);
  xor g_122310_(out[363], _031260_, _031262_);
  xor g_122311_(_004597_, _031260_, _031263_);
  or g_122312_(_031259_, _031262_, _031264_);
  xor g_122313_(out[362], _007799_, _031265_);
  xor g_122314_(_004619_, _007799_, _031266_);
  and g_122315_(_031110_, _031254_, _031267_);
  and g_122316_(_031116_, _031253_, _031268_);
  or g_122317_(_031267_, _031268_, _031269_);
  or g_122318_(_031266_, _031269_, _031270_);
  and g_122319_(_031264_, _031270_, _031271_);
  not g_122320_(_031271_, _031273_);
  and g_122321_(_031266_, _031269_, _031274_);
  and g_122322_(_031259_, _031262_, _031275_);
  or g_122323_(_031274_, _031275_, _031276_);
  or g_122324_(_031273_, _031276_, _031277_);
  or g_122325_(_007682_, _031253_, _031278_);
  not g_122326_(_031278_, _031279_);
  and g_122327_(_031141_, _031253_, _031280_);
  not g_122328_(_031280_, _031281_);
  and g_122329_(_031278_, _031281_, _031282_);
  or g_122330_(_031279_, _031280_, _031284_);
  or g_122331_(_007813_, _031282_, _031285_);
  or g_122332_(_007675_, _031253_, _031286_);
  not g_122333_(_031286_, _031287_);
  and g_122334_(_031134_, _031253_, _031288_);
  not g_122335_(_031288_, _031289_);
  and g_122336_(_031286_, _031289_, _031290_);
  or g_122337_(_031287_, _031288_, _031291_);
  or g_122338_(_007800_, _031290_, _031292_);
  and g_122339_(_031285_, _031292_, _031293_);
  not g_122340_(_031293_, _031295_);
  and g_122341_(_007800_, _031290_, _031296_);
  and g_122342_(_007813_, _031282_, _031297_);
  or g_122343_(_031296_, _031297_, _031298_);
  or g_122344_(_031295_, _031298_, _031299_);
  or g_122345_(_031277_, _031299_, _031300_);
  and g_122346_(_007703_, _031254_, _031301_);
  and g_122347_(_031190_, _031253_, _031302_);
  or g_122348_(_031301_, _031302_, _031303_);
  and g_122349_(_007850_, _031303_, _031304_);
  or g_122350_(_007712_, _031253_, _031306_);
  or g_122351_(_031196_, _031254_, _031307_);
  and g_122352_(_031306_, _031307_, _031308_);
  and g_122353_(_007786_, _031308_, _031309_);
  or g_122354_(_031304_, _031309_, _031310_);
  or g_122355_(_007850_, _031303_, _031311_);
  xor g_122356_(_007785_, _031308_, _031312_);
  xor g_122357_(_007851_, _031303_, _031313_);
  or g_122358_(_031312_, _031313_, _031314_);
  or g_122359_(_007737_, _031253_, _031315_);
  and g_122360_(_031201_, _031253_, _031317_);
  not g_122361_(_031317_, _031318_);
  and g_122362_(_031315_, _031318_, _031319_);
  or g_122363_(_007863_, _031319_, _031320_);
  or g_122364_(_007726_, _031253_, _031321_);
  and g_122365_(_031215_, _031253_, _031322_);
  not g_122366_(_031322_, _031323_);
  and g_122367_(_031321_, _031323_, _031324_);
  or g_122368_(_007836_, _031324_, _031325_);
  and g_122369_(_031320_, _031325_, _031326_);
  and g_122370_(_007863_, _031319_, _031328_);
  xor g_122371_(_007836_, _031324_, _031329_);
  xor g_122372_(_007863_, _031319_, _031330_);
  and g_122373_(_031329_, _031330_, _031331_);
  not g_122374_(_031331_, _031332_);
  or g_122375_(_031314_, _031332_, _031333_);
  or g_122376_(_031300_, _031333_, _031334_);
  or g_122377_(_007616_, _031253_, _031335_);
  not g_122378_(_031335_, _031336_);
  and g_122379_(_031165_, _031253_, _031337_);
  not g_122380_(_031337_, _031339_);
  and g_122381_(_031335_, _031339_, _031340_);
  or g_122382_(_031336_, _031337_, _031341_);
  or g_122383_(_007924_, _031340_, _031342_);
  and g_122384_(_007924_, _031340_, _031343_);
  xor g_122385_(_007923_, _031340_, _031344_);
  and g_122386_(_031160_, _031253_, _031345_);
  and g_122387_(_052354_, _031254_, _031346_);
  or g_122388_(_031345_, _031346_, _031347_);
  or g_122389_(_052549_, _031347_, _031348_);
  xor g_122390_(_052548_, _031347_, _031350_);
  or g_122391_(_031344_, _031350_, _031351_);
  or g_122392_(_053522_, _031253_, _031352_);
  or g_122393_(_031172_, _031254_, _031353_);
  and g_122394_(_031352_, _031353_, _031354_);
  and g_122395_(out[353], _031354_, _031355_);
  not g_122396_(_031355_, _031356_);
  and g_122397_(out[352], _031257_, _031357_);
  xor g_122398_(_053621_, _031354_, _031358_);
  or g_122399_(_031357_, _031358_, _031359_);
  and g_122400_(_031356_, _031359_, _031361_);
  or g_122401_(_031351_, _031361_, _031362_);
  or g_122402_(_031343_, _031348_, _031363_);
  and g_122403_(_031342_, _031363_, _031364_);
  and g_122404_(_031362_, _031364_, _031365_);
  or g_122405_(_031334_, _031365_, _031366_);
  or g_122406_(_031314_, _031328_, _031367_);
  or g_122407_(_031326_, _031367_, _031368_);
  and g_122408_(_031310_, _031311_, _031369_);
  not g_122409_(_031369_, _031370_);
  and g_122410_(_031368_, _031370_, _031372_);
  or g_122411_(_031300_, _031372_, _031373_);
  or g_122412_(_031271_, _031275_, _031374_);
  or g_122413_(_031293_, _031296_, _031375_);
  or g_122414_(_031277_, _031375_, _031376_);
  and g_122415_(_031374_, _031376_, _031377_);
  and g_122416_(_031373_, _031377_, _031378_);
  and g_122417_(_031366_, _031378_, _031379_);
  or g_122418_(out[352], _031257_, _031380_);
  or g_122419_(_031351_, _031359_, _031381_);
  or g_122420_(_031334_, _031381_, _031383_);
  not g_122421_(_031383_, _031384_);
  and g_122422_(_031380_, _031384_, _031385_);
  or g_122423_(_031379_, _031385_, _031386_);
  not g_122424_(_031386_, _031387_);
  and g_122425_(_031257_, _031386_, _031388_);
  not g_122426_(_031388_, _031389_);
  or g_122427_(out[352], _031386_, _031390_);
  not g_122428_(_031390_, _031391_);
  and g_122429_(_031389_, _031390_, _031392_);
  or g_122430_(_031388_, _031391_, _031394_);
  and g_122431_(_031258_, _031262_, _031395_);
  or g_122432_(_031259_, _031263_, _031396_);
  or g_122433_(out[378], _008004_, _031397_);
  xor g_122434_(out[379], _031397_, _031398_);
  xor g_122435_(_004630_, _031397_, _031399_);
  and g_122436_(_031395_, _031399_, _031400_);
  or g_122437_(_031396_, _031398_, _031401_);
  xor g_122438_(out[378], _008004_, _031402_);
  xor g_122439_(_004652_, _008004_, _031403_);
  and g_122440_(_031265_, _031387_, _031405_);
  or g_122441_(_031266_, _031386_, _031406_);
  and g_122442_(_031269_, _031386_, _031407_);
  not g_122443_(_031407_, _031408_);
  and g_122444_(_031406_, _031408_, _031409_);
  or g_122445_(_031405_, _031407_, _031410_);
  and g_122446_(_031402_, _031409_, _031411_);
  or g_122447_(_031403_, _031410_, _031412_);
  and g_122448_(_031401_, _031412_, _031413_);
  or g_122449_(_031400_, _031411_, _031414_);
  and g_122450_(_031396_, _031398_, _031416_);
  or g_122451_(_031395_, _031399_, _031417_);
  and g_122452_(_031403_, _031410_, _031418_);
  or g_122453_(_031402_, _031409_, _031419_);
  and g_122454_(_031417_, _031419_, _031420_);
  or g_122455_(_031416_, _031418_, _031421_);
  and g_122456_(_031413_, _031420_, _031422_);
  or g_122457_(_031414_, _031421_, _031423_);
  and g_122458_(_007813_, _031387_, _031424_);
  and g_122459_(_031284_, _031386_, _031425_);
  or g_122460_(_031424_, _031425_, _031427_);
  and g_122461_(_008024_, _031427_, _031428_);
  not g_122462_(_031428_, _031429_);
  and g_122463_(_007800_, _031387_, _031430_);
  and g_122464_(_031291_, _031386_, _031431_);
  or g_122465_(_031430_, _031431_, _031432_);
  and g_122466_(_008006_, _031432_, _031433_);
  not g_122467_(_031433_, _031434_);
  and g_122468_(_031429_, _031434_, _031435_);
  or g_122469_(_031428_, _031433_, _031436_);
  or g_122470_(_008006_, _031432_, _031438_);
  or g_122471_(_008024_, _031427_, _031439_);
  and g_122472_(_031438_, _031439_, _031440_);
  not g_122473_(_031440_, _031441_);
  and g_122474_(_031435_, _031440_, _031442_);
  or g_122475_(_031436_, _031441_, _031443_);
  and g_122476_(_031422_, _031442_, _031444_);
  or g_122477_(_031423_, _031443_, _031445_);
  and g_122478_(_031308_, _031386_, _031446_);
  not g_122479_(_031446_, _031447_);
  or g_122480_(_007786_, _031386_, _031449_);
  not g_122481_(_031449_, _031450_);
  or g_122482_(_031446_, _031450_, _031451_);
  and g_122483_(_031447_, _031449_, _031452_);
  and g_122484_(_008046_, _031451_, _031453_);
  or g_122485_(_008045_, _031452_, _031454_);
  or g_122486_(_007850_, _031386_, _031455_);
  not g_122487_(_031455_, _031456_);
  and g_122488_(_031303_, _031386_, _031457_);
  not g_122489_(_031457_, _031458_);
  and g_122490_(_031455_, _031458_, _031460_);
  or g_122491_(_031456_, _031457_, _031461_);
  and g_122492_(_008053_, _031461_, _031462_);
  or g_122493_(_008054_, _031460_, _031463_);
  and g_122494_(_008054_, _031460_, _031464_);
  or g_122495_(_008053_, _031461_, _031465_);
  xor g_122496_(_008046_, _031451_, _031466_);
  xor g_122497_(_008045_, _031451_, _031467_);
  and g_122498_(_031463_, _031465_, _031468_);
  or g_122499_(_031462_, _031464_, _031469_);
  and g_122500_(_031466_, _031468_, _031471_);
  or g_122501_(_031467_, _031469_, _031472_);
  and g_122502_(_031319_, _031386_, _031473_);
  not g_122503_(_031473_, _031474_);
  or g_122504_(_007863_, _031386_, _031475_);
  and g_122505_(_031474_, _031475_, _031476_);
  and g_122506_(_008089_, _031476_, _031477_);
  and g_122507_(_031324_, _031386_, _031478_);
  not g_122508_(_031478_, _031479_);
  or g_122509_(_007836_, _031386_, _031480_);
  and g_122510_(_031479_, _031480_, _031482_);
  and g_122511_(_008078_, _031482_, _031483_);
  or g_122512_(_031477_, _031483_, _031484_);
  or g_122513_(_008089_, _031476_, _031485_);
  xor g_122514_(_008089_, _031476_, _031486_);
  xor g_122515_(_008088_, _031476_, _031487_);
  xor g_122516_(_008078_, _031482_, _031488_);
  xor g_122517_(_008077_, _031482_, _031489_);
  and g_122518_(_031486_, _031488_, _031490_);
  or g_122519_(_031487_, _031489_, _031491_);
  and g_122520_(_031471_, _031490_, _031493_);
  or g_122521_(_031472_, _031491_, _031494_);
  and g_122522_(_031444_, _031493_, _031495_);
  or g_122523_(_031445_, _031494_, _031496_);
  and g_122524_(_031354_, _031386_, _031497_);
  not g_122525_(_031497_, _031498_);
  or g_122526_(out[353], _031386_, _031499_);
  not g_122527_(_031499_, _031500_);
  or g_122528_(_031497_, _031500_, _031501_);
  and g_122529_(_031498_, _031499_, _031502_);
  and g_122530_(out[368], _031394_, _031504_);
  or g_122531_(_004641_, _031392_, _031505_);
  and g_122532_(out[369], _031501_, _031506_);
  or g_122533_(_053720_, _031502_, _031507_);
  xor g_122534_(out[369], _031501_, _031508_);
  xor g_122535_(_053720_, _031501_, _031509_);
  and g_122536_(_031505_, _031508_, _031510_);
  or g_122537_(_031504_, _031509_, _031511_);
  and g_122538_(_052548_, _031387_, _031512_);
  and g_122539_(_031347_, _031386_, _031513_);
  or g_122540_(_031512_, _031513_, _031515_);
  or g_122541_(_052743_, _031515_, _031516_);
  not g_122542_(_031516_, _031517_);
  and g_122543_(_007924_, _031387_, _031518_);
  and g_122544_(_031341_, _031386_, _031519_);
  or g_122545_(_031518_, _031519_, _031520_);
  not g_122546_(_031520_, _031521_);
  and g_122547_(_008112_, _031521_, _031522_);
  or g_122548_(_008111_, _031520_, _031523_);
  xor g_122549_(_052743_, _031515_, _031524_);
  xor g_122550_(_052742_, _031515_, _031526_);
  and g_122551_(_031523_, _031524_, _031527_);
  or g_122552_(_031522_, _031526_, _031528_);
  or g_122553_(out[368], _031394_, _031529_);
  not g_122554_(_031529_, _031530_);
  and g_122555_(_008111_, _031520_, _031531_);
  or g_122556_(_008112_, _031521_, _031532_);
  or g_122557_(_031530_, _031531_, _031533_);
  or g_122558_(_031511_, _031533_, _031534_);
  not g_122559_(_031534_, _031535_);
  and g_122560_(_031527_, _031535_, _031537_);
  or g_122561_(_031528_, _031534_, _031538_);
  and g_122562_(_031495_, _031537_, _031539_);
  or g_122563_(_031496_, _031538_, _031540_);
  and g_122564_(_031516_, _031532_, _031541_);
  or g_122565_(_031517_, _031531_, _031542_);
  and g_122566_(_031523_, _031542_, _031543_);
  or g_122567_(_031522_, _031541_, _031544_);
  and g_122568_(_031507_, _031511_, _031545_);
  or g_122569_(_031506_, _031510_, _031546_);
  and g_122570_(_031527_, _031546_, _031548_);
  or g_122571_(_031528_, _031545_, _031549_);
  and g_122572_(_031544_, _031549_, _031550_);
  or g_122573_(_031543_, _031548_, _031551_);
  and g_122574_(_031493_, _031551_, _031552_);
  or g_122575_(_031494_, _031550_, _031553_);
  and g_122576_(_031484_, _031485_, _031554_);
  not g_122577_(_031554_, _031555_);
  and g_122578_(_031471_, _031554_, _031556_);
  or g_122579_(_031472_, _031555_, _031557_);
  and g_122580_(_031453_, _031465_, _031559_);
  or g_122581_(_031454_, _031464_, _031560_);
  and g_122582_(_031463_, _031560_, _031561_);
  or g_122583_(_031462_, _031559_, _031562_);
  and g_122584_(_031557_, _031561_, _031563_);
  or g_122585_(_031556_, _031562_, _031564_);
  and g_122586_(_031553_, _031563_, _031565_);
  or g_122587_(_031552_, _031564_, _031566_);
  and g_122588_(_031444_, _031566_, _031567_);
  or g_122589_(_031445_, _031565_, _031568_);
  and g_122590_(_031414_, _031417_, _031570_);
  or g_122591_(_031413_, _031416_, _031571_);
  and g_122592_(_031436_, _031438_, _031572_);
  and g_122593_(_031422_, _031572_, _031573_);
  not g_122594_(_031573_, _031574_);
  and g_122595_(_031571_, _031574_, _031575_);
  or g_122596_(_031570_, _031573_, _031576_);
  and g_122597_(_031568_, _031575_, _031577_);
  or g_122598_(_031567_, _031576_, _031578_);
  and g_122599_(_031540_, _031578_, _031579_);
  or g_122600_(_031539_, _031577_, _031581_);
  and g_122601_(_031394_, _031581_, _031582_);
  and g_122602_(_004641_, _031579_, _031583_);
  or g_122603_(_031582_, _031583_, _031584_);
  and g_122604_(_031395_, _031398_, _031585_);
  or g_122605_(_031396_, _031399_, _031586_);
  or g_122606_(out[394], _008228_, _031587_);
  xor g_122607_(out[395], _031587_, _031588_);
  xor g_122608_(_004663_, _031587_, _031589_);
  and g_122609_(_031585_, _031589_, _031590_);
  or g_122610_(_031586_, _031588_, _031592_);
  xor g_122611_(out[394], _008228_, _031593_);
  xor g_122612_(_004685_, _008228_, _031594_);
  and g_122613_(_031402_, _031579_, _031595_);
  or g_122614_(_031403_, _031581_, _031596_);
  and g_122615_(_031410_, _031581_, _031597_);
  or g_122616_(_031409_, _031579_, _031598_);
  and g_122617_(_031596_, _031598_, _031599_);
  or g_122618_(_031595_, _031597_, _031600_);
  and g_122619_(_031593_, _031599_, _031601_);
  or g_122620_(_031594_, _031600_, _031603_);
  and g_122621_(_031592_, _031603_, _031604_);
  or g_122622_(_031590_, _031601_, _031605_);
  and g_122623_(_031586_, _031588_, _031606_);
  or g_122624_(_031585_, _031589_, _031607_);
  and g_122625_(_031594_, _031600_, _031608_);
  or g_122626_(_031593_, _031599_, _031609_);
  and g_122627_(_031607_, _031609_, _031610_);
  or g_122628_(_031606_, _031608_, _031611_);
  and g_122629_(_031604_, _031610_, _031612_);
  or g_122630_(_031605_, _031611_, _031614_);
  or g_122631_(_008024_, _031581_, _031615_);
  not g_122632_(_031615_, _031616_);
  and g_122633_(_031427_, _031581_, _031617_);
  not g_122634_(_031617_, _031618_);
  and g_122635_(_031615_, _031618_, _031619_);
  or g_122636_(_031616_, _031617_, _031620_);
  and g_122637_(_008222_, _031620_, _031621_);
  or g_122638_(_008221_, _031619_, _031622_);
  or g_122639_(_008006_, _031581_, _031623_);
  not g_122640_(_031623_, _031625_);
  and g_122641_(_031432_, _031581_, _031626_);
  not g_122642_(_031626_, _031627_);
  and g_122643_(_031623_, _031627_, _031628_);
  or g_122644_(_031625_, _031626_, _031629_);
  and g_122645_(_008230_, _031629_, _031630_);
  or g_122646_(_008229_, _031628_, _031631_);
  and g_122647_(_031622_, _031631_, _031632_);
  or g_122648_(_031621_, _031630_, _031633_);
  and g_122649_(_008221_, _031619_, _031634_);
  or g_122650_(_008222_, _031620_, _031636_);
  and g_122651_(_008229_, _031628_, _031637_);
  or g_122652_(_008230_, _031629_, _031638_);
  and g_122653_(_031636_, _031638_, _031639_);
  or g_122654_(_031634_, _031637_, _031640_);
  and g_122655_(_031632_, _031639_, _031641_);
  or g_122656_(_031633_, _031640_, _031642_);
  and g_122657_(_031612_, _031641_, _031643_);
  or g_122658_(_031614_, _031642_, _031644_);
  and g_122659_(_008054_, _031579_, _031645_);
  or g_122660_(_008053_, _031581_, _031647_);
  and g_122661_(_031461_, _031581_, _031648_);
  or g_122662_(_031460_, _031579_, _031649_);
  and g_122663_(_031647_, _031649_, _031650_);
  or g_122664_(_031645_, _031648_, _031651_);
  and g_122665_(_008251_, _031651_, _031652_);
  or g_122666_(_008252_, _031650_, _031653_);
  and g_122667_(_008046_, _031579_, _031654_);
  or g_122668_(_008045_, _031581_, _031655_);
  and g_122669_(_031452_, _031581_, _031656_);
  or g_122670_(_031451_, _031579_, _031658_);
  and g_122671_(_031655_, _031658_, _031659_);
  or g_122672_(_031654_, _031656_, _031660_);
  or g_122673_(_008262_, _031660_, _031661_);
  not g_122674_(_031661_, _031662_);
  and g_122675_(_031653_, _031661_, _031663_);
  or g_122676_(_031652_, _031662_, _031664_);
  or g_122677_(_008089_, _031581_, _031665_);
  not g_122678_(_031665_, _031666_);
  and g_122679_(_031476_, _031581_, _031667_);
  not g_122680_(_031667_, _031669_);
  and g_122681_(_031665_, _031669_, _031670_);
  or g_122682_(_031666_, _031667_, _031671_);
  and g_122683_(_008295_, _031670_, _031672_);
  or g_122684_(_008296_, _031671_, _031673_);
  and g_122685_(_008252_, _031650_, _031674_);
  or g_122686_(_008251_, _031651_, _031675_);
  and g_122687_(_008262_, _031660_, _031676_);
  or g_122688_(_008263_, _031659_, _031677_);
  and g_122689_(_031675_, _031677_, _031678_);
  or g_122690_(_031674_, _031676_, _031680_);
  and g_122691_(_031673_, _031678_, _031681_);
  or g_122692_(_031672_, _031680_, _031682_);
  and g_122693_(_031663_, _031681_, _031683_);
  or g_122694_(_031664_, _031682_, _031684_);
  and g_122695_(_008296_, _031671_, _031685_);
  or g_122696_(_008295_, _031670_, _031686_);
  or g_122697_(_008078_, _031581_, _031687_);
  not g_122698_(_031687_, _031688_);
  and g_122699_(_031482_, _031581_, _031689_);
  not g_122700_(_031689_, _031691_);
  and g_122701_(_031687_, _031691_, _031692_);
  or g_122702_(_031688_, _031689_, _031693_);
  and g_122703_(_008285_, _031693_, _031694_);
  or g_122704_(_008284_, _031692_, _031695_);
  and g_122705_(_031686_, _031695_, _031696_);
  or g_122706_(_031685_, _031694_, _031697_);
  or g_122707_(_008285_, _031693_, _031698_);
  not g_122708_(_031698_, _031699_);
  and g_122709_(_031696_, _031698_, _031700_);
  or g_122710_(_031697_, _031699_, _031702_);
  and g_122711_(_031683_, _031700_, _031703_);
  or g_122712_(_031684_, _031702_, _031704_);
  and g_122713_(_031643_, _031703_, _031705_);
  or g_122714_(_031644_, _031704_, _031706_);
  and g_122715_(_008112_, _031579_, _031707_);
  and g_122716_(_031520_, _031581_, _031708_);
  or g_122717_(_031707_, _031708_, _031709_);
  not g_122718_(_031709_, _031710_);
  and g_122719_(_008322_, _031710_, _031711_);
  and g_122720_(_031515_, _031581_, _031713_);
  and g_122721_(_052742_, _031579_, _031714_);
  or g_122722_(_031713_, _031714_, _031715_);
  or g_122723_(_052923_, _031715_, _031716_);
  or g_122724_(_008322_, _031710_, _031717_);
  xor g_122725_(_008321_, _031709_, _031718_);
  xor g_122726_(_008322_, _031709_, _031719_);
  xor g_122727_(_052923_, _031715_, _031720_);
  xor g_122728_(_052922_, _031715_, _031721_);
  and g_122729_(_031705_, _031720_, _031722_);
  or g_122730_(_031706_, _031721_, _031724_);
  and g_122731_(_031718_, _031722_, _031725_);
  or g_122732_(_031719_, _031724_, _031726_);
  or g_122733_(_053720_, _031581_, _031727_);
  or g_122734_(_031501_, _031579_, _031728_);
  and g_122735_(_031727_, _031728_, _031729_);
  and g_122736_(out[385], _031729_, _031730_);
  not g_122737_(_031730_, _031731_);
  and g_122738_(out[384], _031584_, _031732_);
  not g_122739_(_031732_, _031733_);
  xor g_122740_(out[385], _031729_, _031735_);
  xor g_122741_(_053819_, _031729_, _031736_);
  and g_122742_(_031733_, _031735_, _031737_);
  or g_122743_(_031732_, _031736_, _031738_);
  and g_122744_(_031731_, _031738_, _031739_);
  or g_122745_(_031730_, _031737_, _031740_);
  and g_122746_(_031725_, _031740_, _031741_);
  or g_122747_(_031726_, _031739_, _031742_);
  or g_122748_(_031663_, _031674_, _031743_);
  or g_122749_(_031684_, _031696_, _031744_);
  and g_122750_(_031743_, _031744_, _031746_);
  not g_122751_(_031746_, _031747_);
  and g_122752_(_031643_, _031747_, _031748_);
  or g_122753_(_031644_, _031746_, _031749_);
  or g_122754_(_031711_, _031716_, _031750_);
  and g_122755_(_031717_, _031750_, _031751_);
  or g_122756_(_031706_, _031751_, _031752_);
  not g_122757_(_031752_, _031753_);
  and g_122758_(_031605_, _031607_, _031754_);
  or g_122759_(_031604_, _031606_, _031755_);
  and g_122760_(_031612_, _031633_, _031757_);
  and g_122761_(_031638_, _031757_, _031758_);
  not g_122762_(_031758_, _031759_);
  and g_122763_(_031755_, _031759_, _031760_);
  or g_122764_(_031754_, _031758_, _031761_);
  and g_122765_(_031752_, _031760_, _031762_);
  or g_122766_(_031753_, _031761_, _031763_);
  and g_122767_(_031749_, _031762_, _031764_);
  or g_122768_(_031741_, _031763_, _031765_);
  and g_122769_(_031742_, _031764_, _031766_);
  or g_122770_(_031748_, _031765_, _031768_);
  or g_122771_(out[384], _031584_, _031769_);
  not g_122772_(_031769_, _031770_);
  or g_122773_(_031726_, _031738_, _031771_);
  not g_122774_(_031771_, _031772_);
  and g_122775_(_031769_, _031772_, _031773_);
  or g_122776_(_031770_, _031771_, _031774_);
  and g_122777_(_031768_, _031774_, _031775_);
  or g_122778_(_031766_, _031773_, _031776_);
  and g_122779_(_031584_, _031776_, _031777_);
  not g_122780_(_031777_, _031779_);
  or g_122781_(out[384], _031776_, _031780_);
  not g_122782_(_031780_, _031781_);
  and g_122783_(_031779_, _031780_, _031782_);
  or g_122784_(_031777_, _031781_, _031783_);
  or g_122785_(_008321_, _031776_, _031784_);
  not g_122786_(_031784_, _031785_);
  and g_122787_(_031709_, _031776_, _031786_);
  not g_122788_(_031786_, _031787_);
  and g_122789_(_031784_, _031787_, _031788_);
  or g_122790_(_031785_, _031786_, _031790_);
  and g_122791_(_008420_, _031788_, _031791_);
  or g_122792_(_008419_, _031790_, _031792_);
  or g_122793_(_052923_, _031776_, _031793_);
  not g_122794_(_031793_, _031794_);
  and g_122795_(_031715_, _031776_, _031795_);
  not g_122796_(_031795_, _031796_);
  and g_122797_(_031793_, _031796_, _031797_);
  or g_122798_(_031794_, _031795_, _031798_);
  and g_122799_(_053010_, _031797_, _031799_);
  or g_122800_(_053011_, _031798_, _031801_);
  and g_122801_(_008419_, _031790_, _031802_);
  or g_122802_(_008420_, _031788_, _031803_);
  and g_122803_(_031801_, _031803_, _031804_);
  or g_122804_(_031799_, _031802_, _031805_);
  or g_122805_(_053819_, _031776_, _031806_);
  or g_122806_(_031729_, _031775_, _031807_);
  and g_122807_(_031806_, _031807_, _031808_);
  and g_122808_(out[401], _031808_, _031809_);
  not g_122809_(_031809_, _031810_);
  and g_122810_(out[400], _031783_, _031812_);
  or g_122811_(_004707_, _031782_, _031813_);
  xor g_122812_(out[401], _031808_, _031814_);
  xor g_122813_(_053918_, _031808_, _031815_);
  and g_122814_(_031813_, _031814_, _031816_);
  or g_122815_(_031812_, _031815_, _031817_);
  and g_122816_(_031810_, _031817_, _031818_);
  or g_122817_(_031809_, _031816_, _031819_);
  xor g_122818_(_053010_, _031797_, _031820_);
  xor g_122819_(_053011_, _031797_, _031821_);
  or g_122820_(_031791_, _031804_, _031823_);
  and g_122821_(_031792_, _031805_, _031824_);
  and g_122822_(_031792_, _031820_, _031825_);
  or g_122823_(_031791_, _031821_, _031826_);
  and g_122824_(_031819_, _031825_, _031827_);
  or g_122825_(_031818_, _031826_, _031828_);
  or g_122826_(_031824_, _031827_, _031829_);
  and g_122827_(_031823_, _031828_, _031830_);
  and g_122828_(_008252_, _031775_, _031831_);
  or g_122829_(_008251_, _031776_, _031832_);
  and g_122830_(_031651_, _031776_, _031834_);
  or g_122831_(_031650_, _031775_, _031835_);
  and g_122832_(_031832_, _031835_, _031836_);
  or g_122833_(_031831_, _031834_, _031837_);
  and g_122834_(_008511_, _031837_, _031838_);
  or g_122835_(_008512_, _031836_, _031839_);
  and g_122836_(_008512_, _031836_, _031840_);
  or g_122837_(_008511_, _031837_, _031841_);
  and g_122838_(_031839_, _031841_, _031842_);
  or g_122839_(_031838_, _031840_, _031843_);
  or g_122840_(_008262_, _031776_, _031845_);
  not g_122841_(_031845_, _031846_);
  and g_122842_(_031660_, _031776_, _031847_);
  not g_122843_(_031847_, _031848_);
  and g_122844_(_031845_, _031848_, _031849_);
  or g_122845_(_031846_, _031847_, _031850_);
  and g_122846_(_008506_, _031849_, _031851_);
  or g_122847_(_008505_, _031850_, _031852_);
  or g_122848_(_008296_, _031776_, _031853_);
  not g_122849_(_031853_, _031854_);
  and g_122850_(_031671_, _031776_, _031856_);
  not g_122851_(_031856_, _031857_);
  and g_122852_(_031853_, _031857_, _031858_);
  or g_122853_(_031854_, _031856_, _031859_);
  and g_122854_(_008540_, _031858_, _031860_);
  or g_122855_(_008541_, _031859_, _031861_);
  xor g_122856_(_008506_, _031849_, _031862_);
  xor g_122857_(_008505_, _031849_, _031863_);
  and g_122858_(_031842_, _031862_, _031864_);
  or g_122859_(_031843_, _031863_, _031865_);
  and g_122860_(_031861_, _031864_, _031867_);
  or g_122861_(_031860_, _031865_, _031868_);
  and g_122862_(_031585_, _031588_, _031869_);
  or g_122863_(_031586_, _031589_, _031870_);
  or g_122864_(out[410], _008479_, _031871_);
  xor g_122865_(out[411], _031871_, _031872_);
  xor g_122866_(_004696_, _031871_, _031873_);
  and g_122867_(_031869_, _031873_, _031874_);
  or g_122868_(_031870_, _031872_, _031875_);
  xor g_122869_(out[410], _008479_, _031876_);
  xor g_122870_(_004718_, _008479_, _031878_);
  and g_122871_(_031593_, _031775_, _031879_);
  or g_122872_(_031594_, _031776_, _031880_);
  and g_122873_(_031600_, _031776_, _031881_);
  or g_122874_(_031599_, _031775_, _031882_);
  and g_122875_(_031880_, _031882_, _031883_);
  or g_122876_(_031879_, _031881_, _031884_);
  and g_122877_(_031876_, _031883_, _031885_);
  or g_122878_(_031878_, _031884_, _031886_);
  and g_122879_(_031875_, _031886_, _031887_);
  or g_122880_(_031874_, _031885_, _031889_);
  and g_122881_(_031878_, _031884_, _031890_);
  or g_122882_(_031876_, _031883_, _031891_);
  and g_122883_(_031870_, _031872_, _031892_);
  or g_122884_(_031869_, _031873_, _031893_);
  and g_122885_(_031891_, _031893_, _031894_);
  or g_122886_(_031890_, _031892_, _031895_);
  and g_122887_(_031887_, _031894_, _031896_);
  or g_122888_(_031889_, _031895_, _031897_);
  or g_122889_(_008222_, _031776_, _031898_);
  not g_122890_(_031898_, _031900_);
  and g_122891_(_031620_, _031776_, _031901_);
  not g_122892_(_031901_, _031902_);
  and g_122893_(_031898_, _031902_, _031903_);
  or g_122894_(_031900_, _031901_, _031904_);
  and g_122895_(_008470_, _031904_, _031905_);
  or g_122896_(_008468_, _031903_, _031906_);
  or g_122897_(_008230_, _031776_, _031907_);
  not g_122898_(_031907_, _031908_);
  and g_122899_(_031629_, _031776_, _031909_);
  not g_122900_(_031909_, _031911_);
  and g_122901_(_031907_, _031911_, _031912_);
  or g_122902_(_031908_, _031909_, _031913_);
  and g_122903_(_008482_, _031913_, _031914_);
  or g_122904_(_008481_, _031912_, _031915_);
  and g_122905_(_031906_, _031915_, _031916_);
  or g_122906_(_031905_, _031914_, _031917_);
  and g_122907_(_008481_, _031912_, _031918_);
  or g_122908_(_008482_, _031913_, _031919_);
  and g_122909_(_008468_, _031903_, _031920_);
  or g_122910_(_008470_, _031904_, _031922_);
  and g_122911_(_031919_, _031922_, _031923_);
  or g_122912_(_031918_, _031920_, _031924_);
  and g_122913_(_031916_, _031923_, _031925_);
  or g_122914_(_031917_, _031924_, _031926_);
  and g_122915_(_031896_, _031925_, _031927_);
  or g_122916_(_031897_, _031926_, _031928_);
  or g_122917_(_008285_, _031776_, _031929_);
  not g_122918_(_031929_, _031930_);
  and g_122919_(_031693_, _031776_, _031931_);
  not g_122920_(_031931_, _031933_);
  and g_122921_(_031929_, _031933_, _031934_);
  or g_122922_(_031930_, _031931_, _031935_);
  and g_122923_(_008530_, _031935_, _031936_);
  or g_122924_(_008529_, _031934_, _031937_);
  and g_122925_(_008541_, _031859_, _031938_);
  or g_122926_(_008540_, _031858_, _031939_);
  and g_122927_(_031937_, _031939_, _031940_);
  or g_122928_(_031936_, _031938_, _031941_);
  and g_122929_(_008529_, _031934_, _031942_);
  or g_122930_(_008530_, _031935_, _031944_);
  and g_122931_(_031940_, _031944_, _031945_);
  or g_122932_(_031941_, _031942_, _031946_);
  and g_122933_(_031867_, _031945_, _031947_);
  or g_122934_(_031868_, _031946_, _031948_);
  and g_122935_(_031927_, _031947_, _031949_);
  or g_122936_(_031928_, _031948_, _031950_);
  and g_122937_(_031829_, _031949_, _031951_);
  or g_122938_(_031830_, _031950_, _031952_);
  and g_122939_(_031867_, _031941_, _031953_);
  or g_122940_(_031868_, _031940_, _031955_);
  and g_122941_(_031841_, _031851_, _031956_);
  or g_122942_(_031840_, _031852_, _031957_);
  and g_122943_(_031839_, _031957_, _031958_);
  or g_122944_(_031838_, _031956_, _031959_);
  and g_122945_(_031955_, _031958_, _031960_);
  or g_122946_(_031953_, _031959_, _031961_);
  and g_122947_(_031927_, _031961_, _031962_);
  or g_122948_(_031928_, _031960_, _031963_);
  and g_122949_(_031889_, _031893_, _031964_);
  or g_122950_(_031887_, _031892_, _031966_);
  and g_122951_(_031896_, _031917_, _031967_);
  or g_122952_(_031897_, _031916_, _031968_);
  and g_122953_(_031919_, _031967_, _031969_);
  or g_122954_(_031918_, _031968_, _031970_);
  and g_122955_(_031966_, _031970_, _031971_);
  or g_122956_(_031964_, _031969_, _031972_);
  and g_122957_(_031952_, _031971_, _031973_);
  or g_122958_(_031951_, _031972_, _031974_);
  and g_122959_(_031963_, _031973_, _031975_);
  or g_122960_(_031962_, _031974_, _031977_);
  and g_122961_(_004707_, _031782_, _031978_);
  or g_122962_(out[400], _031783_, _031979_);
  and g_122963_(_031803_, _031979_, _031980_);
  or g_122964_(_031802_, _031978_, _031981_);
  and g_122965_(_031825_, _031980_, _031982_);
  or g_122966_(_031826_, _031981_, _031983_);
  and g_122967_(_031816_, _031982_, _031984_);
  or g_122968_(_031817_, _031983_, _031985_);
  and g_122969_(_031949_, _031984_, _031986_);
  or g_122970_(_031950_, _031985_, _031988_);
  and g_122971_(_031977_, _031988_, _031989_);
  or g_122972_(_031975_, _031986_, _031990_);
  and g_122973_(_031783_, _031990_, _031991_);
  and g_122974_(_004707_, _031989_, _031992_);
  or g_122975_(_031991_, _031992_, _031993_);
  and g_122976_(_008420_, _031989_, _031994_);
  and g_122977_(_031790_, _031990_, _031995_);
  or g_122978_(_031994_, _031995_, _031996_);
  not g_122979_(_031996_, _031997_);
  and g_122980_(_008728_, _031996_, _031999_);
  or g_122981_(_008729_, _031997_, _032000_);
  and g_122982_(_008729_, _031997_, _032001_);
  or g_122983_(_008728_, _031996_, _032002_);
  and g_122984_(_032000_, _032002_, _032003_);
  or g_122985_(_031999_, _032001_, _032004_);
  and g_122986_(_031798_, _031990_, _032005_);
  and g_122987_(_053010_, _031989_, _032006_);
  or g_122988_(_032005_, _032006_, _032007_);
  not g_122989_(_032007_, _032008_);
  and g_122990_(_053271_, _032008_, _032010_);
  or g_122991_(_053272_, _032007_, _032011_);
  xor g_122992_(_053272_, _032007_, _032012_);
  xor g_122993_(_053271_, _032007_, _032013_);
  and g_122994_(_032003_, _032012_, _032014_);
  or g_122995_(_032004_, _032013_, _032015_);
  and g_122996_(out[401], _031989_, _032016_);
  or g_122997_(_053918_, _031990_, _032017_);
  or g_122998_(_031808_, _031989_, _032018_);
  not g_122999_(_032018_, _032019_);
  and g_123000_(_032017_, _032018_, _032021_);
  or g_123001_(_032016_, _032019_, _032022_);
  and g_123002_(out[417], _032021_, _032023_);
  not g_123003_(_032023_, _032024_);
  and g_123004_(out[416], _031993_, _032025_);
  not g_123005_(_032025_, _032026_);
  xor g_123006_(out[417], _032021_, _032027_);
  xor g_123007_(_054017_, _032021_, _032028_);
  and g_123008_(_032026_, _032027_, _032029_);
  or g_123009_(_032025_, _032028_, _032030_);
  and g_123010_(_032024_, _032030_, _032032_);
  or g_123011_(_032023_, _032029_, _032033_);
  and g_123012_(_032014_, _032033_, _032034_);
  or g_123013_(_032015_, _032032_, _032035_);
  and g_123014_(_032000_, _032011_, _032036_);
  or g_123015_(_031999_, _032010_, _032037_);
  and g_123016_(_032002_, _032037_, _032038_);
  or g_123017_(_032001_, _032036_, _032039_);
  and g_123018_(_032035_, _032039_, _032040_);
  or g_123019_(_032034_, _032038_, _032041_);
  and g_123020_(_031869_, _031872_, _032043_);
  or g_123021_(_031870_, _031873_, _032044_);
  or g_123022_(out[426], _008626_, _032045_);
  xor g_123023_(out[427], _032045_, _032046_);
  xor g_123024_(_004729_, _032045_, _032047_);
  and g_123025_(_032043_, _032047_, _032048_);
  or g_123026_(_032044_, _032046_, _032049_);
  xor g_123027_(out[426], _008626_, _032050_);
  xor g_123028_(_004751_, _008626_, _032051_);
  and g_123029_(_031884_, _031990_, _032052_);
  or g_123030_(_031883_, _031989_, _032054_);
  and g_123031_(_031876_, _031989_, _032055_);
  or g_123032_(_031878_, _031990_, _032056_);
  and g_123033_(_032054_, _032056_, _032057_);
  or g_123034_(_032052_, _032055_, _032058_);
  and g_123035_(_032050_, _032057_, _032059_);
  or g_123036_(_032051_, _032058_, _032060_);
  and g_123037_(_032049_, _032060_, _032061_);
  or g_123038_(_032048_, _032059_, _032062_);
  and g_123039_(_032051_, _032058_, _032063_);
  and g_123040_(_032044_, _032046_, _032065_);
  or g_123041_(_032063_, _032065_, _032066_);
  not g_123042_(_032066_, _032067_);
  and g_123043_(_032061_, _032067_, _032068_);
  or g_123044_(_032062_, _032066_, _032069_);
  and g_123045_(_008468_, _031989_, _032070_);
  and g_123046_(_031904_, _031990_, _032071_);
  or g_123047_(_032070_, _032071_, _032072_);
  not g_123048_(_032072_, _032073_);
  and g_123049_(_008640_, _032072_, _032074_);
  or g_123050_(_008639_, _032073_, _032076_);
  and g_123051_(_008481_, _031989_, _032077_);
  and g_123052_(_031913_, _031990_, _032078_);
  or g_123053_(_032077_, _032078_, _032079_);
  not g_123054_(_032079_, _032080_);
  and g_123055_(_008628_, _032079_, _032081_);
  or g_123056_(_008627_, _032080_, _032082_);
  and g_123057_(_032076_, _032082_, _032083_);
  or g_123058_(_032074_, _032081_, _032084_);
  and g_123059_(_008627_, _032080_, _032085_);
  or g_123060_(_008628_, _032079_, _032087_);
  and g_123061_(_008639_, _032073_, _032088_);
  or g_123062_(_008640_, _032072_, _032089_);
  and g_123063_(_032087_, _032089_, _032090_);
  or g_123064_(_032085_, _032088_, _032091_);
  and g_123065_(_032083_, _032090_, _032092_);
  or g_123066_(_032084_, _032091_, _032093_);
  and g_123067_(_032068_, _032092_, _032094_);
  or g_123068_(_032069_, _032093_, _032095_);
  and g_123069_(_031850_, _031990_, _032096_);
  and g_123070_(_008506_, _031989_, _032098_);
  or g_123071_(_032096_, _032098_, _032099_);
  or g_123072_(_008653_, _032099_, _032100_);
  not g_123073_(_032100_, _032101_);
  xor g_123074_(_008653_, _032099_, _032102_);
  xor g_123075_(_008654_, _032099_, _032103_);
  or g_123076_(_008511_, _031990_, _032104_);
  not g_123077_(_032104_, _032105_);
  and g_123078_(_031837_, _031990_, _032106_);
  not g_123079_(_032106_, _032107_);
  and g_123080_(_032104_, _032107_, _032109_);
  or g_123081_(_032105_, _032106_, _032110_);
  and g_123082_(_008664_, _032110_, _032111_);
  or g_123083_(_008665_, _032109_, _032112_);
  and g_123084_(_008665_, _032109_, _032113_);
  or g_123085_(_008664_, _032110_, _032114_);
  and g_123086_(_032112_, _032114_, _032115_);
  or g_123087_(_032111_, _032113_, _032116_);
  and g_123088_(_032102_, _032115_, _032117_);
  or g_123089_(_032103_, _032116_, _032118_);
  or g_123090_(_008530_, _031990_, _032120_);
  not g_123091_(_032120_, _032121_);
  and g_123092_(_031935_, _031990_, _032122_);
  not g_123093_(_032122_, _032123_);
  and g_123094_(_032120_, _032123_, _032124_);
  or g_123095_(_032121_, _032122_, _032125_);
  and g_123096_(_008687_, _032125_, _032126_);
  or g_123097_(_008686_, _032124_, _032127_);
  xor g_123098_(_008686_, _032124_, _032128_);
  xor g_123099_(_008687_, _032124_, _032129_);
  and g_123100_(_031859_, _031990_, _032131_);
  not g_123101_(_032131_, _032132_);
  or g_123102_(_008541_, _031990_, _032133_);
  not g_123103_(_032133_, _032134_);
  and g_123104_(_032132_, _032133_, _032135_);
  or g_123105_(_032131_, _032134_, _032136_);
  or g_123106_(_008695_, _032136_, _032137_);
  not g_123107_(_032137_, _032138_);
  and g_123108_(_008695_, _032136_, _032139_);
  or g_123109_(_008694_, _032135_, _032140_);
  or g_123110_(_032138_, _032139_, _032142_);
  or g_123111_(_032129_, _032142_, _032143_);
  or g_123112_(_032118_, _032143_, _032144_);
  and g_123113_(_032128_, _032137_, _032145_);
  and g_123114_(_032117_, _032140_, _032146_);
  and g_123115_(_032094_, _032146_, _032147_);
  and g_123116_(_032145_, _032147_, _032148_);
  or g_123117_(_032095_, _032144_, _032149_);
  and g_123118_(_032041_, _032148_, _032150_);
  or g_123119_(_032040_, _032149_, _032151_);
  and g_123120_(_032127_, _032140_, _032153_);
  or g_123121_(_032126_, _032139_, _032154_);
  and g_123122_(_032137_, _032154_, _032155_);
  or g_123123_(_032138_, _032153_, _032156_);
  and g_123124_(_032117_, _032155_, _032157_);
  or g_123125_(_032118_, _032156_, _032158_);
  and g_123126_(_032101_, _032114_, _032159_);
  or g_123127_(_032100_, _032113_, _032160_);
  and g_123128_(_032112_, _032160_, _032161_);
  or g_123129_(_032111_, _032159_, _032162_);
  and g_123130_(_032158_, _032161_, _032164_);
  or g_123131_(_032157_, _032162_, _032165_);
  and g_123132_(_032094_, _032165_, _032166_);
  or g_123133_(_032095_, _032164_, _032167_);
  and g_123134_(_032084_, _032087_, _032168_);
  not g_123135_(_032168_, _032169_);
  and g_123136_(_032068_, _032168_, _032170_);
  or g_123137_(_032069_, _032169_, _032171_);
  or g_123138_(_032061_, _032065_, _032172_);
  not g_123139_(_032172_, _032173_);
  and g_123140_(_032171_, _032172_, _032175_);
  or g_123141_(_032170_, _032173_, _032176_);
  and g_123142_(_032167_, _032175_, _032177_);
  or g_123143_(_032166_, _032176_, _032178_);
  and g_123144_(_032151_, _032177_, _032179_);
  or g_123145_(_032150_, _032178_, _032180_);
  or g_123146_(out[416], _031993_, _032181_);
  not g_123147_(_032181_, _032182_);
  and g_123148_(_032014_, _032181_, _032183_);
  or g_123149_(_032015_, _032182_, _032184_);
  and g_123150_(_032029_, _032183_, _032186_);
  or g_123151_(_032030_, _032184_, _032187_);
  and g_123152_(_032148_, _032186_, _032188_);
  or g_123153_(_032149_, _032187_, _032189_);
  and g_123154_(_032180_, _032189_, _032190_);
  or g_123155_(_032179_, _032188_, _032191_);
  and g_123156_(_031993_, _032191_, _032192_);
  not g_123157_(_032192_, _032193_);
  or g_123158_(out[416], _032191_, _032194_);
  not g_123159_(_032194_, _032195_);
  and g_123160_(_032193_, _032194_, _032197_);
  or g_123161_(_032192_, _032195_, _032198_);
  or g_123162_(_008728_, _032191_, _032199_);
  not g_123163_(_032199_, _032200_);
  and g_123164_(_031996_, _032191_, _032201_);
  not g_123165_(_032201_, _032202_);
  and g_123166_(_032199_, _032202_, _032203_);
  or g_123167_(_032200_, _032201_, _032204_);
  and g_123168_(_008918_, _032204_, _032205_);
  or g_123169_(_008919_, _032203_, _032206_);
  and g_123170_(_008919_, _032203_, _032208_);
  or g_123171_(_008918_, _032204_, _032209_);
  and g_123172_(_032206_, _032209_, _032210_);
  or g_123173_(_032205_, _032208_, _032211_);
  and g_123174_(_032007_, _032191_, _032212_);
  and g_123175_(_053271_, _032190_, _032213_);
  or g_123176_(_032212_, _032213_, _032214_);
  not g_123177_(_032214_, _032215_);
  and g_123178_(_053387_, _032215_, _032216_);
  or g_123179_(_053388_, _032214_, _032217_);
  xor g_123180_(_053388_, _032214_, _032219_);
  xor g_123181_(_053387_, _032214_, _032220_);
  and g_123182_(_032210_, _032219_, _032221_);
  or g_123183_(_032211_, _032220_, _032222_);
  and g_123184_(out[417], _032190_, _032223_);
  and g_123185_(_032022_, _032191_, _032224_);
  or g_123186_(_032223_, _032224_, _032225_);
  or g_123187_(_054116_, _032225_, _032226_);
  not g_123188_(_032226_, _032227_);
  and g_123189_(out[432], _032198_, _032228_);
  or g_123190_(_004773_, _032197_, _032230_);
  xor g_123191_(_054116_, _032225_, _032231_);
  xor g_123192_(out[433], _032225_, _032232_);
  and g_123193_(_032230_, _032231_, _032233_);
  or g_123194_(_032228_, _032232_, _032234_);
  and g_123195_(_032226_, _032234_, _032235_);
  or g_123196_(_032227_, _032233_, _032236_);
  and g_123197_(_032221_, _032236_, _032237_);
  or g_123198_(_032222_, _032235_, _032238_);
  and g_123199_(_032209_, _032216_, _032239_);
  or g_123200_(_032208_, _032217_, _032241_);
  and g_123201_(_032206_, _032241_, _032242_);
  or g_123202_(_032205_, _032239_, _032243_);
  and g_123203_(_032238_, _032242_, _032244_);
  or g_123204_(_032237_, _032243_, _032245_);
  or g_123205_(out[442], _008853_, _032246_);
  xor g_123206_(out[442], _008853_, _032247_);
  not g_123207_(_032247_, _032248_);
  or g_123208_(_032051_, _032191_, _032249_);
  not g_123209_(_032249_, _032250_);
  and g_123210_(_032058_, _032191_, _032252_);
  not g_123211_(_032252_, _032253_);
  and g_123212_(_032249_, _032253_, _032254_);
  or g_123213_(_032250_, _032252_, _032255_);
  and g_123214_(_032247_, _032254_, _032256_);
  or g_123215_(_032248_, _032255_, _032257_);
  and g_123216_(_032248_, _032255_, _032258_);
  or g_123217_(_032247_, _032254_, _032259_);
  and g_123218_(_032043_, _032046_, _032260_);
  or g_123219_(_032044_, _032047_, _032261_);
  xor g_123220_(out[443], _032246_, _032263_);
  xor g_123221_(_004762_, _032246_, _032264_);
  and g_123222_(_032260_, _032264_, _032265_);
  or g_123223_(_032261_, _032263_, _032266_);
  and g_123224_(_032261_, _032263_, _032267_);
  or g_123225_(_032260_, _032264_, _032268_);
  and g_123226_(_032259_, _032266_, _032269_);
  or g_123227_(_032258_, _032265_, _032270_);
  and g_123228_(_032257_, _032268_, _032271_);
  or g_123229_(_032256_, _032267_, _032272_);
  and g_123230_(_032269_, _032271_, _032274_);
  or g_123231_(_032270_, _032272_, _032275_);
  or g_123232_(_008640_, _032191_, _032276_);
  not g_123233_(_032276_, _032277_);
  and g_123234_(_032072_, _032191_, _032278_);
  not g_123235_(_032278_, _032279_);
  and g_123236_(_032276_, _032279_, _032280_);
  or g_123237_(_032277_, _032278_, _032281_);
  and g_123238_(_008846_, _032281_, _032282_);
  or g_123239_(_008845_, _032280_, _032283_);
  or g_123240_(_008628_, _032191_, _032285_);
  not g_123241_(_032285_, _032286_);
  and g_123242_(_032079_, _032191_, _032287_);
  not g_123243_(_032287_, _032288_);
  and g_123244_(_032285_, _032288_, _032289_);
  or g_123245_(_032286_, _032287_, _032290_);
  and g_123246_(_008856_, _032290_, _032291_);
  or g_123247_(_008855_, _032289_, _032292_);
  and g_123248_(_032283_, _032292_, _032293_);
  or g_123249_(_032282_, _032291_, _032294_);
  and g_123250_(_008855_, _032289_, _032296_);
  or g_123251_(_008856_, _032290_, _032297_);
  and g_123252_(_008845_, _032280_, _032298_);
  or g_123253_(_008846_, _032281_, _032299_);
  and g_123254_(_032297_, _032299_, _032300_);
  or g_123255_(_032296_, _032298_, _032301_);
  and g_123256_(_032293_, _032300_, _032302_);
  or g_123257_(_032294_, _032301_, _032303_);
  and g_123258_(_032274_, _032302_, _032304_);
  or g_123259_(_032275_, _032303_, _032305_);
  and g_123260_(_008665_, _032190_, _032307_);
  and g_123261_(_032110_, _032191_, _032308_);
  or g_123262_(_032307_, _032308_, _032309_);
  and g_123263_(_008878_, _032309_, _032310_);
  or g_123264_(_008878_, _032309_, _032311_);
  xor g_123265_(_008878_, _032309_, _032312_);
  xor g_123266_(_008879_, _032309_, _032313_);
  and g_123267_(_008654_, _032190_, _032314_);
  and g_123268_(_032099_, _032191_, _032315_);
  or g_123269_(_032314_, _032315_, _032316_);
  or g_123270_(_008868_, _032316_, _032318_);
  not g_123271_(_032318_, _032319_);
  xor g_123272_(_008868_, _032316_, _032320_);
  xor g_123273_(_008869_, _032316_, _032321_);
  and g_123274_(_032312_, _032320_, _032322_);
  or g_123275_(_032313_, _032321_, _032323_);
  or g_123276_(_008687_, _032191_, _032324_);
  not g_123277_(_032324_, _032325_);
  and g_123278_(_032125_, _032191_, _032326_);
  not g_123279_(_032326_, _032327_);
  and g_123280_(_032324_, _032327_, _032329_);
  or g_123281_(_032325_, _032326_, _032330_);
  and g_123282_(_008893_, _032330_, _032331_);
  or g_123283_(_008892_, _032329_, _032332_);
  or g_123284_(_008695_, _032191_, _032333_);
  not g_123285_(_032333_, _032334_);
  and g_123286_(_032136_, _032191_, _032335_);
  not g_123287_(_032335_, _032336_);
  and g_123288_(_032333_, _032336_, _032337_);
  or g_123289_(_032334_, _032335_, _032338_);
  and g_123290_(_008900_, _032338_, _032340_);
  or g_123291_(_008899_, _032337_, _032341_);
  and g_123292_(_032332_, _032341_, _032342_);
  or g_123293_(_032331_, _032340_, _032343_);
  and g_123294_(_008899_, _032337_, _032344_);
  or g_123295_(_008900_, _032338_, _032345_);
  and g_123296_(_008892_, _032329_, _032346_);
  or g_123297_(_008893_, _032330_, _032347_);
  and g_123298_(_032345_, _032347_, _032348_);
  or g_123299_(_032344_, _032346_, _032349_);
  and g_123300_(_032342_, _032348_, _032351_);
  or g_123301_(_032343_, _032349_, _032352_);
  and g_123302_(_032322_, _032351_, _032353_);
  or g_123303_(_032323_, _032352_, _032354_);
  and g_123304_(_032304_, _032353_, _032355_);
  or g_123305_(_032305_, _032354_, _032356_);
  and g_123306_(_032245_, _032355_, _032357_);
  or g_123307_(_032244_, _032356_, _032358_);
  and g_123308_(_032322_, _032343_, _032359_);
  or g_123309_(_032323_, _032342_, _032360_);
  and g_123310_(_032345_, _032359_, _032362_);
  or g_123311_(_032344_, _032360_, _032363_);
  and g_123312_(_032311_, _032319_, _032364_);
  or g_123313_(_032310_, _032364_, _032365_);
  not g_123314_(_032365_, _032366_);
  and g_123315_(_032363_, _032366_, _032367_);
  or g_123316_(_032362_, _032365_, _032368_);
  and g_123317_(_032304_, _032368_, _032369_);
  or g_123318_(_032305_, _032367_, _032370_);
  and g_123319_(_032294_, _032297_, _032371_);
  or g_123320_(_032293_, _032296_, _032373_);
  and g_123321_(_032274_, _032371_, _032374_);
  or g_123322_(_032275_, _032373_, _032375_);
  and g_123323_(_032257_, _032266_, _032376_);
  or g_123324_(_032256_, _032265_, _032377_);
  and g_123325_(_032268_, _032377_, _032378_);
  or g_123326_(_032267_, _032376_, _032379_);
  and g_123327_(_032375_, _032379_, _032380_);
  or g_123328_(_032374_, _032378_, _032381_);
  and g_123329_(_032358_, _032380_, _032382_);
  or g_123330_(_032357_, _032381_, _032384_);
  and g_123331_(_032370_, _032382_, _032385_);
  or g_123332_(_032369_, _032384_, _032386_);
  or g_123333_(out[432], _032198_, _032387_);
  not g_123334_(_032387_, _032388_);
  or g_123335_(_032234_, _032388_, _032389_);
  not g_123336_(_032389_, _032390_);
  and g_123337_(_032355_, _032390_, _032391_);
  or g_123338_(_032356_, _032389_, _032392_);
  and g_123339_(_032221_, _032391_, _032393_);
  or g_123340_(_032222_, _032392_, _032395_);
  and g_123341_(_032386_, _032395_, _032396_);
  or g_123342_(_032385_, _032393_, _032397_);
  or g_123343_(_032197_, _032396_, _032398_);
  or g_123344_(out[432], _032397_, _032399_);
  and g_123345_(_032398_, _032399_, _032400_);
  not g_123346_(_032400_, _032401_);
  or g_123347_(out[458], _009077_, _032402_);
  xor g_123348_(out[458], _009077_, _032403_);
  not g_123349_(_032403_, _032404_);
  and g_123350_(_032247_, _032396_, _032406_);
  and g_123351_(_032255_, _032397_, _032407_);
  or g_123352_(_032406_, _032407_, _032408_);
  and g_123353_(_032260_, _032263_, _032409_);
  not g_123354_(_032409_, _032410_);
  xor g_123355_(out[459], _032402_, _032411_);
  not g_123356_(_032411_, _032412_);
  and g_123357_(_032409_, _032412_, _032413_);
  or g_123358_(_032410_, _032411_, _032414_);
  and g_123359_(_032410_, _032411_, _032415_);
  or g_123360_(_032409_, _032412_, _032417_);
  and g_123361_(_032414_, _032417_, _032418_);
  or g_123362_(_032404_, _032408_, _032419_);
  not g_123363_(_032419_, _032420_);
  xor g_123364_(_032404_, _032408_, _032421_);
  and g_123365_(_032418_, _032421_, _032422_);
  not g_123366_(_032422_, _032423_);
  and g_123367_(_008845_, _032396_, _032424_);
  or g_123368_(_008846_, _032397_, _032425_);
  and g_123369_(_032281_, _032397_, _032426_);
  or g_123370_(_032280_, _032396_, _032428_);
  and g_123371_(_032425_, _032428_, _032429_);
  or g_123372_(_032424_, _032426_, _032430_);
  and g_123373_(_009067_, _032430_, _032431_);
  or g_123374_(_009066_, _032429_, _032432_);
  and g_123375_(_008855_, _032396_, _032433_);
  or g_123376_(_008856_, _032397_, _032434_);
  and g_123377_(_032290_, _032397_, _032435_);
  or g_123378_(_032289_, _032396_, _032436_);
  and g_123379_(_032434_, _032436_, _032437_);
  or g_123380_(_032433_, _032435_, _032439_);
  and g_123381_(_009079_, _032439_, _032440_);
  or g_123382_(_009078_, _032437_, _032441_);
  and g_123383_(_032432_, _032441_, _032442_);
  or g_123384_(_032431_, _032440_, _032443_);
  and g_123385_(_009078_, _032437_, _032444_);
  or g_123386_(_009079_, _032439_, _032445_);
  and g_123387_(_009066_, _032429_, _032446_);
  or g_123388_(_009067_, _032430_, _032447_);
  and g_123389_(_032445_, _032447_, _032448_);
  or g_123390_(_032444_, _032446_, _032450_);
  and g_123391_(_032442_, _032448_, _032451_);
  or g_123392_(_032443_, _032450_, _032452_);
  and g_123393_(_032422_, _032451_, _032453_);
  or g_123394_(_032423_, _032452_, _032454_);
  or g_123395_(_008868_, _032397_, _032455_);
  not g_123396_(_032455_, _032456_);
  and g_123397_(_032316_, _032397_, _032457_);
  not g_123398_(_032457_, _032458_);
  and g_123399_(_032455_, _032458_, _032459_);
  or g_123400_(_032456_, _032457_, _032461_);
  and g_123401_(_009111_, _032459_, _032462_);
  or g_123402_(_009110_, _032461_, _032463_);
  xor g_123403_(_009111_, _032459_, _032464_);
  xor g_123404_(_009110_, _032459_, _032465_);
  or g_123405_(_008878_, _032397_, _032466_);
  not g_123406_(_032466_, _032467_);
  and g_123407_(_032309_, _032397_, _032468_);
  not g_123408_(_032468_, _032469_);
  and g_123409_(_032466_, _032469_, _032470_);
  or g_123410_(_032467_, _032468_, _032472_);
  or g_123411_(_009101_, _032470_, _032473_);
  not g_123412_(_032473_, _032474_);
  and g_123413_(_009101_, _032470_, _032475_);
  or g_123414_(_009100_, _032472_, _032476_);
  xor g_123415_(_009101_, _032470_, _032477_);
  xor g_123416_(_009100_, _032470_, _032478_);
  and g_123417_(_032464_, _032477_, _032479_);
  or g_123418_(_032465_, _032478_, _032480_);
  and g_123419_(_008892_, _032396_, _032481_);
  or g_123420_(_008893_, _032397_, _032483_);
  and g_123421_(_032330_, _032397_, _032484_);
  or g_123422_(_032329_, _032396_, _032485_);
  and g_123423_(_032483_, _032485_, _032486_);
  or g_123424_(_032481_, _032484_, _032487_);
  and g_123425_(_009125_, _032487_, _032488_);
  or g_123426_(_009124_, _032486_, _032489_);
  xor g_123427_(_009124_, _032486_, _032490_);
  xor g_123428_(_009125_, _032486_, _032491_);
  and g_123429_(_008899_, _032396_, _032492_);
  or g_123430_(_008900_, _032397_, _032494_);
  and g_123431_(_032338_, _032397_, _032495_);
  or g_123432_(_032337_, _032396_, _032496_);
  and g_123433_(_032494_, _032496_, _032497_);
  or g_123434_(_032492_, _032495_, _032498_);
  and g_123435_(_009133_, _032498_, _032499_);
  or g_123436_(_009132_, _032497_, _032500_);
  and g_123437_(_009132_, _032497_, _032501_);
  or g_123438_(_009133_, _032498_, _032502_);
  and g_123439_(_032500_, _032502_, _032503_);
  or g_123440_(_032499_, _032501_, _032505_);
  and g_123441_(_032490_, _032503_, _032506_);
  or g_123442_(_032491_, _032505_, _032507_);
  and g_123443_(_032479_, _032506_, _032508_);
  or g_123444_(_032480_, _032507_, _032509_);
  and g_123445_(_032453_, _032508_, _032510_);
  or g_123446_(_032454_, _032509_, _032511_);
  or g_123447_(_008918_, _032397_, _032512_);
  or g_123448_(_032203_, _032396_, _032513_);
  and g_123449_(_032512_, _032513_, _032514_);
  and g_123450_(_008999_, _032514_, _032516_);
  and g_123451_(_032214_, _032397_, _032517_);
  and g_123452_(_053387_, _032396_, _032518_);
  or g_123453_(_032517_, _032518_, _032519_);
  or g_123454_(_053562_, _032519_, _032520_);
  or g_123455_(_008999_, _032514_, _032521_);
  xor g_123456_(_008999_, _032514_, _032522_);
  xor g_123457_(_008998_, _032514_, _032523_);
  xor g_123458_(_053562_, _032519_, _032524_);
  xor g_123459_(_053561_, _032519_, _032525_);
  and g_123460_(_032510_, _032524_, _032527_);
  or g_123461_(_032511_, _032525_, _032528_);
  and g_123462_(_032522_, _032527_, _032529_);
  or g_123463_(_032523_, _032528_, _032530_);
  and g_123464_(out[433], _032396_, _032531_);
  and g_123465_(_032225_, _032397_, _032532_);
  or g_123466_(_032531_, _032532_, _032533_);
  not g_123467_(_032533_, _032534_);
  and g_123468_(out[449], _032534_, _032535_);
  or g_123469_(_054215_, _032533_, _032536_);
  and g_123470_(out[448], _032401_, _032538_);
  or g_123471_(_004806_, _032400_, _032539_);
  xor g_123472_(_054215_, _032533_, _032540_);
  xor g_123473_(out[449], _032533_, _032541_);
  and g_123474_(_032539_, _032540_, _032542_);
  or g_123475_(_032538_, _032541_, _032543_);
  and g_123476_(_032536_, _032543_, _032544_);
  or g_123477_(_032535_, _032542_, _032545_);
  and g_123478_(_032529_, _032545_, _032546_);
  or g_123479_(_032530_, _032544_, _032547_);
  or g_123480_(_032516_, _032520_, _032549_);
  and g_123481_(_032521_, _032549_, _032550_);
  or g_123482_(_032511_, _032550_, _032551_);
  not g_123483_(_032551_, _032552_);
  and g_123484_(_032489_, _032500_, _032553_);
  or g_123485_(_032488_, _032499_, _032554_);
  and g_123486_(_032502_, _032554_, _032555_);
  or g_123487_(_032501_, _032553_, _032556_);
  and g_123488_(_032479_, _032555_, _032557_);
  or g_123489_(_032480_, _032556_, _032558_);
  and g_123490_(_032462_, _032476_, _032560_);
  or g_123491_(_032463_, _032475_, _032561_);
  and g_123492_(_032473_, _032561_, _032562_);
  or g_123493_(_032474_, _032560_, _032563_);
  and g_123494_(_032558_, _032562_, _032564_);
  or g_123495_(_032557_, _032563_, _032565_);
  and g_123496_(_032453_, _032565_, _032566_);
  or g_123497_(_032454_, _032564_, _032567_);
  and g_123498_(_032422_, _032443_, _032568_);
  and g_123499_(_032445_, _032568_, _032569_);
  not g_123500_(_032569_, _032571_);
  and g_123501_(_032417_, _032420_, _032572_);
  or g_123502_(_032415_, _032419_, _032573_);
  and g_123503_(_032414_, _032573_, _032574_);
  or g_123504_(_032413_, _032572_, _032575_);
  and g_123505_(_032571_, _032574_, _032576_);
  or g_123506_(_032569_, _032575_, _032577_);
  and g_123507_(_032567_, _032576_, _032578_);
  or g_123508_(_032566_, _032577_, _032579_);
  and g_123509_(_032551_, _032578_, _032580_);
  or g_123510_(_032552_, _032579_, _032582_);
  and g_123511_(_032547_, _032580_, _032583_);
  or g_123512_(_032546_, _032582_, _032584_);
  and g_123513_(_004806_, _032400_, _032585_);
  or g_123514_(_032543_, _032585_, _032586_);
  or g_123515_(_032530_, _032586_, _032587_);
  not g_123516_(_032587_, _032588_);
  and g_123517_(_032584_, _032587_, _032589_);
  or g_123518_(_032583_, _032588_, _032590_);
  or g_123519_(_032400_, _032589_, _032591_);
  or g_123520_(out[448], _032590_, _032593_);
  and g_123521_(_032591_, _032593_, _032594_);
  not g_123522_(_032594_, _032595_);
  and g_123523_(_009078_, _032589_, _032596_);
  and g_123524_(_032439_, _032590_, _032597_);
  or g_123525_(_032596_, _032597_, _032598_);
  not g_123526_(_032598_, _032599_);
  and g_123527_(_009192_, _032598_, _032600_);
  or g_123528_(_009191_, _032599_, _032601_);
  or g_123529_(_009066_, _032590_, _032602_);
  not g_123530_(_032602_, _032604_);
  and g_123531_(_032429_, _032590_, _032605_);
  not g_123532_(_032605_, _032606_);
  and g_123533_(_032602_, _032606_, _032607_);
  or g_123534_(_032604_, _032605_, _032608_);
  and g_123535_(_009204_, _032608_, _032609_);
  or g_123536_(_009205_, _032607_, _032610_);
  and g_123537_(_032601_, _032610_, _032611_);
  or g_123538_(_032600_, _032609_, _032612_);
  or g_123539_(out[474], _009190_, _032613_);
  xor g_123540_(out[474], _009190_, _032615_);
  not g_123541_(_032615_, _032616_);
  and g_123542_(_032403_, _032589_, _032617_);
  and g_123543_(_032408_, _032590_, _032618_);
  or g_123544_(_032617_, _032618_, _032619_);
  not g_123545_(_032619_, _032620_);
  and g_123546_(_032616_, _032619_, _032621_);
  or g_123547_(_032615_, _032620_, _032622_);
  and g_123548_(_009205_, _032607_, _032623_);
  or g_123549_(_009204_, _032608_, _032624_);
  or g_123550_(_032621_, _032623_, _032626_);
  or g_123551_(_032612_, _032626_, _032627_);
  and g_123552_(_032409_, _032411_, _032628_);
  not g_123553_(_032628_, _032629_);
  xor g_123554_(out[475], _032613_, _032630_);
  not g_123555_(_032630_, _032631_);
  and g_123556_(_032628_, _032631_, _032632_);
  or g_123557_(_032629_, _032630_, _032633_);
  and g_123558_(_032615_, _032620_, _032634_);
  or g_123559_(_032616_, _032619_, _032635_);
  and g_123560_(_032633_, _032635_, _032637_);
  or g_123561_(_032632_, _032634_, _032638_);
  and g_123562_(_032629_, _032630_, _032639_);
  or g_123563_(_032628_, _032631_, _032640_);
  and g_123564_(_009191_, _032599_, _032641_);
  or g_123565_(_009192_, _032598_, _032642_);
  or g_123566_(_032639_, _032641_, _032643_);
  or g_123567_(_032638_, _032643_, _032644_);
  and g_123568_(_032622_, _032637_, _032645_);
  and g_123569_(_032640_, _032645_, _032646_);
  and g_123570_(_032624_, _032642_, _032648_);
  and g_123571_(_032611_, _032648_, _032649_);
  and g_123572_(_032646_, _032649_, _032650_);
  or g_123573_(_032627_, _032644_, _032651_);
  or g_123574_(_009110_, _032590_, _032652_);
  or g_123575_(_032459_, _032589_, _032653_);
  and g_123576_(_032652_, _032653_, _032654_);
  not g_123577_(_032654_, _032655_);
  or g_123578_(_009233_, _032655_, _032656_);
  xor g_123579_(_009233_, _032654_, _032657_);
  or g_123580_(_009100_, _032590_, _032659_);
  or g_123581_(_032470_, _032589_, _032660_);
  and g_123582_(_032659_, _032660_, _032661_);
  or g_123583_(_003130_, _032661_, _032662_);
  and g_123584_(_003130_, _032661_, _032663_);
  xor g_123585_(_003129_, _032661_, _032664_);
  or g_123586_(_032657_, _032664_, _032665_);
  not g_123587_(_032665_, _032666_);
  and g_123588_(_009132_, _032589_, _032667_);
  or g_123589_(_009133_, _032590_, _032668_);
  and g_123590_(_032498_, _032590_, _032670_);
  or g_123591_(_032497_, _032589_, _032671_);
  and g_123592_(_032668_, _032671_, _032672_);
  or g_123593_(_032667_, _032670_, _032673_);
  and g_123594_(_009265_, _032673_, _032674_);
  or g_123595_(_009264_, _032672_, _032675_);
  and g_123596_(_009125_, _032589_, _032676_);
  or g_123597_(_009124_, _032590_, _032677_);
  and g_123598_(_032486_, _032590_, _032678_);
  or g_123599_(_032487_, _032589_, _032679_);
  and g_123600_(_032677_, _032679_, _032681_);
  or g_123601_(_032676_, _032678_, _032682_);
  and g_123602_(_009255_, _032681_, _032683_);
  or g_123603_(_009254_, _032682_, _032684_);
  and g_123604_(_032675_, _032684_, _032685_);
  or g_123605_(_032674_, _032683_, _032686_);
  or g_123606_(_009255_, _032681_, _032687_);
  not g_123607_(_032687_, _032688_);
  and g_123608_(_009264_, _032672_, _032689_);
  not g_123609_(_032689_, _032690_);
  or g_123610_(_032686_, _032688_, _032692_);
  or g_123611_(_032689_, _032692_, _032693_);
  or g_123612_(_032665_, _032693_, _032694_);
  not g_123613_(_032694_, _032695_);
  and g_123614_(_032650_, _032695_, _032696_);
  or g_123615_(_032651_, _032694_, _032697_);
  or g_123616_(_008998_, _032590_, _032698_);
  or g_123617_(_032514_, _032589_, _032699_);
  and g_123618_(_032698_, _032699_, _032700_);
  or g_123619_(_009291_, _032700_, _032701_);
  and g_123620_(_032519_, _032590_, _032703_);
  and g_123621_(_053561_, _032589_, _032704_);
  or g_123622_(_032703_, _032704_, _032705_);
  or g_123623_(_053882_, _032705_, _032706_);
  and g_123624_(_032701_, _032706_, _032707_);
  and g_123625_(_009291_, _032700_, _032708_);
  xor g_123626_(_009290_, _032700_, _032709_);
  xor g_123627_(_053881_, _032705_, _032710_);
  or g_123628_(_032709_, _032710_, _032711_);
  and g_123629_(out[449], _032589_, _032712_);
  and g_123630_(_032533_, _032590_, _032714_);
  or g_123631_(_032712_, _032714_, _032715_);
  or g_123632_(_054314_, _032715_, _032716_);
  and g_123633_(out[464], _032595_, _032717_);
  xor g_123634_(out[465], _032715_, _032718_);
  or g_123635_(_032717_, _032718_, _032719_);
  and g_123636_(_032716_, _032719_, _032720_);
  or g_123637_(_032711_, _032720_, _032721_);
  or g_123638_(_032707_, _032708_, _032722_);
  and g_123639_(_032721_, _032722_, _032723_);
  not g_123640_(_032723_, _032725_);
  and g_123641_(_032696_, _032725_, _032726_);
  or g_123642_(_032697_, _032723_, _032727_);
  and g_123643_(_032686_, _032690_, _032728_);
  or g_123644_(_032685_, _032689_, _032729_);
  and g_123645_(_032666_, _032728_, _032730_);
  or g_123646_(_032665_, _032729_, _032731_);
  or g_123647_(_032656_, _032663_, _032732_);
  and g_123648_(_032662_, _032732_, _032733_);
  not g_123649_(_032733_, _032734_);
  and g_123650_(_032731_, _032733_, _032736_);
  or g_123651_(_032730_, _032734_, _032737_);
  and g_123652_(_032650_, _032737_, _032738_);
  or g_123653_(_032651_, _032736_, _032739_);
  and g_123654_(_032601_, _032624_, _032740_);
  or g_123655_(_032600_, _032623_, _032741_);
  and g_123656_(_032622_, _032642_, _032742_);
  or g_123657_(_032621_, _032641_, _032743_);
  and g_123658_(_032741_, _032742_, _032744_);
  or g_123659_(_032740_, _032743_, _032745_);
  and g_123660_(_032637_, _032745_, _032747_);
  or g_123661_(_032638_, _032744_, _032748_);
  and g_123662_(_032640_, _032748_, _032749_);
  or g_123663_(_032639_, _032747_, _032750_);
  and g_123664_(_032739_, _032750_, _032751_);
  or g_123665_(_032738_, _032749_, _032752_);
  and g_123666_(_032727_, _032751_, _032753_);
  or g_123667_(_032726_, _032752_, _032754_);
  and g_123668_(_004839_, _032594_, _032755_);
  or g_123669_(_032711_, _032755_, _032756_);
  or g_123670_(_032719_, _032756_, _032758_);
  not g_123671_(_032758_, _032759_);
  and g_123672_(_032696_, _032759_, _032760_);
  or g_123673_(_032697_, _032758_, _032761_);
  and g_123674_(_032754_, _032761_, _032762_);
  or g_123675_(_032753_, _032760_, _032763_);
  or g_123676_(_032594_, _032762_, _032764_);
  or g_123677_(out[464], _032763_, _032765_);
  and g_123678_(_032764_, _032765_, _032766_);
  or g_123679_(out[490], _009872_, _032767_);
  xor g_123680_(out[491], _032767_, _032769_);
  xor g_123681_(_054358_, _032767_, _032770_);
  or g_123682_(out[506], _009875_, _032771_);
  xor g_123683_(out[507], _032771_, _032772_);
  xor g_123684_(_054479_, _032771_, _032773_);
  and g_123685_(_032770_, _032772_, _032774_);
  or g_123686_(_032769_, _032773_, _032775_);
  xor g_123687_(out[490], _009872_, _032776_);
  xor g_123688_(_054468_, _009872_, _032777_);
  xor g_123689_(out[506], _009875_, _032778_);
  xor g_123690_(_054600_, _009875_, _032780_);
  and g_123691_(_032777_, _032778_, _032781_);
  or g_123692_(_032776_, _032780_, _032782_);
  and g_123693_(_032776_, _032780_, _032783_);
  or g_123694_(_032777_, _032778_, _032784_);
  and g_123695_(_009880_, _010001_, _032785_);
  or g_123696_(_009879_, _010000_, _032786_);
  and g_123697_(_032784_, _032786_, _032787_);
  or g_123698_(_032783_, _032785_, _032788_);
  and g_123699_(_032782_, _032788_, _032789_);
  or g_123700_(_032781_, _032787_, _032791_);
  and g_123701_(_032775_, _032791_, _032792_);
  or g_123702_(_032774_, _032789_, _032793_);
  and g_123703_(_032769_, _032773_, _032794_);
  or g_123704_(_032770_, _032772_, _032795_);
  or g_123705_(_032792_, _032794_, _032796_);
  and g_123706_(_032793_, _032795_, _032797_);
  and g_123707_(_009996_, _032797_, _032798_);
  or g_123708_(_009995_, _032796_, _032799_);
  and g_123709_(_009966_, _032799_, _032800_);
  or g_123710_(_009964_, _032798_, _032802_);
  and g_123711_(_054347_, _032802_, _032803_);
  or g_123712_(out[480], _032800_, _032804_);
  and g_123713_(_054545_, _032800_, _032805_);
  or g_123714_(out[496], _032802_, _032806_);
  and g_123715_(_032804_, _032806_, _032807_);
  or g_123716_(_032803_, _032805_, _032808_);
  and g_123717_(_009967_, _032800_, _032809_);
  or g_123718_(_009968_, _032802_, _032810_);
  and g_123719_(_009969_, _032802_, _032811_);
  or g_123720_(_009970_, _032800_, _032813_);
  and g_123721_(_032810_, _032813_, _032814_);
  or g_123722_(_032809_, _032811_, _032815_);
  and g_123723_(_010133_, _032815_, _032816_);
  or g_123724_(_010132_, _032814_, _032817_);
  and g_123725_(_009939_, _032800_, _032818_);
  or g_123726_(_009938_, _032802_, _032819_);
  and g_123727_(_009935_, _032802_, _032820_);
  or g_123728_(_009934_, _032800_, _032821_);
  and g_123729_(_032819_, _032821_, _032822_);
  or g_123730_(_032818_, _032820_, _032824_);
  and g_123731_(_010094_, _032824_, _032825_);
  or g_123732_(_010095_, _032822_, _032826_);
  and g_123733_(_032817_, _032826_, _032827_);
  or g_123734_(_032816_, _032825_, _032828_);
  and g_123735_(_016367_, _032800_, _032829_);
  or g_123736_(_016378_, _032802_, _032830_);
  and g_123737_(_016400_, _032802_, _032831_);
  or g_123738_(_016411_, _032800_, _032832_);
  and g_123739_(_032830_, _032832_, _032833_);
  or g_123740_(_032829_, _032831_, _032835_);
  and g_123741_(_010132_, _032814_, _032836_);
  or g_123742_(_010133_, _032815_, _032837_);
  and g_123743_(_019084_, _032833_, _032838_);
  or g_123744_(_019095_, _032835_, _032839_);
  and g_123745_(_032837_, _032839_, _032840_);
  or g_123746_(_032836_, _032838_, _032841_);
  and g_123747_(_032817_, _032837_, _032842_);
  or g_123748_(_032816_, _032836_, _032843_);
  xor g_123749_(_019084_, _032833_, _032844_);
  xor g_123750_(_019095_, _032833_, _032846_);
  and g_123751_(_032826_, _032844_, _032847_);
  or g_123752_(_032825_, _032846_, _032848_);
  and g_123753_(_032842_, _032847_, _032849_);
  or g_123754_(_032843_, _032848_, _032850_);
  and g_123755_(out[497], _032800_, _032851_);
  or g_123756_(_054534_, _032802_, _032852_);
  and g_123757_(out[481], _032802_, _032853_);
  or g_123758_(_054413_, _032800_, _032854_);
  and g_123759_(_032852_, _032854_, _032855_);
  or g_123760_(_032851_, _032853_, _032857_);
  and g_123761_(out[512], _032808_, _032858_);
  or g_123762_(_054677_, _032807_, _032859_);
  and g_123763_(out[513], _032855_, _032860_);
  or g_123764_(_054666_, _032857_, _032861_);
  xor g_123765_(out[513], _032855_, _032862_);
  xor g_123766_(_054666_, _032855_, _032863_);
  and g_123767_(_032859_, _032862_, _032864_);
  or g_123768_(_032858_, _032863_, _032865_);
  and g_123769_(_010095_, _032822_, _032866_);
  or g_123770_(_010094_, _032824_, _032868_);
  and g_123771_(_009944_, _032800_, _032869_);
  or g_123772_(_009942_, _032802_, _032870_);
  and g_123773_(_009946_, _032802_, _032871_);
  or g_123774_(_009945_, _032800_, _032872_);
  and g_123775_(_032870_, _032872_, _032873_);
  or g_123776_(_032869_, _032871_, _032874_);
  and g_123777_(_010106_, _032873_, _032875_);
  or g_123778_(_010105_, _032874_, _032876_);
  and g_123779_(_032868_, _032876_, _032877_);
  or g_123780_(_032866_, _032875_, _032879_);
  and g_123781_(_054677_, _032807_, _032880_);
  or g_123782_(out[512], _032808_, _032881_);
  and g_123783_(_032877_, _032881_, _032882_);
  or g_123784_(_032879_, _032880_, _032883_);
  and g_123785_(_032864_, _032882_, _032884_);
  or g_123786_(_032865_, _032883_, _032885_);
  and g_123787_(_032849_, _032884_, _032886_);
  or g_123788_(_032850_, _032885_, _032887_);
  and g_123789_(_032778_, _032800_, _032888_);
  or g_123790_(_032780_, _032802_, _032890_);
  and g_123791_(_032776_, _032802_, _032891_);
  or g_123792_(_032777_, _032800_, _032892_);
  and g_123793_(_032890_, _032892_, _032893_);
  or g_123794_(_032888_, _032891_, _032894_);
  or g_123795_(out[522], _010035_, _032895_);
  xor g_123796_(out[522], _010035_, _032896_);
  xor g_123797_(_054732_, _010035_, _032897_);
  and g_123798_(_032893_, _032896_, _032898_);
  or g_123799_(_032894_, _032897_, _032899_);
  xor g_123800_(out[523], _032895_, _032901_);
  xor g_123801_(_054611_, _032895_, _032902_);
  and g_123802_(_032773_, _032800_, _032903_);
  or g_123803_(_032772_, _032802_, _032904_);
  and g_123804_(_032770_, _032802_, _032905_);
  or g_123805_(_032769_, _032800_, _032906_);
  and g_123806_(_032904_, _032906_, _032907_);
  or g_123807_(_032903_, _032905_, _032908_);
  and g_123808_(_032902_, _032907_, _032909_);
  or g_123809_(_032901_, _032908_, _032910_);
  and g_123810_(_032899_, _032910_, _032912_);
  or g_123811_(_032898_, _032909_, _032913_);
  and g_123812_(_032894_, _032897_, _032914_);
  or g_123813_(_032893_, _032896_, _032915_);
  and g_123814_(_032901_, _032908_, _032916_);
  or g_123815_(_032902_, _032907_, _032917_);
  and g_123816_(_032915_, _032917_, _032918_);
  or g_123817_(_032914_, _032916_, _032919_);
  and g_123818_(_032912_, _032918_, _032920_);
  or g_123819_(_032913_, _032919_, _032921_);
  or g_123820_(_009887_, _032802_, _032923_);
  or g_123821_(_009885_, _032800_, _032924_);
  and g_123822_(_032923_, _032924_, _032925_);
  not g_123823_(_032925_, _032926_);
  or g_123824_(_010054_, _032926_, _032927_);
  and g_123825_(_009876_, _032800_, _032928_);
  and g_123826_(_009873_, _032802_, _032929_);
  or g_123827_(_032928_, _032929_, _032930_);
  not g_123828_(_032930_, _032931_);
  or g_123829_(_010036_, _032931_, _032932_);
  and g_123830_(_032927_, _032932_, _032934_);
  not g_123831_(_032934_, _032935_);
  and g_123832_(_010054_, _032926_, _032936_);
  or g_123833_(_010055_, _032925_, _032937_);
  and g_123834_(_010036_, _032931_, _032938_);
  or g_123835_(_010037_, _032930_, _032939_);
  and g_123836_(_032937_, _032939_, _032940_);
  or g_123837_(_032936_, _032938_, _032941_);
  and g_123838_(_032934_, _032940_, _032942_);
  or g_123839_(_032935_, _032941_, _032943_);
  and g_123840_(_032920_, _032942_, _032945_);
  or g_123841_(_032921_, _032943_, _032946_);
  and g_123842_(_009909_, _032800_, _032947_);
  and g_123843_(_009907_, _032802_, _032948_);
  or g_123844_(_032947_, _032948_, _032949_);
  not g_123845_(_032949_, _032950_);
  and g_123846_(_010080_, _032950_, _032951_);
  or g_123847_(_010081_, _032949_, _032952_);
  or g_123848_(_009916_, _032802_, _032953_);
  or g_123849_(_009914_, _032800_, _032954_);
  and g_123850_(_032953_, _032954_, _032956_);
  not g_123851_(_032956_, _032957_);
  and g_123852_(_010071_, _032957_, _032958_);
  or g_123853_(_010072_, _032956_, _032959_);
  and g_123854_(_032952_, _032959_, _032960_);
  or g_123855_(_032951_, _032958_, _032961_);
  and g_123856_(_010072_, _032956_, _032962_);
  or g_123857_(_010071_, _032957_, _032963_);
  and g_123858_(_010105_, _032874_, _032964_);
  or g_123859_(_010106_, _032873_, _032965_);
  and g_123860_(_010081_, _032949_, _032967_);
  or g_123861_(_010080_, _032950_, _032968_);
  and g_123862_(_032965_, _032968_, _032969_);
  or g_123863_(_032964_, _032967_, _032970_);
  and g_123864_(_032963_, _032969_, _032971_);
  or g_123865_(_032962_, _032970_, _032972_);
  and g_123866_(_032960_, _032971_, _032973_);
  or g_123867_(_032961_, _032972_, _032974_);
  and g_123868_(_032945_, _032973_, _032975_);
  or g_123869_(_032946_, _032974_, _032976_);
  and g_123870_(_032886_, _032975_, _032978_);
  or g_123871_(_032887_, _032976_, _032979_);
  and g_123872_(_032861_, _032865_, _032980_);
  or g_123873_(_032860_, _032864_, _032981_);
  and g_123874_(_032849_, _032981_, _032982_);
  or g_123875_(_032850_, _032980_, _032983_);
  and g_123876_(_032827_, _032841_, _032984_);
  or g_123877_(_032828_, _032840_, _032985_);
  and g_123878_(_032877_, _032985_, _032986_);
  or g_123879_(_032879_, _032984_, _032987_);
  and g_123880_(_032983_, _032986_, _032989_);
  or g_123881_(_032982_, _032987_, _032990_);
  and g_123882_(_032973_, _032990_, _032991_);
  or g_123883_(_032974_, _032989_, _032992_);
  and g_123884_(_032962_, _032968_, _032993_);
  or g_123885_(_032963_, _032967_, _032994_);
  and g_123886_(_032952_, _032994_, _032995_);
  or g_123887_(_032951_, _032993_, _032996_);
  and g_123888_(_032992_, _032995_, _032997_);
  or g_123889_(_032991_, _032996_, _032998_);
  and g_123890_(_032945_, _032998_, _033000_);
  or g_123891_(_032946_, _032997_, _033001_);
  and g_123892_(_032913_, _032917_, _033002_);
  or g_123893_(_032912_, _032916_, _033003_);
  and g_123894_(_032920_, _032939_, _033004_);
  not g_123895_(_033004_, _033005_);
  and g_123896_(_032935_, _033004_, _033006_);
  or g_123897_(_032934_, _033005_, _033007_);
  and g_123898_(_033003_, _033007_, _033008_);
  or g_123899_(_033002_, _033006_, _033009_);
  and g_123900_(_033001_, _033008_, _033011_);
  or g_123901_(_033000_, _033009_, _033012_);
  and g_123902_(_032979_, _033012_, _033013_);
  or g_123903_(_032978_, _033011_, _033014_);
  and g_123904_(_032808_, _033014_, _033015_);
  or g_123905_(_032807_, _033013_, _033016_);
  and g_123906_(_054677_, _033013_, _033017_);
  or g_123907_(out[512], _033014_, _033018_);
  and g_123908_(_033016_, _033018_, _033019_);
  or g_123909_(_033015_, _033017_, _033020_);
  and g_123910_(_032901_, _032907_, _033022_);
  or g_123911_(_032902_, _032908_, _033023_);
  or g_123912_(out[538], _010255_, _033024_);
  xor g_123913_(out[539], _033024_, _033025_);
  xor g_123914_(_054743_, _033024_, _033026_);
  and g_123915_(_033023_, _033025_, _033027_);
  or g_123916_(_033022_, _033026_, _033028_);
  and g_123917_(_033022_, _033026_, _033029_);
  or g_123918_(_033023_, _033025_, _033030_);
  and g_123919_(_032894_, _033014_, _033031_);
  or g_123920_(_032893_, _033013_, _033033_);
  and g_123921_(_032896_, _033013_, _033034_);
  or g_123922_(_032897_, _033014_, _033035_);
  and g_123923_(_033033_, _033035_, _033036_);
  or g_123924_(_033031_, _033034_, _033037_);
  xor g_123925_(out[538], _010255_, _033038_);
  xor g_123926_(_054864_, _010255_, _033039_);
  and g_123927_(_033036_, _033038_, _033040_);
  or g_123928_(_033037_, _033039_, _033041_);
  and g_123929_(_033030_, _033041_, _033042_);
  or g_123930_(_033029_, _033040_, _033044_);
  and g_123931_(_033028_, _033044_, _033045_);
  or g_123932_(_033027_, _033042_, _033046_);
  and g_123933_(_033037_, _033039_, _033047_);
  or g_123934_(_033036_, _033038_, _033048_);
  and g_123935_(_033028_, _033048_, _033049_);
  or g_123936_(_033027_, _033047_, _033050_);
  and g_123937_(_033042_, _033049_, _033051_);
  or g_123938_(_033044_, _033050_, _033052_);
  and g_123939_(_010036_, _033013_, _033053_);
  or g_123940_(_010037_, _033014_, _033055_);
  and g_123941_(_032930_, _033014_, _033056_);
  not g_123942_(_033056_, _033057_);
  and g_123943_(_033055_, _033057_, _033058_);
  or g_123944_(_033053_, _033056_, _033059_);
  and g_123945_(_010256_, _033058_, _033060_);
  or g_123946_(_010257_, _033059_, _033061_);
  or g_123947_(_033052_, _033060_, _033062_);
  and g_123948_(_010257_, _033059_, _033063_);
  or g_123949_(_010256_, _033058_, _033064_);
  and g_123950_(_010054_, _033013_, _033066_);
  or g_123951_(_010055_, _033014_, _033067_);
  and g_123952_(_032925_, _033014_, _033068_);
  not g_123953_(_033068_, _033069_);
  and g_123954_(_033067_, _033069_, _033070_);
  or g_123955_(_033066_, _033068_, _033071_);
  and g_123956_(_010252_, _033071_, _033072_);
  or g_123957_(_010250_, _033070_, _033073_);
  and g_123958_(_033064_, _033073_, _033074_);
  or g_123959_(_033063_, _033072_, _033075_);
  or g_123960_(_032949_, _033013_, _033077_);
  or g_123961_(_010080_, _033014_, _033078_);
  and g_123962_(_033077_, _033078_, _033079_);
  not g_123963_(_033079_, _033080_);
  and g_123964_(_010297_, _033079_, _033081_);
  or g_123965_(_010296_, _033080_, _033082_);
  and g_123966_(_010296_, _033080_, _033083_);
  or g_123967_(_010297_, _033079_, _033084_);
  or g_123968_(_032956_, _033013_, _033085_);
  or g_123969_(_010071_, _033014_, _033086_);
  and g_123970_(_033085_, _033086_, _033088_);
  not g_123971_(_033088_, _033089_);
  and g_123972_(_010288_, _033088_, _033090_);
  or g_123973_(_010287_, _033089_, _033091_);
  and g_123974_(_033084_, _033091_, _033092_);
  or g_123975_(_033083_, _033090_, _033093_);
  and g_123976_(_033082_, _033093_, _033094_);
  or g_123977_(_033081_, _033092_, _033095_);
  and g_123978_(_010094_, _033013_, _033096_);
  or g_123979_(_010095_, _033014_, _033097_);
  and g_123980_(_032822_, _033014_, _033099_);
  or g_123981_(_032824_, _033013_, _033100_);
  and g_123982_(_033097_, _033100_, _033101_);
  or g_123983_(_033096_, _033099_, _033102_);
  and g_123984_(_010312_, _033101_, _033103_);
  or g_123985_(_010313_, _033102_, _033104_);
  or g_123986_(_010132_, _033014_, _033105_);
  or g_123987_(_032815_, _033013_, _033106_);
  and g_123988_(_033105_, _033106_, _033107_);
  or g_123989_(_010351_, _033107_, _033108_);
  and g_123990_(_032835_, _033014_, _033110_);
  or g_123991_(_032833_, _033013_, _033111_);
  and g_123992_(_019084_, _033013_, _033112_);
  or g_123993_(_019095_, _033014_, _033113_);
  and g_123994_(_033111_, _033113_, _033114_);
  or g_123995_(_033110_, _033112_, _033115_);
  or g_123996_(_020998_, _033115_, _033116_);
  and g_123997_(_010351_, _033107_, _033117_);
  xor g_123998_(_010351_, _033107_, _033118_);
  xor g_123999_(_010349_, _033107_, _033119_);
  xor g_124000_(_020987_, _033114_, _033121_);
  xor g_124001_(_020998_, _033114_, _033122_);
  and g_124002_(_033118_, _033121_, _033123_);
  or g_124003_(_033119_, _033122_, _033124_);
  and g_124004_(out[513], _033013_, _033125_);
  or g_124005_(_054666_, _033014_, _033126_);
  and g_124006_(_032857_, _033014_, _033127_);
  or g_124007_(_032855_, _033013_, _033128_);
  and g_124008_(_033126_, _033128_, _033129_);
  or g_124009_(_033125_, _033127_, _033130_);
  and g_124010_(out[529], _033129_, _033132_);
  not g_124011_(_033132_, _033133_);
  and g_124012_(out[528], _033020_, _033134_);
  or g_124013_(_054809_, _033019_, _033135_);
  and g_124014_(_054798_, _033130_, _033136_);
  or g_124015_(out[529], _033129_, _033137_);
  and g_124016_(_033135_, _033137_, _033138_);
  or g_124017_(_033134_, _033136_, _033139_);
  and g_124018_(_033133_, _033139_, _033140_);
  or g_124019_(_033132_, _033138_, _033141_);
  and g_124020_(_033123_, _033141_, _033143_);
  or g_124021_(_033124_, _033140_, _033144_);
  or g_124022_(_033116_, _033117_, _033145_);
  and g_124023_(_033108_, _033145_, _033146_);
  not g_124024_(_033146_, _033147_);
  and g_124025_(_033144_, _033146_, _033148_);
  or g_124026_(_033143_, _033147_, _033149_);
  and g_124027_(_033104_, _033149_, _033150_);
  or g_124028_(_033103_, _033148_, _033151_);
  and g_124029_(_032873_, _033014_, _033152_);
  or g_124030_(_032874_, _033013_, _033154_);
  and g_124031_(_010105_, _033013_, _033155_);
  or g_124032_(_010106_, _033014_, _033156_);
  and g_124033_(_033154_, _033156_, _033157_);
  or g_124034_(_033152_, _033155_, _033158_);
  and g_124035_(_010324_, _033158_, _033159_);
  or g_124036_(_010323_, _033157_, _033160_);
  and g_124037_(_010313_, _033102_, _033161_);
  or g_124038_(_010312_, _033101_, _033162_);
  and g_124039_(_033160_, _033162_, _033163_);
  or g_124040_(_033159_, _033161_, _033165_);
  and g_124041_(_033151_, _033163_, _033166_);
  or g_124042_(_033150_, _033165_, _033167_);
  and g_124043_(_010323_, _033157_, _033168_);
  or g_124044_(_010324_, _033158_, _033169_);
  and g_124045_(_010287_, _033089_, _033170_);
  or g_124046_(_010288_, _033088_, _033171_);
  and g_124047_(_033082_, _033171_, _033172_);
  or g_124048_(_033081_, _033170_, _033173_);
  and g_124049_(_033092_, _033172_, _033174_);
  or g_124050_(_033093_, _033173_, _033176_);
  and g_124051_(_033169_, _033174_, _033177_);
  or g_124052_(_033168_, _033176_, _033178_);
  and g_124053_(_033167_, _033177_, _033179_);
  or g_124054_(_033166_, _033178_, _033180_);
  and g_124055_(_033095_, _033180_, _033181_);
  or g_124056_(_033094_, _033179_, _033182_);
  and g_124057_(_010250_, _033070_, _033183_);
  or g_124058_(_010252_, _033071_, _033184_);
  and g_124059_(_033061_, _033184_, _033185_);
  or g_124060_(_033060_, _033183_, _033187_);
  and g_124061_(_033074_, _033185_, _033188_);
  or g_124062_(_033075_, _033187_, _033189_);
  and g_124063_(_033051_, _033188_, _033190_);
  or g_124064_(_033052_, _033189_, _033191_);
  and g_124065_(_033182_, _033190_, _033192_);
  or g_124066_(_033181_, _033191_, _033193_);
  and g_124067_(_033061_, _033075_, _033194_);
  and g_124068_(_033051_, _033194_, _033195_);
  or g_124069_(_033062_, _033074_, _033196_);
  and g_124070_(_033046_, _033196_, _033198_);
  or g_124071_(_033045_, _033195_, _033199_);
  and g_124072_(_033193_, _033198_, _033200_);
  or g_124073_(_033192_, _033199_, _033201_);
  and g_124074_(_054809_, _033019_, _033202_);
  or g_124075_(out[528], _033020_, _033203_);
  and g_124076_(_033138_, _033169_, _033204_);
  and g_124077_(_033160_, _033204_, _033205_);
  and g_124078_(_033174_, _033205_, _033206_);
  not g_124079_(_033206_, _033207_);
  and g_124080_(_033104_, _033162_, _033209_);
  or g_124081_(_033103_, _033161_, _033210_);
  and g_124082_(_033133_, _033203_, _033211_);
  or g_124083_(_033132_, _033202_, _033212_);
  and g_124084_(_033209_, _033211_, _033213_);
  or g_124085_(_033210_, _033212_, _033214_);
  and g_124086_(_033123_, _033213_, _033215_);
  or g_124087_(_033124_, _033214_, _033216_);
  and g_124088_(_033190_, _033215_, _033217_);
  or g_124089_(_033191_, _033216_, _033218_);
  and g_124090_(_033206_, _033217_, _033220_);
  or g_124091_(_033207_, _033218_, _033221_);
  and g_124092_(_033201_, _033221_, _033222_);
  or g_124093_(_033200_, _033220_, _033223_);
  and g_124094_(_033020_, _033223_, _033224_);
  or g_124095_(_033019_, _033222_, _033225_);
  or g_124096_(out[528], _033223_, _033226_);
  not g_124097_(_033226_, _033227_);
  and g_124098_(_033225_, _033226_, _033228_);
  or g_124099_(_033224_, _033227_, _033229_);
  and g_124100_(_033107_, _033223_, _033231_);
  not g_124101_(_033231_, _033232_);
  and g_124102_(_010349_, _033222_, _033233_);
  or g_124103_(_010351_, _033223_, _033234_);
  or g_124104_(_033231_, _033233_, _033235_);
  and g_124105_(_033232_, _033234_, _033236_);
  or g_124106_(_010566_, _033236_, _033237_);
  or g_124107_(_033114_, _033222_, _033238_);
  or g_124108_(_020998_, _033223_, _033239_);
  and g_124109_(_033238_, _033239_, _033240_);
  and g_124110_(_054004_, _033240_, _033242_);
  and g_124111_(_010566_, _033236_, _033243_);
  xor g_124112_(_010567_, _033235_, _033244_);
  xor g_124113_(_054004_, _033240_, _033245_);
  and g_124114_(_033244_, _033245_, _033246_);
  or g_124115_(_054798_, _033223_, _033247_);
  or g_124116_(_033129_, _033222_, _033248_);
  and g_124117_(_033247_, _033248_, _033249_);
  and g_124118_(out[545], _033249_, _033250_);
  or g_124119_(_054941_, _033228_, _033251_);
  xor g_124120_(out[545], _033249_, _033253_);
  and g_124121_(_033251_, _033253_, _033254_);
  and g_124122_(_033246_, _033254_, _033255_);
  or g_124123_(_033242_, _033243_, _033256_);
  and g_124124_(_033237_, _033256_, _033257_);
  or g_124125_(_033250_, _033254_, _033258_);
  and g_124126_(_033246_, _033258_, _033259_);
  or g_124127_(_033257_, _033259_, _033260_);
  not g_124128_(_033260_, _033261_);
  or g_124129_(_010296_, _033223_, _033262_);
  or g_124130_(_033079_, _033222_, _033264_);
  and g_124131_(_033262_, _033264_, _033265_);
  not g_124132_(_033265_, _033266_);
  and g_124133_(_010470_, _033266_, _033267_);
  or g_124134_(_010472_, _033265_, _033268_);
  or g_124135_(_010287_, _033223_, _033269_);
  or g_124136_(_033088_, _033222_, _033270_);
  and g_124137_(_033269_, _033270_, _033271_);
  not g_124138_(_033271_, _033272_);
  and g_124139_(_010455_, _033271_, _033273_);
  or g_124140_(_010454_, _033272_, _033275_);
  and g_124141_(_010472_, _033265_, _033276_);
  or g_124142_(_010470_, _033266_, _033277_);
  and g_124143_(_010323_, _033222_, _033278_);
  or g_124144_(_010324_, _033223_, _033279_);
  and g_124145_(_033158_, _033223_, _033280_);
  not g_124146_(_033280_, _033281_);
  and g_124147_(_033279_, _033281_, _033282_);
  or g_124148_(_033278_, _033280_, _033283_);
  and g_124149_(_010459_, _033282_, _033284_);
  or g_124150_(_010461_, _033283_, _033286_);
  xor g_124151_(_010472_, _033265_, _033287_);
  xor g_124152_(_010470_, _033265_, _033288_);
  xor g_124153_(_010455_, _033271_, _033289_);
  xor g_124154_(_010454_, _033271_, _033290_);
  and g_124155_(_033287_, _033289_, _033291_);
  or g_124156_(_033288_, _033290_, _033292_);
  and g_124157_(_033286_, _033291_, _033293_);
  or g_124158_(_033284_, _033292_, _033294_);
  and g_124159_(_033022_, _033025_, _033295_);
  or g_124160_(_033023_, _033026_, _033297_);
  or g_124161_(out[554], _010525_, _033298_);
  xor g_124162_(out[555], _033298_, _033299_);
  xor g_124163_(_054875_, _033298_, _033300_);
  and g_124164_(_033295_, _033300_, _033301_);
  or g_124165_(_033297_, _033299_, _033302_);
  xor g_124166_(out[554], _010525_, _033303_);
  xor g_124167_(_054996_, _010525_, _033304_);
  and g_124168_(_033038_, _033222_, _033305_);
  or g_124169_(_033039_, _033223_, _033306_);
  and g_124170_(_033037_, _033223_, _033308_);
  or g_124171_(_033036_, _033222_, _033309_);
  and g_124172_(_033306_, _033309_, _033310_);
  or g_124173_(_033305_, _033308_, _033311_);
  and g_124174_(_033303_, _033310_, _033312_);
  or g_124175_(_033304_, _033311_, _033313_);
  and g_124176_(_033302_, _033313_, _033314_);
  or g_124177_(_033301_, _033312_, _033315_);
  and g_124178_(_033297_, _033299_, _033316_);
  or g_124179_(_033295_, _033300_, _033317_);
  and g_124180_(_033304_, _033311_, _033319_);
  or g_124181_(_033303_, _033310_, _033320_);
  and g_124182_(_033317_, _033320_, _033321_);
  or g_124183_(_033316_, _033319_, _033322_);
  and g_124184_(_033314_, _033321_, _033323_);
  or g_124185_(_033315_, _033322_, _033324_);
  and g_124186_(_010256_, _033222_, _033325_);
  or g_124187_(_010257_, _033223_, _033326_);
  and g_124188_(_033059_, _033223_, _033327_);
  or g_124189_(_033058_, _033222_, _033328_);
  and g_124190_(_033326_, _033328_, _033330_);
  or g_124191_(_033325_, _033327_, _033331_);
  and g_124192_(_010528_, _033331_, _033332_);
  or g_124193_(_010527_, _033330_, _033333_);
  and g_124194_(_010250_, _033222_, _033334_);
  or g_124195_(_010252_, _033223_, _033335_);
  and g_124196_(_033071_, _033223_, _033336_);
  or g_124197_(_033070_, _033222_, _033337_);
  and g_124198_(_033335_, _033337_, _033338_);
  or g_124199_(_033334_, _033336_, _033339_);
  and g_124200_(_010545_, _033339_, _033341_);
  or g_124201_(_010544_, _033338_, _033342_);
  and g_124202_(_033333_, _033342_, _033343_);
  or g_124203_(_033332_, _033341_, _033344_);
  and g_124204_(_010527_, _033330_, _033345_);
  or g_124205_(_010528_, _033331_, _033346_);
  and g_124206_(_010544_, _033338_, _033347_);
  or g_124207_(_010545_, _033339_, _033348_);
  and g_124208_(_033346_, _033348_, _033349_);
  or g_124209_(_033345_, _033347_, _033350_);
  and g_124210_(_033343_, _033349_, _033352_);
  or g_124211_(_033344_, _033350_, _033353_);
  and g_124212_(_033323_, _033352_, _033354_);
  or g_124213_(_033324_, _033353_, _033355_);
  and g_124214_(_010312_, _033222_, _033356_);
  or g_124215_(_010313_, _033223_, _033357_);
  and g_124216_(_033102_, _033223_, _033358_);
  not g_124217_(_033358_, _033359_);
  and g_124218_(_033357_, _033359_, _033360_);
  or g_124219_(_033356_, _033358_, _033361_);
  and g_124220_(_010491_, _033361_, _033363_);
  or g_124221_(_010490_, _033360_, _033364_);
  and g_124222_(_010461_, _033283_, _033365_);
  or g_124223_(_010459_, _033282_, _033366_);
  and g_124224_(_033364_, _033366_, _033367_);
  or g_124225_(_033363_, _033365_, _033368_);
  and g_124226_(_010490_, _033360_, _033369_);
  or g_124227_(_010491_, _033361_, _033370_);
  and g_124228_(_033367_, _033370_, _033371_);
  or g_124229_(_033368_, _033369_, _033372_);
  and g_124230_(_033354_, _033371_, _033374_);
  or g_124231_(_033355_, _033372_, _033375_);
  and g_124232_(_033293_, _033374_, _033376_);
  or g_124233_(_033294_, _033375_, _033377_);
  and g_124234_(_033260_, _033376_, _033378_);
  or g_124235_(_033261_, _033377_, _033379_);
  and g_124236_(_033315_, _033317_, _033380_);
  or g_124237_(_033314_, _033316_, _033381_);
  and g_124238_(_033344_, _033346_, _033382_);
  or g_124239_(_033343_, _033345_, _033383_);
  and g_124240_(_033323_, _033382_, _033385_);
  or g_124241_(_033324_, _033383_, _033386_);
  and g_124242_(_033381_, _033386_, _033387_);
  or g_124243_(_033380_, _033385_, _033388_);
  and g_124244_(_033293_, _033368_, _033389_);
  or g_124245_(_033294_, _033367_, _033390_);
  and g_124246_(_033273_, _033277_, _033391_);
  or g_124247_(_033275_, _033276_, _033392_);
  and g_124248_(_033268_, _033392_, _033393_);
  or g_124249_(_033267_, _033391_, _033394_);
  and g_124250_(_033390_, _033393_, _033396_);
  or g_124251_(_033389_, _033394_, _033397_);
  and g_124252_(_033354_, _033397_, _033398_);
  or g_124253_(_033355_, _033396_, _033399_);
  and g_124254_(_033387_, _033399_, _033400_);
  or g_124255_(_033388_, _033398_, _033401_);
  and g_124256_(_033379_, _033400_, _033402_);
  or g_124257_(_033378_, _033401_, _033403_);
  or g_124258_(out[544], _033229_, _033404_);
  and g_124259_(_033255_, _033404_, _033405_);
  not g_124260_(_033405_, _033407_);
  and g_124261_(_033376_, _033405_, _033408_);
  or g_124262_(_033377_, _033407_, _033409_);
  and g_124263_(_033403_, _033409_, _033410_);
  or g_124264_(_033402_, _033408_, _033411_);
  and g_124265_(_033229_, _033411_, _033412_);
  or g_124266_(_033228_, _033410_, _033413_);
  and g_124267_(_054941_, _033410_, _033414_);
  or g_124268_(out[544], _033411_, _033415_);
  and g_124269_(_033413_, _033415_, _033416_);
  or g_124270_(_033412_, _033414_, _033418_);
  and g_124271_(_033295_, _033299_, _033419_);
  or g_124272_(_033297_, _033300_, _033420_);
  or g_124273_(out[570], _010677_, _033421_);
  xor g_124274_(out[571], _033421_, _033422_);
  xor g_124275_(_055007_, _033421_, _033423_);
  and g_124276_(_033419_, _033423_, _033424_);
  or g_124277_(_033420_, _033422_, _033425_);
  and g_124278_(_033311_, _033411_, _033426_);
  or g_124279_(_033310_, _033410_, _033427_);
  and g_124280_(_033303_, _033410_, _033429_);
  or g_124281_(_033304_, _033411_, _033430_);
  and g_124282_(_033427_, _033430_, _033431_);
  or g_124283_(_033426_, _033429_, _033432_);
  xor g_124284_(out[570], _010677_, _033433_);
  xor g_124285_(_055128_, _010677_, _033434_);
  and g_124286_(_033431_, _033433_, _033435_);
  or g_124287_(_033432_, _033434_, _033436_);
  and g_124288_(_033425_, _033436_, _033437_);
  or g_124289_(_033424_, _033435_, _033438_);
  and g_124290_(_033432_, _033434_, _033440_);
  or g_124291_(_033431_, _033433_, _033441_);
  and g_124292_(_033420_, _033422_, _033442_);
  or g_124293_(_033419_, _033423_, _033443_);
  and g_124294_(_033441_, _033443_, _033444_);
  or g_124295_(_033440_, _033442_, _033445_);
  and g_124296_(_033437_, _033444_, _033446_);
  or g_124297_(_033438_, _033445_, _033447_);
  and g_124298_(_010544_, _033410_, _033448_);
  or g_124299_(_010545_, _033411_, _033449_);
  and g_124300_(_033339_, _033411_, _033451_);
  or g_124301_(_033338_, _033410_, _033452_);
  and g_124302_(_033449_, _033452_, _033453_);
  or g_124303_(_033448_, _033451_, _033454_);
  and g_124304_(_010701_, _033454_, _033455_);
  or g_124305_(_010700_, _033453_, _033456_);
  and g_124306_(_010527_, _033410_, _033457_);
  or g_124307_(_010528_, _033411_, _033458_);
  and g_124308_(_033331_, _033411_, _033459_);
  or g_124309_(_033330_, _033410_, _033460_);
  and g_124310_(_033458_, _033460_, _033462_);
  or g_124311_(_033457_, _033459_, _033463_);
  and g_124312_(_010679_, _033463_, _033464_);
  or g_124313_(_010678_, _033462_, _033465_);
  and g_124314_(_033456_, _033465_, _033466_);
  or g_124315_(_033455_, _033464_, _033467_);
  and g_124316_(_010678_, _033462_, _033468_);
  or g_124317_(_010679_, _033463_, _033469_);
  and g_124318_(_010700_, _033453_, _033470_);
  or g_124319_(_010701_, _033454_, _033471_);
  and g_124320_(_033469_, _033471_, _033473_);
  or g_124321_(_033468_, _033470_, _033474_);
  and g_124322_(_033466_, _033473_, _033475_);
  or g_124323_(_033467_, _033474_, _033476_);
  and g_124324_(_033446_, _033475_, _033477_);
  or g_124325_(_033447_, _033476_, _033478_);
  or g_124326_(_010454_, _033411_, _033479_);
  or g_124327_(_033271_, _033410_, _033480_);
  and g_124328_(_033479_, _033480_, _033481_);
  and g_124329_(_010727_, _033481_, _033482_);
  not g_124330_(_033482_, _033484_);
  xor g_124331_(_010727_, _033481_, _033485_);
  xor g_124332_(_010726_, _033481_, _033486_);
  or g_124333_(_010470_, _033411_, _033487_);
  or g_124334_(_033265_, _033410_, _033488_);
  and g_124335_(_033487_, _033488_, _033489_);
  not g_124336_(_033489_, _033490_);
  and g_124337_(_010716_, _033490_, _033491_);
  not g_124338_(_033491_, _033492_);
  and g_124339_(_010717_, _033489_, _033493_);
  not g_124340_(_033493_, _033495_);
  and g_124341_(_033485_, _033495_, _033496_);
  or g_124342_(_033486_, _033493_, _033497_);
  and g_124343_(_033492_, _033496_, _033498_);
  or g_124344_(_033491_, _033497_, _033499_);
  and g_124345_(_010490_, _033410_, _033500_);
  or g_124346_(_010491_, _033411_, _033501_);
  and g_124347_(_033361_, _033411_, _033502_);
  or g_124348_(_033360_, _033410_, _033503_);
  and g_124349_(_033501_, _033503_, _033504_);
  or g_124350_(_033500_, _033502_, _033506_);
  and g_124351_(_010740_, _033506_, _033507_);
  or g_124352_(_010739_, _033504_, _033508_);
  and g_124353_(_010459_, _033410_, _033509_);
  or g_124354_(_010461_, _033411_, _033510_);
  and g_124355_(_033283_, _033411_, _033511_);
  or g_124356_(_033282_, _033410_, _033512_);
  and g_124357_(_033510_, _033512_, _033513_);
  or g_124358_(_033509_, _033511_, _033514_);
  and g_124359_(_010751_, _033514_, _033515_);
  or g_124360_(_010750_, _033513_, _033517_);
  and g_124361_(_033508_, _033517_, _033518_);
  or g_124362_(_033507_, _033515_, _033519_);
  and g_124363_(_010750_, _033513_, _033520_);
  or g_124364_(_010751_, _033514_, _033521_);
  and g_124365_(_010739_, _033504_, _033522_);
  or g_124366_(_010740_, _033506_, _033523_);
  and g_124367_(_033521_, _033523_, _033524_);
  or g_124368_(_033520_, _033522_, _033525_);
  and g_124369_(_033518_, _033524_, _033526_);
  or g_124370_(_033519_, _033525_, _033528_);
  and g_124371_(_033498_, _033526_, _033529_);
  or g_124372_(_033499_, _033528_, _033530_);
  and g_124373_(_033477_, _033529_, _033531_);
  or g_124374_(_033478_, _033530_, _033532_);
  or g_124375_(_010566_, _033411_, _033533_);
  or g_124376_(_033235_, _033410_, _033534_);
  and g_124377_(_033533_, _033534_, _033535_);
  not g_124378_(_033535_, _033536_);
  and g_124379_(_010776_, _033536_, _033537_);
  or g_124380_(_010777_, _033535_, _033539_);
  or g_124381_(_033240_, _033410_, _033540_);
  or g_124382_(_054005_, _033411_, _033541_);
  and g_124383_(_033540_, _033541_, _033542_);
  not g_124384_(_033542_, _033543_);
  and g_124385_(_054261_, _033542_, _033544_);
  or g_124386_(_054262_, _033543_, _033545_);
  and g_124387_(_033539_, _033545_, _033546_);
  or g_124388_(_033537_, _033544_, _033547_);
  and g_124389_(_010777_, _033535_, _033548_);
  or g_124390_(_010776_, _033536_, _033550_);
  and g_124391_(_054262_, _033543_, _033551_);
  or g_124392_(_054261_, _033542_, _033552_);
  and g_124393_(_033550_, _033552_, _033553_);
  or g_124394_(_033548_, _033551_, _033554_);
  and g_124395_(_033546_, _033553_, _033555_);
  or g_124396_(_033547_, _033554_, _033556_);
  or g_124397_(_054930_, _033411_, _033557_);
  or g_124398_(_033249_, _033410_, _033558_);
  and g_124399_(_033557_, _033558_, _033559_);
  and g_124400_(out[561], _033559_, _033561_);
  not g_124401_(_033561_, _033562_);
  and g_124402_(out[560], _033418_, _033563_);
  or g_124403_(_055073_, _033416_, _033564_);
  xor g_124404_(out[561], _033559_, _033565_);
  xor g_124405_(_055062_, _033559_, _033566_);
  and g_124406_(_033564_, _033565_, _033567_);
  or g_124407_(_033563_, _033566_, _033568_);
  and g_124408_(_033562_, _033568_, _033569_);
  or g_124409_(_033561_, _033567_, _033570_);
  and g_124410_(_033555_, _033570_, _033572_);
  or g_124411_(_033556_, _033569_, _033573_);
  and g_124412_(_033547_, _033550_, _033574_);
  or g_124413_(_033546_, _033548_, _033575_);
  and g_124414_(_033573_, _033575_, _033576_);
  or g_124415_(_033572_, _033574_, _033577_);
  and g_124416_(_033531_, _033577_, _033578_);
  or g_124417_(_033532_, _033576_, _033579_);
  or g_124418_(_033518_, _033520_, _033580_);
  and g_124419_(_033498_, _033519_, _033581_);
  and g_124420_(_033521_, _033581_, _033583_);
  or g_124421_(_033499_, _033580_, _033584_);
  and g_124422_(_033482_, _033495_, _033585_);
  or g_124423_(_033484_, _033493_, _033586_);
  and g_124424_(_033492_, _033586_, _033587_);
  or g_124425_(_033491_, _033585_, _033588_);
  and g_124426_(_033584_, _033587_, _033589_);
  or g_124427_(_033583_, _033588_, _033590_);
  and g_124428_(_033477_, _033590_, _033591_);
  or g_124429_(_033478_, _033589_, _033592_);
  and g_124430_(_033438_, _033443_, _033594_);
  or g_124431_(_033437_, _033442_, _033595_);
  and g_124432_(_033467_, _033469_, _033596_);
  or g_124433_(_033466_, _033468_, _033597_);
  and g_124434_(_033446_, _033596_, _033598_);
  or g_124435_(_033447_, _033597_, _033599_);
  and g_124436_(_033595_, _033599_, _033600_);
  or g_124437_(_033594_, _033598_, _033601_);
  and g_124438_(_033579_, _033600_, _033602_);
  or g_124439_(_033578_, _033601_, _033603_);
  and g_124440_(_033592_, _033602_, _033605_);
  or g_124441_(_033591_, _033603_, _033606_);
  and g_124442_(_055073_, _033416_, _033607_);
  or g_124443_(out[560], _033418_, _033608_);
  and g_124444_(_033555_, _033608_, _033609_);
  or g_124445_(_033556_, _033607_, _033610_);
  and g_124446_(_033567_, _033609_, _033611_);
  or g_124447_(_033568_, _033610_, _033612_);
  and g_124448_(_033531_, _033611_, _033613_);
  or g_124449_(_033532_, _033612_, _033614_);
  and g_124450_(_033606_, _033614_, _033616_);
  or g_124451_(_033605_, _033613_, _033617_);
  and g_124452_(_033418_, _033617_, _033618_);
  not g_124453_(_033618_, _033619_);
  or g_124454_(out[560], _033617_, _033620_);
  not g_124455_(_033620_, _033621_);
  and g_124456_(_033619_, _033620_, _033622_);
  or g_124457_(_033618_, _033621_, _033623_);
  or g_124458_(_010726_, _033617_, _033624_);
  or g_124459_(_033481_, _033616_, _033625_);
  and g_124460_(_033624_, _033625_, _033627_);
  not g_124461_(_033627_, _033628_);
  and g_124462_(_010940_, _033628_, _033629_);
  or g_124463_(_010941_, _033627_, _033630_);
  and g_124464_(_010750_, _033616_, _033631_);
  or g_124465_(_010751_, _033617_, _033632_);
  and g_124466_(_033514_, _033617_, _033633_);
  or g_124467_(_033513_, _033616_, _033634_);
  and g_124468_(_033632_, _033634_, _033635_);
  or g_124469_(_033631_, _033633_, _033636_);
  and g_124470_(_010954_, _033635_, _033638_);
  or g_124471_(_010956_, _033636_, _033639_);
  and g_124472_(_033630_, _033639_, _033640_);
  or g_124473_(_033629_, _033638_, _033641_);
  or g_124474_(_010716_, _033617_, _033642_);
  or g_124475_(_033489_, _033616_, _033643_);
  and g_124476_(_033642_, _033643_, _033644_);
  not g_124477_(_033644_, _033645_);
  and g_124478_(_010934_, _033645_, _033646_);
  or g_124479_(_010935_, _033644_, _033647_);
  and g_124480_(_010941_, _033627_, _033649_);
  or g_124481_(_010940_, _033628_, _033650_);
  and g_124482_(_010935_, _033644_, _033651_);
  or g_124483_(_010934_, _033645_, _033652_);
  and g_124484_(_033650_, _033652_, _033653_);
  or g_124485_(_033649_, _033651_, _033654_);
  and g_124486_(_033647_, _033653_, _033655_);
  or g_124487_(_033646_, _033654_, _033656_);
  and g_124488_(_033640_, _033655_, _033657_);
  or g_124489_(_033641_, _033656_, _033658_);
  and g_124490_(_010739_, _033616_, _033660_);
  or g_124491_(_010740_, _033617_, _033661_);
  and g_124492_(_033506_, _033617_, _033662_);
  or g_124493_(_033504_, _033616_, _033663_);
  and g_124494_(_033661_, _033663_, _033664_);
  or g_124495_(_033660_, _033662_, _033665_);
  and g_124496_(_010969_, _033665_, _033666_);
  or g_124497_(_010968_, _033664_, _033667_);
  and g_124498_(_010956_, _033636_, _033668_);
  or g_124499_(_010954_, _033635_, _033669_);
  and g_124500_(_033667_, _033669_, _033671_);
  or g_124501_(_033666_, _033668_, _033672_);
  and g_124502_(_010968_, _033664_, _033673_);
  or g_124503_(_010969_, _033665_, _033674_);
  and g_124504_(_033671_, _033674_, _033675_);
  or g_124505_(_033672_, _033673_, _033676_);
  and g_124506_(_033657_, _033675_, _033677_);
  or g_124507_(_033658_, _033676_, _033678_);
  or g_124508_(_010776_, _033617_, _033679_);
  or g_124509_(_033535_, _033616_, _033680_);
  and g_124510_(_033679_, _033680_, _033682_);
  not g_124511_(_033682_, _033683_);
  and g_124512_(_011003_, _033682_, _033684_);
  or g_124513_(_011002_, _033683_, _033685_);
  or g_124514_(_054262_, _033617_, _033686_);
  not g_124515_(_033686_, _033687_);
  and g_124516_(_033543_, _033617_, _033688_);
  not g_124517_(_033688_, _033689_);
  and g_124518_(_033686_, _033689_, _033690_);
  or g_124519_(_033687_, _033688_, _033691_);
  and g_124520_(_054572_, _033691_, _033693_);
  or g_124521_(_054571_, _033690_, _033694_);
  and g_124522_(_033685_, _033694_, _033695_);
  or g_124523_(_033684_, _033693_, _033696_);
  and g_124524_(_011002_, _033683_, _033697_);
  or g_124525_(_011003_, _033682_, _033698_);
  and g_124526_(_054571_, _033690_, _033699_);
  or g_124527_(_054572_, _033691_, _033700_);
  and g_124528_(_033698_, _033700_, _033701_);
  or g_124529_(_033697_, _033699_, _033702_);
  and g_124530_(_033695_, _033701_, _033704_);
  or g_124531_(_033696_, _033702_, _033705_);
  and g_124532_(_033677_, _033704_, _033706_);
  or g_124533_(_033678_, _033705_, _033707_);
  or g_124534_(_055205_, _033622_, _033708_);
  or g_124535_(_055062_, _033617_, _033709_);
  or g_124536_(_033559_, _033616_, _033710_);
  and g_124537_(_033709_, _033710_, _033711_);
  and g_124538_(out[577], _033711_, _033712_);
  xor g_124539_(out[577], _033711_, _033713_);
  and g_124540_(_033708_, _033713_, _033715_);
  and g_124541_(_033706_, _033715_, _033716_);
  or g_124542_(out[576], _033623_, _033717_);
  or g_124543_(_033434_, _033617_, _033718_);
  not g_124544_(_033718_, _033719_);
  and g_124545_(_033432_, _033617_, _033720_);
  not g_124546_(_033720_, _033721_);
  and g_124547_(_033718_, _033721_, _033722_);
  or g_124548_(_033719_, _033720_, _033723_);
  or g_124549_(out[586], _010888_, _033724_);
  xor g_124550_(out[586], _010888_, _033726_);
  xor g_124551_(_055260_, _010888_, _033727_);
  and g_124552_(_033722_, _033726_, _033728_);
  or g_124553_(_033723_, _033727_, _033729_);
  and g_124554_(_033419_, _033422_, _033730_);
  or g_124555_(_033420_, _033423_, _033731_);
  xor g_124556_(out[587], _033724_, _033732_);
  xor g_124557_(_055139_, _033724_, _033733_);
  and g_124558_(_033730_, _033733_, _033734_);
  or g_124559_(_033731_, _033732_, _033735_);
  and g_124560_(_033729_, _033735_, _033737_);
  or g_124561_(_033728_, _033734_, _033738_);
  and g_124562_(_033731_, _033732_, _033739_);
  or g_124563_(_033730_, _033733_, _033740_);
  and g_124564_(_033723_, _033727_, _033741_);
  or g_124565_(_033722_, _033726_, _033742_);
  and g_124566_(_033740_, _033742_, _033743_);
  or g_124567_(_033739_, _033741_, _033744_);
  and g_124568_(_033737_, _033743_, _033745_);
  or g_124569_(_033738_, _033744_, _033746_);
  or g_124570_(_010679_, _033617_, _033748_);
  not g_124571_(_033748_, _033749_);
  and g_124572_(_033463_, _033617_, _033750_);
  not g_124573_(_033750_, _033751_);
  and g_124574_(_033748_, _033751_, _033752_);
  or g_124575_(_033749_, _033750_, _033753_);
  and g_124576_(_010891_, _033753_, _033754_);
  or g_124577_(_010890_, _033752_, _033755_);
  or g_124578_(_010701_, _033617_, _033756_);
  not g_124579_(_033756_, _033757_);
  and g_124580_(_033454_, _033617_, _033759_);
  not g_124581_(_033759_, _033760_);
  and g_124582_(_033756_, _033760_, _033761_);
  or g_124583_(_033757_, _033759_, _033762_);
  and g_124584_(_010908_, _033762_, _033763_);
  or g_124585_(_010907_, _033761_, _033764_);
  and g_124586_(_033755_, _033764_, _033765_);
  or g_124587_(_033754_, _033763_, _033766_);
  and g_124588_(_010890_, _033752_, _033767_);
  or g_124589_(_010891_, _033753_, _033768_);
  and g_124590_(_010907_, _033761_, _033770_);
  or g_124591_(_010908_, _033762_, _033771_);
  and g_124592_(_033768_, _033771_, _033772_);
  or g_124593_(_033767_, _033770_, _033773_);
  and g_124594_(_033765_, _033772_, _033774_);
  or g_124595_(_033766_, _033773_, _033775_);
  and g_124596_(_033745_, _033774_, _033776_);
  or g_124597_(_033746_, _033775_, _033777_);
  and g_124598_(_033717_, _033776_, _033778_);
  and g_124599_(_033716_, _033778_, _033779_);
  not g_124600_(_033779_, _033781_);
  and g_124601_(_033685_, _033702_, _033782_);
  or g_124602_(_033684_, _033701_, _033783_);
  and g_124603_(_033677_, _033782_, _033784_);
  or g_124604_(_033678_, _033783_, _033785_);
  and g_124605_(_033657_, _033672_, _033786_);
  or g_124606_(_033658_, _033671_, _033787_);
  and g_124607_(_033649_, _033652_, _033788_);
  or g_124608_(_033650_, _033651_, _033789_);
  and g_124609_(_033647_, _033789_, _033790_);
  or g_124610_(_033646_, _033788_, _033792_);
  and g_124611_(_033787_, _033790_, _033793_);
  or g_124612_(_033786_, _033792_, _033794_);
  and g_124613_(_033785_, _033793_, _033795_);
  or g_124614_(_033784_, _033794_, _033796_);
  or g_124615_(_033712_, _033715_, _033797_);
  not g_124616_(_033797_, _033798_);
  and g_124617_(_033706_, _033797_, _033799_);
  or g_124618_(_033707_, _033798_, _033800_);
  and g_124619_(_033795_, _033800_, _033801_);
  or g_124620_(_033796_, _033799_, _033803_);
  and g_124621_(_033776_, _033803_, _033804_);
  or g_124622_(_033777_, _033801_, _033805_);
  and g_124623_(_033766_, _033768_, _033806_);
  or g_124624_(_033765_, _033767_, _033807_);
  and g_124625_(_033745_, _033806_, _033808_);
  or g_124626_(_033746_, _033807_, _033809_);
  and g_124627_(_033738_, _033740_, _033810_);
  or g_124628_(_033737_, _033739_, _033811_);
  and g_124629_(_033809_, _033811_, _033812_);
  or g_124630_(_033808_, _033810_, _033814_);
  and g_124631_(_033805_, _033812_, _033815_);
  or g_124632_(_033804_, _033814_, _033816_);
  and g_124633_(_033781_, _033816_, _033817_);
  or g_124634_(_033779_, _033815_, _033818_);
  and g_124635_(_033623_, _033818_, _033819_);
  or g_124636_(_033622_, _033817_, _033820_);
  and g_124637_(_055205_, _033817_, _033821_);
  or g_124638_(out[576], _033818_, _033822_);
  and g_124639_(_033820_, _033822_, _033823_);
  or g_124640_(_033819_, _033821_, _033825_);
  and g_124641_(_033730_, _033732_, _033826_);
  or g_124642_(_033731_, _033733_, _033827_);
  or g_124643_(out[602], _011111_, _033828_);
  xor g_124644_(out[603], _033828_, _033829_);
  xor g_124645_(_055271_, _033828_, _033830_);
  and g_124646_(_033826_, _033830_, _033831_);
  or g_124647_(_033827_, _033829_, _033832_);
  and g_124648_(_033726_, _033817_, _033833_);
  or g_124649_(_033727_, _033818_, _033834_);
  and g_124650_(_033723_, _033818_, _033836_);
  or g_124651_(_033722_, _033817_, _033837_);
  and g_124652_(_033834_, _033837_, _033838_);
  or g_124653_(_033833_, _033836_, _033839_);
  xor g_124654_(out[602], _011111_, _033840_);
  xor g_124655_(_055392_, _011111_, _033841_);
  and g_124656_(_033838_, _033840_, _033842_);
  or g_124657_(_033839_, _033841_, _033843_);
  and g_124658_(_033832_, _033843_, _033844_);
  or g_124659_(_033831_, _033842_, _033845_);
  and g_124660_(_033839_, _033841_, _033847_);
  or g_124661_(_033838_, _033840_, _033848_);
  and g_124662_(_033827_, _033829_, _033849_);
  or g_124663_(_033826_, _033830_, _033850_);
  and g_124664_(_033848_, _033850_, _033851_);
  or g_124665_(_033847_, _033849_, _033852_);
  and g_124666_(_033844_, _033851_, _033853_);
  or g_124667_(_033845_, _033852_, _033854_);
  and g_124668_(_010907_, _033817_, _033855_);
  or g_124669_(_010908_, _033818_, _033856_);
  and g_124670_(_033762_, _033818_, _033858_);
  or g_124671_(_033761_, _033817_, _033859_);
  and g_124672_(_033856_, _033859_, _033860_);
  or g_124673_(_033855_, _033858_, _033861_);
  and g_124674_(_011133_, _033861_, _033862_);
  or g_124675_(_011132_, _033860_, _033863_);
  and g_124676_(_010890_, _033817_, _033864_);
  or g_124677_(_010891_, _033818_, _033865_);
  and g_124678_(_033753_, _033818_, _033866_);
  or g_124679_(_033752_, _033817_, _033867_);
  and g_124680_(_033865_, _033867_, _033869_);
  or g_124681_(_033864_, _033866_, _033870_);
  and g_124682_(_011113_, _033870_, _033871_);
  or g_124683_(_011112_, _033869_, _033872_);
  and g_124684_(_033863_, _033872_, _033873_);
  or g_124685_(_033862_, _033871_, _033874_);
  and g_124686_(_011112_, _033869_, _033875_);
  or g_124687_(_011113_, _033870_, _033876_);
  and g_124688_(_011132_, _033860_, _033877_);
  or g_124689_(_011133_, _033861_, _033878_);
  and g_124690_(_033876_, _033878_, _033880_);
  or g_124691_(_033875_, _033877_, _033881_);
  and g_124692_(_033873_, _033880_, _033882_);
  or g_124693_(_033874_, _033881_, _033883_);
  and g_124694_(_033853_, _033882_, _033884_);
  or g_124695_(_033854_, _033883_, _033885_);
  and g_124696_(_010935_, _033817_, _033886_);
  or g_124697_(_010934_, _033818_, _033887_);
  and g_124698_(_033645_, _033818_, _033888_);
  or g_124699_(_033644_, _033817_, _033889_);
  and g_124700_(_033887_, _033889_, _033891_);
  or g_124701_(_033886_, _033888_, _033892_);
  and g_124702_(_011146_, _033892_, _033893_);
  or g_124703_(_010940_, _033818_, _033894_);
  or g_124704_(_033627_, _033817_, _033895_);
  and g_124705_(_033894_, _033895_, _033896_);
  or g_124706_(_011146_, _033892_, _033897_);
  and g_124707_(_011154_, _033896_, _033898_);
  xor g_124708_(_011147_, _033891_, _033899_);
  xor g_124709_(_011146_, _033891_, _033900_);
  xor g_124710_(_011154_, _033896_, _033902_);
  xor g_124711_(_011152_, _033896_, _033903_);
  and g_124712_(_033899_, _033902_, _033904_);
  or g_124713_(_033900_, _033903_, _033905_);
  and g_124714_(_010968_, _033817_, _033906_);
  or g_124715_(_010969_, _033818_, _033907_);
  and g_124716_(_033665_, _033818_, _033908_);
  or g_124717_(_033664_, _033817_, _033909_);
  and g_124718_(_033907_, _033909_, _033910_);
  or g_124719_(_033906_, _033908_, _033911_);
  and g_124720_(_010954_, _033817_, _033913_);
  or g_124721_(_010956_, _033818_, _033914_);
  and g_124722_(_033636_, _033818_, _033915_);
  or g_124723_(_033635_, _033817_, _033916_);
  and g_124724_(_033914_, _033916_, _033917_);
  or g_124725_(_033913_, _033915_, _033918_);
  and g_124726_(_011168_, _033918_, _033919_);
  or g_124727_(_011167_, _033917_, _033920_);
  and g_124728_(_011167_, _033917_, _033921_);
  or g_124729_(_011168_, _033918_, _033922_);
  and g_124730_(_011181_, _033911_, _033924_);
  or g_124731_(_011180_, _033910_, _033925_);
  and g_124732_(_033920_, _033922_, _033926_);
  or g_124733_(_033919_, _033921_, _033927_);
  xor g_124734_(_011180_, _033910_, _033928_);
  xor g_124735_(_011181_, _033910_, _033929_);
  and g_124736_(_033926_, _033928_, _033930_);
  or g_124737_(_033927_, _033929_, _033931_);
  and g_124738_(_033904_, _033930_, _033932_);
  or g_124739_(_033905_, _033931_, _033933_);
  or g_124740_(_011002_, _033818_, _033935_);
  or g_124741_(_033682_, _033817_, _033936_);
  and g_124742_(_033935_, _033936_, _033937_);
  or g_124743_(_011232_, _033937_, _033938_);
  and g_124744_(_033691_, _033818_, _033939_);
  and g_124745_(_054571_, _033817_, _033940_);
  or g_124746_(_033939_, _033940_, _033941_);
  and g_124747_(_011232_, _033937_, _033942_);
  or g_124748_(_054793_, _033941_, _033943_);
  xor g_124749_(_011232_, _033937_, _033944_);
  xor g_124750_(_011231_, _033937_, _033946_);
  xor g_124751_(_054793_, _033941_, _033947_);
  xor g_124752_(_054792_, _033941_, _033948_);
  and g_124753_(_033944_, _033947_, _033949_);
  or g_124754_(_033946_, _033948_, _033950_);
  or g_124755_(_055194_, _033818_, _033951_);
  or g_124756_(_033711_, _033817_, _033952_);
  and g_124757_(_033951_, _033952_, _033953_);
  and g_124758_(out[593], _033953_, _033954_);
  not g_124759_(_033954_, _033955_);
  and g_124760_(out[592], _033825_, _033957_);
  or g_124761_(_055337_, _033823_, _033958_);
  xor g_124762_(out[593], _033953_, _033959_);
  xor g_124763_(_055326_, _033953_, _033960_);
  and g_124764_(_033958_, _033959_, _033961_);
  or g_124765_(_033957_, _033960_, _033962_);
  and g_124766_(_033955_, _033962_, _033963_);
  or g_124767_(_033954_, _033961_, _033964_);
  and g_124768_(_033949_, _033964_, _033965_);
  or g_124769_(_033950_, _033963_, _033966_);
  or g_124770_(_033942_, _033943_, _033968_);
  and g_124771_(_033938_, _033968_, _033969_);
  not g_124772_(_033969_, _033970_);
  and g_124773_(_033966_, _033969_, _033971_);
  or g_124774_(_033965_, _033970_, _033972_);
  and g_124775_(_033932_, _033972_, _033973_);
  or g_124776_(_033933_, _033971_, _033974_);
  and g_124777_(_033920_, _033925_, _033975_);
  or g_124778_(_033919_, _033924_, _033976_);
  and g_124779_(_033922_, _033976_, _033977_);
  or g_124780_(_033921_, _033975_, _033979_);
  and g_124781_(_033904_, _033977_, _033980_);
  or g_124782_(_033905_, _033979_, _033981_);
  and g_124783_(_033897_, _033898_, _033982_);
  or g_124784_(_033893_, _033982_, _033983_);
  not g_124785_(_033983_, _033984_);
  and g_124786_(_033981_, _033984_, _033985_);
  or g_124787_(_033980_, _033983_, _033986_);
  and g_124788_(_033974_, _033985_, _033987_);
  or g_124789_(_033973_, _033986_, _033988_);
  and g_124790_(_033884_, _033988_, _033990_);
  or g_124791_(_033885_, _033987_, _033991_);
  and g_124792_(_033874_, _033876_, _033992_);
  or g_124793_(_033873_, _033875_, _033993_);
  and g_124794_(_033853_, _033992_, _033994_);
  or g_124795_(_033854_, _033993_, _033995_);
  and g_124796_(_033845_, _033850_, _033996_);
  or g_124797_(_033844_, _033849_, _033997_);
  and g_124798_(_033995_, _033997_, _033998_);
  or g_124799_(_033994_, _033996_, _033999_);
  and g_124800_(_033991_, _033998_, _034001_);
  or g_124801_(_033990_, _033999_, _034002_);
  and g_124802_(_055337_, _033823_, _034003_);
  or g_124803_(out[592], _033825_, _034004_);
  and g_124804_(_033961_, _034004_, _034005_);
  or g_124805_(_033962_, _034003_, _034006_);
  and g_124806_(_033949_, _034005_, _034007_);
  or g_124807_(_033950_, _034006_, _034008_);
  and g_124808_(_033932_, _034007_, _034009_);
  or g_124809_(_033933_, _034008_, _034010_);
  and g_124810_(_033884_, _034009_, _034012_);
  or g_124811_(_033885_, _034010_, _034013_);
  and g_124812_(_034002_, _034013_, _034014_);
  or g_124813_(_034001_, _034012_, _034015_);
  and g_124814_(_033825_, _034015_, _034016_);
  or g_124815_(_033823_, _034014_, _034017_);
  and g_124816_(_055337_, _034014_, _034018_);
  or g_124817_(out[592], _034015_, _034019_);
  and g_124818_(_034017_, _034019_, _034020_);
  or g_124819_(_034016_, _034018_, _034021_);
  and g_124820_(_033826_, _033829_, _034023_);
  or g_124821_(_033827_, _033830_, _034024_);
  or g_124822_(out[618], _011321_, _034025_);
  xor g_124823_(out[619], _034025_, _034026_);
  xor g_124824_(_055403_, _034025_, _034027_);
  and g_124825_(_034023_, _034027_, _034028_);
  or g_124826_(_034024_, _034026_, _034029_);
  and g_124827_(_033840_, _034014_, _034030_);
  not g_124828_(_034030_, _034031_);
  or g_124829_(_033838_, _034014_, _034032_);
  not g_124830_(_034032_, _034034_);
  and g_124831_(_034031_, _034032_, _034035_);
  or g_124832_(_034030_, _034034_, _034036_);
  xor g_124833_(out[618], _011321_, _034037_);
  xor g_124834_(_055524_, _011321_, _034038_);
  and g_124835_(_034035_, _034037_, _034039_);
  or g_124836_(_034036_, _034038_, _034040_);
  and g_124837_(_034029_, _034040_, _034041_);
  or g_124838_(_034028_, _034039_, _034042_);
  and g_124839_(_034024_, _034026_, _034043_);
  or g_124840_(_034023_, _034027_, _034045_);
  and g_124841_(_034036_, _034038_, _034046_);
  or g_124842_(_034035_, _034037_, _034047_);
  and g_124843_(_034045_, _034047_, _034048_);
  or g_124844_(_034043_, _034046_, _034049_);
  and g_124845_(_011112_, _034014_, _034050_);
  not g_124846_(_034050_, _034051_);
  or g_124847_(_033869_, _034014_, _034052_);
  not g_124848_(_034052_, _034053_);
  and g_124849_(_034051_, _034052_, _034054_);
  or g_124850_(_034050_, _034053_, _034056_);
  and g_124851_(_011322_, _034054_, _034057_);
  or g_124852_(_011323_, _034056_, _034058_);
  and g_124853_(_034048_, _034058_, _034059_);
  or g_124854_(_034049_, _034057_, _034060_);
  and g_124855_(_034041_, _034059_, _034061_);
  or g_124856_(_034042_, _034060_, _034062_);
  and g_124857_(_011323_, _034056_, _034063_);
  or g_124858_(_011322_, _034054_, _034064_);
  and g_124859_(_011132_, _034014_, _034065_);
  not g_124860_(_034065_, _034067_);
  or g_124861_(_033860_, _034014_, _034068_);
  not g_124862_(_034068_, _034069_);
  and g_124863_(_034067_, _034068_, _034070_);
  or g_124864_(_034065_, _034069_, _034071_);
  and g_124865_(_011320_, _034071_, _034072_);
  or g_124866_(_011319_, _034070_, _034073_);
  and g_124867_(_034064_, _034073_, _034074_);
  or g_124868_(_034063_, _034072_, _034075_);
  and g_124869_(_011319_, _034070_, _034076_);
  or g_124870_(_011320_, _034071_, _034078_);
  and g_124871_(_034074_, _034078_, _034079_);
  or g_124872_(_034075_, _034076_, _034080_);
  and g_124873_(_034061_, _034079_, _034081_);
  or g_124874_(_034062_, _034080_, _034082_);
  and g_124875_(_011147_, _034014_, _034083_);
  or g_124876_(_011146_, _034015_, _034084_);
  and g_124877_(_033892_, _034015_, _034085_);
  or g_124878_(_033891_, _034014_, _034086_);
  and g_124879_(_034084_, _034086_, _034087_);
  or g_124880_(_034083_, _034085_, _034089_);
  and g_124881_(_011341_, _034089_, _034090_);
  or g_124882_(_011342_, _034087_, _034091_);
  and g_124883_(_011154_, _034014_, _034092_);
  not g_124884_(_034092_, _034093_);
  or g_124885_(_033896_, _034014_, _034094_);
  not g_124886_(_034094_, _034095_);
  and g_124887_(_034093_, _034094_, _034096_);
  or g_124888_(_034092_, _034095_, _034097_);
  and g_124889_(_011350_, _034097_, _034098_);
  or g_124890_(_034090_, _034098_, _034100_);
  and g_124891_(_011352_, _034096_, _034101_);
  or g_124892_(_011350_, _034097_, _034102_);
  and g_124893_(_011342_, _034087_, _034103_);
  or g_124894_(_011341_, _034089_, _034104_);
  and g_124895_(_011167_, _034014_, _034105_);
  not g_124896_(_034105_, _034106_);
  or g_124897_(_033917_, _034014_, _034107_);
  not g_124898_(_034107_, _034108_);
  and g_124899_(_034106_, _034107_, _034109_);
  or g_124900_(_034105_, _034108_, _034111_);
  and g_124901_(_011375_, _034109_, _034112_);
  or g_124902_(_011376_, _034111_, _034113_);
  or g_124903_(_034103_, _034112_, _034114_);
  or g_124904_(_034101_, _034114_, _034115_);
  and g_124905_(_034091_, _034104_, _034116_);
  xor g_124906_(_011352_, _034096_, _034117_);
  and g_124907_(_034116_, _034117_, _034118_);
  and g_124908_(_034113_, _034118_, _034119_);
  or g_124909_(_034100_, _034115_, _034120_);
  and g_124910_(_011180_, _034014_, _034122_);
  not g_124911_(_034122_, _034123_);
  or g_124912_(_033910_, _034014_, _034124_);
  not g_124913_(_034124_, _034125_);
  and g_124914_(_034123_, _034124_, _034126_);
  or g_124915_(_034122_, _034125_, _034127_);
  and g_124916_(_011365_, _034127_, _034128_);
  or g_124917_(_011364_, _034126_, _034129_);
  and g_124918_(_011376_, _034111_, _034130_);
  or g_124919_(_011375_, _034109_, _034131_);
  and g_124920_(_034129_, _034131_, _034133_);
  or g_124921_(_034128_, _034130_, _034134_);
  and g_124922_(_011364_, _034126_, _034135_);
  or g_124923_(_011365_, _034127_, _034136_);
  and g_124924_(_034133_, _034136_, _034137_);
  or g_124925_(_034134_, _034135_, _034138_);
  and g_124926_(_034119_, _034137_, _034139_);
  or g_124927_(_034120_, _034138_, _034140_);
  or g_124928_(_011231_, _034015_, _034141_);
  or g_124929_(_033937_, _034014_, _034142_);
  and g_124930_(_034141_, _034142_, _034144_);
  or g_124931_(_011402_, _034144_, _034145_);
  and g_124932_(_011402_, _034144_, _034146_);
  xor g_124933_(_011402_, _034144_, _034147_);
  xor g_124934_(_011401_, _034144_, _034148_);
  and g_124935_(_033941_, _034015_, _034149_);
  and g_124936_(_054792_, _034014_, _034150_);
  or g_124937_(_034149_, _034150_, _034151_);
  or g_124938_(_054979_, _034151_, _034152_);
  xor g_124939_(_054979_, _034151_, _034153_);
  xor g_124940_(_054978_, _034151_, _034155_);
  and g_124941_(_034147_, _034153_, _034156_);
  or g_124942_(_034148_, _034155_, _034157_);
  or g_124943_(_055326_, _034015_, _034158_);
  or g_124944_(_033953_, _034014_, _034159_);
  and g_124945_(_034158_, _034159_, _034160_);
  and g_124946_(out[609], _034160_, _034161_);
  not g_124947_(_034161_, _034162_);
  and g_124948_(out[608], _034021_, _034163_);
  or g_124949_(_055469_, _034020_, _034164_);
  xor g_124950_(out[609], _034160_, _034166_);
  xor g_124951_(_055458_, _034160_, _034167_);
  and g_124952_(_034164_, _034166_, _034168_);
  or g_124953_(_034163_, _034167_, _034169_);
  and g_124954_(_034162_, _034169_, _034170_);
  or g_124955_(_034161_, _034168_, _034171_);
  and g_124956_(_034156_, _034171_, _034172_);
  or g_124957_(_034157_, _034170_, _034173_);
  and g_124958_(_034145_, _034152_, _034174_);
  or g_124959_(_034146_, _034174_, _034175_);
  not g_124960_(_034175_, _034177_);
  and g_124961_(_034173_, _034175_, _034178_);
  or g_124962_(_034172_, _034177_, _034179_);
  and g_124963_(_034139_, _034179_, _034180_);
  or g_124964_(_034140_, _034178_, _034181_);
  and g_124965_(_034119_, _034134_, _034182_);
  or g_124966_(_034120_, _034133_, _034183_);
  and g_124967_(_034101_, _034104_, _034184_);
  or g_124968_(_034102_, _034103_, _034185_);
  and g_124969_(_034091_, _034185_, _034186_);
  or g_124970_(_034090_, _034184_, _034188_);
  and g_124971_(_034183_, _034186_, _034189_);
  or g_124972_(_034182_, _034188_, _034190_);
  and g_124973_(_034181_, _034189_, _034191_);
  or g_124974_(_034180_, _034190_, _034192_);
  and g_124975_(_034081_, _034192_, _034193_);
  or g_124976_(_034082_, _034191_, _034194_);
  and g_124977_(_034061_, _034075_, _034195_);
  or g_124978_(_034062_, _034074_, _034196_);
  and g_124979_(_034042_, _034045_, _034197_);
  or g_124980_(_034041_, _034043_, _034199_);
  and g_124981_(_034196_, _034199_, _034200_);
  or g_124982_(_034195_, _034197_, _034201_);
  and g_124983_(_034194_, _034200_, _034202_);
  or g_124984_(_034193_, _034201_, _034203_);
  and g_124985_(_055469_, _034020_, _034204_);
  or g_124986_(out[608], _034021_, _034205_);
  and g_124987_(_034156_, _034205_, _034206_);
  or g_124988_(_034157_, _034204_, _034207_);
  and g_124989_(_034168_, _034206_, _034208_);
  or g_124990_(_034169_, _034207_, _034210_);
  and g_124991_(_034139_, _034208_, _034211_);
  or g_124992_(_034140_, _034210_, _034212_);
  and g_124993_(_034081_, _034211_, _034213_);
  or g_124994_(_034082_, _034212_, _034214_);
  and g_124995_(_034203_, _034214_, _034215_);
  or g_124996_(_034202_, _034213_, _034216_);
  and g_124997_(_034021_, _034216_, _034217_);
  or g_124998_(_034020_, _034215_, _034218_);
  and g_124999_(_055469_, _034215_, _034219_);
  or g_125000_(out[608], _034216_, _034221_);
  and g_125001_(_034218_, _034221_, _034222_);
  or g_125002_(_034217_, _034219_, _034223_);
  and g_125003_(_011322_, _034215_, _034224_);
  or g_125004_(_011323_, _034216_, _034225_);
  and g_125005_(_034056_, _034216_, _034226_);
  or g_125006_(_034054_, _034215_, _034227_);
  and g_125007_(_034225_, _034227_, _034228_);
  or g_125008_(_034224_, _034226_, _034229_);
  and g_125009_(_011507_, _034229_, _034230_);
  or g_125010_(_011506_, _034228_, _034232_);
  and g_125011_(_011319_, _034215_, _034233_);
  or g_125012_(_011320_, _034216_, _034234_);
  and g_125013_(_034071_, _034216_, _034235_);
  or g_125014_(_034070_, _034215_, _034236_);
  and g_125015_(_034234_, _034236_, _034237_);
  or g_125016_(_034233_, _034235_, _034238_);
  and g_125017_(_011529_, _034238_, _034239_);
  or g_125018_(_011528_, _034237_, _034240_);
  and g_125019_(_034232_, _034240_, _034241_);
  or g_125020_(_034230_, _034239_, _034243_);
  and g_125021_(_034151_, _034216_, _034244_);
  not g_125022_(_034244_, _034245_);
  and g_125023_(_054978_, _034215_, _034246_);
  or g_125024_(_054979_, _034216_, _034247_);
  and g_125025_(_034245_, _034247_, _034248_);
  or g_125026_(_034244_, _034246_, _034249_);
  and g_125027_(_055091_, _034248_, _034250_);
  or g_125028_(_055092_, _034249_, _034251_);
  or g_125029_(_011401_, _034216_, _034252_);
  or g_125030_(_034144_, _034215_, _034254_);
  and g_125031_(_034252_, _034254_, _034255_);
  not g_125032_(_034255_, _034256_);
  and g_125033_(_011613_, _034256_, _034257_);
  or g_125034_(_011614_, _034255_, _034258_);
  and g_125035_(_034251_, _034258_, _034259_);
  or g_125036_(_034250_, _034257_, _034260_);
  or g_125037_(_055458_, _034216_, _034261_);
  or g_125038_(_034160_, _034215_, _034262_);
  and g_125039_(_034261_, _034262_, _034263_);
  and g_125040_(out[625], _034263_, _034265_);
  not g_125041_(_034265_, _034266_);
  and g_125042_(out[624], _034223_, _034267_);
  or g_125043_(_055601_, _034222_, _034268_);
  xor g_125044_(out[625], _034263_, _034269_);
  xor g_125045_(_055590_, _034263_, _034270_);
  and g_125046_(_034268_, _034269_, _034271_);
  or g_125047_(_034267_, _034270_, _034272_);
  and g_125048_(_034266_, _034272_, _034273_);
  or g_125049_(_034265_, _034271_, _034274_);
  and g_125050_(_055092_, _034249_, _034276_);
  or g_125051_(_055091_, _034248_, _034277_);
  and g_125052_(_034274_, _034277_, _034278_);
  or g_125053_(_034273_, _034276_, _034279_);
  and g_125054_(_034259_, _034277_, _034280_);
  and g_125055_(_034259_, _034279_, _034281_);
  or g_125056_(_034260_, _034278_, _034282_);
  and g_125057_(_011342_, _034215_, _034283_);
  or g_125058_(_011341_, _034216_, _034284_);
  and g_125059_(_034089_, _034216_, _034285_);
  or g_125060_(_034087_, _034215_, _034287_);
  and g_125061_(_034284_, _034287_, _034288_);
  or g_125062_(_034283_, _034285_, _034289_);
  and g_125063_(_011556_, _034289_, _034290_);
  or g_125064_(_011557_, _034288_, _034291_);
  and g_125065_(_011352_, _034215_, _034292_);
  or g_125066_(_011350_, _034216_, _034293_);
  and g_125067_(_034097_, _034216_, _034294_);
  or g_125068_(_034096_, _034215_, _034295_);
  and g_125069_(_034293_, _034295_, _034296_);
  or g_125070_(_034292_, _034294_, _034298_);
  and g_125071_(_011543_, _034298_, _034299_);
  or g_125072_(_011544_, _034296_, _034300_);
  and g_125073_(_034291_, _034300_, _034301_);
  or g_125074_(_034290_, _034299_, _034302_);
  and g_125075_(_011557_, _034288_, _034303_);
  or g_125076_(_011556_, _034289_, _034304_);
  and g_125077_(_011544_, _034296_, _034305_);
  or g_125078_(_011543_, _034298_, _034306_);
  and g_125079_(_034304_, _034306_, _034307_);
  or g_125080_(_034303_, _034305_, _034309_);
  and g_125081_(_034301_, _034307_, _034310_);
  or g_125082_(_034302_, _034309_, _034311_);
  and g_125083_(_011375_, _034215_, _034312_);
  or g_125084_(_011376_, _034216_, _034313_);
  and g_125085_(_034111_, _034216_, _034314_);
  or g_125086_(_034109_, _034215_, _034315_);
  and g_125087_(_034313_, _034315_, _034316_);
  or g_125088_(_034312_, _034314_, _034317_);
  and g_125089_(_011588_, _034317_, _034318_);
  or g_125090_(_011587_, _034316_, _034320_);
  and g_125091_(_011364_, _034215_, _034321_);
  or g_125092_(_011365_, _034216_, _034322_);
  and g_125093_(_034127_, _034216_, _034323_);
  or g_125094_(_034126_, _034215_, _034324_);
  and g_125095_(_034322_, _034324_, _034325_);
  or g_125096_(_034321_, _034323_, _034326_);
  and g_125097_(_011577_, _034326_, _034327_);
  or g_125098_(_011576_, _034325_, _034328_);
  and g_125099_(_034320_, _034328_, _034329_);
  or g_125100_(_034318_, _034327_, _034331_);
  and g_125101_(_011576_, _034325_, _034332_);
  or g_125102_(_011577_, _034326_, _034333_);
  and g_125103_(_011587_, _034316_, _034334_);
  or g_125104_(_011588_, _034317_, _034335_);
  and g_125105_(_011614_, _034255_, _034336_);
  or g_125106_(_011613_, _034256_, _034337_);
  and g_125107_(_034333_, _034335_, _034338_);
  or g_125108_(_034332_, _034334_, _034339_);
  and g_125109_(_034329_, _034338_, _034340_);
  or g_125110_(_034331_, _034339_, _034342_);
  and g_125111_(_034310_, _034340_, _034343_);
  or g_125112_(_034311_, _034342_, _034344_);
  and g_125113_(_034337_, _034343_, _034345_);
  or g_125114_(_034336_, _034344_, _034346_);
  and g_125115_(_034282_, _034345_, _034347_);
  or g_125116_(_034281_, _034346_, _034348_);
  and g_125117_(_034331_, _034335_, _034349_);
  or g_125118_(_034329_, _034334_, _034350_);
  and g_125119_(_034310_, _034349_, _034351_);
  or g_125120_(_034311_, _034350_, _034353_);
  and g_125121_(_034304_, _034305_, _034354_);
  or g_125122_(_034303_, _034306_, _034355_);
  and g_125123_(_034291_, _034355_, _034356_);
  or g_125124_(_034290_, _034354_, _034357_);
  and g_125125_(_034353_, _034356_, _034358_);
  or g_125126_(_034351_, _034357_, _034359_);
  and g_125127_(_034348_, _034358_, _034360_);
  or g_125128_(_034347_, _034359_, _034361_);
  and g_125129_(_011528_, _034237_, _034362_);
  or g_125130_(_011529_, _034238_, _034364_);
  and g_125131_(_034361_, _034364_, _034365_);
  or g_125132_(_034360_, _034362_, _034366_);
  and g_125133_(_034241_, _034364_, _034367_);
  and g_125134_(_034241_, _034366_, _034368_);
  or g_125135_(_034243_, _034365_, _034369_);
  and g_125136_(_034037_, _034215_, _034370_);
  or g_125137_(_034038_, _034216_, _034371_);
  and g_125138_(_034036_, _034216_, _034372_);
  or g_125139_(_034035_, _034215_, _034373_);
  and g_125140_(_034371_, _034373_, _034375_);
  or g_125141_(_034370_, _034372_, _034376_);
  or g_125142_(out[634], _011504_, _034377_);
  xor g_125143_(out[634], _011504_, _034378_);
  xor g_125144_(_055656_, _011504_, _034379_);
  and g_125145_(_034375_, _034378_, _034380_);
  or g_125146_(_034376_, _034379_, _034381_);
  and g_125147_(_034023_, _034026_, _034382_);
  or g_125148_(_034024_, _034027_, _034383_);
  xor g_125149_(out[635], _034377_, _034384_);
  xor g_125150_(_055535_, _034377_, _034386_);
  and g_125151_(_034382_, _034386_, _034387_);
  or g_125152_(_034383_, _034384_, _034388_);
  and g_125153_(_034381_, _034388_, _034389_);
  or g_125154_(_034380_, _034387_, _034390_);
  and g_125155_(_034383_, _034384_, _034391_);
  or g_125156_(_034382_, _034386_, _034392_);
  and g_125157_(_034376_, _034379_, _034393_);
  or g_125158_(_034375_, _034378_, _034394_);
  and g_125159_(_034392_, _034394_, _034395_);
  or g_125160_(_034391_, _034393_, _034397_);
  and g_125161_(_034389_, _034395_, _034398_);
  or g_125162_(_034390_, _034397_, _034399_);
  and g_125163_(_011506_, _034228_, _034400_);
  or g_125164_(_011507_, _034229_, _034401_);
  and g_125165_(_034398_, _034401_, _034402_);
  or g_125166_(_034399_, _034400_, _034403_);
  and g_125167_(_034369_, _034402_, _034404_);
  or g_125168_(_034368_, _034403_, _034405_);
  and g_125169_(_034390_, _034392_, _034406_);
  or g_125170_(_034389_, _034391_, _034408_);
  and g_125171_(_034405_, _034408_, _034409_);
  or g_125172_(_034404_, _034406_, _034410_);
  or g_125173_(out[624], _034223_, _034411_);
  and g_125174_(_034280_, _034401_, _034412_);
  and g_125175_(_034411_, _034412_, _034413_);
  and g_125176_(_034271_, _034367_, _034414_);
  and g_125177_(_034398_, _034414_, _034415_);
  and g_125178_(_034413_, _034415_, _034416_);
  not g_125179_(_034416_, _034417_);
  and g_125180_(_034345_, _034416_, _034419_);
  or g_125181_(_034346_, _034417_, _034420_);
  and g_125182_(_034410_, _034420_, _034421_);
  or g_125183_(_034409_, _034419_, _034422_);
  and g_125184_(_034223_, _034422_, _034423_);
  or g_125185_(_034222_, _034421_, _034424_);
  or g_125186_(out[624], _034422_, _034425_);
  not g_125187_(_034425_, _034426_);
  and g_125188_(_034424_, _034425_, _034427_);
  or g_125189_(_034423_, _034426_, _034428_);
  or g_125190_(_034379_, _034422_, _034430_);
  not g_125191_(_034430_, _034431_);
  and g_125192_(_034376_, _034422_, _034432_);
  not g_125193_(_034432_, _034433_);
  and g_125194_(_034430_, _034433_, _034434_);
  or g_125195_(_034431_, _034432_, _034435_);
  or g_125196_(out[650], _011798_, _034436_);
  xor g_125197_(out[650], _011798_, _034437_);
  xor g_125198_(_055788_, _011798_, _034438_);
  and g_125199_(_034434_, _034437_, _034439_);
  or g_125200_(_034435_, _034438_, _034441_);
  and g_125201_(_034382_, _034384_, _034442_);
  or g_125202_(_034383_, _034386_, _034443_);
  xor g_125203_(out[651], _034436_, _034444_);
  xor g_125204_(_055667_, _034436_, _034445_);
  and g_125205_(_034442_, _034445_, _034446_);
  or g_125206_(_034443_, _034444_, _034447_);
  and g_125207_(_034441_, _034447_, _034448_);
  or g_125208_(_034439_, _034446_, _034449_);
  or g_125209_(_011507_, _034422_, _034450_);
  not g_125210_(_034450_, _034452_);
  and g_125211_(_034229_, _034422_, _034453_);
  not g_125212_(_034453_, _034454_);
  and g_125213_(_034450_, _034454_, _034455_);
  or g_125214_(_034452_, _034453_, _034456_);
  and g_125215_(_011800_, _034456_, _034457_);
  or g_125216_(_011799_, _034455_, _034458_);
  and g_125217_(_034238_, _034422_, _034459_);
  not g_125218_(_034459_, _034460_);
  or g_125219_(_011529_, _034422_, _034461_);
  not g_125220_(_034461_, _034463_);
  and g_125221_(_034460_, _034461_, _034464_);
  or g_125222_(_034459_, _034463_, _034465_);
  and g_125223_(_011788_, _034465_, _034466_);
  or g_125224_(_011787_, _034464_, _034467_);
  and g_125225_(_034458_, _034467_, _034468_);
  or g_125226_(_034457_, _034466_, _034469_);
  or g_125227_(_011543_, _034422_, _034470_);
  or g_125228_(_034296_, _034421_, _034471_);
  and g_125229_(_034470_, _034471_, _034472_);
  and g_125230_(_011825_, _034472_, _034474_);
  and g_125231_(_034289_, _034422_, _034475_);
  or g_125232_(_034288_, _034421_, _034476_);
  and g_125233_(_011557_, _034421_, _034477_);
  or g_125234_(_011556_, _034422_, _034478_);
  and g_125235_(_034476_, _034478_, _034479_);
  or g_125236_(_034475_, _034477_, _034480_);
  and g_125237_(_011832_, _034480_, _034481_);
  or g_125238_(_034474_, _034481_, _034482_);
  or g_125239_(_011825_, _034472_, _034483_);
  not g_125240_(_034483_, _034485_);
  and g_125241_(_034317_, _034422_, _034486_);
  not g_125242_(_034486_, _034487_);
  or g_125243_(_011588_, _034422_, _034488_);
  not g_125244_(_034488_, _034489_);
  and g_125245_(_034487_, _034488_, _034490_);
  or g_125246_(_034486_, _034489_, _034491_);
  and g_125247_(_011856_, _034490_, _034492_);
  or g_125248_(_011858_, _034491_, _034493_);
  and g_125249_(_034483_, _034493_, _034494_);
  or g_125250_(_011577_, _034422_, _034496_);
  not g_125251_(_034496_, _034497_);
  and g_125252_(_034326_, _034422_, _034498_);
  not g_125253_(_034498_, _034499_);
  and g_125254_(_034496_, _034499_, _034500_);
  or g_125255_(_034497_, _034498_, _034501_);
  and g_125256_(_011848_, _034501_, _034502_);
  or g_125257_(_011847_, _034500_, _034503_);
  and g_125258_(_011858_, _034491_, _034504_);
  or g_125259_(_011856_, _034490_, _034505_);
  and g_125260_(_034503_, _034505_, _034507_);
  or g_125261_(_034502_, _034504_, _034508_);
  and g_125262_(_011847_, _034500_, _034509_);
  or g_125263_(_011848_, _034501_, _034510_);
  or g_125264_(_011613_, _034422_, _034511_);
  or g_125265_(_034255_, _034421_, _034512_);
  and g_125266_(_034511_, _034512_, _034513_);
  not g_125267_(_034513_, _034514_);
  and g_125268_(_011711_, _034514_, _034515_);
  or g_125269_(_011712_, _034513_, _034516_);
  or g_125270_(_055092_, _034422_, _034518_);
  not g_125271_(_034518_, _034519_);
  and g_125272_(_034249_, _034422_, _034520_);
  not g_125273_(_034520_, _034521_);
  and g_125274_(_034518_, _034521_, _034522_);
  or g_125275_(_034519_, _034520_, _034523_);
  and g_125276_(_055357_, _034522_, _034524_);
  or g_125277_(_055358_, _034523_, _034525_);
  and g_125278_(_011712_, _034513_, _034526_);
  or g_125279_(_011711_, _034514_, _034527_);
  and g_125280_(_034524_, _034527_, _034529_);
  or g_125281_(_034525_, _034526_, _034530_);
  and g_125282_(_034516_, _034530_, _034531_);
  or g_125283_(_034515_, _034529_, _034532_);
  and g_125284_(_055358_, _034523_, _034533_);
  or g_125285_(_034526_, _034533_, _034534_);
  or g_125286_(_034524_, _034534_, _034535_);
  or g_125287_(_055590_, _034422_, _034536_);
  or g_125288_(_034263_, _034421_, _034537_);
  and g_125289_(_034536_, _034537_, _034538_);
  and g_125290_(out[641], _034538_, _034540_);
  or g_125291_(_055733_, _034427_, _034541_);
  xor g_125292_(out[641], _034538_, _034542_);
  and g_125293_(_034541_, _034542_, _034543_);
  or g_125294_(_034540_, _034543_, _034544_);
  not g_125295_(_034544_, _034545_);
  or g_125296_(_034535_, _034545_, _034546_);
  xor g_125297_(_055357_, _034522_, _034547_);
  and g_125298_(_034516_, _034547_, _034548_);
  and g_125299_(_034527_, _034548_, _034549_);
  and g_125300_(_034541_, _034549_, _034551_);
  and g_125301_(_034542_, _034551_, _034552_);
  and g_125302_(_034544_, _034549_, _034553_);
  and g_125303_(_034531_, _034546_, _034554_);
  or g_125304_(_034532_, _034553_, _034555_);
  and g_125305_(_034510_, _034555_, _034556_);
  or g_125306_(_034508_, _034556_, _034557_);
  and g_125307_(_034494_, _034557_, _034558_);
  or g_125308_(_034482_, _034558_, _034559_);
  or g_125309_(_011832_, _034480_, _034560_);
  not g_125310_(_034560_, _034562_);
  and g_125311_(_011787_, _034464_, _034563_);
  or g_125312_(_011788_, _034465_, _034564_);
  and g_125313_(_034560_, _034564_, _034565_);
  and g_125314_(_034559_, _034565_, _034566_);
  or g_125315_(_034469_, _034566_, _034567_);
  and g_125316_(_034435_, _034438_, _034568_);
  or g_125317_(_034434_, _034437_, _034569_);
  and g_125318_(_011799_, _034455_, _034570_);
  or g_125319_(_011800_, _034456_, _034571_);
  and g_125320_(_034569_, _034571_, _034573_);
  and g_125321_(_034567_, _034573_, _034574_);
  and g_125322_(_034448_, _034569_, _034575_);
  or g_125323_(_034449_, _034568_, _034576_);
  or g_125324_(_034563_, _034570_, _034577_);
  or g_125325_(_034469_, _034577_, _034578_);
  or g_125326_(_034508_, _034509_, _034579_);
  or g_125327_(_034482_, _034485_, _034580_);
  or g_125328_(_034562_, _034580_, _034581_);
  or g_125329_(_034492_, _034581_, _034582_);
  or g_125330_(_034579_, _034582_, _034584_);
  or g_125331_(_034554_, _034584_, _034585_);
  and g_125332_(_034482_, _034560_, _034586_);
  not g_125333_(_034586_, _034587_);
  or g_125334_(_034507_, _034582_, _034588_);
  and g_125335_(_034587_, _034588_, _034589_);
  and g_125336_(_034585_, _034589_, _034590_);
  or g_125337_(_034578_, _034590_, _034591_);
  or g_125338_(_034468_, _034570_, _034592_);
  and g_125339_(_034591_, _034592_, _034593_);
  or g_125340_(_034576_, _034593_, _034595_);
  and g_125341_(_034448_, _034595_, _034596_);
  or g_125342_(_034449_, _034574_, _034597_);
  and g_125343_(_034443_, _034444_, _034598_);
  or g_125344_(_034442_, _034445_, _034599_);
  or g_125345_(out[640], _034428_, _034600_);
  and g_125346_(_034575_, _034600_, _034601_);
  and g_125347_(_034599_, _034601_, _034602_);
  and g_125348_(_034552_, _034602_, _034603_);
  not g_125349_(_034603_, _034604_);
  or g_125350_(_034578_, _034584_, _034606_);
  not g_125351_(_034606_, _034607_);
  and g_125352_(_034603_, _034607_, _034608_);
  or g_125353_(_034604_, _034606_, _034609_);
  and g_125354_(_034599_, _034609_, _034610_);
  or g_125355_(_034598_, _034608_, _034611_);
  and g_125356_(_034597_, _034610_, _034612_);
  or g_125357_(_034596_, _034611_, _034613_);
  and g_125358_(_034428_, _034613_, _034614_);
  not g_125359_(_034614_, _034615_);
  and g_125360_(_055733_, _034612_, _034617_);
  or g_125361_(out[640], _034613_, _034618_);
  and g_125362_(_034615_, _034618_, _034619_);
  or g_125363_(_034614_, _034617_, _034620_);
  and g_125364_(_034442_, _034444_, _034621_);
  or g_125365_(_034443_, _034445_, _034622_);
  or g_125366_(out[666], _011942_, _034623_);
  xor g_125367_(out[667], _034623_, _034624_);
  xor g_125368_(_055799_, _034623_, _034625_);
  and g_125369_(_034622_, _034624_, _034626_);
  or g_125370_(_034621_, _034625_, _034628_);
  and g_125371_(_034621_, _034625_, _034629_);
  or g_125372_(_034622_, _034624_, _034630_);
  and g_125373_(_034435_, _034613_, _034631_);
  or g_125374_(_034434_, _034612_, _034632_);
  and g_125375_(_034437_, _034612_, _034633_);
  or g_125376_(_034438_, _034613_, _034634_);
  and g_125377_(_034632_, _034634_, _034635_);
  or g_125378_(_034631_, _034633_, _034636_);
  xor g_125379_(out[666], _011942_, _034637_);
  xor g_125380_(_055920_, _011942_, _034639_);
  and g_125381_(_034635_, _034637_, _034640_);
  or g_125382_(_034636_, _034639_, _034641_);
  and g_125383_(_034630_, _034641_, _034642_);
  or g_125384_(_034629_, _034640_, _034643_);
  and g_125385_(_034628_, _034643_, _034644_);
  or g_125386_(_034626_, _034642_, _034645_);
  and g_125387_(_034636_, _034639_, _034646_);
  or g_125388_(_034635_, _034637_, _034647_);
  and g_125389_(_034628_, _034647_, _034648_);
  or g_125390_(_034626_, _034646_, _034650_);
  and g_125391_(_011799_, _034612_, _034651_);
  or g_125392_(_011800_, _034613_, _034652_);
  and g_125393_(_034456_, _034613_, _034653_);
  or g_125394_(_034455_, _034612_, _034654_);
  and g_125395_(_034652_, _034654_, _034655_);
  or g_125396_(_034651_, _034653_, _034656_);
  and g_125397_(_011943_, _034655_, _034657_);
  or g_125398_(_011944_, _034656_, _034658_);
  and g_125399_(_034465_, _034613_, _034659_);
  or g_125400_(_034464_, _034612_, _034661_);
  and g_125401_(_011787_, _034612_, _034662_);
  or g_125402_(_011788_, _034613_, _034663_);
  and g_125403_(_034661_, _034663_, _034664_);
  or g_125404_(_034659_, _034662_, _034665_);
  and g_125405_(_011933_, _034665_, _034666_);
  or g_125406_(_011932_, _034664_, _034667_);
  and g_125407_(_011944_, _034656_, _034668_);
  or g_125408_(_011943_, _034655_, _034669_);
  and g_125409_(_034667_, _034669_, _034670_);
  or g_125410_(_034666_, _034668_, _034672_);
  and g_125411_(_011932_, _034664_, _034673_);
  or g_125412_(_011933_, _034665_, _034674_);
  or g_125413_(_034472_, _034612_, _034675_);
  or g_125414_(_011823_, _034613_, _034676_);
  and g_125415_(_034675_, _034676_, _034677_);
  not g_125416_(_034677_, _034678_);
  or g_125417_(_011966_, _034678_, _034679_);
  or g_125418_(_011832_, _034613_, _034680_);
  or g_125419_(_034479_, _034612_, _034681_);
  and g_125420_(_034680_, _034681_, _034683_);
  and g_125421_(_011974_, _034683_, _034684_);
  or g_125422_(_011974_, _034683_, _034685_);
  not g_125423_(_034685_, _034686_);
  xor g_125424_(_011968_, _034677_, _034687_);
  xor g_125425_(_011966_, _034677_, _034688_);
  or g_125426_(_034684_, _034688_, _034689_);
  xor g_125427_(_011974_, _034683_, _034690_);
  and g_125428_(_034687_, _034690_, _034691_);
  or g_125429_(_034686_, _034689_, _034692_);
  and g_125430_(_034491_, _034613_, _034694_);
  or g_125431_(_034490_, _034612_, _034695_);
  and g_125432_(_011856_, _034612_, _034696_);
  or g_125433_(_011858_, _034613_, _034697_);
  and g_125434_(_034695_, _034697_, _034698_);
  or g_125435_(_034694_, _034696_, _034699_);
  and g_125436_(_012001_, _034698_, _034700_);
  or g_125437_(_012002_, _034699_, _034701_);
  and g_125438_(_012002_, _034699_, _034702_);
  or g_125439_(_012001_, _034698_, _034703_);
  and g_125440_(_011847_, _034612_, _034705_);
  or g_125441_(_011848_, _034613_, _034706_);
  and g_125442_(_034501_, _034613_, _034707_);
  or g_125443_(_034500_, _034612_, _034708_);
  and g_125444_(_034706_, _034708_, _034709_);
  or g_125445_(_034705_, _034707_, _034710_);
  and g_125446_(_011991_, _034710_, _034711_);
  or g_125447_(_011990_, _034709_, _034712_);
  and g_125448_(_034703_, _034712_, _034713_);
  or g_125449_(_034702_, _034711_, _034714_);
  and g_125450_(_034701_, _034714_, _034716_);
  or g_125451_(_034700_, _034713_, _034717_);
  or g_125452_(_011711_, _034613_, _034718_);
  or g_125453_(_034513_, _034612_, _034719_);
  and g_125454_(_034718_, _034719_, _034720_);
  or g_125455_(_012048_, _034720_, _034721_);
  and g_125456_(_012048_, _034720_, _034722_);
  xor g_125457_(_012048_, _034720_, _034723_);
  xor g_125458_(_012047_, _034720_, _034724_);
  and g_125459_(_034523_, _034613_, _034725_);
  and g_125460_(_055357_, _034612_, _034727_);
  or g_125461_(_034725_, _034727_, _034728_);
  or g_125462_(_055439_, _034728_, _034729_);
  xor g_125463_(_055439_, _034728_, _034730_);
  xor g_125464_(_055438_, _034728_, _034731_);
  and g_125465_(_034723_, _034730_, _034732_);
  or g_125466_(_034724_, _034731_, _034733_);
  or g_125467_(_055722_, _034613_, _034734_);
  or g_125468_(_034538_, _034612_, _034735_);
  and g_125469_(_034734_, _034735_, _034736_);
  and g_125470_(out[657], _034736_, _034738_);
  not g_125471_(_034738_, _034739_);
  and g_125472_(out[656], _034620_, _034740_);
  or g_125473_(_055865_, _034619_, _034741_);
  xor g_125474_(out[657], _034736_, _034742_);
  xor g_125475_(_055854_, _034736_, _034743_);
  and g_125476_(_034741_, _034742_, _034744_);
  or g_125477_(_034740_, _034743_, _034745_);
  and g_125478_(_034739_, _034745_, _034746_);
  or g_125479_(_034738_, _034744_, _034747_);
  and g_125480_(_034732_, _034747_, _034749_);
  or g_125481_(_034733_, _034746_, _034750_);
  or g_125482_(_034722_, _034729_, _034751_);
  and g_125483_(_034721_, _034751_, _034752_);
  not g_125484_(_034752_, _034753_);
  and g_125485_(_034750_, _034752_, _034754_);
  or g_125486_(_034749_, _034753_, _034755_);
  and g_125487_(_011990_, _034709_, _034756_);
  or g_125488_(_011991_, _034710_, _034757_);
  and g_125489_(_034701_, _034757_, _034758_);
  or g_125490_(_034700_, _034756_, _034760_);
  and g_125491_(_034713_, _034758_, _034761_);
  or g_125492_(_034714_, _034760_, _034762_);
  or g_125493_(_034679_, _034684_, _034763_);
  not g_125494_(_034763_, _034764_);
  and g_125495_(_034642_, _034648_, _034765_);
  or g_125496_(_034643_, _034650_, _034766_);
  and g_125497_(_034658_, _034674_, _034767_);
  or g_125498_(_034657_, _034673_, _034768_);
  and g_125499_(_034670_, _034767_, _034769_);
  or g_125500_(_034672_, _034768_, _034771_);
  and g_125501_(_034765_, _034769_, _034772_);
  or g_125502_(_034766_, _034771_, _034773_);
  and g_125503_(_034691_, _034716_, _034774_);
  or g_125504_(_034692_, _034717_, _034775_);
  and g_125505_(_034763_, _034775_, _034776_);
  or g_125506_(_034764_, _034774_, _034777_);
  and g_125507_(_034685_, _034776_, _034778_);
  or g_125508_(_034686_, _034777_, _034779_);
  and g_125509_(_034772_, _034779_, _034780_);
  or g_125510_(_034773_, _034778_, _034782_);
  and g_125511_(_034691_, _034761_, _034783_);
  or g_125512_(_034692_, _034762_, _034784_);
  and g_125513_(_034772_, _034783_, _034785_);
  or g_125514_(_034773_, _034784_, _034786_);
  and g_125515_(_034755_, _034785_, _034787_);
  or g_125516_(_034754_, _034786_, _034788_);
  and g_125517_(_034658_, _034672_, _034789_);
  or g_125518_(_034657_, _034670_, _034790_);
  and g_125519_(_034765_, _034789_, _034791_);
  or g_125520_(_034766_, _034790_, _034793_);
  and g_125521_(_034645_, _034788_, _034794_);
  or g_125522_(_034644_, _034787_, _034795_);
  and g_125523_(_034782_, _034793_, _034796_);
  or g_125524_(_034780_, _034791_, _034797_);
  and g_125525_(_034794_, _034796_, _034798_);
  or g_125526_(_034795_, _034797_, _034799_);
  and g_125527_(_034732_, _034744_, _034800_);
  or g_125528_(_034733_, _034745_, _034801_);
  and g_125529_(_055865_, _034619_, _034802_);
  or g_125530_(out[656], _034620_, _034804_);
  and g_125531_(_034785_, _034800_, _034805_);
  or g_125532_(_034786_, _034801_, _034806_);
  and g_125533_(_034804_, _034805_, _034807_);
  or g_125534_(_034802_, _034806_, _034808_);
  and g_125535_(_034799_, _034808_, _034809_);
  or g_125536_(_034798_, _034807_, _034810_);
  and g_125537_(_034620_, _034810_, _034811_);
  or g_125538_(_034619_, _034809_, _034812_);
  and g_125539_(_055865_, _034809_, _034813_);
  or g_125540_(out[656], _034810_, _034815_);
  and g_125541_(_034812_, _034815_, _034816_);
  or g_125542_(_034811_, _034813_, _034817_);
  and g_125543_(_034621_, _034624_, _034818_);
  or g_125544_(_034622_, _034625_, _034819_);
  or g_125545_(out[682], _012127_, _034820_);
  xor g_125546_(out[683], _034820_, _034821_);
  xor g_125547_(_055931_, _034820_, _034822_);
  and g_125548_(_034818_, _034822_, _034823_);
  or g_125549_(_034819_, _034821_, _034824_);
  and g_125550_(_034637_, _034809_, _034826_);
  or g_125551_(_034639_, _034810_, _034827_);
  and g_125552_(_034636_, _034810_, _034828_);
  or g_125553_(_034635_, _034809_, _034829_);
  and g_125554_(_034827_, _034829_, _034830_);
  or g_125555_(_034826_, _034828_, _034831_);
  xor g_125556_(out[682], _012127_, _034832_);
  xor g_125557_(_000087_, _012127_, _034833_);
  and g_125558_(_034830_, _034832_, _034834_);
  or g_125559_(_034831_, _034833_, _034835_);
  and g_125560_(_034824_, _034835_, _034837_);
  or g_125561_(_034823_, _034834_, _034838_);
  and g_125562_(_034831_, _034833_, _034839_);
  or g_125563_(_034830_, _034832_, _034840_);
  and g_125564_(_034819_, _034821_, _034841_);
  or g_125565_(_034818_, _034822_, _034842_);
  and g_125566_(_034840_, _034842_, _034843_);
  or g_125567_(_034839_, _034841_, _034844_);
  and g_125568_(_034837_, _034843_, _034845_);
  or g_125569_(_034838_, _034844_, _034846_);
  and g_125570_(_011932_, _034809_, _034848_);
  and g_125571_(_034665_, _034810_, _034849_);
  or g_125572_(_034848_, _034849_, _034850_);
  not g_125573_(_034850_, _034851_);
  and g_125574_(_012118_, _034850_, _034852_);
  or g_125575_(_012117_, _034851_, _034853_);
  and g_125576_(_011943_, _034809_, _034854_);
  and g_125577_(_034656_, _034810_, _034855_);
  or g_125578_(_034854_, _034855_, _034856_);
  not g_125579_(_034856_, _034857_);
  and g_125580_(_012129_, _034856_, _034859_);
  or g_125581_(_012128_, _034857_, _034860_);
  and g_125582_(_034853_, _034860_, _034861_);
  or g_125583_(_034852_, _034859_, _034862_);
  and g_125584_(_012128_, _034857_, _034863_);
  or g_125585_(_012129_, _034856_, _034864_);
  and g_125586_(_012117_, _034851_, _034865_);
  or g_125587_(_012118_, _034850_, _034866_);
  and g_125588_(_034864_, _034866_, _034867_);
  or g_125589_(_034863_, _034865_, _034868_);
  and g_125590_(_034861_, _034867_, _034870_);
  or g_125591_(_034862_, _034868_, _034871_);
  and g_125592_(_034845_, _034870_, _034872_);
  or g_125593_(_034846_, _034871_, _034873_);
  or g_125594_(_011966_, _034810_, _034874_);
  or g_125595_(_034677_, _034809_, _034875_);
  and g_125596_(_034874_, _034875_, _034876_);
  not g_125597_(_034876_, _034877_);
  and g_125598_(_012152_, _034876_, _034878_);
  or g_125599_(_012151_, _034877_, _034879_);
  or g_125600_(_011973_, _034810_, _034881_);
  or g_125601_(_034683_, _034809_, _034882_);
  and g_125602_(_034881_, _034882_, _034883_);
  not g_125603_(_034883_, _034884_);
  and g_125604_(_012159_, _034884_, _034885_);
  not g_125605_(_034885_, _034886_);
  and g_125606_(_012160_, _034883_, _034887_);
  not g_125607_(_034887_, _034888_);
  xor g_125608_(_012152_, _034876_, _034889_);
  xor g_125609_(_012151_, _034876_, _034890_);
  and g_125610_(_034888_, _034889_, _034892_);
  or g_125611_(_034887_, _034890_, _034893_);
  and g_125612_(_034886_, _034892_, _034894_);
  or g_125613_(_034885_, _034893_, _034895_);
  and g_125614_(_012001_, _034809_, _034896_);
  or g_125615_(_012002_, _034810_, _034897_);
  and g_125616_(_034699_, _034810_, _034898_);
  or g_125617_(_034698_, _034809_, _034899_);
  and g_125618_(_034897_, _034899_, _034900_);
  or g_125619_(_034896_, _034898_, _034901_);
  and g_125620_(_012192_, _034901_, _034903_);
  or g_125621_(_012191_, _034900_, _034904_);
  and g_125622_(_011990_, _034809_, _034905_);
  or g_125623_(_011991_, _034810_, _034906_);
  and g_125624_(_034710_, _034810_, _034907_);
  or g_125625_(_034709_, _034809_, _034908_);
  and g_125626_(_034906_, _034908_, _034909_);
  or g_125627_(_034905_, _034907_, _034910_);
  and g_125628_(_012181_, _034910_, _034911_);
  or g_125629_(_012180_, _034909_, _034912_);
  and g_125630_(_034904_, _034912_, _034914_);
  or g_125631_(_034903_, _034911_, _034915_);
  or g_125632_(_012192_, _034901_, _034916_);
  not g_125633_(_034916_, _034917_);
  or g_125634_(_012181_, _034910_, _034918_);
  and g_125635_(_034916_, _034918_, _034919_);
  not g_125636_(_034919_, _034920_);
  and g_125637_(_034914_, _034919_, _034921_);
  or g_125638_(_034915_, _034920_, _034922_);
  and g_125639_(_034894_, _034921_, _034923_);
  or g_125640_(_034895_, _034922_, _034925_);
  and g_125641_(_034872_, _034923_, _034926_);
  or g_125642_(_034873_, _034925_, _034927_);
  or g_125643_(_012047_, _034810_, _034928_);
  or g_125644_(_034720_, _034809_, _034929_);
  and g_125645_(_034928_, _034929_, _034930_);
  not g_125646_(_034930_, _034931_);
  or g_125647_(_012216_, _034930_, _034932_);
  and g_125648_(_034728_, _034810_, _034933_);
  and g_125649_(_055438_, _034809_, _034934_);
  or g_125650_(_034933_, _034934_, _034936_);
  and g_125651_(_012216_, _034930_, _034937_);
  or g_125652_(_055742_, _034936_, _034938_);
  xor g_125653_(_012216_, _034930_, _034939_);
  xor g_125654_(_012215_, _034930_, _034940_);
  xor g_125655_(_055742_, _034936_, _034941_);
  xor g_125656_(_055743_, _034936_, _034942_);
  and g_125657_(_034939_, _034941_, _034943_);
  or g_125658_(_034940_, _034942_, _034944_);
  or g_125659_(_055854_, _034810_, _034945_);
  or g_125660_(_034736_, _034809_, _034947_);
  and g_125661_(_034945_, _034947_, _034948_);
  and g_125662_(out[673], _034948_, _034949_);
  not g_125663_(_034949_, _034950_);
  and g_125664_(out[672], _034817_, _034951_);
  or g_125665_(_000032_, _034816_, _034952_);
  xor g_125666_(out[673], _034948_, _034953_);
  xor g_125667_(_000021_, _034948_, _034954_);
  and g_125668_(_034952_, _034953_, _034955_);
  or g_125669_(_034951_, _034954_, _034956_);
  and g_125670_(_034950_, _034956_, _034958_);
  or g_125671_(_034949_, _034955_, _034959_);
  and g_125672_(_034943_, _034959_, _034960_);
  or g_125673_(_034944_, _034958_, _034961_);
  or g_125674_(_034937_, _034938_, _034962_);
  and g_125675_(_034932_, _034962_, _034963_);
  not g_125676_(_034963_, _034964_);
  and g_125677_(_034961_, _034963_, _034965_);
  or g_125678_(_034960_, _034964_, _034966_);
  and g_125679_(_034926_, _034966_, _034967_);
  or g_125680_(_034927_, _034965_, _034969_);
  and g_125681_(_034915_, _034916_, _034970_);
  or g_125682_(_034914_, _034917_, _034971_);
  and g_125683_(_034894_, _034970_, _034972_);
  or g_125684_(_034895_, _034971_, _034973_);
  and g_125685_(_034878_, _034888_, _034974_);
  or g_125686_(_034879_, _034887_, _034975_);
  and g_125687_(_034886_, _034975_, _034976_);
  or g_125688_(_034885_, _034974_, _034977_);
  and g_125689_(_034973_, _034976_, _034978_);
  or g_125690_(_034972_, _034977_, _034980_);
  and g_125691_(_034872_, _034980_, _034981_);
  or g_125692_(_034873_, _034978_, _034982_);
  or g_125693_(_034837_, _034841_, _034983_);
  not g_125694_(_034983_, _034984_);
  and g_125695_(_034862_, _034864_, _034985_);
  or g_125696_(_034846_, _034861_, _034986_);
  and g_125697_(_034845_, _034985_, _034987_);
  or g_125698_(_034863_, _034986_, _034988_);
  and g_125699_(_034983_, _034988_, _034989_);
  or g_125700_(_034984_, _034987_, _034991_);
  and g_125701_(_034982_, _034989_, _034992_);
  or g_125702_(_034981_, _034991_, _034993_);
  and g_125703_(_034969_, _034992_, _034994_);
  or g_125704_(_034967_, _034993_, _034995_);
  and g_125705_(_000032_, _034816_, _034996_);
  or g_125706_(_034956_, _034996_, _034997_);
  or g_125707_(_034944_, _034997_, _034998_);
  or g_125708_(_034927_, _034998_, _034999_);
  not g_125709_(_034999_, _035000_);
  and g_125710_(_034995_, _034999_, _035002_);
  or g_125711_(_034994_, _035000_, _035003_);
  and g_125712_(_034817_, _035003_, _035004_);
  not g_125713_(_035004_, _035005_);
  or g_125714_(out[672], _035003_, _035006_);
  not g_125715_(_035006_, _035007_);
  and g_125716_(_035005_, _035006_, _035008_);
  or g_125717_(_035004_, _035007_, _035009_);
  or g_125718_(_034833_, _035003_, _035010_);
  not g_125719_(_035010_, _035011_);
  and g_125720_(_034831_, _035003_, _035013_);
  not g_125721_(_035013_, _035014_);
  and g_125722_(_035010_, _035014_, _035015_);
  or g_125723_(_035011_, _035013_, _035016_);
  or g_125724_(out[698], _012333_, _035017_);
  xor g_125725_(out[698], _012333_, _035018_);
  xor g_125726_(_000219_, _012333_, _035019_);
  and g_125727_(_035015_, _035018_, _035020_);
  or g_125728_(_035016_, _035019_, _035021_);
  and g_125729_(_034818_, _034821_, _035022_);
  or g_125730_(_034819_, _034822_, _035024_);
  xor g_125731_(out[699], _035017_, _035025_);
  xor g_125732_(_000098_, _035017_, _035026_);
  and g_125733_(_035022_, _035026_, _035027_);
  or g_125734_(_035024_, _035025_, _035028_);
  and g_125735_(_035021_, _035028_, _035029_);
  or g_125736_(_035020_, _035027_, _035030_);
  and g_125737_(_035016_, _035019_, _035031_);
  or g_125738_(_035015_, _035018_, _035032_);
  or g_125739_(_012129_, _035003_, _035033_);
  not g_125740_(_035033_, _035035_);
  and g_125741_(_034856_, _035003_, _035036_);
  not g_125742_(_035036_, _035037_);
  and g_125743_(_035033_, _035037_, _035038_);
  or g_125744_(_035035_, _035036_, _035039_);
  and g_125745_(_012335_, _035039_, _035040_);
  or g_125746_(_012334_, _035038_, _035041_);
  or g_125747_(_012118_, _035003_, _035042_);
  not g_125748_(_035042_, _035043_);
  and g_125749_(_034850_, _035003_, _035044_);
  not g_125750_(_035044_, _035046_);
  and g_125751_(_035042_, _035046_, _035047_);
  or g_125752_(_035043_, _035044_, _035048_);
  and g_125753_(_012343_, _035048_, _035049_);
  or g_125754_(_012342_, _035047_, _035050_);
  and g_125755_(_035041_, _035050_, _035051_);
  or g_125756_(_035040_, _035049_, _035052_);
  and g_125757_(_012334_, _035038_, _035053_);
  or g_125758_(_012335_, _035039_, _035054_);
  and g_125759_(_035052_, _035054_, _035055_);
  or g_125760_(_035051_, _035053_, _035057_);
  and g_125761_(_012342_, _035047_, _035058_);
  or g_125762_(_035053_, _035058_, _035059_);
  not g_125763_(_035059_, _035060_);
  and g_125764_(_035051_, _035060_, _035061_);
  or g_125765_(_035052_, _035059_, _035062_);
  and g_125766_(_012160_, _035002_, _035063_);
  or g_125767_(_012159_, _035003_, _035064_);
  and g_125768_(_034884_, _035003_, _035065_);
  or g_125769_(_034883_, _035002_, _035066_);
  and g_125770_(_035064_, _035066_, _035068_);
  or g_125771_(_035063_, _035065_, _035069_);
  or g_125772_(_012364_, _035068_, _035070_);
  or g_125773_(_012151_, _035003_, _035071_);
  or g_125774_(_034876_, _035002_, _035072_);
  and g_125775_(_035071_, _035072_, _035073_);
  not g_125776_(_035073_, _035074_);
  or g_125777_(_012373_, _035074_, _035075_);
  and g_125778_(_012364_, _035068_, _035076_);
  or g_125779_(_035075_, _035076_, _035077_);
  and g_125780_(_035070_, _035077_, _035079_);
  or g_125781_(_012192_, _035003_, _035080_);
  not g_125782_(_035080_, _035081_);
  and g_125783_(_034901_, _035003_, _035082_);
  not g_125784_(_035082_, _035083_);
  and g_125785_(_035080_, _035083_, _035084_);
  or g_125786_(_035081_, _035082_, _035085_);
  and g_125787_(_012403_, _035084_, _035086_);
  or g_125788_(_012404_, _035085_, _035087_);
  xor g_125789_(_012375_, _035073_, _035088_);
  xor g_125790_(_012373_, _035073_, _035090_);
  xor g_125791_(_012364_, _035068_, _035091_);
  xor g_125792_(_012362_, _035068_, _035092_);
  and g_125793_(_035088_, _035091_, _035093_);
  or g_125794_(_035090_, _035092_, _035094_);
  and g_125795_(_035087_, _035093_, _035095_);
  or g_125796_(_035086_, _035094_, _035096_);
  or g_125797_(_012181_, _035003_, _035097_);
  not g_125798_(_035097_, _035098_);
  and g_125799_(_034910_, _035003_, _035099_);
  not g_125800_(_035099_, _035101_);
  and g_125801_(_035097_, _035101_, _035102_);
  or g_125802_(_035098_, _035099_, _035103_);
  and g_125803_(_012393_, _035103_, _035104_);
  or g_125804_(_012392_, _035102_, _035105_);
  and g_125805_(_012404_, _035085_, _035106_);
  or g_125806_(_012403_, _035084_, _035107_);
  and g_125807_(_035105_, _035107_, _035108_);
  or g_125808_(_035104_, _035106_, _035109_);
  and g_125809_(_012392_, _035102_, _035110_);
  or g_125810_(_012393_, _035103_, _035112_);
  or g_125811_(_012215_, _035003_, _035113_);
  not g_125812_(_035113_, _035114_);
  and g_125813_(_034931_, _035003_, _035115_);
  not g_125814_(_035115_, _035116_);
  and g_125815_(_035113_, _035116_, _035117_);
  or g_125816_(_035114_, _035115_, _035118_);
  and g_125817_(_012424_, _035118_, _035119_);
  or g_125818_(_012425_, _035117_, _035120_);
  and g_125819_(_012425_, _035117_, _035121_);
  or g_125820_(_012424_, _035118_, _035123_);
  and g_125821_(_034936_, _035003_, _035124_);
  not g_125822_(_035124_, _035125_);
  or g_125823_(_055742_, _035003_, _035126_);
  not g_125824_(_035126_, _035127_);
  and g_125825_(_035125_, _035126_, _035128_);
  or g_125826_(_035124_, _035127_, _035129_);
  and g_125827_(_055930_, _035128_, _035130_);
  or g_125828_(_055932_, _035129_, _035131_);
  and g_125829_(_035123_, _035130_, _035132_);
  or g_125830_(_035121_, _035131_, _035134_);
  and g_125831_(_035120_, _035134_, _035135_);
  or g_125832_(_035119_, _035132_, _035136_);
  and g_125833_(_055932_, _035129_, _035137_);
  or g_125834_(_035121_, _035130_, _035138_);
  or g_125835_(_035137_, _035138_, _035139_);
  and g_125836_(_034948_, _035003_, _035140_);
  not g_125837_(_035140_, _035141_);
  and g_125838_(_000021_, _035002_, _035142_);
  or g_125839_(out[673], _035003_, _035143_);
  or g_125840_(_035140_, _035142_, _035145_);
  and g_125841_(_035141_, _035143_, _035146_);
  and g_125842_(out[689], _035145_, _035147_);
  or g_125843_(_000153_, _035146_, _035148_);
  and g_125844_(out[688], _035009_, _035149_);
  and g_125845_(_000153_, _035146_, _035150_);
  or g_125846_(_035149_, _035150_, _035151_);
  or g_125847_(_035147_, _035150_, _035152_);
  or g_125848_(_035149_, _035152_, _035153_);
  not g_125849_(_035153_, _035154_);
  and g_125850_(_035148_, _035151_, _035156_);
  or g_125851_(_035147_, _035154_, _035157_);
  or g_125852_(_035139_, _035156_, _035158_);
  and g_125853_(_035135_, _035158_, _035159_);
  or g_125854_(_035110_, _035159_, _035160_);
  and g_125855_(_035108_, _035160_, _035161_);
  or g_125856_(_035096_, _035161_, _035162_);
  and g_125857_(_035108_, _035112_, _035163_);
  and g_125858_(_035095_, _035163_, _035164_);
  and g_125859_(_035136_, _035164_, _035165_);
  and g_125860_(_035120_, _035123_, _035167_);
  xor g_125861_(_055930_, _035128_, _035168_);
  and g_125862_(_035164_, _035168_, _035169_);
  and g_125863_(_035167_, _035169_, _035170_);
  and g_125864_(_035157_, _035170_, _035171_);
  or g_125865_(_035096_, _035108_, _035172_);
  and g_125866_(_035079_, _035172_, _035173_);
  not g_125867_(_035173_, _035174_);
  or g_125868_(_035171_, _035174_, _035175_);
  and g_125869_(_035079_, _035162_, _035176_);
  or g_125870_(_035165_, _035175_, _035178_);
  and g_125871_(_035061_, _035178_, _035179_);
  or g_125872_(_035062_, _035176_, _035180_);
  and g_125873_(_035057_, _035180_, _035181_);
  or g_125874_(_035055_, _035179_, _035182_);
  and g_125875_(_035032_, _035182_, _035183_);
  or g_125876_(_035031_, _035181_, _035184_);
  and g_125877_(_035029_, _035184_, _035185_);
  or g_125878_(_035030_, _035183_, _035186_);
  and g_125879_(_035024_, _035025_, _035187_);
  or g_125880_(_035022_, _035026_, _035189_);
  or g_125881_(_035110_, _035147_, _035190_);
  and g_125882_(_000164_, _035008_, _035191_);
  or g_125883_(out[688], _035009_, _035192_);
  or g_125884_(_035119_, _035191_, _035193_);
  or g_125885_(_035190_, _035193_, _035194_);
  or g_125886_(_035062_, _035194_, _035195_);
  or g_125887_(_035139_, _035195_, _035196_);
  and g_125888_(_035032_, _035189_, _035197_);
  or g_125889_(_035031_, _035187_, _035198_);
  and g_125890_(_035029_, _035197_, _035200_);
  or g_125891_(_035030_, _035198_, _035201_);
  or g_125892_(_035109_, _035151_, _035202_);
  or g_125893_(_035201_, _035202_, _035203_);
  or g_125894_(_035096_, _035203_, _035204_);
  and g_125895_(_035154_, _035192_, _035205_);
  and g_125896_(_035061_, _035205_, _035206_);
  and g_125897_(_035200_, _035206_, _035207_);
  and g_125898_(_035170_, _035207_, _035208_);
  or g_125899_(_035196_, _035204_, _035209_);
  and g_125900_(_035189_, _035209_, _035211_);
  or g_125901_(_035187_, _035208_, _035212_);
  and g_125902_(_035186_, _035211_, _035213_);
  or g_125903_(_035185_, _035212_, _035214_);
  and g_125904_(_035009_, _035214_, _035215_);
  not g_125905_(_035215_, _035216_);
  or g_125906_(out[688], _035214_, _035217_);
  not g_125907_(_035217_, _035218_);
  and g_125908_(_035216_, _035217_, _035219_);
  or g_125909_(_035215_, _035218_, _035220_);
  and g_125910_(_035022_, _035025_, _035222_);
  or g_125911_(_035024_, _035026_, _035223_);
  or g_125912_(out[714], _012532_, _035224_);
  xor g_125913_(out[715], _035224_, _035225_);
  not g_125914_(_035225_, _035226_);
  or g_125915_(_035223_, _035225_, _035227_);
  xor g_125916_(out[714], _012532_, _035228_);
  not g_125917_(_035228_, _035229_);
  and g_125918_(_035016_, _035214_, _035230_);
  not g_125919_(_035230_, _035231_);
  or g_125920_(_035019_, _035214_, _035233_);
  not g_125921_(_035233_, _035234_);
  and g_125922_(_035231_, _035233_, _035235_);
  or g_125923_(_035230_, _035234_, _035236_);
  or g_125924_(_035229_, _035236_, _035237_);
  and g_125925_(_035227_, _035237_, _035238_);
  and g_125926_(_035223_, _035225_, _035239_);
  or g_125927_(_035222_, _035226_, _035240_);
  or g_125928_(_035228_, _035235_, _035241_);
  and g_125929_(_035240_, _035241_, _035242_);
  xor g_125930_(_035222_, _035225_, _035244_);
  xor g_125931_(_035229_, _035235_, _035245_);
  and g_125932_(_035238_, _035242_, _035246_);
  or g_125933_(_035244_, _035245_, _035247_);
  or g_125934_(_012335_, _035214_, _035248_);
  not g_125935_(_035248_, _035249_);
  and g_125936_(_035039_, _035214_, _035250_);
  not g_125937_(_035250_, _035251_);
  and g_125938_(_035248_, _035251_, _035252_);
  or g_125939_(_035249_, _035250_, _035253_);
  and g_125940_(_012534_, _035253_, _035255_);
  or g_125941_(_012533_, _035252_, _035256_);
  and g_125942_(_035048_, _035214_, _035257_);
  not g_125943_(_035257_, _035258_);
  or g_125944_(_012343_, _035214_, _035259_);
  not g_125945_(_035259_, _035260_);
  and g_125946_(_035258_, _035259_, _035261_);
  or g_125947_(_035257_, _035260_, _035262_);
  and g_125948_(_012522_, _035262_, _035263_);
  or g_125949_(_012521_, _035261_, _035264_);
  and g_125950_(_035256_, _035264_, _035266_);
  or g_125951_(_035255_, _035263_, _035267_);
  and g_125952_(_012533_, _035252_, _035268_);
  or g_125953_(_012534_, _035253_, _035269_);
  and g_125954_(_012521_, _035261_, _035270_);
  or g_125955_(_012522_, _035262_, _035271_);
  and g_125956_(_035269_, _035271_, _035272_);
  or g_125957_(_035268_, _035270_, _035273_);
  and g_125958_(_035266_, _035272_, _035274_);
  or g_125959_(_035267_, _035273_, _035275_);
  and g_125960_(_035246_, _035274_, _035277_);
  or g_125961_(_035247_, _035275_, _035278_);
  and g_125962_(_035069_, _035214_, _035279_);
  or g_125963_(_035068_, _035213_, _035280_);
  and g_125964_(_012364_, _035213_, _035281_);
  or g_125965_(_012362_, _035214_, _035282_);
  and g_125966_(_035280_, _035282_, _035283_);
  or g_125967_(_035279_, _035281_, _035284_);
  and g_125968_(_012557_, _035284_, _035285_);
  or g_125969_(_012558_, _035283_, _035286_);
  or g_125970_(_035073_, _035213_, _035288_);
  or g_125971_(_012373_, _035214_, _035289_);
  and g_125972_(_035288_, _035289_, _035290_);
  not g_125973_(_035290_, _035291_);
  and g_125974_(_012574_, _035290_, _035292_);
  or g_125975_(_012573_, _035291_, _035293_);
  and g_125976_(_012558_, _035283_, _035294_);
  or g_125977_(_012557_, _035284_, _035295_);
  and g_125978_(_035085_, _035214_, _035296_);
  not g_125979_(_035296_, _035297_);
  or g_125980_(_012404_, _035214_, _035299_);
  not g_125981_(_035299_, _035300_);
  and g_125982_(_035297_, _035299_, _035301_);
  or g_125983_(_035296_, _035300_, _035302_);
  and g_125984_(_012598_, _035301_, _035303_);
  or g_125985_(_012599_, _035302_, _035304_);
  and g_125986_(_035286_, _035295_, _035305_);
  or g_125987_(_035285_, _035294_, _035306_);
  xor g_125988_(_012574_, _035290_, _035307_);
  xor g_125989_(_012573_, _035290_, _035308_);
  and g_125990_(_035305_, _035307_, _035310_);
  or g_125991_(_035306_, _035308_, _035311_);
  and g_125992_(_035304_, _035310_, _035312_);
  or g_125993_(_035303_, _035311_, _035313_);
  or g_125994_(_012393_, _035214_, _035314_);
  not g_125995_(_035314_, _035315_);
  and g_125996_(_035103_, _035214_, _035316_);
  not g_125997_(_035316_, _035317_);
  and g_125998_(_035314_, _035317_, _035318_);
  or g_125999_(_035315_, _035316_, _035319_);
  and g_126000_(_012588_, _035319_, _035321_);
  or g_126001_(_012587_, _035318_, _035322_);
  and g_126002_(_012599_, _035302_, _035323_);
  or g_126003_(_012598_, _035301_, _035324_);
  and g_126004_(_035322_, _035324_, _035325_);
  or g_126005_(_035321_, _035323_, _035326_);
  and g_126006_(_012587_, _035318_, _035327_);
  or g_126007_(_012588_, _035319_, _035328_);
  and g_126008_(_035325_, _035328_, _035329_);
  or g_126009_(_035326_, _035327_, _035330_);
  and g_126010_(_035312_, _035329_, _035332_);
  or g_126011_(_035313_, _035330_, _035333_);
  and g_126012_(_035118_, _035214_, _035334_);
  not g_126013_(_035334_, _035335_);
  or g_126014_(_012424_, _035214_, _035336_);
  not g_126015_(_035336_, _035337_);
  and g_126016_(_035335_, _035336_, _035338_);
  or g_126017_(_035334_, _035337_, _035339_);
  and g_126018_(_012622_, _035338_, _035340_);
  or g_126019_(_012621_, _035339_, _035341_);
  and g_126020_(_012621_, _035339_, _035343_);
  or g_126021_(_012622_, _035338_, _035344_);
  and g_126022_(_035341_, _035344_, _035345_);
  or g_126023_(_035340_, _035343_, _035346_);
  and g_126024_(_035129_, _035214_, _035347_);
  not g_126025_(_035347_, _035348_);
  or g_126026_(_055932_, _035214_, _035349_);
  not g_126027_(_035349_, _035350_);
  and g_126028_(_035348_, _035349_, _035351_);
  or g_126029_(_035347_, _035350_, _035352_);
  and g_126030_(_000141_, _035351_, _035354_);
  or g_126031_(_000143_, _035352_, _035355_);
  xor g_126032_(_000141_, _035351_, _035356_);
  xor g_126033_(_000143_, _035351_, _035357_);
  and g_126034_(_035345_, _035356_, _035358_);
  or g_126035_(_035346_, _035357_, _035359_);
  and g_126036_(_035146_, _035214_, _035360_);
  not g_126037_(_035360_, _035361_);
  or g_126038_(_000153_, _035214_, _035362_);
  not g_126039_(_035362_, _035363_);
  and g_126040_(_035361_, _035362_, _035365_);
  or g_126041_(_035360_, _035363_, _035366_);
  and g_126042_(out[705], _035365_, _035367_);
  or g_126043_(_000285_, _035366_, _035368_);
  and g_126044_(out[704], _035220_, _035369_);
  or g_126045_(_000296_, _035219_, _035370_);
  xor g_126046_(out[705], _035365_, _035371_);
  xor g_126047_(_000285_, _035365_, _035372_);
  and g_126048_(_035370_, _035371_, _035373_);
  or g_126049_(_035369_, _035372_, _035374_);
  and g_126050_(_035368_, _035374_, _035376_);
  or g_126051_(_035367_, _035373_, _035377_);
  and g_126052_(_035358_, _035377_, _035378_);
  or g_126053_(_035359_, _035376_, _035379_);
  and g_126054_(_035344_, _035355_, _035380_);
  or g_126055_(_035343_, _035354_, _035381_);
  and g_126056_(_035341_, _035381_, _035382_);
  or g_126057_(_035340_, _035380_, _035383_);
  and g_126058_(_035379_, _035383_, _035384_);
  or g_126059_(_035378_, _035382_, _035385_);
  and g_126060_(_035332_, _035385_, _035387_);
  or g_126061_(_035333_, _035384_, _035388_);
  and g_126062_(_035312_, _035326_, _035389_);
  or g_126063_(_035313_, _035325_, _035390_);
  and g_126064_(_035292_, _035295_, _035391_);
  or g_126065_(_035293_, _035294_, _035392_);
  and g_126066_(_035286_, _035392_, _035393_);
  or g_126067_(_035285_, _035391_, _035394_);
  and g_126068_(_035390_, _035393_, _035395_);
  or g_126069_(_035389_, _035394_, _035396_);
  and g_126070_(_035388_, _035395_, _035398_);
  or g_126071_(_035387_, _035396_, _035399_);
  and g_126072_(_035277_, _035399_, _035400_);
  or g_126073_(_035278_, _035398_, _035401_);
  or g_126074_(_035238_, _035239_, _035402_);
  or g_126075_(_035247_, _035268_, _035403_);
  or g_126076_(_035266_, _035403_, _035404_);
  and g_126077_(_035402_, _035404_, _035405_);
  not g_126078_(_035405_, _035406_);
  and g_126079_(_035401_, _035405_, _035407_);
  or g_126080_(_035400_, _035406_, _035409_);
  and g_126081_(_000296_, _035219_, _035410_);
  or g_126082_(out[704], _035220_, _035411_);
  and g_126083_(_035373_, _035411_, _035412_);
  or g_126084_(_035374_, _035410_, _035413_);
  and g_126085_(_035358_, _035412_, _035414_);
  or g_126086_(_035359_, _035413_, _035415_);
  and g_126087_(_035277_, _035414_, _035416_);
  or g_126088_(_035278_, _035415_, _035417_);
  and g_126089_(_035332_, _035416_, _035418_);
  or g_126090_(_035333_, _035417_, _035420_);
  and g_126091_(_035409_, _035420_, _035421_);
  or g_126092_(_035407_, _035418_, _035422_);
  and g_126093_(_035220_, _035422_, _035423_);
  or g_126094_(_035219_, _035421_, _035424_);
  or g_126095_(out[704], _035422_, _035425_);
  not g_126096_(_035425_, _035426_);
  and g_126097_(_035424_, _035425_, _035427_);
  or g_126098_(_035423_, _035426_, _035428_);
  and g_126099_(_035222_, _035225_, _035429_);
  or g_126100_(_035223_, _035226_, _035431_);
  or g_126101_(out[730], _012732_, _035432_);
  xor g_126102_(out[731], _035432_, _035433_);
  xor g_126103_(_000362_, _035432_, _035434_);
  and g_126104_(_035429_, _035434_, _035435_);
  or g_126105_(_035431_, _035433_, _035436_);
  and g_126106_(_035236_, _035422_, _035437_);
  not g_126107_(_035437_, _035438_);
  or g_126108_(_035229_, _035422_, _035439_);
  not g_126109_(_035439_, _035440_);
  and g_126110_(_035438_, _035439_, _035442_);
  or g_126111_(_035437_, _035440_, _035443_);
  xor g_126112_(out[730], _012732_, _035444_);
  xor g_126113_(_000483_, _012732_, _035445_);
  and g_126114_(_035442_, _035444_, _035446_);
  or g_126115_(_035443_, _035445_, _035447_);
  and g_126116_(_035436_, _035447_, _035448_);
  or g_126117_(_035435_, _035446_, _035449_);
  and g_126118_(_035443_, _035445_, _035450_);
  or g_126119_(_035442_, _035444_, _035451_);
  and g_126120_(_035431_, _035433_, _035453_);
  or g_126121_(_035429_, _035434_, _035454_);
  and g_126122_(_035451_, _035454_, _035455_);
  or g_126123_(_035450_, _035453_, _035456_);
  and g_126124_(_035448_, _035455_, _035457_);
  or g_126125_(_035449_, _035456_, _035458_);
  or g_126126_(_012522_, _035422_, _035459_);
  not g_126127_(_035459_, _035460_);
  and g_126128_(_035262_, _035422_, _035461_);
  not g_126129_(_035461_, _035462_);
  and g_126130_(_035459_, _035462_, _035464_);
  or g_126131_(_035460_, _035461_, _035465_);
  and g_126132_(_012718_, _035465_, _035466_);
  or g_126133_(_012717_, _035464_, _035467_);
  or g_126134_(_012534_, _035422_, _035468_);
  not g_126135_(_035468_, _035469_);
  and g_126136_(_035253_, _035422_, _035470_);
  not g_126137_(_035470_, _035471_);
  and g_126138_(_035468_, _035471_, _035472_);
  or g_126139_(_035469_, _035470_, _035473_);
  and g_126140_(_012734_, _035473_, _035475_);
  or g_126141_(_012733_, _035472_, _035476_);
  and g_126142_(_035467_, _035476_, _035477_);
  or g_126143_(_035466_, _035475_, _035478_);
  and g_126144_(_012733_, _035472_, _035479_);
  or g_126145_(_012734_, _035473_, _035480_);
  and g_126146_(_012717_, _035464_, _035481_);
  or g_126147_(_012718_, _035465_, _035482_);
  and g_126148_(_035480_, _035482_, _035483_);
  or g_126149_(_035479_, _035481_, _035484_);
  and g_126150_(_035477_, _035483_, _035486_);
  or g_126151_(_035478_, _035484_, _035487_);
  and g_126152_(_035457_, _035486_, _035488_);
  or g_126153_(_035458_, _035487_, _035489_);
  or g_126154_(_012557_, _035422_, _035490_);
  not g_126155_(_035490_, _035491_);
  and g_126156_(_035284_, _035422_, _035492_);
  not g_126157_(_035492_, _035493_);
  and g_126158_(_035490_, _035493_, _035494_);
  or g_126159_(_035491_, _035492_, _035495_);
  and g_126160_(_012760_, _035495_, _035497_);
  or g_126161_(_012573_, _035422_, _035498_);
  or g_126162_(_035290_, _035421_, _035499_);
  and g_126163_(_035498_, _035499_, _035500_);
  and g_126164_(_012767_, _035500_, _035501_);
  or g_126165_(_012760_, _035495_, _035502_);
  or g_126166_(_012599_, _035422_, _035503_);
  not g_126167_(_035503_, _035504_);
  and g_126168_(_035302_, _035422_, _035505_);
  not g_126169_(_035505_, _035506_);
  and g_126170_(_035503_, _035506_, _035508_);
  or g_126171_(_035504_, _035505_, _035509_);
  and g_126172_(_012794_, _035508_, _035510_);
  or g_126173_(_012795_, _035509_, _035511_);
  xor g_126174_(_012761_, _035494_, _035512_);
  xor g_126175_(_012760_, _035494_, _035513_);
  xor g_126176_(_012767_, _035500_, _035514_);
  xor g_126177_(_012766_, _035500_, _035515_);
  and g_126178_(_035512_, _035514_, _035516_);
  or g_126179_(_035513_, _035515_, _035517_);
  and g_126180_(_035511_, _035516_, _035519_);
  or g_126181_(_035510_, _035517_, _035520_);
  or g_126182_(_012588_, _035422_, _035521_);
  not g_126183_(_035521_, _035522_);
  and g_126184_(_035319_, _035422_, _035523_);
  not g_126185_(_035523_, _035524_);
  and g_126186_(_035521_, _035524_, _035525_);
  or g_126187_(_035522_, _035523_, _035526_);
  and g_126188_(_012784_, _035526_, _035527_);
  or g_126189_(_012783_, _035525_, _035528_);
  and g_126190_(_012795_, _035509_, _035530_);
  or g_126191_(_012794_, _035508_, _035531_);
  and g_126192_(_035528_, _035531_, _035532_);
  or g_126193_(_035527_, _035530_, _035533_);
  and g_126194_(_012783_, _035525_, _035534_);
  or g_126195_(_012784_, _035526_, _035535_);
  and g_126196_(_035532_, _035535_, _035536_);
  or g_126197_(_035533_, _035534_, _035537_);
  and g_126198_(_035519_, _035536_, _035538_);
  or g_126199_(_035520_, _035537_, _035539_);
  and g_126200_(_012622_, _035421_, _035541_);
  or g_126201_(_012621_, _035422_, _035542_);
  and g_126202_(_035339_, _035422_, _035543_);
  or g_126203_(_035338_, _035421_, _035544_);
  and g_126204_(_035542_, _035544_, _035545_);
  or g_126205_(_035541_, _035543_, _035546_);
  and g_126206_(_012820_, _035546_, _035547_);
  and g_126207_(_035352_, _035422_, _035548_);
  not g_126208_(_035548_, _035549_);
  or g_126209_(_000143_, _035422_, _035550_);
  not g_126210_(_035550_, _035552_);
  and g_126211_(_035549_, _035550_, _035553_);
  or g_126212_(_035548_, _035552_, _035554_);
  or g_126213_(_012820_, _035546_, _035555_);
  and g_126214_(_000240_, _035553_, _035556_);
  xor g_126215_(_012821_, _035545_, _035557_);
  xor g_126216_(_012820_, _035545_, _035558_);
  xor g_126217_(_000240_, _035553_, _035559_);
  xor g_126218_(_000242_, _035553_, _035560_);
  and g_126219_(_035557_, _035559_, _035561_);
  or g_126220_(_035558_, _035560_, _035563_);
  or g_126221_(_000285_, _035422_, _035564_);
  not g_126222_(_035564_, _035565_);
  and g_126223_(_035366_, _035422_, _035566_);
  or g_126224_(_035365_, _035421_, _035567_);
  and g_126225_(_035564_, _035567_, _035568_);
  or g_126226_(_035565_, _035566_, _035569_);
  and g_126227_(out[721], _035568_, _035570_);
  and g_126228_(out[720], _035428_, _035571_);
  or g_126229_(_000428_, _035427_, _035572_);
  xor g_126230_(out[721], _035568_, _035574_);
  xor g_126231_(_000417_, _035568_, _035575_);
  and g_126232_(_035572_, _035574_, _035576_);
  or g_126233_(_035571_, _035575_, _035577_);
  or g_126234_(_035570_, _035576_, _035578_);
  and g_126235_(_035561_, _035578_, _035579_);
  and g_126236_(_035555_, _035556_, _035580_);
  or g_126237_(_035547_, _035580_, _035581_);
  or g_126238_(_035579_, _035581_, _035582_);
  and g_126239_(_035538_, _035582_, _035583_);
  and g_126240_(_035519_, _035533_, _035585_);
  and g_126241_(_035501_, _035502_, _035586_);
  or g_126242_(_035497_, _035586_, _035587_);
  or g_126243_(_035585_, _035587_, _035588_);
  or g_126244_(_035583_, _035588_, _035589_);
  and g_126245_(_035488_, _035589_, _035590_);
  and g_126246_(_035478_, _035480_, _035591_);
  and g_126247_(_035457_, _035591_, _035592_);
  and g_126248_(_035449_, _035454_, _035593_);
  or g_126249_(_035592_, _035593_, _035594_);
  or g_126250_(_035590_, _035594_, _035596_);
  or g_126251_(out[720], _035428_, _035597_);
  not g_126252_(_035597_, _035598_);
  or g_126253_(_035577_, _035598_, _035599_);
  or g_126254_(_035563_, _035599_, _035600_);
  or g_126255_(_035489_, _035600_, _035601_);
  or g_126256_(_035539_, _035601_, _035602_);
  and g_126257_(_035596_, _035602_, _035603_);
  not g_126258_(_035603_, _035604_);
  and g_126259_(_035428_, _035604_, _035605_);
  and g_126260_(_000428_, _035603_, _035607_);
  or g_126261_(_035605_, _035607_, _035608_);
  and g_126262_(_035429_, _035433_, _035609_);
  or g_126263_(_035431_, _035434_, _035610_);
  or g_126264_(out[746], _012918_, _035611_);
  xor g_126265_(out[747], _035611_, _035612_);
  xor g_126266_(_000494_, _035611_, _035613_);
  and g_126267_(_035609_, _035613_, _035614_);
  or g_126268_(_035610_, _035612_, _035615_);
  and g_126269_(_035444_, _035603_, _035616_);
  not g_126270_(_035616_, _035618_);
  and g_126271_(_035443_, _035604_, _035619_);
  or g_126272_(_035442_, _035603_, _035620_);
  and g_126273_(_035618_, _035620_, _035621_);
  or g_126274_(_035616_, _035619_, _035622_);
  xor g_126275_(out[746], _012918_, _035623_);
  xor g_126276_(_000615_, _012918_, _035624_);
  and g_126277_(_035621_, _035623_, _035625_);
  or g_126278_(_035622_, _035624_, _035626_);
  and g_126279_(_035615_, _035626_, _035627_);
  or g_126280_(_035614_, _035625_, _035629_);
  and g_126281_(_035610_, _035612_, _035630_);
  or g_126282_(_035627_, _035630_, _035631_);
  and g_126283_(_012733_, _035603_, _035632_);
  and g_126284_(_035473_, _035604_, _035633_);
  or g_126285_(_035632_, _035633_, _035634_);
  not g_126286_(_035634_, _035635_);
  and g_126287_(_012919_, _035635_, _035636_);
  or g_126288_(_012920_, _035634_, _035637_);
  and g_126289_(_035622_, _035624_, _035638_);
  or g_126290_(_035630_, _035638_, _035640_);
  not g_126291_(_035640_, _035641_);
  and g_126292_(_035627_, _035641_, _035642_);
  or g_126293_(_035629_, _035640_, _035643_);
  or g_126294_(_035636_, _035643_, _035644_);
  and g_126295_(_012717_, _035603_, _035645_);
  and g_126296_(_035465_, _035604_, _035646_);
  or g_126297_(_035645_, _035646_, _035647_);
  not g_126298_(_035647_, _035648_);
  or g_126299_(_012931_, _035648_, _035649_);
  or g_126300_(_012919_, _035635_, _035651_);
  and g_126301_(_035649_, _035651_, _035652_);
  and g_126302_(_035495_, _035604_, _035653_);
  and g_126303_(_012761_, _035603_, _035654_);
  or g_126304_(_035653_, _035654_, _035655_);
  and g_126305_(_012950_, _035655_, _035656_);
  or g_126306_(_035500_, _035603_, _035657_);
  or g_126307_(_012766_, _035604_, _035658_);
  and g_126308_(_035657_, _035658_, _035659_);
  not g_126309_(_035659_, _035660_);
  and g_126310_(_012958_, _035659_, _035662_);
  or g_126311_(_035656_, _035662_, _035663_);
  and g_126312_(_035509_, _035604_, _035664_);
  and g_126313_(_012794_, _035603_, _035665_);
  or g_126314_(_035664_, _035665_, _035666_);
  not g_126315_(_035666_, _035667_);
  and g_126316_(_012982_, _035666_, _035668_);
  or g_126317_(_012981_, _035667_, _035669_);
  and g_126318_(_012783_, _035603_, _035670_);
  and g_126319_(_035526_, _035604_, _035671_);
  or g_126320_(_035670_, _035671_, _035673_);
  not g_126321_(_035673_, _035674_);
  and g_126322_(_012971_, _035673_, _035675_);
  or g_126323_(_012970_, _035674_, _035676_);
  and g_126324_(_035669_, _035676_, _035677_);
  or g_126325_(_035668_, _035675_, _035678_);
  and g_126326_(_035545_, _035604_, _035679_);
  or g_126327_(_035546_, _035603_, _035680_);
  and g_126328_(_012820_, _035603_, _035681_);
  not g_126329_(_035681_, _035682_);
  or g_126330_(_035679_, _035681_, _035684_);
  and g_126331_(_035680_, _035682_, _035685_);
  or g_126332_(_013006_, _035684_, _035686_);
  and g_126333_(_013006_, _035684_, _035687_);
  xor g_126334_(_013006_, _035684_, _035688_);
  xor g_126335_(_013005_, _035684_, _035689_);
  and g_126336_(_035554_, _035604_, _035690_);
  and g_126337_(_000240_, _035603_, _035691_);
  or g_126338_(_035690_, _035691_, _035692_);
  not g_126339_(_035692_, _035693_);
  or g_126340_(_000363_, _035692_, _035695_);
  xor g_126341_(_000363_, _035692_, _035696_);
  xor g_126342_(_000363_, _035693_, _035697_);
  and g_126343_(_035688_, _035696_, _035698_);
  or g_126344_(_035689_, _035697_, _035699_);
  and g_126345_(_035569_, _035604_, _035700_);
  or g_126346_(_035568_, _035603_, _035701_);
  and g_126347_(out[721], _035603_, _035702_);
  not g_126348_(_035702_, _035703_);
  and g_126349_(_035701_, _035703_, _035704_);
  or g_126350_(_035700_, _035702_, _035706_);
  or g_126351_(_000549_, _035706_, _035707_);
  and g_126352_(out[736], _035608_, _035708_);
  xor g_126353_(_000549_, _035704_, _035709_);
  or g_126354_(_035708_, _035709_, _035710_);
  and g_126355_(_035707_, _035710_, _035711_);
  or g_126356_(_035699_, _035711_, _035712_);
  and g_126357_(_035686_, _035695_, _035713_);
  or g_126358_(_035687_, _035713_, _035714_);
  and g_126359_(_035712_, _035714_, _035715_);
  and g_126360_(_012970_, _035674_, _035717_);
  or g_126361_(_012971_, _035673_, _035718_);
  or g_126362_(_035715_, _035717_, _035719_);
  and g_126363_(_035677_, _035719_, _035720_);
  or g_126364_(_012982_, _035666_, _035721_);
  and g_126365_(_012956_, _035660_, _035722_);
  or g_126366_(_012932_, _035647_, _035723_);
  or g_126367_(_012950_, _035655_, _035724_);
  and g_126368_(_035637_, _035723_, _035725_);
  and g_126369_(_035652_, _035725_, _035726_);
  and g_126370_(_035642_, _035726_, _035728_);
  not g_126371_(_035728_, _035729_);
  xor g_126372_(_012950_, _035655_, _035730_);
  and g_126373_(_035721_, _035730_, _035731_);
  not g_126374_(_035731_, _035732_);
  or g_126375_(_035722_, _035732_, _035733_);
  xor g_126376_(_012958_, _035659_, _035734_);
  and g_126377_(_035721_, _035734_, _035735_);
  and g_126378_(_035730_, _035735_, _035736_);
  or g_126379_(_035662_, _035733_, _035737_);
  and g_126380_(_035728_, _035736_, _035739_);
  or g_126381_(_035729_, _035737_, _035740_);
  or g_126382_(_035720_, _035740_, _035741_);
  or g_126383_(_035644_, _035652_, _035742_);
  and g_126384_(_035631_, _035742_, _035743_);
  and g_126385_(_035663_, _035724_, _035744_);
  and g_126386_(_035728_, _035744_, _035745_);
  not g_126387_(_035745_, _035746_);
  and g_126388_(_035743_, _035746_, _035747_);
  and g_126389_(_035741_, _035747_, _035748_);
  or g_126390_(out[736], _035608_, _035750_);
  and g_126391_(_035718_, _035750_, _035751_);
  and g_126392_(_035698_, _035751_, _035752_);
  or g_126393_(_035678_, _035710_, _035753_);
  not g_126394_(_035753_, _035754_);
  and g_126395_(_035739_, _035754_, _035755_);
  and g_126396_(_035752_, _035755_, _035756_);
  or g_126397_(_035748_, _035756_, _035757_);
  not g_126398_(_035757_, _035758_);
  and g_126399_(_035608_, _035757_, _035759_);
  and g_126400_(_000560_, _035758_, _035761_);
  or g_126401_(_035759_, _035761_, _035762_);
  and g_126402_(out[737], _035758_, _035763_);
  or g_126403_(_000549_, _035757_, _035764_);
  and g_126404_(_035706_, _035757_, _035765_);
  or g_126405_(_035704_, _035758_, _035766_);
  and g_126406_(_035764_, _035766_, _035767_);
  or g_126407_(_035763_, _035765_, _035768_);
  and g_126408_(out[752], _035762_, _035769_);
  or g_126409_(_000681_, _035768_, _035770_);
  xor g_126410_(_000681_, _035767_, _035772_);
  or g_126411_(_035769_, _035772_, _035773_);
  not g_126412_(_035773_, _035774_);
  or g_126413_(out[752], _035762_, _035775_);
  and g_126414_(_035774_, _035775_, _035776_);
  or g_126415_(_013005_, _035757_, _035777_);
  not g_126416_(_035777_, _035778_);
  and g_126417_(_035685_, _035757_, _035779_);
  or g_126418_(_035684_, _035758_, _035780_);
  and g_126419_(_035777_, _035780_, _035781_);
  or g_126420_(_035778_, _035779_, _035783_);
  or g_126421_(_013146_, _035781_, _035784_);
  and g_126422_(_035692_, _035757_, _035785_);
  or g_126423_(_000363_, _035757_, _035786_);
  not g_126424_(_035786_, _035787_);
  or g_126425_(_035785_, _035787_, _035788_);
  and g_126426_(_013146_, _035781_, _035789_);
  or g_126427_(_000652_, _035788_, _035790_);
  xor g_126428_(_013146_, _035781_, _035791_);
  xor g_126429_(_013145_, _035781_, _035792_);
  xor g_126430_(_000652_, _035788_, _035794_);
  xor g_126431_(_000651_, _035788_, _035795_);
  and g_126432_(_035791_, _035794_, _035796_);
  or g_126433_(_035792_, _035795_, _035797_);
  and g_126434_(_035776_, _035796_, _035798_);
  or g_126435_(_012956_, _035757_, _035799_);
  not g_126436_(_035799_, _035800_);
  and g_126437_(_035660_, _035757_, _035801_);
  not g_126438_(_035801_, _035802_);
  and g_126439_(_035799_, _035802_, _035803_);
  or g_126440_(_035800_, _035801_, _035805_);
  and g_126441_(_013103_, _035803_, _035806_);
  or g_126442_(_013102_, _035805_, _035807_);
  or g_126443_(_012950_, _035757_, _035808_);
  not g_126444_(_035808_, _035809_);
  and g_126445_(_035655_, _035757_, _035810_);
  not g_126446_(_035810_, _035811_);
  and g_126447_(_035808_, _035811_, _035812_);
  or g_126448_(_035809_, _035810_, _035813_);
  and g_126449_(_013095_, _035813_, _035814_);
  or g_126450_(_013096_, _035812_, _035816_);
  and g_126451_(_035807_, _035816_, _035817_);
  or g_126452_(_035806_, _035814_, _035818_);
  and g_126453_(_013102_, _035805_, _035819_);
  and g_126454_(_013096_, _035812_, _035820_);
  or g_126455_(_035819_, _035820_, _035821_);
  or g_126456_(_035818_, _035821_, _035822_);
  not g_126457_(_035822_, _035823_);
  or g_126458_(_012982_, _035757_, _035824_);
  or g_126459_(_035667_, _035758_, _035825_);
  and g_126460_(_035824_, _035825_, _035827_);
  or g_126461_(_013109_, _035827_, _035828_);
  or g_126462_(_012971_, _035757_, _035829_);
  or g_126463_(_035674_, _035758_, _035830_);
  and g_126464_(_035829_, _035830_, _035831_);
  or g_126465_(_013127_, _035831_, _035832_);
  and g_126466_(_035828_, _035832_, _035833_);
  and g_126467_(_013109_, _035827_, _035834_);
  xor g_126468_(_013127_, _035831_, _035835_);
  xor g_126469_(_013109_, _035827_, _035836_);
  and g_126470_(_035835_, _035836_, _035838_);
  not g_126471_(_035838_, _035839_);
  and g_126472_(_035823_, _035838_, _035840_);
  or g_126473_(_035822_, _035839_, _035841_);
  and g_126474_(_035623_, _035758_, _035842_);
  and g_126475_(_035622_, _035757_, _035843_);
  or g_126476_(_035842_, _035843_, _035844_);
  or g_126477_(out[762], _013075_, _035845_);
  xor g_126478_(out[762], _013075_, _035846_);
  not g_126479_(_035846_, _035847_);
  and g_126480_(_035609_, _035612_, _035849_);
  or g_126481_(_035610_, _035613_, _035850_);
  xor g_126482_(out[763], _035845_, _035851_);
  xor g_126483_(_000626_, _035845_, _035852_);
  or g_126484_(_035850_, _035851_, _035853_);
  and g_126485_(_035850_, _035851_, _035854_);
  xor g_126486_(_035849_, _035851_, _035855_);
  or g_126487_(_035844_, _035847_, _035856_);
  xor g_126488_(_035844_, _035846_, _035857_);
  or g_126489_(_035855_, _035857_, _035858_);
  not g_126490_(_035858_, _035860_);
  or g_126491_(_012932_, _035757_, _035861_);
  not g_126492_(_035861_, _035862_);
  and g_126493_(_035647_, _035757_, _035863_);
  not g_126494_(_035863_, _035864_);
  and g_126495_(_035861_, _035864_, _035865_);
  or g_126496_(_035862_, _035863_, _035866_);
  or g_126497_(_013086_, _035865_, _035867_);
  or g_126498_(_012920_, _035757_, _035868_);
  not g_126499_(_035868_, _035869_);
  and g_126500_(_035634_, _035757_, _035871_);
  not g_126501_(_035871_, _035872_);
  and g_126502_(_035868_, _035872_, _035873_);
  or g_126503_(_035869_, _035871_, _035874_);
  or g_126504_(_013076_, _035873_, _035875_);
  and g_126505_(_035867_, _035875_, _035876_);
  not g_126506_(_035876_, _035877_);
  and g_126507_(_013076_, _035873_, _035878_);
  and g_126508_(_013086_, _035865_, _035879_);
  or g_126509_(_035878_, _035879_, _035880_);
  not g_126510_(_035880_, _035882_);
  and g_126511_(_035876_, _035882_, _035883_);
  or g_126512_(_035877_, _035880_, _035884_);
  and g_126513_(_035860_, _035883_, _035885_);
  or g_126514_(_035858_, _035884_, _035886_);
  and g_126515_(_035840_, _035885_, _035887_);
  and g_126516_(_035798_, _035887_, _035888_);
  and g_126517_(_035770_, _035773_, _035889_);
  or g_126518_(_035797_, _035889_, _035890_);
  or g_126519_(_035789_, _035790_, _035891_);
  and g_126520_(_035784_, _035891_, _035893_);
  and g_126521_(_035890_, _035893_, _035894_);
  or g_126522_(_035858_, _035876_, _035895_);
  or g_126523_(_035878_, _035895_, _035896_);
  or g_126524_(_035854_, _035856_, _035897_);
  and g_126525_(_035853_, _035897_, _035898_);
  and g_126526_(_035896_, _035898_, _035899_);
  or g_126527_(_035833_, _035834_, _035900_);
  or g_126528_(_035822_, _035900_, _035901_);
  or g_126529_(_035817_, _035820_, _035902_);
  or g_126530_(_035841_, _035894_, _035904_);
  and g_126531_(_035901_, _035904_, _035905_);
  and g_126532_(_035902_, _035905_, _035906_);
  or g_126533_(_035886_, _035906_, _035907_);
  and g_126534_(_035899_, _035907_, _035908_);
  or g_126535_(_035888_, _035908_, _035909_);
  not g_126536_(_035909_, _035910_);
  and g_126537_(_035762_, _035909_, _035911_);
  not g_126538_(_035911_, _035912_);
  or g_126539_(out[752], _035909_, _035913_);
  not g_126540_(_035913_, _035915_);
  and g_126541_(_035912_, _035913_, _035916_);
  or g_126542_(_035911_, _035915_, _035917_);
  or g_126543_(_013145_, _035909_, _035918_);
  not g_126544_(_035918_, _035919_);
  and g_126545_(_035783_, _035909_, _035920_);
  or g_126546_(_035781_, _035910_, _035921_);
  and g_126547_(_035918_, _035921_, _035922_);
  or g_126548_(_035919_, _035920_, _035923_);
  and g_126549_(_013303_, _035923_, _035924_);
  or g_126550_(_013304_, _035922_, _035926_);
  and g_126551_(_013304_, _035922_, _035927_);
  or g_126552_(_013303_, _035923_, _035928_);
  and g_126553_(_035926_, _035928_, _035929_);
  or g_126554_(_035924_, _035927_, _035930_);
  and g_126555_(_035788_, _035909_, _035931_);
  and g_126556_(_000651_, _035910_, _035932_);
  or g_126557_(_035931_, _035932_, _035933_);
  or g_126558_(_000829_, _035933_, _035934_);
  not g_126559_(_035934_, _035935_);
  xor g_126560_(_000829_, _035933_, _035937_);
  xor g_126561_(_000828_, _035933_, _035938_);
  and g_126562_(_035929_, _035937_, _035939_);
  or g_126563_(_035930_, _035938_, _035940_);
  and g_126564_(_035767_, _035909_, _035941_);
  not g_126565_(_035941_, _035942_);
  or g_126566_(out[753], _035909_, _035943_);
  not g_126567_(_035943_, _035944_);
  or g_126568_(_035941_, _035944_, _035945_);
  and g_126569_(_035942_, _035943_, _035946_);
  and g_126570_(out[769], _035945_, _035948_);
  or g_126571_(_000813_, _035946_, _035949_);
  and g_126572_(out[768], _035917_, _035950_);
  or g_126573_(_000824_, _035916_, _035951_);
  xor g_126574_(out[769], _035945_, _035952_);
  xor g_126575_(_000813_, _035945_, _035953_);
  and g_126576_(_035951_, _035952_, _035954_);
  or g_126577_(_035950_, _035953_, _035955_);
  and g_126578_(_035949_, _035955_, _035956_);
  or g_126579_(_035948_, _035954_, _035957_);
  and g_126580_(_035939_, _035957_, _035959_);
  or g_126581_(_035940_, _035956_, _035960_);
  and g_126582_(_035926_, _035934_, _035961_);
  or g_126583_(_035924_, _035935_, _035962_);
  and g_126584_(_035928_, _035962_, _035963_);
  or g_126585_(_035927_, _035961_, _035964_);
  and g_126586_(_035960_, _035964_, _035965_);
  or g_126587_(_035959_, _035963_, _035966_);
  and g_126588_(_035849_, _035851_, _035967_);
  or g_126589_(_035850_, _035852_, _035968_);
  or g_126590_(out[778], _013223_, _035970_);
  xor g_126591_(out[779], _035970_, _035971_);
  xor g_126592_(_000758_, _035970_, _035972_);
  and g_126593_(_035967_, _035972_, _035973_);
  or g_126594_(_035968_, _035971_, _035974_);
  and g_126595_(_035846_, _035910_, _035975_);
  and g_126596_(_035844_, _035909_, _035976_);
  or g_126597_(_035975_, _035976_, _035977_);
  xor g_126598_(_000879_, _013223_, _035978_);
  or g_126599_(_035977_, _035978_, _035979_);
  not g_126600_(_035979_, _035981_);
  and g_126601_(_035974_, _035979_, _035982_);
  or g_126602_(_035973_, _035981_, _035983_);
  and g_126603_(_035968_, _035971_, _035984_);
  or g_126604_(_035967_, _035972_, _035985_);
  and g_126605_(_035977_, _035978_, _035986_);
  or g_126606_(_035984_, _035986_, _035987_);
  not g_126607_(_035987_, _035988_);
  and g_126608_(_035982_, _035988_, _035989_);
  or g_126609_(_035983_, _035987_, _035990_);
  and g_126610_(_013086_, _035910_, _035992_);
  and g_126611_(_035866_, _035909_, _035993_);
  or g_126612_(_035992_, _035993_, _035994_);
  not g_126613_(_035994_, _035995_);
  and g_126614_(_013233_, _035994_, _035996_);
  or g_126615_(_013231_, _035995_, _035997_);
  and g_126616_(_013076_, _035910_, _035998_);
  and g_126617_(_035874_, _035909_, _035999_);
  or g_126618_(_035998_, _035999_, _036000_);
  not g_126619_(_036000_, _036001_);
  and g_126620_(_013225_, _036000_, _036003_);
  or g_126621_(_013224_, _036001_, _036004_);
  and g_126622_(_035997_, _036004_, _036005_);
  or g_126623_(_035996_, _036003_, _036006_);
  or g_126624_(_013225_, _036000_, _036007_);
  or g_126625_(_013233_, _035994_, _036008_);
  and g_126626_(_036007_, _036008_, _036009_);
  not g_126627_(_036009_, _036010_);
  and g_126628_(_036005_, _036009_, _036011_);
  or g_126629_(_036006_, _036010_, _036012_);
  and g_126630_(_035989_, _036011_, _036014_);
  or g_126631_(_035990_, _036012_, _036015_);
  or g_126632_(_013095_, _035909_, _036016_);
  not g_126633_(_036016_, _036017_);
  and g_126634_(_035813_, _035909_, _036018_);
  or g_126635_(_035812_, _035910_, _036019_);
  and g_126636_(_036016_, _036019_, _036020_);
  or g_126637_(_036017_, _036018_, _036021_);
  and g_126638_(_013259_, _036021_, _036022_);
  or g_126639_(_013260_, _036020_, _036023_);
  or g_126640_(_013102_, _035909_, _036025_);
  not g_126641_(_036025_, _036026_);
  and g_126642_(_035805_, _035909_, _036027_);
  or g_126643_(_035803_, _035910_, _036028_);
  and g_126644_(_036025_, _036028_, _036029_);
  or g_126645_(_036026_, _036027_, _036030_);
  and g_126646_(_013260_, _036020_, _036031_);
  or g_126647_(_013259_, _036021_, _036032_);
  and g_126648_(_013250_, _036029_, _036033_);
  or g_126649_(_013249_, _036030_, _036034_);
  and g_126650_(_036023_, _036032_, _036036_);
  or g_126651_(_036022_, _036031_, _036037_);
  xor g_126652_(_013250_, _036029_, _036038_);
  xor g_126653_(_013249_, _036029_, _036039_);
  and g_126654_(_036036_, _036038_, _036040_);
  or g_126655_(_036037_, _036039_, _036041_);
  and g_126656_(_035827_, _035909_, _036042_);
  not g_126657_(_036042_, _036043_);
  or g_126658_(_013109_, _035909_, _036044_);
  and g_126659_(_036043_, _036044_, _036045_);
  or g_126660_(_013281_, _036045_, _036047_);
  and g_126661_(_035831_, _035909_, _036048_);
  not g_126662_(_036048_, _036049_);
  or g_126663_(_013127_, _035909_, _036050_);
  and g_126664_(_036049_, _036050_, _036051_);
  and g_126665_(_013273_, _036051_, _036052_);
  and g_126666_(_013281_, _036045_, _036053_);
  xor g_126667_(_013281_, _036045_, _036054_);
  xor g_126668_(_013280_, _036045_, _036055_);
  xor g_126669_(_013273_, _036051_, _036056_);
  xor g_126670_(_013272_, _036051_, _036058_);
  and g_126671_(_036054_, _036056_, _036059_);
  or g_126672_(_036055_, _036058_, _036060_);
  and g_126673_(_036040_, _036059_, _036061_);
  or g_126674_(_036041_, _036060_, _036062_);
  and g_126675_(_036014_, _036061_, _036063_);
  or g_126676_(_036015_, _036062_, _036064_);
  and g_126677_(_035966_, _036063_, _036065_);
  and g_126678_(_035983_, _035985_, _036066_);
  or g_126679_(_035982_, _035984_, _036067_);
  and g_126680_(_036006_, _036007_, _036069_);
  not g_126681_(_036069_, _036070_);
  and g_126682_(_035989_, _036069_, _036071_);
  or g_126683_(_035990_, _036070_, _036072_);
  and g_126684_(_036067_, _036072_, _036073_);
  or g_126685_(_036066_, _036071_, _036074_);
  or g_126686_(_036052_, _036053_, _036075_);
  and g_126687_(_036047_, _036075_, _036076_);
  not g_126688_(_036076_, _036077_);
  and g_126689_(_036040_, _036076_, _036078_);
  or g_126690_(_036041_, _036077_, _036080_);
  and g_126691_(_036032_, _036033_, _036081_);
  or g_126692_(_036031_, _036034_, _036082_);
  and g_126693_(_036023_, _036082_, _036083_);
  or g_126694_(_036022_, _036081_, _036084_);
  and g_126695_(_036080_, _036083_, _036085_);
  or g_126696_(_036078_, _036084_, _036086_);
  and g_126697_(_036014_, _036086_, _036087_);
  or g_126698_(_036074_, _036087_, _036088_);
  or g_126699_(_035965_, _036062_, _036089_);
  and g_126700_(_036085_, _036089_, _036091_);
  or g_126701_(_036015_, _036091_, _036092_);
  and g_126702_(_036073_, _036092_, _036093_);
  or g_126703_(_036065_, _036088_, _036094_);
  or g_126704_(out[768], _035917_, _036095_);
  not g_126705_(_036095_, _036096_);
  or g_126706_(_035955_, _036096_, _036097_);
  not g_126707_(_036097_, _036098_);
  and g_126708_(_035939_, _036098_, _036099_);
  or g_126709_(_035940_, _036097_, _036100_);
  and g_126710_(_036063_, _036099_, _036102_);
  or g_126711_(_036064_, _036100_, _036103_);
  and g_126712_(_036094_, _036103_, _036104_);
  or g_126713_(_036093_, _036102_, _036105_);
  and g_126714_(_035917_, _036105_, _036106_);
  not g_126715_(_036106_, _036107_);
  or g_126716_(out[768], _036105_, _036108_);
  not g_126717_(_036108_, _036109_);
  and g_126718_(_036107_, _036108_, _036110_);
  or g_126719_(_036106_, _036109_, _036111_);
  and g_126720_(_035967_, _035971_, _036113_);
  or g_126721_(_035968_, _035972_, _036114_);
  or g_126722_(out[794], _013421_, _036115_);
  xor g_126723_(out[795], _036115_, _036116_);
  xor g_126724_(_000890_, _036115_, _036117_);
  and g_126725_(_036113_, _036117_, _036118_);
  or g_126726_(_036114_, _036116_, _036119_);
  xor g_126727_(out[794], _013421_, _036120_);
  xor g_126728_(_001011_, _013421_, _036121_);
  or g_126729_(_035978_, _036105_, _036122_);
  not g_126730_(_036122_, _036124_);
  and g_126731_(_035977_, _036105_, _036125_);
  not g_126732_(_036125_, _036126_);
  and g_126733_(_036122_, _036126_, _036127_);
  or g_126734_(_036124_, _036125_, _036128_);
  and g_126735_(_036120_, _036127_, _036129_);
  or g_126736_(_036121_, _036128_, _036130_);
  and g_126737_(_036119_, _036130_, _036131_);
  or g_126738_(_036118_, _036129_, _036132_);
  and g_126739_(_036121_, _036128_, _036133_);
  or g_126740_(_036120_, _036127_, _036135_);
  or g_126741_(_013233_, _036105_, _036136_);
  not g_126742_(_036136_, _036137_);
  and g_126743_(_035994_, _036105_, _036138_);
  not g_126744_(_036138_, _036139_);
  and g_126745_(_036136_, _036139_, _036140_);
  or g_126746_(_036137_, _036138_, _036141_);
  and g_126747_(_013431_, _036141_, _036142_);
  or g_126748_(_013429_, _036140_, _036143_);
  or g_126749_(_013225_, _036105_, _036144_);
  not g_126750_(_036144_, _036146_);
  and g_126751_(_036000_, _036105_, _036147_);
  not g_126752_(_036147_, _036148_);
  and g_126753_(_036144_, _036148_, _036149_);
  or g_126754_(_036146_, _036147_, _036150_);
  and g_126755_(_013423_, _036150_, _036151_);
  or g_126756_(_013422_, _036149_, _036152_);
  and g_126757_(_036143_, _036152_, _036153_);
  or g_126758_(_036142_, _036151_, _036154_);
  and g_126759_(_013422_, _036149_, _036155_);
  and g_126760_(_036114_, _036116_, _036157_);
  or g_126761_(_036113_, _036117_, _036158_);
  and g_126762_(_013429_, _036140_, _036159_);
  and g_126763_(_036135_, _036158_, _036160_);
  or g_126764_(_036133_, _036157_, _036161_);
  and g_126765_(_036131_, _036160_, _036162_);
  or g_126766_(_036132_, _036161_, _036163_);
  or g_126767_(_036155_, _036159_, _036164_);
  not g_126768_(_036164_, _036165_);
  and g_126769_(_036153_, _036165_, _036166_);
  or g_126770_(_036154_, _036164_, _036168_);
  and g_126771_(_036162_, _036166_, _036169_);
  or g_126772_(_036163_, _036168_, _036170_);
  or g_126773_(_013249_, _036105_, _036171_);
  or g_126774_(_036029_, _036104_, _036172_);
  and g_126775_(_036171_, _036172_, _036173_);
  and g_126776_(_013456_, _036173_, _036174_);
  xor g_126777_(_013455_, _036173_, _036175_);
  and g_126778_(_013260_, _036104_, _036176_);
  or g_126779_(_013259_, _036105_, _036177_);
  and g_126780_(_036021_, _036105_, _036179_);
  or g_126781_(_036020_, _036104_, _036180_);
  and g_126782_(_036177_, _036180_, _036181_);
  or g_126783_(_036176_, _036179_, _036182_);
  and g_126784_(_013462_, _036182_, _036183_);
  or g_126785_(_013462_, _036182_, _036184_);
  xor g_126786_(_013462_, _036181_, _036185_);
  or g_126787_(_036175_, _036185_, _036186_);
  and g_126788_(_036045_, _036105_, _036187_);
  not g_126789_(_036187_, _036188_);
  or g_126790_(_013281_, _036105_, _036190_);
  not g_126791_(_036190_, _036191_);
  and g_126792_(_036188_, _036190_, _036192_);
  or g_126793_(_036187_, _036191_, _036193_);
  and g_126794_(_013381_, _036193_, _036194_);
  or g_126795_(_013380_, _036192_, _036195_);
  or g_126796_(_013273_, _036105_, _036196_);
  not g_126797_(_036196_, _036197_);
  and g_126798_(_036051_, _036105_, _036198_);
  not g_126799_(_036198_, _036199_);
  and g_126800_(_036196_, _036199_, _036201_);
  or g_126801_(_036197_, _036198_, _036202_);
  and g_126802_(_013371_, _036202_, _036203_);
  or g_126803_(_013370_, _036201_, _036204_);
  and g_126804_(_036195_, _036204_, _036205_);
  or g_126805_(_036194_, _036203_, _036206_);
  and g_126806_(_013380_, _036192_, _036207_);
  or g_126807_(_013381_, _036193_, _036208_);
  and g_126808_(_013370_, _036201_, _036209_);
  or g_126809_(_036186_, _036209_, _036210_);
  not g_126810_(_036210_, _036212_);
  and g_126811_(_036205_, _036208_, _036213_);
  or g_126812_(_036206_, _036207_, _036214_);
  and g_126813_(_036169_, _036213_, _036215_);
  or g_126814_(_036170_, _036214_, _036216_);
  and g_126815_(_036212_, _036215_, _036217_);
  or g_126816_(_036210_, _036216_, _036218_);
  or g_126817_(_000829_, _036105_, _036219_);
  not g_126818_(_036219_, _036220_);
  and g_126819_(_035933_, _036105_, _036221_);
  not g_126820_(_036221_, _036223_);
  and g_126821_(_036219_, _036223_, _036224_);
  or g_126822_(_036220_, _036221_, _036225_);
  and g_126823_(_001010_, _036224_, _036226_);
  xor g_126824_(_001010_, _036224_, _036227_);
  or g_126825_(_013303_, _036105_, _036228_);
  not g_126826_(_036228_, _036229_);
  and g_126827_(_035923_, _036105_, _036230_);
  not g_126828_(_036230_, _036231_);
  and g_126829_(_036228_, _036231_, _036232_);
  or g_126830_(_036229_, _036230_, _036234_);
  and g_126831_(_013385_, _036234_, _036235_);
  or g_126832_(_013385_, _036234_, _036236_);
  xor g_126833_(_013387_, _036232_, _036237_);
  and g_126834_(_036227_, _036237_, _036238_);
  or g_126835_(_000813_, _036105_, _036239_);
  or g_126836_(_035945_, _036104_, _036240_);
  and g_126837_(_036239_, _036240_, _036241_);
  and g_126838_(out[785], _036241_, _036242_);
  or g_126839_(_000956_, _036110_, _036243_);
  xor g_126840_(out[785], _036241_, _036245_);
  and g_126841_(_036243_, _036245_, _036246_);
  and g_126842_(_036238_, _036246_, _036247_);
  and g_126843_(_036238_, _036242_, _036248_);
  and g_126844_(_036226_, _036236_, _036249_);
  or g_126845_(_036235_, _036249_, _036250_);
  or g_126846_(_036247_, _036248_, _036251_);
  or g_126847_(_036250_, _036251_, _036252_);
  not g_126848_(_036252_, _036253_);
  or g_126849_(_036218_, _036253_, _036254_);
  or g_126850_(_036186_, _036205_, _036256_);
  or g_126851_(_036207_, _036256_, _036257_);
  and g_126852_(_036174_, _036184_, _036258_);
  or g_126853_(_036183_, _036258_, _036259_);
  not g_126854_(_036259_, _036260_);
  and g_126855_(_036257_, _036260_, _036261_);
  or g_126856_(_036170_, _036261_, _036262_);
  or g_126857_(_036153_, _036155_, _036263_);
  or g_126858_(_036131_, _036157_, _036264_);
  or g_126859_(_036163_, _036263_, _036265_);
  and g_126860_(_036262_, _036265_, _036267_);
  and g_126861_(_036264_, _036267_, _036268_);
  and g_126862_(_036254_, _036268_, _036269_);
  or g_126863_(out[784], _036111_, _036270_);
  and g_126864_(_036247_, _036270_, _036271_);
  and g_126865_(_036217_, _036271_, _036272_);
  or g_126866_(_036269_, _036272_, _036273_);
  not g_126867_(_036273_, _036274_);
  and g_126868_(_036111_, _036273_, _036275_);
  and g_126869_(_000956_, _036274_, _036276_);
  or g_126870_(_036275_, _036276_, _036278_);
  and g_126871_(_036113_, _036116_, _036279_);
  or g_126872_(_036114_, _036117_, _036280_);
  or g_126873_(out[810], _013545_, _036281_);
  xor g_126874_(out[811], _036281_, _036282_);
  xor g_126875_(_001022_, _036281_, _036283_);
  or g_126876_(_036280_, _036282_, _036284_);
  xor g_126877_(out[810], _013545_, _036285_);
  not g_126878_(_036285_, _036286_);
  and g_126879_(_036128_, _036273_, _036287_);
  or g_126880_(_036127_, _036274_, _036289_);
  and g_126881_(_036120_, _036274_, _036290_);
  or g_126882_(_036121_, _036273_, _036291_);
  and g_126883_(_036289_, _036291_, _036292_);
  or g_126884_(_036287_, _036290_, _036293_);
  or g_126885_(_036286_, _036293_, _036294_);
  and g_126886_(_036284_, _036294_, _036295_);
  or g_126887_(_036285_, _036292_, _036296_);
  and g_126888_(_036295_, _036296_, _036297_);
  not g_126889_(_036297_, _036298_);
  and g_126890_(_013429_, _036274_, _036300_);
  or g_126891_(_013431_, _036273_, _036301_);
  and g_126892_(_036141_, _036273_, _036302_);
  or g_126893_(_036140_, _036274_, _036303_);
  and g_126894_(_036301_, _036303_, _036304_);
  or g_126895_(_036300_, _036302_, _036305_);
  or g_126896_(_013537_, _036304_, _036306_);
  and g_126897_(_013422_, _036274_, _036307_);
  or g_126898_(_013423_, _036273_, _036308_);
  and g_126899_(_036150_, _036273_, _036309_);
  or g_126900_(_036149_, _036274_, _036311_);
  and g_126901_(_036308_, _036311_, _036312_);
  or g_126902_(_036307_, _036309_, _036313_);
  or g_126903_(_013546_, _036312_, _036314_);
  and g_126904_(_036306_, _036314_, _036315_);
  not g_126905_(_036315_, _036316_);
  and g_126906_(_013546_, _036312_, _036317_);
  and g_126907_(_036280_, _036282_, _036318_);
  and g_126908_(_013537_, _036304_, _036319_);
  or g_126909_(_036318_, _036319_, _036320_);
  or g_126910_(_036317_, _036320_, _036322_);
  or g_126911_(_036316_, _036322_, _036323_);
  or g_126912_(_036298_, _036323_, _036324_);
  or g_126913_(_013462_, _036273_, _036325_);
  not g_126914_(_036325_, _036326_);
  and g_126915_(_036182_, _036273_, _036327_);
  or g_126916_(_036181_, _036274_, _036328_);
  and g_126917_(_036325_, _036328_, _036329_);
  or g_126918_(_036326_, _036327_, _036330_);
  or g_126919_(_013506_, _036329_, _036331_);
  and g_126920_(_013506_, _036329_, _036333_);
  xor g_126921_(_013505_, _036329_, _036334_);
  or g_126922_(_013455_, _036273_, _036335_);
  or g_126923_(_036173_, _036274_, _036336_);
  and g_126924_(_036335_, _036336_, _036337_);
  not g_126925_(_036337_, _036338_);
  or g_126926_(_013497_, _036338_, _036339_);
  xor g_126927_(_013497_, _036337_, _036340_);
  or g_126928_(_036334_, _036340_, _036341_);
  and g_126929_(_013370_, _036274_, _036342_);
  or g_126930_(_013371_, _036273_, _036344_);
  and g_126931_(_036202_, _036273_, _036345_);
  or g_126932_(_036201_, _036274_, _036346_);
  and g_126933_(_036344_, _036346_, _036347_);
  or g_126934_(_036342_, _036345_, _036348_);
  or g_126935_(_013578_, _036347_, _036349_);
  and g_126936_(_013380_, _036274_, _036350_);
  or g_126937_(_013381_, _036273_, _036351_);
  and g_126938_(_036193_, _036273_, _036352_);
  or g_126939_(_036192_, _036274_, _036353_);
  and g_126940_(_036351_, _036353_, _036355_);
  or g_126941_(_036350_, _036352_, _036356_);
  or g_126942_(_013516_, _036355_, _036357_);
  and g_126943_(_036349_, _036357_, _036358_);
  not g_126944_(_036358_, _036359_);
  and g_126945_(_013516_, _036355_, _036360_);
  and g_126946_(_013578_, _036347_, _036361_);
  or g_126947_(_036360_, _036361_, _036362_);
  or g_126948_(_036359_, _036362_, _036363_);
  or g_126949_(_036341_, _036363_, _036364_);
  or g_126950_(_036324_, _036364_, _036366_);
  or g_126951_(_013385_, _036273_, _036367_);
  not g_126952_(_036367_, _036368_);
  and g_126953_(_036234_, _036273_, _036369_);
  or g_126954_(_036232_, _036274_, _036370_);
  and g_126955_(_036367_, _036370_, _036371_);
  or g_126956_(_036368_, _036369_, _036372_);
  or g_126957_(_013599_, _036371_, _036373_);
  and g_126958_(_013599_, _036371_, _036374_);
  xor g_126959_(_013598_, _036371_, _036375_);
  and g_126960_(_036225_, _036273_, _036377_);
  and g_126961_(_001010_, _036274_, _036378_);
  or g_126962_(_036377_, _036378_, _036379_);
  or g_126963_(_001212_, _036379_, _036380_);
  xor g_126964_(_001211_, _036379_, _036381_);
  or g_126965_(_036375_, _036381_, _036382_);
  or g_126966_(out[785], _036273_, _036383_);
  and g_126967_(_036241_, _036273_, _036384_);
  not g_126968_(_036384_, _036385_);
  and g_126969_(_036383_, _036385_, _036386_);
  or g_126970_(_001077_, _036386_, _036388_);
  and g_126971_(out[800], _036278_, _036389_);
  xor g_126972_(out[801], _036386_, _036390_);
  or g_126973_(_036389_, _036390_, _036391_);
  and g_126974_(_036388_, _036391_, _036392_);
  or g_126975_(_036382_, _036392_, _036393_);
  or g_126976_(_036374_, _036380_, _036394_);
  and g_126977_(_036373_, _036394_, _036395_);
  and g_126978_(_036393_, _036395_, _036396_);
  or g_126979_(_036366_, _036396_, _036397_);
  or g_126980_(_036341_, _036358_, _036399_);
  or g_126981_(_036360_, _036399_, _036400_);
  or g_126982_(_036333_, _036339_, _036401_);
  and g_126983_(_036331_, _036401_, _036402_);
  and g_126984_(_036400_, _036402_, _036403_);
  or g_126985_(_036324_, _036403_, _036404_);
  or g_126986_(_036315_, _036317_, _036405_);
  or g_126987_(_036298_, _036405_, _036406_);
  and g_126988_(_036295_, _036406_, _036407_);
  or g_126989_(_036318_, _036407_, _036408_);
  and g_126990_(_036404_, _036408_, _036410_);
  and g_126991_(_036397_, _036410_, _036411_);
  or g_126992_(out[800], _036278_, _036412_);
  or g_126993_(_036382_, _036391_, _036413_);
  or g_126994_(_036366_, _036413_, _036414_);
  not g_126995_(_036414_, _036415_);
  and g_126996_(_036412_, _036415_, _036416_);
  or g_126997_(_036411_, _036416_, _036417_);
  not g_126998_(_036417_, _036418_);
  and g_126999_(_036278_, _036417_, _036419_);
  and g_127000_(_001088_, _036418_, _036421_);
  or g_127001_(_036419_, _036421_, _036422_);
  or g_127002_(_013598_, _036417_, _036423_);
  not g_127003_(_036423_, _036424_);
  and g_127004_(_036372_, _036417_, _036425_);
  or g_127005_(_036371_, _036418_, _036426_);
  and g_127006_(_036423_, _036426_, _036427_);
  or g_127007_(_036424_, _036425_, _036428_);
  or g_127008_(_013803_, _036427_, _036429_);
  and g_127009_(_013803_, _036427_, _036430_);
  xor g_127010_(_013803_, _036427_, _036432_);
  xor g_127011_(_013802_, _036427_, _036433_);
  and g_127012_(_036379_, _036417_, _036434_);
  and g_127013_(_001211_, _036418_, _036435_);
  or g_127014_(_036434_, _036435_, _036436_);
  or g_127015_(_001340_, _036436_, _036437_);
  xor g_127016_(_001340_, _036436_, _036438_);
  xor g_127017_(_001339_, _036436_, _036439_);
  and g_127018_(_036432_, _036438_, _036440_);
  or g_127019_(_036433_, _036439_, _036441_);
  and g_127020_(out[801], _036418_, _036443_);
  or g_127021_(_001077_, _036417_, _036444_);
  and g_127022_(_036386_, _036417_, _036445_);
  not g_127023_(_036445_, _036446_);
  and g_127024_(_036444_, _036446_, _036447_);
  or g_127025_(_036443_, _036445_, _036448_);
  or g_127026_(_001209_, _036448_, _036449_);
  and g_127027_(out[816], _036422_, _036450_);
  not g_127028_(_036450_, _036451_);
  xor g_127029_(out[817], _036447_, _036452_);
  xor g_127030_(_001209_, _036447_, _036454_);
  and g_127031_(_036451_, _036452_, _036455_);
  or g_127032_(_036450_, _036454_, _036456_);
  and g_127033_(_036449_, _036456_, _036457_);
  or g_127034_(_036441_, _036457_, _036458_);
  and g_127035_(_036429_, _036437_, _036459_);
  or g_127036_(_036430_, _036459_, _036460_);
  and g_127037_(_036458_, _036460_, _036461_);
  and g_127038_(_036279_, _036282_, _036462_);
  or g_127039_(_036280_, _036283_, _036463_);
  or g_127040_(out[826], _013698_, _036465_);
  xor g_127041_(out[827], _036465_, _036466_);
  xor g_127042_(_001154_, _036465_, _036467_);
  and g_127043_(_036462_, _036467_, _036468_);
  or g_127044_(_036463_, _036466_, _036469_);
  xor g_127045_(out[826], _013698_, _036470_);
  xor g_127046_(_001275_, _013698_, _036471_);
  and g_127047_(_036285_, _036418_, _036472_);
  or g_127048_(_036286_, _036417_, _036473_);
  and g_127049_(_036293_, _036417_, _036474_);
  or g_127050_(_036292_, _036418_, _036476_);
  and g_127051_(_036473_, _036476_, _036477_);
  or g_127052_(_036472_, _036474_, _036478_);
  and g_127053_(_036470_, _036477_, _036479_);
  or g_127054_(_036471_, _036478_, _036480_);
  and g_127055_(_036469_, _036480_, _036481_);
  or g_127056_(_036468_, _036479_, _036482_);
  and g_127057_(_036471_, _036478_, _036483_);
  and g_127058_(_036463_, _036466_, _036484_);
  or g_127059_(_036483_, _036484_, _036485_);
  not g_127060_(_036485_, _036487_);
  and g_127061_(_036481_, _036487_, _036488_);
  or g_127062_(_036482_, _036485_, _036489_);
  and g_127063_(_036304_, _036417_, _036490_);
  or g_127064_(_036305_, _036418_, _036491_);
  or g_127065_(_013537_, _036417_, _036492_);
  not g_127066_(_036492_, _036493_);
  or g_127067_(_036490_, _036493_, _036494_);
  and g_127068_(_036491_, _036492_, _036495_);
  and g_127069_(_013718_, _036495_, _036496_);
  not g_127070_(_036496_, _036498_);
  and g_127071_(_013546_, _036418_, _036499_);
  or g_127072_(_013547_, _036417_, _036500_);
  and g_127073_(_036313_, _036417_, _036501_);
  or g_127074_(_036312_, _036418_, _036502_);
  and g_127075_(_036500_, _036502_, _036503_);
  or g_127076_(_036499_, _036501_, _036504_);
  and g_127077_(_013700_, _036504_, _036505_);
  not g_127078_(_036505_, _036506_);
  and g_127079_(_036498_, _036506_, _036507_);
  or g_127080_(_036496_, _036505_, _036509_);
  and g_127081_(_013699_, _036503_, _036510_);
  or g_127082_(_013700_, _036504_, _036511_);
  and g_127083_(_013717_, _036494_, _036512_);
  or g_127084_(_013718_, _036495_, _036513_);
  and g_127085_(_036511_, _036513_, _036514_);
  or g_127086_(_036510_, _036512_, _036515_);
  and g_127087_(_036507_, _036514_, _036516_);
  or g_127088_(_036509_, _036515_, _036517_);
  and g_127089_(_036488_, _036516_, _036518_);
  or g_127090_(_036489_, _036517_, _036520_);
  and g_127091_(_013506_, _036418_, _036521_);
  and g_127092_(_036330_, _036417_, _036522_);
  or g_127093_(_036521_, _036522_, _036523_);
  and g_127094_(_013739_, _036523_, _036524_);
  or g_127095_(_013739_, _036523_, _036525_);
  xor g_127096_(_013739_, _036523_, _036526_);
  xor g_127097_(_013740_, _036523_, _036527_);
  and g_127098_(_013498_, _036418_, _036528_);
  and g_127099_(_036338_, _036417_, _036529_);
  or g_127100_(_036528_, _036529_, _036531_);
  or g_127101_(_013750_, _036531_, _036532_);
  not g_127102_(_036532_, _036533_);
  xor g_127103_(_013750_, _036531_, _036534_);
  xor g_127104_(_013751_, _036531_, _036535_);
  and g_127105_(_036526_, _036534_, _036536_);
  or g_127106_(_036527_, _036535_, _036537_);
  and g_127107_(_036355_, _036417_, _036538_);
  or g_127108_(_036356_, _036418_, _036539_);
  or g_127109_(_013516_, _036417_, _036540_);
  not g_127110_(_036540_, _036542_);
  or g_127111_(_036538_, _036542_, _036543_);
  and g_127112_(_036539_, _036540_, _036544_);
  or g_127113_(_013779_, _036543_, _036545_);
  and g_127114_(_036347_, _036417_, _036546_);
  or g_127115_(_036348_, _036418_, _036547_);
  or g_127116_(_013578_, _036417_, _036548_);
  not g_127117_(_036548_, _036549_);
  or g_127118_(_036546_, _036549_, _036550_);
  and g_127119_(_036547_, _036548_, _036551_);
  or g_127120_(_013768_, _036550_, _036553_);
  and g_127121_(_036545_, _036553_, _036554_);
  or g_127122_(_013780_, _036544_, _036555_);
  not g_127123_(_036555_, _036556_);
  or g_127124_(_013769_, _036551_, _036557_);
  and g_127125_(_036555_, _036557_, _036558_);
  xor g_127126_(_013780_, _036543_, _036559_);
  xor g_127127_(_013769_, _036550_, _036560_);
  and g_127128_(_036554_, _036558_, _036561_);
  or g_127129_(_036559_, _036560_, _036562_);
  and g_127130_(_036536_, _036561_, _036564_);
  or g_127131_(_036537_, _036562_, _036565_);
  and g_127132_(_036518_, _036564_, _036566_);
  or g_127133_(_036520_, _036565_, _036567_);
  or g_127134_(_036461_, _036567_, _036568_);
  or g_127135_(_036554_, _036556_, _036569_);
  or g_127136_(_036537_, _036569_, _036570_);
  and g_127137_(_036525_, _036533_, _036571_);
  or g_127138_(_036524_, _036571_, _036572_);
  not g_127139_(_036572_, _036573_);
  and g_127140_(_036570_, _036573_, _036575_);
  or g_127141_(_036520_, _036575_, _036576_);
  or g_127142_(_036489_, _036507_, _036577_);
  or g_127143_(_036510_, _036577_, _036578_);
  or g_127144_(_036481_, _036484_, _036579_);
  and g_127145_(_036578_, _036579_, _036580_);
  and g_127146_(_036568_, _036580_, _036581_);
  and g_127147_(_036576_, _036581_, _036582_);
  or g_127148_(out[816], _036422_, _036583_);
  and g_127149_(_036440_, _036583_, _036584_);
  and g_127150_(_036455_, _036584_, _036586_);
  and g_127151_(_036566_, _036586_, _036587_);
  or g_127152_(_036582_, _036587_, _036588_);
  and g_127153_(_036422_, _036588_, _036589_);
  not g_127154_(_036589_, _036590_);
  or g_127155_(out[816], _036588_, _036591_);
  not g_127156_(_036591_, _036592_);
  and g_127157_(_036590_, _036591_, _036593_);
  or g_127158_(_036589_, _036592_, _036594_);
  or g_127159_(out[842], _013956_, _036595_);
  xor g_127160_(out[842], _013956_, _036597_);
  xor g_127161_(_001407_, _013956_, _036598_);
  or g_127162_(_036471_, _036588_, _036599_);
  not g_127163_(_036599_, _036600_);
  and g_127164_(_036478_, _036588_, _036601_);
  not g_127165_(_036601_, _036602_);
  and g_127166_(_036599_, _036602_, _036603_);
  or g_127167_(_036600_, _036601_, _036604_);
  and g_127168_(_036598_, _036604_, _036605_);
  not g_127169_(_036605_, _036606_);
  and g_127170_(_036462_, _036466_, _036608_);
  or g_127171_(_036463_, _036467_, _036609_);
  xor g_127172_(out[843], _036595_, _036610_);
  xor g_127173_(_001286_, _036595_, _036611_);
  and g_127174_(_036609_, _036610_, _036612_);
  or g_127175_(_036608_, _036611_, _036613_);
  or g_127176_(_036605_, _036612_, _036614_);
  or g_127177_(_013718_, _036588_, _036615_);
  not g_127178_(_036615_, _036616_);
  and g_127179_(_036495_, _036588_, _036617_);
  or g_127180_(_036616_, _036617_, _036619_);
  not g_127181_(_036619_, _036620_);
  and g_127182_(_013949_, _036620_, _036621_);
  or g_127183_(_013950_, _036619_, _036622_);
  or g_127184_(_013700_, _036588_, _036623_);
  not g_127185_(_036623_, _036624_);
  and g_127186_(_036504_, _036588_, _036625_);
  or g_127187_(_036624_, _036625_, _036626_);
  not g_127188_(_036626_, _036627_);
  and g_127189_(_013957_, _036627_, _036628_);
  or g_127190_(_013959_, _036626_, _036630_);
  and g_127191_(_036622_, _036630_, _036631_);
  or g_127192_(_036621_, _036628_, _036632_);
  and g_127193_(_036608_, _036611_, _036633_);
  or g_127194_(_036609_, _036610_, _036634_);
  and g_127195_(_036597_, _036603_, _036635_);
  or g_127196_(_036598_, _036604_, _036636_);
  and g_127197_(_036634_, _036636_, _036637_);
  or g_127198_(_036633_, _036635_, _036638_);
  and g_127199_(_013950_, _036619_, _036639_);
  or g_127200_(_013949_, _036620_, _036641_);
  and g_127201_(_013959_, _036626_, _036642_);
  or g_127202_(_013957_, _036627_, _036643_);
  and g_127203_(_036641_, _036643_, _036644_);
  or g_127204_(_036639_, _036642_, _036645_);
  and g_127205_(_036606_, _036637_, _036646_);
  and g_127206_(_036613_, _036646_, _036647_);
  or g_127207_(_036614_, _036638_, _036648_);
  and g_127208_(_036631_, _036644_, _036649_);
  or g_127209_(_036632_, _036645_, _036650_);
  and g_127210_(_036647_, _036649_, _036652_);
  or g_127211_(_036648_, _036650_, _036653_);
  or g_127212_(_013750_, _036588_, _036654_);
  not g_127213_(_036654_, _036655_);
  and g_127214_(_036531_, _036588_, _036656_);
  or g_127215_(_036655_, _036656_, _036657_);
  or g_127216_(_013992_, _036657_, _036658_);
  not g_127217_(_036658_, _036659_);
  xor g_127218_(_013992_, _036657_, _036660_);
  xor g_127219_(_013993_, _036657_, _036661_);
  or g_127220_(_013739_, _036588_, _036663_);
  not g_127221_(_036663_, _036664_);
  and g_127222_(_036523_, _036588_, _036665_);
  not g_127223_(_036665_, _036666_);
  and g_127224_(_036663_, _036666_, _036667_);
  or g_127225_(_036664_, _036665_, _036668_);
  and g_127226_(_013981_, _036668_, _036669_);
  or g_127227_(_013982_, _036667_, _036670_);
  and g_127228_(_013982_, _036667_, _036671_);
  or g_127229_(_013981_, _036668_, _036672_);
  and g_127230_(_036670_, _036672_, _036674_);
  or g_127231_(_036669_, _036671_, _036675_);
  and g_127232_(_036660_, _036674_, _036676_);
  or g_127233_(_036661_, _036675_, _036677_);
  or g_127234_(_013780_, _036588_, _036678_);
  not g_127235_(_036678_, _036679_);
  and g_127236_(_036544_, _036588_, _036680_);
  not g_127237_(_036680_, _036681_);
  and g_127238_(_036678_, _036681_, _036682_);
  or g_127239_(_036679_, _036680_, _036683_);
  and g_127240_(_014022_, _036683_, _036685_);
  or g_127241_(_014021_, _036682_, _036686_);
  or g_127242_(_013769_, _036588_, _036687_);
  not g_127243_(_036687_, _036688_);
  and g_127244_(_036551_, _036588_, _036689_);
  not g_127245_(_036689_, _036690_);
  and g_127246_(_036687_, _036690_, _036691_);
  or g_127247_(_036688_, _036689_, _036692_);
  and g_127248_(_014011_, _036692_, _036693_);
  or g_127249_(_014010_, _036691_, _036694_);
  and g_127250_(_036686_, _036694_, _036696_);
  or g_127251_(_036685_, _036693_, _036697_);
  or g_127252_(_014011_, _036692_, _036698_);
  or g_127253_(_014022_, _036683_, _036699_);
  not g_127254_(_036699_, _036700_);
  and g_127255_(_036698_, _036699_, _036701_);
  not g_127256_(_036701_, _036702_);
  and g_127257_(_036696_, _036701_, _036703_);
  or g_127258_(_036697_, _036702_, _036704_);
  and g_127259_(_036676_, _036703_, _036705_);
  or g_127260_(_036677_, _036704_, _036707_);
  and g_127261_(_036652_, _036705_, _036708_);
  or g_127262_(_036653_, _036707_, _036709_);
  or g_127263_(_013802_, _036588_, _036710_);
  not g_127264_(_036710_, _036711_);
  and g_127265_(_036428_, _036588_, _036712_);
  or g_127266_(_036711_, _036712_, _036713_);
  or g_127267_(_013888_, _036713_, _036714_);
  and g_127268_(_036436_, _036588_, _036715_);
  or g_127269_(_001340_, _036588_, _036716_);
  not g_127270_(_036716_, _036718_);
  or g_127271_(_036715_, _036718_, _036719_);
  not g_127272_(_036719_, _036720_);
  and g_127273_(_013888_, _036713_, _036721_);
  and g_127274_(_001515_, _036720_, _036722_);
  xor g_127275_(_013888_, _036713_, _036723_);
  xor g_127276_(_013889_, _036713_, _036724_);
  xor g_127277_(_001516_, _036719_, _036725_);
  xor g_127278_(_001515_, _036719_, _036726_);
  and g_127279_(_036723_, _036725_, _036727_);
  or g_127280_(_036724_, _036726_, _036729_);
  and g_127281_(_036447_, _036588_, _036730_);
  or g_127282_(out[817], _036588_, _036731_);
  not g_127283_(_036731_, _036732_);
  or g_127284_(_036730_, _036732_, _036733_);
  and g_127285_(out[832], _036594_, _036734_);
  or g_127286_(_001352_, _036593_, _036735_);
  and g_127287_(out[833], _036733_, _036736_);
  not g_127288_(_036736_, _036737_);
  xor g_127289_(out[833], _036733_, _036738_);
  xor g_127290_(_001341_, _036733_, _036740_);
  and g_127291_(_036735_, _036738_, _036741_);
  or g_127292_(_036734_, _036740_, _036742_);
  and g_127293_(_001352_, _036593_, _036743_);
  or g_127294_(_036742_, _036743_, _036744_);
  or g_127295_(_036729_, _036744_, _036745_);
  or g_127296_(_036709_, _036745_, _036746_);
  not g_127297_(_036746_, _036747_);
  and g_127298_(_036737_, _036742_, _036748_);
  or g_127299_(_036736_, _036741_, _036749_);
  and g_127300_(_036727_, _036749_, _036751_);
  or g_127301_(_036729_, _036748_, _036752_);
  and g_127302_(_036714_, _036722_, _036753_);
  or g_127303_(_036721_, _036753_, _036754_);
  not g_127304_(_036754_, _036755_);
  and g_127305_(_036752_, _036755_, _036756_);
  or g_127306_(_036751_, _036754_, _036757_);
  and g_127307_(_036708_, _036757_, _036758_);
  or g_127308_(_036709_, _036756_, _036759_);
  and g_127309_(_036697_, _036699_, _036760_);
  or g_127310_(_036696_, _036700_, _036762_);
  and g_127311_(_036676_, _036760_, _036763_);
  or g_127312_(_036677_, _036762_, _036764_);
  and g_127313_(_036659_, _036672_, _036765_);
  or g_127314_(_036658_, _036671_, _036766_);
  and g_127315_(_036670_, _036766_, _036767_);
  or g_127316_(_036669_, _036765_, _036768_);
  and g_127317_(_036764_, _036767_, _036769_);
  or g_127318_(_036763_, _036768_, _036770_);
  and g_127319_(_036652_, _036770_, _036771_);
  or g_127320_(_036653_, _036769_, _036773_);
  and g_127321_(_036606_, _036630_, _036774_);
  or g_127322_(_036605_, _036628_, _036775_);
  and g_127323_(_036645_, _036774_, _036776_);
  or g_127324_(_036644_, _036775_, _036777_);
  and g_127325_(_036637_, _036777_, _036778_);
  or g_127326_(_036638_, _036776_, _036779_);
  and g_127327_(_036613_, _036779_, _036780_);
  or g_127328_(_036612_, _036778_, _036781_);
  and g_127329_(_036773_, _036781_, _036782_);
  or g_127330_(_036771_, _036780_, _036784_);
  and g_127331_(_036759_, _036782_, _036785_);
  or g_127332_(_036758_, _036784_, _036786_);
  and g_127333_(_036746_, _036786_, _036787_);
  or g_127334_(_036747_, _036785_, _036788_);
  and g_127335_(_036594_, _036788_, _036789_);
  and g_127336_(_001352_, _036787_, _036790_);
  or g_127337_(_036789_, _036790_, _036791_);
  or g_127338_(_013950_, _036788_, _036792_);
  not g_127339_(_036792_, _036793_);
  and g_127340_(_036619_, _036788_, _036795_);
  not g_127341_(_036795_, _036796_);
  and g_127342_(_036792_, _036796_, _036797_);
  or g_127343_(_036793_, _036795_, _036798_);
  and g_127344_(_014118_, _036798_, _036799_);
  or g_127345_(_014117_, _036797_, _036800_);
  or g_127346_(_013959_, _036788_, _036801_);
  not g_127347_(_036801_, _036802_);
  and g_127348_(_036626_, _036788_, _036803_);
  not g_127349_(_036803_, _036804_);
  and g_127350_(_036801_, _036804_, _036806_);
  or g_127351_(_036802_, _036803_, _036807_);
  and g_127352_(_014108_, _036807_, _036808_);
  or g_127353_(_014107_, _036806_, _036809_);
  and g_127354_(_036800_, _036809_, _036810_);
  or g_127355_(_036799_, _036808_, _036811_);
  and g_127356_(_036608_, _036610_, _036812_);
  or g_127357_(_036609_, _036611_, _036813_);
  or g_127358_(out[858], _014106_, _036814_);
  xor g_127359_(out[859], _036814_, _036815_);
  xor g_127360_(_001418_, _036814_, _036817_);
  and g_127361_(_036813_, _036815_, _036818_);
  and g_127362_(_014117_, _036797_, _036819_);
  or g_127363_(_014118_, _036798_, _036820_);
  and g_127364_(_036812_, _036817_, _036821_);
  or g_127365_(_036813_, _036815_, _036822_);
  xor g_127366_(out[858], _014106_, _036823_);
  xor g_127367_(_001539_, _014106_, _036824_);
  and g_127368_(_036604_, _036788_, _036825_);
  not g_127369_(_036825_, _036826_);
  or g_127370_(_036598_, _036788_, _036828_);
  not g_127371_(_036828_, _036829_);
  and g_127372_(_036826_, _036828_, _036830_);
  or g_127373_(_036825_, _036829_, _036831_);
  and g_127374_(_036823_, _036830_, _036832_);
  or g_127375_(_036824_, _036831_, _036833_);
  and g_127376_(_036822_, _036833_, _036834_);
  or g_127377_(_036821_, _036832_, _036835_);
  and g_127378_(_036824_, _036831_, _036836_);
  and g_127379_(_014107_, _036806_, _036837_);
  or g_127380_(_014108_, _036807_, _036839_);
  or g_127381_(_036836_, _036837_, _036840_);
  or g_127382_(_036818_, _036836_, _036841_);
  not g_127383_(_036841_, _036842_);
  and g_127384_(_036834_, _036842_, _036843_);
  or g_127385_(_036835_, _036841_, _036844_);
  and g_127386_(_036820_, _036839_, _036845_);
  or g_127387_(_036819_, _036837_, _036846_);
  and g_127388_(_036810_, _036845_, _036847_);
  or g_127389_(_036811_, _036846_, _036848_);
  and g_127390_(_036843_, _036847_, _036850_);
  or g_127391_(_036844_, _036848_, _036851_);
  and g_127392_(_013982_, _036787_, _036852_);
  or g_127393_(_013981_, _036788_, _036853_);
  and g_127394_(_036668_, _036788_, _036854_);
  or g_127395_(_036667_, _036787_, _036855_);
  and g_127396_(_036853_, _036855_, _036856_);
  or g_127397_(_036852_, _036854_, _036857_);
  and g_127398_(_014147_, _036857_, _036858_);
  or g_127399_(_014147_, _036857_, _036859_);
  xor g_127400_(_014148_, _036856_, _036861_);
  xor g_127401_(_014147_, _036856_, _036862_);
  or g_127402_(_013992_, _036788_, _036863_);
  not g_127403_(_036863_, _036864_);
  and g_127404_(_036657_, _036788_, _036865_);
  not g_127405_(_036865_, _036866_);
  and g_127406_(_036863_, _036866_, _036867_);
  or g_127407_(_036864_, _036865_, _036868_);
  and g_127408_(_014154_, _036867_, _036869_);
  xor g_127409_(_014154_, _036867_, _036870_);
  xor g_127410_(_014153_, _036867_, _036872_);
  and g_127411_(_036861_, _036870_, _036873_);
  or g_127412_(_036862_, _036872_, _036874_);
  and g_127413_(_014010_, _036787_, _036875_);
  and g_127414_(_036692_, _036788_, _036876_);
  or g_127415_(_036875_, _036876_, _036877_);
  and g_127416_(_014182_, _036877_, _036878_);
  and g_127417_(_014021_, _036787_, _036879_);
  and g_127418_(_036683_, _036788_, _036880_);
  or g_127419_(_036879_, _036880_, _036881_);
  and g_127420_(_014169_, _036881_, _036883_);
  or g_127421_(_036878_, _036883_, _036884_);
  or g_127422_(_014169_, _036881_, _036885_);
  not g_127423_(_036885_, _036886_);
  or g_127424_(_014182_, _036877_, _036887_);
  and g_127425_(_036885_, _036887_, _036888_);
  not g_127426_(_036888_, _036889_);
  or g_127427_(_036884_, _036886_, _036890_);
  not g_127428_(_036890_, _036891_);
  and g_127429_(_036887_, _036891_, _036892_);
  or g_127430_(_036884_, _036889_, _036894_);
  and g_127431_(_036873_, _036892_, _036895_);
  or g_127432_(_036874_, _036894_, _036896_);
  and g_127433_(_036850_, _036895_, _036897_);
  or g_127434_(_036851_, _036896_, _036898_);
  and g_127435_(_013889_, _036787_, _036899_);
  and g_127436_(_036713_, _036788_, _036900_);
  or g_127437_(_036899_, _036900_, _036901_);
  not g_127438_(_036901_, _036902_);
  and g_127439_(_014206_, _036901_, _036903_);
  or g_127440_(_014207_, _036902_, _036905_);
  and g_127441_(_036719_, _036788_, _036906_);
  and g_127442_(_001515_, _036787_, _036907_);
  or g_127443_(_036906_, _036907_, _036908_);
  and g_127444_(_001846_, _036908_, _036909_);
  or g_127445_(_036903_, _036909_, _036910_);
  and g_127446_(_014207_, _036902_, _036911_);
  or g_127447_(_014206_, _036901_, _036912_);
  or g_127448_(_001846_, _036908_, _036913_);
  not g_127449_(_036913_, _036914_);
  or g_127450_(_036911_, _036914_, _036916_);
  and g_127451_(_036905_, _036912_, _036917_);
  xor g_127452_(_001846_, _036908_, _036918_);
  and g_127453_(_036917_, _036918_, _036919_);
  or g_127454_(_036910_, _036916_, _036920_);
  or g_127455_(_001341_, _036788_, _036921_);
  or g_127456_(_036733_, _036787_, _036922_);
  and g_127457_(_036921_, _036922_, _036923_);
  and g_127458_(out[849], _036923_, _036924_);
  not g_127459_(_036924_, _036925_);
  and g_127460_(out[848], _036791_, _036927_);
  not g_127461_(_036927_, _036928_);
  xor g_127462_(out[849], _036923_, _036929_);
  xor g_127463_(_001473_, _036923_, _036930_);
  and g_127464_(_036928_, _036929_, _036931_);
  or g_127465_(_036927_, _036930_, _036932_);
  and g_127466_(_036925_, _036932_, _036933_);
  or g_127467_(_036924_, _036931_, _036934_);
  and g_127468_(_036919_, _036934_, _036935_);
  or g_127469_(_036920_, _036933_, _036936_);
  and g_127470_(_036912_, _036914_, _036938_);
  or g_127471_(_036911_, _036913_, _036939_);
  and g_127472_(_036905_, _036939_, _036940_);
  or g_127473_(_036903_, _036938_, _036941_);
  and g_127474_(_036936_, _036940_, _036942_);
  or g_127475_(_036935_, _036941_, _036943_);
  and g_127476_(_036897_, _036943_, _036944_);
  or g_127477_(_036898_, _036942_, _036945_);
  and g_127478_(_036884_, _036885_, _036946_);
  and g_127479_(_036873_, _036946_, _036947_);
  and g_127480_(_036859_, _036869_, _036949_);
  or g_127481_(_036947_, _036949_, _036950_);
  or g_127482_(_036858_, _036950_, _036951_);
  and g_127483_(_036850_, _036951_, _036952_);
  not g_127484_(_036952_, _036953_);
  or g_127485_(_036810_, _036840_, _036954_);
  and g_127486_(_036834_, _036954_, _036955_);
  or g_127487_(_036818_, _036955_, _036956_);
  not g_127488_(_036956_, _036957_);
  or g_127489_(_036952_, _036957_, _036958_);
  and g_127490_(_036945_, _036956_, _036960_);
  and g_127491_(_036953_, _036960_, _036961_);
  or g_127492_(_036944_, _036958_, _036962_);
  or g_127493_(out[848], _036791_, _036963_);
  and g_127494_(_036919_, _036963_, _036964_);
  not g_127495_(_036964_, _036965_);
  and g_127496_(_036931_, _036964_, _036966_);
  or g_127497_(_036932_, _036965_, _036967_);
  and g_127498_(_036897_, _036966_, _036968_);
  or g_127499_(_036898_, _036967_, _036969_);
  and g_127500_(_036962_, _036969_, _036971_);
  or g_127501_(_036961_, _036968_, _036972_);
  and g_127502_(_036791_, _036972_, _036973_);
  not g_127503_(_036973_, _036974_);
  or g_127504_(out[848], _036972_, _036975_);
  not g_127505_(_036975_, _036976_);
  and g_127506_(_036974_, _036975_, _036977_);
  or g_127507_(_036973_, _036976_, _036978_);
  or g_127508_(_014206_, _036972_, _036979_);
  not g_127509_(_036979_, _036980_);
  and g_127510_(_036901_, _036972_, _036982_);
  not g_127511_(_036982_, _036983_);
  and g_127512_(_036979_, _036983_, _036984_);
  or g_127513_(_036980_, _036982_, _036985_);
  and g_127514_(_014399_, _036985_, _036986_);
  or g_127515_(_014400_, _036984_, _036987_);
  and g_127516_(_014400_, _036984_, _036988_);
  or g_127517_(_014399_, _036985_, _036989_);
  and g_127518_(_036987_, _036989_, _036990_);
  or g_127519_(_036986_, _036988_, _036991_);
  and g_127520_(_036908_, _036972_, _036993_);
  and g_127521_(_001845_, _036971_, _036994_);
  or g_127522_(_036993_, _036994_, _036995_);
  and g_127523_(_002017_, _036995_, _036996_);
  or g_127524_(_002017_, _036995_, _036997_);
  not g_127525_(_036997_, _036998_);
  xor g_127526_(_002017_, _036995_, _036999_);
  or g_127527_(_036991_, _036998_, _037000_);
  and g_127528_(_036990_, _036999_, _037001_);
  or g_127529_(_036996_, _037000_, _037002_);
  or g_127530_(_001473_, _036972_, _037004_);
  or g_127531_(_036923_, _036971_, _037005_);
  and g_127532_(_037004_, _037005_, _037006_);
  and g_127533_(out[865], _037006_, _037007_);
  not g_127534_(_037007_, _037008_);
  and g_127535_(out[864], _036978_, _037009_);
  or g_127536_(_001616_, _036977_, _037010_);
  xor g_127537_(out[865], _037006_, _037011_);
  xor g_127538_(_001605_, _037006_, _037012_);
  and g_127539_(_037010_, _037011_, _037013_);
  or g_127540_(_037009_, _037012_, _037015_);
  and g_127541_(_037008_, _037015_, _037016_);
  or g_127542_(_037007_, _037013_, _037017_);
  and g_127543_(_037001_, _037017_, _037018_);
  or g_127544_(_037002_, _037016_, _037019_);
  and g_127545_(_036987_, _036997_, _037020_);
  or g_127546_(_036986_, _036998_, _037021_);
  and g_127547_(_036989_, _037021_, _037022_);
  or g_127548_(_036988_, _037020_, _037023_);
  and g_127549_(_037019_, _037023_, _037024_);
  or g_127550_(_037018_, _037022_, _037026_);
  and g_127551_(_036812_, _036815_, _037027_);
  or g_127552_(_036813_, _036817_, _037028_);
  or g_127553_(out[874], _014314_, _037029_);
  xor g_127554_(out[875], _037029_, _037030_);
  xor g_127555_(_001550_, _037029_, _037031_);
  and g_127556_(_037027_, _037031_, _037032_);
  or g_127557_(_037028_, _037030_, _037033_);
  xor g_127558_(out[874], _014314_, _037034_);
  xor g_127559_(_001671_, _014314_, _037035_);
  or g_127560_(_036824_, _036972_, _037037_);
  not g_127561_(_037037_, _037038_);
  and g_127562_(_036831_, _036972_, _037039_);
  not g_127563_(_037039_, _037040_);
  and g_127564_(_037037_, _037040_, _037041_);
  or g_127565_(_037038_, _037039_, _037042_);
  and g_127566_(_037034_, _037041_, _037043_);
  or g_127567_(_037035_, _037042_, _037044_);
  and g_127568_(_037033_, _037044_, _037045_);
  or g_127569_(_037032_, _037043_, _037046_);
  and g_127570_(_037035_, _037042_, _037048_);
  or g_127571_(_037034_, _037041_, _037049_);
  and g_127572_(_014117_, _036971_, _037050_);
  or g_127573_(_014118_, _036972_, _037051_);
  and g_127574_(_036798_, _036972_, _037052_);
  or g_127575_(_036797_, _036971_, _037053_);
  and g_127576_(_037051_, _037053_, _037054_);
  or g_127577_(_037050_, _037052_, _037055_);
  and g_127578_(_014323_, _037055_, _037056_);
  or g_127579_(_014322_, _037054_, _037057_);
  and g_127580_(_014107_, _036971_, _037059_);
  or g_127581_(_014108_, _036972_, _037060_);
  and g_127582_(_036807_, _036972_, _037061_);
  or g_127583_(_036806_, _036971_, _037062_);
  and g_127584_(_037060_, _037062_, _037063_);
  or g_127585_(_037059_, _037061_, _037064_);
  and g_127586_(_014316_, _037064_, _037065_);
  or g_127587_(_014315_, _037063_, _037066_);
  and g_127588_(_037057_, _037066_, _037067_);
  or g_127589_(_037056_, _037065_, _037068_);
  or g_127590_(_014316_, _037064_, _037070_);
  and g_127591_(_037028_, _037030_, _037071_);
  or g_127592_(_037027_, _037031_, _037072_);
  or g_127593_(_014323_, _037055_, _037073_);
  and g_127594_(_037049_, _037072_, _037074_);
  or g_127595_(_037048_, _037071_, _037075_);
  and g_127596_(_037045_, _037074_, _037076_);
  or g_127597_(_037046_, _037075_, _037077_);
  and g_127598_(_037070_, _037073_, _037078_);
  not g_127599_(_037078_, _037079_);
  and g_127600_(_037067_, _037078_, _037081_);
  or g_127601_(_037068_, _037079_, _037082_);
  and g_127602_(_037076_, _037081_, _037083_);
  or g_127603_(_037077_, _037082_, _037084_);
  and g_127604_(_014154_, _036971_, _037085_);
  or g_127605_(_014153_, _036972_, _037086_);
  and g_127606_(_036868_, _036972_, _037087_);
  or g_127607_(_036867_, _036971_, _037088_);
  and g_127608_(_037086_, _037088_, _037089_);
  or g_127609_(_037085_, _037087_, _037090_);
  and g_127610_(_014353_, _037089_, _037092_);
  or g_127611_(_014352_, _037090_, _037093_);
  and g_127612_(_014148_, _036971_, _037094_);
  or g_127613_(_014147_, _036972_, _037095_);
  and g_127614_(_036857_, _036972_, _037096_);
  or g_127615_(_036856_, _036971_, _037097_);
  and g_127616_(_037095_, _037097_, _037098_);
  or g_127617_(_037094_, _037096_, _037099_);
  and g_127618_(_014339_, _037099_, _037100_);
  or g_127619_(_014340_, _037098_, _037101_);
  and g_127620_(_037093_, _037101_, _037103_);
  or g_127621_(_037092_, _037100_, _037104_);
  and g_127622_(_014340_, _037098_, _037105_);
  or g_127623_(_014339_, _037099_, _037106_);
  and g_127624_(_014352_, _037090_, _037107_);
  or g_127625_(_014353_, _037089_, _037108_);
  and g_127626_(_037106_, _037108_, _037109_);
  or g_127627_(_037105_, _037107_, _037110_);
  and g_127628_(_037103_, _037109_, _037111_);
  or g_127629_(_037104_, _037110_, _037112_);
  or g_127630_(_014182_, _036972_, _037114_);
  not g_127631_(_037114_, _037115_);
  and g_127632_(_036877_, _036972_, _037116_);
  not g_127633_(_037116_, _037117_);
  and g_127634_(_037114_, _037117_, _037118_);
  or g_127635_(_037115_, _037116_, _037119_);
  and g_127636_(_014368_, _037119_, _037120_);
  or g_127637_(_014367_, _037118_, _037121_);
  or g_127638_(_014169_, _036972_, _037122_);
  not g_127639_(_037122_, _037123_);
  and g_127640_(_036881_, _036972_, _037125_);
  not g_127641_(_037125_, _037126_);
  and g_127642_(_037122_, _037126_, _037127_);
  or g_127643_(_037123_, _037125_, _037128_);
  and g_127644_(_014375_, _037128_, _037129_);
  or g_127645_(_014374_, _037127_, _037130_);
  and g_127646_(_037121_, _037130_, _037131_);
  or g_127647_(_037120_, _037129_, _037132_);
  and g_127648_(_014374_, _037127_, _037133_);
  or g_127649_(_014375_, _037128_, _037134_);
  and g_127650_(_014367_, _037118_, _037136_);
  or g_127651_(_014368_, _037119_, _037137_);
  and g_127652_(_037134_, _037137_, _037138_);
  or g_127653_(_037133_, _037136_, _037139_);
  and g_127654_(_037131_, _037138_, _037140_);
  or g_127655_(_037132_, _037139_, _037141_);
  and g_127656_(_037111_, _037140_, _037142_);
  or g_127657_(_037112_, _037141_, _037143_);
  and g_127658_(_037083_, _037142_, _037144_);
  or g_127659_(_037084_, _037143_, _037145_);
  and g_127660_(_037026_, _037144_, _037147_);
  or g_127661_(_037024_, _037145_, _037148_);
  and g_127662_(_037104_, _037106_, _037149_);
  or g_127663_(_037103_, _037105_, _037150_);
  and g_127664_(_037111_, _037134_, _037151_);
  and g_127665_(_037132_, _037151_, _037152_);
  not g_127666_(_037152_, _037153_);
  and g_127667_(_037150_, _037153_, _037154_);
  or g_127668_(_037149_, _037152_, _037155_);
  and g_127669_(_037083_, _037155_, _037156_);
  or g_127670_(_037084_, _037154_, _037158_);
  and g_127671_(_037068_, _037070_, _037159_);
  not g_127672_(_037159_, _037160_);
  or g_127673_(_037045_, _037071_, _037161_);
  or g_127674_(_037077_, _037160_, _037162_);
  and g_127675_(_037161_, _037162_, _037163_);
  not g_127676_(_037163_, _037164_);
  and g_127677_(_037158_, _037163_, _037165_);
  or g_127678_(_037156_, _037164_, _037166_);
  and g_127679_(_037148_, _037165_, _037167_);
  or g_127680_(_037147_, _037166_, _037169_);
  and g_127681_(_001616_, _036977_, _037170_);
  or g_127682_(_037002_, _037015_, _037171_);
  or g_127683_(_037170_, _037171_, _037172_);
  or g_127684_(_037145_, _037172_, _037173_);
  not g_127685_(_037173_, _037174_);
  and g_127686_(_037169_, _037173_, _037175_);
  or g_127687_(_037167_, _037174_, _037176_);
  and g_127688_(_036978_, _037176_, _037177_);
  and g_127689_(_001616_, _037175_, _037178_);
  or g_127690_(_037177_, _037178_, _037180_);
  and g_127691_(_036995_, _037176_, _037181_);
  or g_127692_(_002017_, _037176_, _037182_);
  not g_127693_(_037182_, _037183_);
  or g_127694_(_037181_, _037183_, _037184_);
  or g_127695_(_002077_, _037184_, _037185_);
  not g_127696_(_037185_, _037186_);
  and g_127697_(_036985_, _037176_, _037187_);
  not g_127698_(_037187_, _037188_);
  or g_127699_(_014399_, _037176_, _037189_);
  not g_127700_(_037189_, _037191_);
  and g_127701_(_037188_, _037189_, _037192_);
  or g_127702_(_037187_, _037191_, _037193_);
  and g_127703_(_014615_, _037193_, _037194_);
  or g_127704_(_014616_, _037192_, _037195_);
  and g_127705_(_037185_, _037195_, _037196_);
  or g_127706_(_037186_, _037194_, _037197_);
  and g_127707_(_002077_, _037184_, _037198_);
  not g_127708_(_037198_, _037199_);
  and g_127709_(_014616_, _037192_, _037200_);
  or g_127710_(_014615_, _037193_, _037202_);
  or g_127711_(_037198_, _037200_, _037203_);
  and g_127712_(_037196_, _037199_, _037204_);
  and g_127713_(_037202_, _037204_, _037205_);
  or g_127714_(_037197_, _037203_, _037206_);
  or g_127715_(_001605_, _037176_, _037207_);
  or g_127716_(_037006_, _037175_, _037208_);
  and g_127717_(_037207_, _037208_, _037209_);
  and g_127718_(out[881], _037209_, _037210_);
  not g_127719_(_037210_, _037211_);
  and g_127720_(out[880], _037180_, _037213_);
  not g_127721_(_037213_, _037214_);
  xor g_127722_(out[881], _037209_, _037215_);
  xor g_127723_(_001737_, _037209_, _037216_);
  and g_127724_(_037214_, _037215_, _037217_);
  or g_127725_(_037213_, _037216_, _037218_);
  and g_127726_(_037211_, _037218_, _037219_);
  or g_127727_(_037206_, _037219_, _037220_);
  or g_127728_(_037196_, _037200_, _037221_);
  and g_127729_(_037220_, _037221_, _037222_);
  or g_127730_(out[890], _014483_, _037224_);
  xor g_127731_(out[890], _014483_, _037225_);
  xor g_127732_(_001803_, _014483_, _037226_);
  or g_127733_(_037035_, _037176_, _037227_);
  not g_127734_(_037227_, _037228_);
  and g_127735_(_037042_, _037176_, _037229_);
  not g_127736_(_037229_, _037230_);
  and g_127737_(_037227_, _037230_, _037231_);
  or g_127738_(_037228_, _037229_, _037232_);
  and g_127739_(_037226_, _037232_, _037233_);
  not g_127740_(_037233_, _037235_);
  and g_127741_(_037027_, _037030_, _037236_);
  or g_127742_(_037028_, _037031_, _037237_);
  xor g_127743_(out[891], _037224_, _037238_);
  xor g_127744_(_001682_, _037224_, _037239_);
  and g_127745_(_037237_, _037238_, _037240_);
  or g_127746_(_037236_, _037239_, _037241_);
  or g_127747_(_037233_, _037240_, _037242_);
  and g_127748_(_014322_, _037175_, _037243_);
  and g_127749_(_037055_, _037176_, _037244_);
  or g_127750_(_037243_, _037244_, _037246_);
  or g_127751_(_014503_, _037246_, _037247_);
  and g_127752_(_014315_, _037175_, _037248_);
  and g_127753_(_037064_, _037176_, _037249_);
  or g_127754_(_037248_, _037249_, _037250_);
  or g_127755_(_014485_, _037250_, _037251_);
  and g_127756_(_037247_, _037251_, _037252_);
  not g_127757_(_037252_, _037253_);
  and g_127758_(_037225_, _037231_, _037254_);
  or g_127759_(_037226_, _037232_, _037255_);
  and g_127760_(_037236_, _037239_, _037257_);
  or g_127761_(_037237_, _037238_, _037258_);
  and g_127762_(_037255_, _037258_, _037259_);
  or g_127763_(_037254_, _037257_, _037260_);
  and g_127764_(_014485_, _037250_, _037261_);
  not g_127765_(_037261_, _037262_);
  and g_127766_(_014503_, _037246_, _037263_);
  not g_127767_(_037263_, _037264_);
  and g_127768_(_037262_, _037264_, _037265_);
  or g_127769_(_037261_, _037263_, _037266_);
  and g_127770_(_037235_, _037259_, _037268_);
  and g_127771_(_037241_, _037268_, _037269_);
  or g_127772_(_037242_, _037260_, _037270_);
  and g_127773_(_037252_, _037265_, _037271_);
  or g_127774_(_037253_, _037266_, _037272_);
  and g_127775_(_037269_, _037271_, _037273_);
  or g_127776_(_037270_, _037272_, _037274_);
  and g_127777_(_014340_, _037175_, _037275_);
  or g_127778_(_014339_, _037176_, _037276_);
  and g_127779_(_037099_, _037176_, _037277_);
  not g_127780_(_037277_, _037279_);
  and g_127781_(_037276_, _037279_, _037280_);
  or g_127782_(_037275_, _037277_, _037281_);
  and g_127783_(_014533_, _037281_, _037282_);
  or g_127784_(_014534_, _037280_, _037283_);
  or g_127785_(_014352_, _037176_, _037284_);
  not g_127786_(_037284_, _037285_);
  and g_127787_(_037090_, _037176_, _037286_);
  or g_127788_(_037089_, _037175_, _037287_);
  and g_127789_(_037284_, _037287_, _037288_);
  or g_127790_(_037285_, _037286_, _037290_);
  and g_127791_(_014525_, _037288_, _037291_);
  or g_127792_(_014524_, _037290_, _037292_);
  and g_127793_(_037283_, _037292_, _037293_);
  or g_127794_(_037282_, _037291_, _037294_);
  and g_127795_(_014534_, _037280_, _037295_);
  and g_127796_(_014524_, _037290_, _037296_);
  or g_127797_(_037295_, _037296_, _037297_);
  not g_127798_(_037297_, _037298_);
  and g_127799_(_037293_, _037298_, _037299_);
  or g_127800_(_037294_, _037297_, _037301_);
  and g_127801_(_014374_, _037175_, _037302_);
  and g_127802_(_037128_, _037176_, _037303_);
  or g_127803_(_037302_, _037303_, _037304_);
  and g_127804_(_014567_, _037304_, _037305_);
  not g_127805_(_037305_, _037306_);
  and g_127806_(_014367_, _037175_, _037307_);
  and g_127807_(_037119_, _037176_, _037308_);
  or g_127808_(_037307_, _037308_, _037309_);
  and g_127809_(_014556_, _037309_, _037310_);
  or g_127810_(_037305_, _037310_, _037312_);
  or g_127811_(_014567_, _037304_, _037313_);
  xor g_127812_(_014556_, _037309_, _037314_);
  and g_127813_(_037313_, _037314_, _037315_);
  and g_127814_(_037306_, _037315_, _037316_);
  and g_127815_(_037299_, _037316_, _037317_);
  not g_127816_(_037317_, _037318_);
  and g_127817_(_037273_, _037317_, _037319_);
  or g_127818_(_037274_, _037318_, _037320_);
  or g_127819_(_037222_, _037320_, _037321_);
  or g_127820_(_037293_, _037295_, _037323_);
  and g_127821_(_037312_, _037313_, _037324_);
  not g_127822_(_037324_, _037325_);
  or g_127823_(_037301_, _037325_, _037326_);
  and g_127824_(_037323_, _037326_, _037327_);
  or g_127825_(_037274_, _037327_, _037328_);
  and g_127826_(_037251_, _037266_, _037329_);
  and g_127827_(_037268_, _037329_, _037330_);
  not g_127828_(_037330_, _037331_);
  and g_127829_(_037259_, _037331_, _037332_);
  or g_127830_(_037240_, _037332_, _037334_);
  and g_127831_(_037328_, _037334_, _037335_);
  and g_127832_(_037321_, _037335_, _037336_);
  or g_127833_(out[880], _037180_, _037337_);
  and g_127834_(_037205_, _037337_, _037338_);
  and g_127835_(_037217_, _037338_, _037339_);
  and g_127836_(_037319_, _037339_, _037340_);
  or g_127837_(_037336_, _037340_, _037341_);
  and g_127838_(_037180_, _037341_, _037342_);
  not g_127839_(_037342_, _037343_);
  or g_127840_(out[880], _037341_, _037345_);
  not g_127841_(_037345_, _037346_);
  and g_127842_(_037343_, _037345_, _037347_);
  or g_127843_(_037342_, _037346_, _037348_);
  or g_127844_(_014503_, _037341_, _037349_);
  not g_127845_(_037349_, _037350_);
  and g_127846_(_037246_, _037341_, _037351_);
  or g_127847_(_037350_, _037351_, _037352_);
  not g_127848_(_037352_, _037353_);
  and g_127849_(_014713_, _037352_, _037354_);
  or g_127850_(_014712_, _037353_, _037356_);
  or g_127851_(_014485_, _037341_, _037357_);
  not g_127852_(_037357_, _037358_);
  and g_127853_(_037250_, _037341_, _037359_);
  or g_127854_(_037358_, _037359_, _037360_);
  not g_127855_(_037360_, _037361_);
  and g_127856_(_014707_, _037360_, _037362_);
  or g_127857_(_014705_, _037361_, _037363_);
  and g_127858_(_037356_, _037363_, _037364_);
  or g_127859_(_037354_, _037362_, _037365_);
  and g_127860_(_037236_, _037238_, _037367_);
  or g_127861_(_037237_, _037239_, _037368_);
  or g_127862_(out[906], _014704_, _037369_);
  xor g_127863_(out[907], _037369_, _037370_);
  xor g_127864_(_001814_, _037369_, _037371_);
  and g_127865_(_037368_, _037370_, _037372_);
  or g_127866_(_037367_, _037371_, _037373_);
  or g_127867_(_014713_, _037352_, _037374_);
  and g_127868_(_037367_, _037371_, _037375_);
  or g_127869_(_037368_, _037370_, _037376_);
  xor g_127870_(out[906], _014704_, _037378_);
  xor g_127871_(_001935_, _014704_, _037379_);
  or g_127872_(_037226_, _037341_, _037380_);
  not g_127873_(_037380_, _037381_);
  and g_127874_(_037232_, _037341_, _037382_);
  not g_127875_(_037382_, _037383_);
  and g_127876_(_037380_, _037383_, _037384_);
  or g_127877_(_037381_, _037382_, _037385_);
  and g_127878_(_037378_, _037384_, _037386_);
  or g_127879_(_037379_, _037385_, _037387_);
  and g_127880_(_037376_, _037387_, _037389_);
  or g_127881_(_037375_, _037386_, _037390_);
  and g_127882_(_037379_, _037385_, _037391_);
  not g_127883_(_037391_, _037392_);
  and g_127884_(_014705_, _037361_, _037393_);
  or g_127885_(_014707_, _037360_, _037394_);
  and g_127886_(_037392_, _037394_, _037395_);
  or g_127887_(_037391_, _037393_, _037396_);
  and g_127888_(_037389_, _037392_, _037397_);
  or g_127889_(_037372_, _037391_, _037398_);
  and g_127890_(_037373_, _037397_, _037400_);
  or g_127891_(_037390_, _037398_, _037401_);
  and g_127892_(_037374_, _037394_, _037402_);
  not g_127893_(_037402_, _037403_);
  and g_127894_(_037364_, _037402_, _037404_);
  or g_127895_(_037365_, _037403_, _037405_);
  and g_127896_(_037400_, _037404_, _037406_);
  or g_127897_(_037401_, _037405_, _037407_);
  or g_127898_(_014524_, _037341_, _037408_);
  not g_127899_(_037408_, _037409_);
  and g_127900_(_037290_, _037341_, _037411_);
  or g_127901_(_037409_, _037411_, _037412_);
  not g_127902_(_037412_, _037413_);
  or g_127903_(_014746_, _037412_, _037414_);
  not g_127904_(_037414_, _037415_);
  xor g_127905_(_014746_, _037412_, _037416_);
  xor g_127906_(_014746_, _037413_, _037417_);
  or g_127907_(_014533_, _037341_, _037418_);
  not g_127908_(_037418_, _037419_);
  and g_127909_(_037281_, _037341_, _037420_);
  not g_127910_(_037420_, _037422_);
  and g_127911_(_037418_, _037422_, _037423_);
  or g_127912_(_037419_, _037420_, _037424_);
  and g_127913_(_014735_, _037424_, _037425_);
  or g_127914_(_014736_, _037423_, _037426_);
  and g_127915_(_014736_, _037423_, _037427_);
  or g_127916_(_014735_, _037424_, _037428_);
  and g_127917_(_037426_, _037428_, _037429_);
  or g_127918_(_037425_, _037427_, _037430_);
  and g_127919_(_037416_, _037429_, _037431_);
  or g_127920_(_037417_, _037430_, _037433_);
  and g_127921_(_037304_, _037341_, _037434_);
  not g_127922_(_037434_, _037435_);
  or g_127923_(_014567_, _037341_, _037436_);
  not g_127924_(_037436_, _037437_);
  and g_127925_(_037435_, _037436_, _037438_);
  or g_127926_(_037434_, _037437_, _037439_);
  and g_127927_(_014774_, _037439_, _037440_);
  or g_127928_(_014773_, _037438_, _037441_);
  or g_127929_(_014556_, _037341_, _037442_);
  not g_127930_(_037442_, _037444_);
  and g_127931_(_037309_, _037341_, _037445_);
  not g_127932_(_037445_, _037446_);
  and g_127933_(_037442_, _037446_, _037447_);
  or g_127934_(_037444_, _037445_, _037448_);
  and g_127935_(_014766_, _037448_, _037449_);
  or g_127936_(_014765_, _037447_, _037450_);
  and g_127937_(_037441_, _037450_, _037451_);
  or g_127938_(_037440_, _037449_, _037452_);
  and g_127939_(_014765_, _037447_, _037453_);
  or g_127940_(_014766_, _037448_, _037455_);
  and g_127941_(_014773_, _037438_, _037456_);
  or g_127942_(_014774_, _037439_, _037457_);
  and g_127943_(_037455_, _037457_, _037458_);
  or g_127944_(_037453_, _037456_, _037459_);
  and g_127945_(_037451_, _037458_, _037460_);
  or g_127946_(_037452_, _037459_, _037461_);
  and g_127947_(_037431_, _037460_, _037462_);
  or g_127948_(_037433_, _037461_, _037463_);
  and g_127949_(_037406_, _037462_, _037464_);
  or g_127950_(_037407_, _037463_, _037466_);
  or g_127951_(_014615_, _037341_, _037467_);
  not g_127952_(_037467_, _037468_);
  and g_127953_(_037193_, _037341_, _037469_);
  or g_127954_(_037468_, _037469_, _037470_);
  and g_127955_(_014798_, _037470_, _037471_);
  and g_127956_(_037184_, _037341_, _037472_);
  or g_127957_(_002077_, _037341_, _037473_);
  not g_127958_(_037473_, _037474_);
  or g_127959_(_037472_, _037474_, _037475_);
  or g_127960_(_014798_, _037470_, _037477_);
  or g_127961_(_002334_, _037475_, _037478_);
  not g_127962_(_037478_, _037479_);
  xor g_127963_(_014798_, _037470_, _037480_);
  xor g_127964_(_014799_, _037470_, _037481_);
  xor g_127965_(_002334_, _037475_, _037482_);
  xor g_127966_(_002333_, _037475_, _037483_);
  and g_127967_(_037480_, _037482_, _037484_);
  or g_127968_(_037481_, _037483_, _037485_);
  and g_127969_(_037209_, _037341_, _037486_);
  or g_127970_(out[881], _037341_, _037488_);
  not g_127971_(_037488_, _037489_);
  or g_127972_(_037486_, _037489_, _037490_);
  and g_127973_(out[897], _037490_, _037491_);
  not g_127974_(_037491_, _037492_);
  and g_127975_(out[896], _037348_, _037493_);
  or g_127976_(_001880_, _037347_, _037494_);
  xor g_127977_(out[897], _037490_, _037495_);
  xor g_127978_(_001869_, _037490_, _037496_);
  and g_127979_(_037494_, _037495_, _037497_);
  or g_127980_(_037493_, _037496_, _037499_);
  and g_127981_(_037492_, _037499_, _037500_);
  or g_127982_(_037491_, _037497_, _037501_);
  and g_127983_(_037484_, _037501_, _037502_);
  or g_127984_(_037485_, _037500_, _037503_);
  or g_127985_(_037471_, _037479_, _037504_);
  and g_127986_(_037477_, _037504_, _037505_);
  not g_127987_(_037505_, _037506_);
  and g_127988_(_037503_, _037506_, _037507_);
  or g_127989_(_037502_, _037505_, _037508_);
  and g_127990_(_037464_, _037508_, _037510_);
  or g_127991_(_037466_, _037507_, _037511_);
  and g_127992_(_037452_, _037457_, _037512_);
  or g_127993_(_037451_, _037456_, _037513_);
  and g_127994_(_037431_, _037512_, _037514_);
  or g_127995_(_037433_, _037513_, _037515_);
  and g_127996_(_037415_, _037428_, _037516_);
  or g_127997_(_037414_, _037427_, _037517_);
  and g_127998_(_037426_, _037517_, _037518_);
  or g_127999_(_037425_, _037516_, _037519_);
  and g_128000_(_037515_, _037518_, _037521_);
  or g_128001_(_037514_, _037519_, _037522_);
  and g_128002_(_037406_, _037522_, _037523_);
  or g_128003_(_037407_, _037521_, _037524_);
  and g_128004_(_037365_, _037395_, _037525_);
  or g_128005_(_037364_, _037396_, _037526_);
  and g_128006_(_037389_, _037526_, _037527_);
  or g_128007_(_037390_, _037525_, _037528_);
  and g_128008_(_037373_, _037528_, _037529_);
  or g_128009_(_037372_, _037527_, _037530_);
  and g_128010_(_037524_, _037530_, _037532_);
  or g_128011_(_037523_, _037529_, _037533_);
  and g_128012_(_037511_, _037532_, _037534_);
  or g_128013_(_037510_, _037533_, _037535_);
  or g_128014_(out[896], _037348_, _037536_);
  and g_128015_(_037484_, _037536_, _037537_);
  not g_128016_(_037537_, _037538_);
  and g_128017_(_037497_, _037537_, _037539_);
  or g_128018_(_037499_, _037538_, _037540_);
  and g_128019_(_037464_, _037539_, _037541_);
  or g_128020_(_037466_, _037540_, _037543_);
  and g_128021_(_037535_, _037543_, _037544_);
  or g_128022_(_037534_, _037541_, _037545_);
  and g_128023_(_037348_, _037545_, _037546_);
  and g_128024_(_001880_, _037544_, _037547_);
  or g_128025_(_037546_, _037547_, _037548_);
  and g_128026_(_037367_, _037370_, _037549_);
  or g_128027_(_037368_, _037371_, _037550_);
  or g_128028_(out[922], _014962_, _037551_);
  xor g_128029_(out[923], _037551_, _037552_);
  xor g_128030_(_001946_, _037551_, _037554_);
  and g_128031_(_037550_, _037552_, _037555_);
  or g_128032_(_037549_, _037554_, _037556_);
  xor g_128033_(_002067_, _014962_, _037557_);
  and g_128034_(_037378_, _037544_, _037558_);
  and g_128035_(_037385_, _037545_, _037559_);
  or g_128036_(_037558_, _037559_, _037560_);
  or g_128037_(_037557_, _037560_, _037561_);
  not g_128038_(_037561_, _037562_);
  and g_128039_(_037549_, _037554_, _037563_);
  or g_128040_(_037550_, _037552_, _037565_);
  and g_128041_(_037561_, _037565_, _037566_);
  or g_128042_(_037562_, _037563_, _037567_);
  and g_128043_(_037556_, _037567_, _037568_);
  or g_128044_(_037555_, _037566_, _037569_);
  and g_128045_(_014705_, _037544_, _037570_);
  and g_128046_(_037360_, _037545_, _037571_);
  or g_128047_(_037570_, _037571_, _037572_);
  not g_128048_(_037572_, _037573_);
  and g_128049_(_014964_, _037572_, _037574_);
  or g_128050_(_014963_, _037573_, _037576_);
  and g_128051_(_014712_, _037544_, _037577_);
  and g_128052_(_037352_, _037545_, _037578_);
  or g_128053_(_037577_, _037578_, _037579_);
  not g_128054_(_037579_, _037580_);
  and g_128055_(_014972_, _037579_, _037581_);
  or g_128056_(_014971_, _037580_, _037582_);
  and g_128057_(_037576_, _037582_, _037583_);
  or g_128058_(_037574_, _037581_, _037584_);
  and g_128059_(_014971_, _037580_, _037585_);
  or g_128060_(_014972_, _037579_, _037587_);
  and g_128061_(_014963_, _037573_, _037588_);
  or g_128062_(_014964_, _037572_, _037589_);
  and g_128063_(_037587_, _037589_, _037590_);
  or g_128064_(_037585_, _037588_, _037591_);
  and g_128065_(_037583_, _037590_, _037592_);
  or g_128066_(_037584_, _037591_, _037593_);
  or g_128067_(_001869_, _037545_, _037594_);
  or g_128068_(_037490_, _037544_, _037595_);
  and g_128069_(_037594_, _037595_, _037596_);
  not g_128070_(_037596_, _037598_);
  and g_128071_(out[913], _037596_, _037599_);
  and g_128072_(out[912], _037548_, _037600_);
  not g_128073_(_037600_, _037601_);
  xor g_128074_(out[913], _037596_, _037602_);
  xor g_128075_(_002001_, _037596_, _037603_);
  and g_128076_(_037601_, _037602_, _037604_);
  or g_128077_(_037600_, _037603_, _037605_);
  or g_128078_(_037599_, _037604_, _037606_);
  and g_128079_(_014736_, _037544_, _037607_);
  or g_128080_(_014735_, _037545_, _037609_);
  and g_128081_(_037424_, _037545_, _037610_);
  or g_128082_(_037423_, _037544_, _037611_);
  and g_128083_(_037609_, _037611_, _037612_);
  or g_128084_(_037607_, _037610_, _037613_);
  and g_128085_(_014991_, _037613_, _037614_);
  or g_128086_(_014991_, _037613_, _037615_);
  xor g_128087_(_014993_, _037612_, _037616_);
  xor g_128088_(_014991_, _037612_, _037617_);
  or g_128089_(_014746_, _037545_, _037618_);
  not g_128090_(_037618_, _037620_);
  and g_128091_(_037412_, _037545_, _037621_);
  or g_128092_(_037620_, _037621_, _037622_);
  or g_128093_(_015002_, _037622_, _037623_);
  not g_128094_(_037623_, _037624_);
  xor g_128095_(_015002_, _037622_, _037625_);
  xor g_128096_(_015004_, _037622_, _037626_);
  and g_128097_(_037616_, _037625_, _037627_);
  or g_128098_(_037617_, _037626_, _037628_);
  and g_128099_(_014765_, _037544_, _037629_);
  or g_128100_(_014766_, _037545_, _037631_);
  and g_128101_(_037448_, _037545_, _037632_);
  or g_128102_(_037447_, _037544_, _037633_);
  and g_128103_(_037631_, _037633_, _037634_);
  or g_128104_(_037629_, _037632_, _037635_);
  and g_128105_(_015041_, _037635_, _037636_);
  or g_128106_(_015040_, _037634_, _037637_);
  and g_128107_(_014773_, _037544_, _037638_);
  or g_128108_(_014774_, _037545_, _037639_);
  and g_128109_(_037439_, _037545_, _037640_);
  or g_128110_(_037438_, _037544_, _037642_);
  and g_128111_(_037639_, _037642_, _037643_);
  or g_128112_(_037638_, _037640_, _037644_);
  and g_128113_(_015019_, _037644_, _037645_);
  or g_128114_(_015018_, _037643_, _037646_);
  and g_128115_(_037637_, _037646_, _037647_);
  or g_128116_(_037636_, _037645_, _037648_);
  and g_128117_(_015040_, _037634_, _037649_);
  or g_128118_(_015041_, _037635_, _037650_);
  and g_128119_(_015018_, _037643_, _037651_);
  or g_128120_(_015019_, _037644_, _037653_);
  and g_128121_(_037650_, _037653_, _037654_);
  or g_128122_(_037649_, _037651_, _037655_);
  and g_128123_(_037647_, _037654_, _037656_);
  or g_128124_(_037648_, _037655_, _037657_);
  and g_128125_(_037627_, _037656_, _037658_);
  or g_128126_(_037628_, _037657_, _037659_);
  and g_128127_(_037470_, _037545_, _037660_);
  not g_128128_(_037660_, _037661_);
  or g_128129_(_014798_, _037545_, _037662_);
  not g_128130_(_037662_, _037664_);
  and g_128131_(_037661_, _037662_, _037665_);
  or g_128132_(_037660_, _037664_, _037666_);
  and g_128133_(_014899_, _037666_, _037667_);
  or g_128134_(_014900_, _037665_, _037668_);
  or g_128135_(_014899_, _037666_, _037669_);
  not g_128136_(_037669_, _037670_);
  or g_128137_(_002334_, _037545_, _037671_);
  not g_128138_(_037671_, _037672_);
  and g_128139_(_037475_, _037545_, _037673_);
  not g_128140_(_037673_, _037675_);
  and g_128141_(_037671_, _037675_, _037676_);
  or g_128142_(_037672_, _037673_, _037677_);
  and g_128143_(_002530_, _037676_, _037678_);
  or g_128144_(_002531_, _037677_, _037679_);
  xor g_128145_(_002530_, _037676_, _037680_);
  and g_128146_(_037669_, _037680_, _037681_);
  and g_128147_(_037668_, _037681_, _037682_);
  and g_128148_(_037658_, _037682_, _037683_);
  and g_128149_(_037606_, _037683_, _037684_);
  not g_128150_(_037684_, _037686_);
  and g_128151_(_037668_, _037679_, _037687_);
  or g_128152_(_037667_, _037678_, _037688_);
  and g_128153_(_037669_, _037688_, _037689_);
  or g_128154_(_037670_, _037687_, _037690_);
  and g_128155_(_037658_, _037689_, _037691_);
  or g_128156_(_037659_, _037690_, _037692_);
  and g_128157_(_037627_, _037648_, _037693_);
  and g_128158_(_037653_, _037693_, _037694_);
  and g_128159_(_037615_, _037624_, _037695_);
  or g_128160_(_037614_, _037695_, _037697_);
  or g_128161_(_037694_, _037697_, _037698_);
  not g_128162_(_037698_, _037699_);
  and g_128163_(_037692_, _037699_, _037700_);
  or g_128164_(_037691_, _037698_, _037701_);
  and g_128165_(_037686_, _037700_, _037702_);
  or g_128166_(_037684_, _037701_, _037703_);
  and g_128167_(_037592_, _037703_, _037704_);
  or g_128168_(_037593_, _037702_, _037705_);
  and g_128169_(_037584_, _037589_, _037706_);
  or g_128170_(_037583_, _037588_, _037708_);
  and g_128171_(_037705_, _037708_, _037709_);
  or g_128172_(_037704_, _037706_, _037710_);
  and g_128173_(_037557_, _037560_, _037711_);
  not g_128174_(_037711_, _037712_);
  and g_128175_(_037556_, _037712_, _037713_);
  or g_128176_(_037555_, _037711_, _037714_);
  and g_128177_(_037710_, _037713_, _037715_);
  or g_128178_(_037709_, _037714_, _037716_);
  and g_128179_(_037569_, _037716_, _037717_);
  or g_128180_(_037568_, _037715_, _037719_);
  or g_128181_(out[912], _037548_, _037720_);
  and g_128182_(_037566_, _037720_, _037721_);
  and g_128183_(_037713_, _037721_, _037722_);
  and g_128184_(_037592_, _037722_, _037723_);
  and g_128185_(_037683_, _037723_, _037724_);
  not g_128186_(_037724_, _037725_);
  and g_128187_(_037604_, _037724_, _037726_);
  or g_128188_(_037605_, _037725_, _037727_);
  and g_128189_(_037719_, _037727_, _037728_);
  or g_128190_(_037717_, _037726_, _037730_);
  and g_128191_(_037548_, _037730_, _037731_);
  not g_128192_(_037731_, _037732_);
  or g_128193_(out[912], _037730_, _037733_);
  and g_128194_(_037732_, _037733_, _037734_);
  not g_128195_(_037734_, _037735_);
  and g_128196_(_014900_, _037728_, _037736_);
  and g_128197_(_037666_, _037730_, _037737_);
  or g_128198_(_037736_, _037737_, _037738_);
  and g_128199_(_015196_, _037738_, _037739_);
  and g_128200_(_037677_, _037730_, _037741_);
  not g_128201_(_037741_, _037742_);
  or g_128202_(_002531_, _037730_, _037743_);
  not g_128203_(_037743_, _037744_);
  and g_128204_(_037742_, _037743_, _037745_);
  or g_128205_(_037741_, _037744_, _037746_);
  or g_128206_(_015196_, _037738_, _037747_);
  and g_128207_(_002720_, _037745_, _037748_);
  xor g_128208_(_015196_, _037738_, _037749_);
  xor g_128209_(_002720_, _037745_, _037750_);
  and g_128210_(_037749_, _037750_, _037752_);
  or g_128211_(_002001_, _037730_, _037753_);
  not g_128212_(_037753_, _037754_);
  and g_128213_(_037598_, _037730_, _037755_);
  or g_128214_(_037596_, _037728_, _037756_);
  and g_128215_(_037753_, _037756_, _037757_);
  or g_128216_(_037754_, _037755_, _037758_);
  and g_128217_(out[929], _037757_, _037759_);
  or g_128218_(_002122_, _037734_, _037760_);
  xor g_128219_(out[929], _037757_, _037761_);
  and g_128220_(_037760_, _037761_, _037763_);
  or g_128221_(_037759_, _037763_, _037764_);
  and g_128222_(_037752_, _037764_, _037765_);
  or g_128223_(_037739_, _037748_, _037766_);
  and g_128224_(_037747_, _037766_, _037767_);
  or g_128225_(_037765_, _037767_, _037768_);
  not g_128226_(_037768_, _037769_);
  or g_128227_(out[938], _015118_, _037770_);
  xor g_128228_(_002177_, _015118_, _037771_);
  and g_128229_(_037560_, _037730_, _037772_);
  or g_128230_(_037557_, _037730_, _037774_);
  not g_128231_(_037774_, _037775_);
  or g_128232_(_037772_, _037775_, _037776_);
  or g_128233_(_037771_, _037776_, _037777_);
  not g_128234_(_037777_, _037778_);
  and g_128235_(_037549_, _037552_, _037779_);
  not g_128236_(_037779_, _037780_);
  xor g_128237_(out[939], _037770_, _037781_);
  not g_128238_(_037781_, _037782_);
  and g_128239_(_037779_, _037782_, _037783_);
  or g_128240_(_037780_, _037781_, _037785_);
  and g_128241_(_037777_, _037785_, _037786_);
  or g_128242_(_037778_, _037783_, _037787_);
  and g_128243_(_037771_, _037776_, _037788_);
  not g_128244_(_037788_, _037789_);
  and g_128245_(_037780_, _037781_, _037790_);
  or g_128246_(_037779_, _037782_, _037791_);
  and g_128247_(_037789_, _037791_, _037792_);
  or g_128248_(_037788_, _037790_, _037793_);
  and g_128249_(_037786_, _037792_, _037794_);
  or g_128250_(_037787_, _037793_, _037796_);
  or g_128251_(_014964_, _037730_, _037797_);
  not g_128252_(_037797_, _037798_);
  and g_128253_(_037572_, _037730_, _037799_);
  not g_128254_(_037799_, _037800_);
  and g_128255_(_037797_, _037800_, _037801_);
  or g_128256_(_037798_, _037799_, _037802_);
  and g_128257_(_015120_, _037802_, _037803_);
  or g_128258_(_015119_, _037801_, _037804_);
  or g_128259_(_014972_, _037730_, _037805_);
  not g_128260_(_037805_, _037807_);
  and g_128261_(_037579_, _037730_, _037808_);
  not g_128262_(_037808_, _037809_);
  and g_128263_(_037805_, _037809_, _037810_);
  or g_128264_(_037807_, _037808_, _037811_);
  and g_128265_(_015129_, _037811_, _037812_);
  or g_128266_(_015128_, _037810_, _037813_);
  and g_128267_(_037804_, _037813_, _037814_);
  or g_128268_(_037803_, _037812_, _037815_);
  and g_128269_(_015128_, _037810_, _037816_);
  not g_128270_(_037816_, _037818_);
  or g_128271_(_015120_, _037802_, _037819_);
  not g_128272_(_037819_, _037820_);
  and g_128273_(_037814_, _037819_, _037821_);
  or g_128274_(_037815_, _037820_, _037822_);
  and g_128275_(_037818_, _037821_, _037823_);
  or g_128276_(_037816_, _037822_, _037824_);
  and g_128277_(_037794_, _037823_, _037825_);
  or g_128278_(_037796_, _037824_, _037826_);
  or g_128279_(_015002_, _037730_, _037827_);
  not g_128280_(_037827_, _037829_);
  and g_128281_(_037622_, _037730_, _037830_);
  not g_128282_(_037830_, _037831_);
  and g_128283_(_037827_, _037831_, _037832_);
  or g_128284_(_037829_, _037830_, _037833_);
  and g_128285_(_015156_, _037832_, _037834_);
  or g_128286_(_015155_, _037833_, _037835_);
  xor g_128287_(_015156_, _037832_, _037836_);
  xor g_128288_(_015155_, _037832_, _037837_);
  and g_128289_(_014993_, _037728_, _037838_);
  or g_128290_(_014991_, _037730_, _037840_);
  and g_128291_(_037613_, _037730_, _037841_);
  or g_128292_(_037612_, _037728_, _037842_);
  and g_128293_(_037840_, _037842_, _037843_);
  or g_128294_(_037838_, _037841_, _037844_);
  and g_128295_(_015149_, _037844_, _037845_);
  or g_128296_(_015150_, _037843_, _037846_);
  and g_128297_(_015150_, _037843_, _037847_);
  or g_128298_(_015149_, _037844_, _037848_);
  and g_128299_(_037846_, _037848_, _037849_);
  or g_128300_(_037845_, _037847_, _037851_);
  and g_128301_(_037836_, _037849_, _037852_);
  or g_128302_(_037837_, _037851_, _037853_);
  or g_128303_(_015041_, _037730_, _037854_);
  not g_128304_(_037854_, _037855_);
  and g_128305_(_037635_, _037730_, _037856_);
  not g_128306_(_037856_, _037857_);
  and g_128307_(_037854_, _037857_, _037858_);
  or g_128308_(_037855_, _037856_, _037859_);
  and g_128309_(_015173_, _037859_, _037860_);
  or g_128310_(_015172_, _037858_, _037862_);
  or g_128311_(_015019_, _037730_, _037863_);
  not g_128312_(_037863_, _037864_);
  and g_128313_(_037644_, _037730_, _037865_);
  not g_128314_(_037865_, _037866_);
  and g_128315_(_037863_, _037866_, _037867_);
  or g_128316_(_037864_, _037865_, _037868_);
  and g_128317_(_015180_, _037868_, _037869_);
  or g_128318_(_015178_, _037867_, _037870_);
  and g_128319_(_037862_, _037870_, _037871_);
  or g_128320_(_037860_, _037869_, _037873_);
  or g_128321_(_015180_, _037868_, _037874_);
  not g_128322_(_037874_, _037875_);
  or g_128323_(_015173_, _037859_, _037876_);
  not g_128324_(_037876_, _037877_);
  or g_128325_(_037873_, _037877_, _037878_);
  not g_128326_(_037878_, _037879_);
  and g_128327_(_037874_, _037879_, _037880_);
  or g_128328_(_037875_, _037878_, _037881_);
  or g_128329_(_037853_, _037881_, _037882_);
  and g_128330_(_037825_, _037880_, _037884_);
  and g_128331_(_037852_, _037884_, _037885_);
  or g_128332_(_037826_, _037882_, _037886_);
  and g_128333_(_037768_, _037885_, _037887_);
  or g_128334_(_037769_, _037886_, _037888_);
  and g_128335_(_037852_, _037873_, _037889_);
  or g_128336_(_037853_, _037871_, _037890_);
  and g_128337_(_037874_, _037889_, _037891_);
  or g_128338_(_037875_, _037890_, _037892_);
  and g_128339_(_037834_, _037848_, _037893_);
  or g_128340_(_037835_, _037847_, _037895_);
  and g_128341_(_037846_, _037895_, _037896_);
  or g_128342_(_037845_, _037893_, _037897_);
  and g_128343_(_037892_, _037896_, _037898_);
  or g_128344_(_037891_, _037897_, _037899_);
  and g_128345_(_037825_, _037899_, _037900_);
  or g_128346_(_037826_, _037898_, _037901_);
  and g_128347_(_037815_, _037819_, _037902_);
  or g_128348_(_037814_, _037820_, _037903_);
  and g_128349_(_037794_, _037902_, _037904_);
  or g_128350_(_037796_, _037903_, _037906_);
  and g_128351_(_037787_, _037791_, _037907_);
  or g_128352_(_037786_, _037790_, _037908_);
  and g_128353_(_037906_, _037908_, _037909_);
  or g_128354_(_037904_, _037907_, _037910_);
  and g_128355_(_037901_, _037909_, _037911_);
  or g_128356_(_037900_, _037910_, _037912_);
  and g_128357_(_037888_, _037911_, _037913_);
  or g_128358_(_037887_, _037912_, _037914_);
  and g_128359_(_002122_, _037734_, _037915_);
  or g_128360_(out[928], _037735_, _037917_);
  and g_128361_(_037752_, _037763_, _037918_);
  not g_128362_(_037918_, _037919_);
  and g_128363_(_037885_, _037918_, _037920_);
  or g_128364_(_037886_, _037919_, _037921_);
  and g_128365_(_037917_, _037920_, _037922_);
  or g_128366_(_037915_, _037921_, _037923_);
  and g_128367_(_037914_, _037923_, _037924_);
  or g_128368_(_037913_, _037922_, _037925_);
  or g_128369_(_037734_, _037924_, _037926_);
  or g_128370_(out[928], _037925_, _037928_);
  and g_128371_(_037926_, _037928_, _037929_);
  not g_128372_(_037929_, _037930_);
  and g_128373_(_037779_, _037781_, _037931_);
  not g_128374_(_037931_, _037932_);
  or g_128375_(out[954], _015303_, _037933_);
  xor g_128376_(out[955], _037933_, _037934_);
  not g_128377_(_037934_, _037935_);
  and g_128378_(_037932_, _037934_, _037936_);
  or g_128379_(_037931_, _037935_, _037937_);
  or g_128380_(_015128_, _037925_, _037939_);
  not g_128381_(_037939_, _037940_);
  and g_128382_(_037810_, _037925_, _037941_);
  not g_128383_(_037941_, _037942_);
  and g_128384_(_037939_, _037942_, _037943_);
  or g_128385_(_037940_, _037941_, _037944_);
  and g_128386_(_015296_, _037944_, _037945_);
  or g_128387_(_015297_, _037943_, _037946_);
  xor g_128388_(out[954], _015303_, _037947_);
  not g_128389_(_037947_, _037948_);
  or g_128390_(_037771_, _037925_, _037950_);
  not g_128391_(_037950_, _037951_);
  and g_128392_(_037776_, _037925_, _037952_);
  or g_128393_(_037951_, _037952_, _037953_);
  not g_128394_(_037953_, _037954_);
  and g_128395_(_037948_, _037953_, _037955_);
  or g_128396_(_037947_, _037954_, _037956_);
  and g_128397_(_015119_, _037924_, _037957_);
  and g_128398_(_037802_, _037925_, _037958_);
  or g_128399_(_037957_, _037958_, _037959_);
  not g_128400_(_037959_, _037961_);
  and g_128401_(_015304_, _037961_, _037962_);
  or g_128402_(_015305_, _037959_, _037963_);
  and g_128403_(_037931_, _037935_, _037964_);
  or g_128404_(_037932_, _037934_, _037965_);
  and g_128405_(_037947_, _037954_, _037966_);
  or g_128406_(_037948_, _037953_, _037967_);
  and g_128407_(_037965_, _037967_, _037968_);
  or g_128408_(_037964_, _037966_, _037969_);
  and g_128409_(_015305_, _037959_, _037970_);
  or g_128410_(_015304_, _037961_, _037972_);
  and g_128411_(_015297_, _037943_, _037973_);
  or g_128412_(_015296_, _037944_, _037974_);
  and g_128413_(_037972_, _037974_, _037975_);
  or g_128414_(_037970_, _037973_, _037976_);
  and g_128415_(_037937_, _037956_, _037977_);
  or g_128416_(_037936_, _037955_, _037978_);
  and g_128417_(_037968_, _037977_, _037979_);
  or g_128418_(_037969_, _037978_, _037980_);
  and g_128419_(_037946_, _037972_, _037981_);
  or g_128420_(_037945_, _037970_, _037983_);
  and g_128421_(_037963_, _037974_, _037984_);
  or g_128422_(_037962_, _037973_, _037985_);
  and g_128423_(_037981_, _037984_, _037986_);
  or g_128424_(_037983_, _037985_, _037987_);
  and g_128425_(_037979_, _037986_, _037988_);
  or g_128426_(_037980_, _037987_, _037989_);
  and g_128427_(_015156_, _037924_, _037990_);
  or g_128428_(_015155_, _037925_, _037991_);
  and g_128429_(_037833_, _037925_, _037992_);
  or g_128430_(_037832_, _037924_, _037994_);
  and g_128431_(_037991_, _037994_, _037995_);
  or g_128432_(_037990_, _037992_, _037996_);
  and g_128433_(_015320_, _037995_, _037997_);
  or g_128434_(_015319_, _037996_, _037998_);
  and g_128435_(_015150_, _037924_, _037999_);
  or g_128436_(_015149_, _037925_, _038000_);
  and g_128437_(_037844_, _037925_, _038001_);
  or g_128438_(_037843_, _037924_, _038002_);
  and g_128439_(_038000_, _038002_, _038003_);
  or g_128440_(_037999_, _038001_, _038005_);
  and g_128441_(_009389_, _038005_, _038006_);
  or g_128442_(_009390_, _038003_, _038007_);
  and g_128443_(_037998_, _038007_, _038008_);
  or g_128444_(_037997_, _038006_, _038009_);
  or g_128445_(_015320_, _037995_, _038010_);
  not g_128446_(_038010_, _038011_);
  and g_128447_(_009390_, _038003_, _038012_);
  not g_128448_(_038012_, _038013_);
  and g_128449_(_038008_, _038013_, _038014_);
  or g_128450_(_038009_, _038012_, _038016_);
  and g_128451_(_038010_, _038014_, _038017_);
  or g_128452_(_038011_, _038016_, _038018_);
  or g_128453_(_015172_, _037925_, _038019_);
  or g_128454_(_037859_, _037924_, _038020_);
  and g_128455_(_038019_, _038020_, _038021_);
  not g_128456_(_038021_, _038022_);
  and g_128457_(_015337_, _038022_, _038023_);
  or g_128458_(_015338_, _038021_, _038024_);
  or g_128459_(_015180_, _037925_, _038025_);
  not g_128460_(_038025_, _038027_);
  and g_128461_(_037868_, _037925_, _038028_);
  not g_128462_(_038028_, _038029_);
  and g_128463_(_038025_, _038029_, _038030_);
  or g_128464_(_038027_, _038028_, _038031_);
  and g_128465_(_015346_, _038031_, _038032_);
  or g_128466_(_015345_, _038030_, _038033_);
  and g_128467_(_038024_, _038033_, _038034_);
  or g_128468_(_038023_, _038032_, _038035_);
  and g_128469_(_015338_, _038021_, _038036_);
  or g_128470_(_015337_, _038022_, _038038_);
  and g_128471_(_015345_, _038030_, _038039_);
  or g_128472_(_015346_, _038031_, _038040_);
  and g_128473_(_038038_, _038040_, _038041_);
  or g_128474_(_038036_, _038039_, _038042_);
  and g_128475_(_038034_, _038041_, _038043_);
  or g_128476_(_038035_, _038042_, _038044_);
  and g_128477_(_038017_, _038043_, _038045_);
  or g_128478_(_038018_, _038044_, _038046_);
  and g_128479_(_037988_, _038045_, _038047_);
  or g_128480_(_037989_, _038046_, _038049_);
  or g_128481_(_015196_, _037925_, _038050_);
  and g_128482_(_037738_, _037925_, _038051_);
  not g_128483_(_038051_, _038052_);
  and g_128484_(_038050_, _038052_, _038053_);
  or g_128485_(_015361_, _038053_, _038054_);
  and g_128486_(_002720_, _037924_, _038055_);
  and g_128487_(_037746_, _037925_, _038056_);
  or g_128488_(_038055_, _038056_, _038057_);
  or g_128489_(_002906_, _038057_, _038058_);
  and g_128490_(_038054_, _038058_, _038060_);
  and g_128491_(_015361_, _038053_, _038061_);
  not g_128492_(_038061_, _038062_);
  xor g_128493_(_002906_, _038057_, _038063_);
  xor g_128494_(_002905_, _038057_, _038064_);
  and g_128495_(_038054_, _038063_, _038065_);
  xor g_128496_(_015360_, _038053_, _038066_);
  and g_128497_(_038062_, _038065_, _038067_);
  or g_128498_(_038064_, _038066_, _038068_);
  and g_128499_(out[929], _037924_, _038069_);
  and g_128500_(_037758_, _037925_, _038071_);
  or g_128501_(_038069_, _038071_, _038072_);
  or g_128502_(_054336_, _038072_, _038073_);
  and g_128503_(out[944], _037930_, _038074_);
  or g_128504_(_002232_, _037929_, _038075_);
  xor g_128505_(_054336_, _038072_, _038076_);
  xor g_128506_(out[945], _038072_, _038077_);
  and g_128507_(_038075_, _038076_, _038078_);
  or g_128508_(_038074_, _038077_, _038079_);
  and g_128509_(_038073_, _038079_, _038080_);
  not g_128510_(_038080_, _038082_);
  and g_128511_(_038067_, _038082_, _038083_);
  or g_128512_(_038068_, _038080_, _038084_);
  or g_128513_(_038060_, _038061_, _038085_);
  not g_128514_(_038085_, _038086_);
  and g_128515_(_038084_, _038085_, _038087_);
  or g_128516_(_038083_, _038086_, _038088_);
  and g_128517_(_038047_, _038088_, _038089_);
  or g_128518_(_038049_, _038087_, _038090_);
  or g_128519_(_038008_, _038012_, _038091_);
  not g_128520_(_038091_, _038093_);
  and g_128521_(_038033_, _038038_, _038094_);
  or g_128522_(_038032_, _038036_, _038095_);
  and g_128523_(_038040_, _038095_, _038096_);
  or g_128524_(_038039_, _038094_, _038097_);
  and g_128525_(_038017_, _038096_, _038098_);
  or g_128526_(_038018_, _038097_, _038099_);
  and g_128527_(_038091_, _038099_, _038100_);
  or g_128528_(_038093_, _038098_, _038101_);
  and g_128529_(_037988_, _038101_, _038102_);
  or g_128530_(_037989_, _038100_, _038104_);
  and g_128531_(_037963_, _037976_, _038105_);
  or g_128532_(_037962_, _037975_, _038106_);
  and g_128533_(_037979_, _038105_, _038107_);
  or g_128534_(_037980_, _038106_, _038108_);
  and g_128535_(_037937_, _037969_, _038109_);
  or g_128536_(_037936_, _037968_, _038110_);
  and g_128537_(_038108_, _038110_, _038111_);
  or g_128538_(_038107_, _038109_, _038112_);
  and g_128539_(_038104_, _038111_, _038113_);
  or g_128540_(_038102_, _038112_, _038115_);
  and g_128541_(_038090_, _038113_, _038116_);
  or g_128542_(_038089_, _038115_, _038117_);
  or g_128543_(out[944], _037930_, _038118_);
  and g_128544_(_038067_, _038078_, _038119_);
  and g_128545_(_038118_, _038119_, _038120_);
  and g_128546_(_038047_, _038120_, _038121_);
  not g_128547_(_038121_, _038122_);
  and g_128548_(_038117_, _038122_, _038123_);
  or g_128549_(_038116_, _038121_, _038124_);
  or g_128550_(_037929_, _038123_, _038126_);
  or g_128551_(out[944], _038124_, _038127_);
  and g_128552_(_038126_, _038127_, _038128_);
  xor g_128553_(_032766_, _038128_, _038129_);
  or g_128554_(_009233_, _032763_, _038130_);
  or g_128555_(_032654_, _032762_, _038131_);
  and g_128556_(_038130_, _038131_, _038132_);
  or g_128557_(_037995_, _038123_, _038133_);
  or g_128558_(_015319_, _038124_, _038134_);
  and g_128559_(_038133_, _038134_, _038135_);
  xor g_128560_(_038132_, _038135_, _038137_);
  and g_128561_(_009205_, _032762_, _038138_);
  not g_128562_(_038138_, _038139_);
  and g_128563_(_032608_, _032763_, _038140_);
  or g_128564_(_032607_, _032762_, _038141_);
  and g_128565_(_038139_, _038141_, _038142_);
  or g_128566_(_038138_, _038140_, _038143_);
  and g_128567_(_015297_, _038123_, _038144_);
  or g_128568_(_015296_, _038124_, _038145_);
  or g_128569_(_037943_, _038123_, _038146_);
  not g_128570_(_038146_, _038148_);
  and g_128571_(_038145_, _038146_, _038149_);
  or g_128572_(_038144_, _038148_, _038150_);
  and g_128573_(_038142_, _038150_, _038151_);
  and g_128574_(_032628_, _032630_, _038152_);
  and g_128575_(_037931_, _037934_, _038153_);
  xor g_128576_(_038152_, _038153_, _038154_);
  or g_128577_(_038151_, _038154_, _038155_);
  or g_128578_(_003129_, _032763_, _038156_);
  or g_128579_(_032661_, _032762_, _038157_);
  and g_128580_(_038156_, _038157_, _038159_);
  and g_128581_(_009389_, _038123_, _038160_);
  and g_128582_(_038003_, _038124_, _038161_);
  or g_128583_(_038160_, _038161_, _038162_);
  xor g_128584_(_038159_, _038162_, _038163_);
  and g_128585_(_009255_, _032762_, _038164_);
  and g_128586_(_032682_, _032763_, _038165_);
  or g_128587_(_038164_, _038165_, _038166_);
  or g_128588_(_015338_, _038124_, _038167_);
  or g_128589_(_038022_, _038123_, _038168_);
  and g_128590_(_038167_, _038168_, _038170_);
  and g_128591_(out[465], _032762_, _038171_);
  and g_128592_(_032715_, _032763_, _038172_);
  or g_128593_(_038171_, _038172_, _038173_);
  and g_128594_(out[945], _038123_, _038174_);
  and g_128595_(_038072_, _038124_, _038175_);
  or g_128596_(_038174_, _038175_, _038176_);
  and g_128597_(_009264_, _032762_, _038177_);
  not g_128598_(_038177_, _038178_);
  and g_128599_(_032673_, _032763_, _038179_);
  or g_128600_(_032672_, _032762_, _038181_);
  and g_128601_(_038178_, _038181_, _038182_);
  or g_128602_(_038177_, _038179_, _038183_);
  and g_128603_(_015345_, _038123_, _038184_);
  or g_128604_(_015346_, _038124_, _038185_);
  or g_128605_(_038030_, _038123_, _038186_);
  not g_128606_(_038186_, _038187_);
  and g_128607_(_038185_, _038186_, _038188_);
  or g_128608_(_038184_, _038187_, _038189_);
  and g_128609_(_038182_, _038189_, _038190_);
  or g_128610_(_009192_, _032763_, _038192_);
  or g_128611_(_032599_, _032762_, _038193_);
  and g_128612_(_038192_, _038193_, _038194_);
  or g_128613_(_015305_, _038124_, _038195_);
  or g_128614_(_037961_, _038123_, _038196_);
  and g_128615_(_038195_, _038196_, _038197_);
  or g_128616_(_032620_, _032762_, _038198_);
  or g_128617_(_032616_, _032763_, _038199_);
  and g_128618_(_038198_, _038199_, _038200_);
  or g_128619_(_037954_, _038123_, _038201_);
  or g_128620_(_037948_, _038124_, _038203_);
  and g_128621_(_038201_, _038203_, _038204_);
  and g_128622_(_038183_, _038188_, _038205_);
  or g_128623_(_009290_, _032763_, _038206_);
  or g_128624_(_032700_, _032762_, _038207_);
  and g_128625_(_038206_, _038207_, _038208_);
  or g_128626_(_015360_, _038124_, _038209_);
  or g_128627_(_038053_, _038123_, _038210_);
  and g_128628_(_038209_, _038210_, _038211_);
  and g_128629_(_032705_, _032763_, _038212_);
  and g_128630_(_053881_, _032762_, _038214_);
  or g_128631_(_038212_, _038214_, _038215_);
  and g_128632_(_038057_, _038124_, _038216_);
  and g_128633_(_002905_, _038123_, _038217_);
  or g_128634_(_038216_, _038217_, _038218_);
  and g_128635_(_038143_, _038149_, _038219_);
  xor g_128636_(_038215_, _038218_, _038220_);
  or g_128637_(_038155_, _038220_, _038221_);
  or g_128638_(_038163_, _038190_, _038222_);
  or g_128639_(_038221_, _038222_, _038223_);
  not g_128640_(_038223_, _038225_);
  xor g_128641_(_038173_, _038176_, _038226_);
  or g_128642_(_038137_, _038226_, _038227_);
  xor g_128643_(_038208_, _038211_, _038228_);
  or g_128644_(_038129_, _038228_, _038229_);
  or g_128645_(_038227_, _038229_, _038230_);
  xor g_128646_(_038194_, _038197_, _038231_);
  xor g_128647_(_038166_, _038170_, _038232_);
  or g_128648_(_038231_, _038232_, _038233_);
  xor g_128649_(_038200_, _038204_, _038234_);
  or g_128650_(_038205_, _038219_, _038236_);
  or g_128651_(_038234_, _038236_, _038237_);
  or g_128652_(_038233_, _038237_, _038238_);
  or g_128653_(_038230_, _038238_, _038239_);
  not g_128654_(_038239_, _038240_);
  and g_128655_(_038225_, _038240_, _038241_);
  or g_128656_(out[465], out[464], _038242_);
  or g_128657_(out[464], _053880_, _038243_);
  and g_128658_(out[467], _038243_, _038244_);
  and g_128659_(_021300_, _038243_, _038245_);
  and g_128660_(out[469], _038245_, _038247_);
  or g_128661_(out[470], _038247_, _038248_);
  and g_128662_(out[471], _038248_, _038249_);
  and g_128663_(out[472], _038249_, _038250_);
  or g_128664_(out[473], _038250_, _038251_);
  and g_128665_(out[474], _038251_, _038252_);
  xor g_128666_(out[475], _038252_, _038253_);
  xor g_128667_(_004828_, _038252_, _038254_);
  or g_128668_(out[449], out[448], _038255_);
  or g_128669_(out[448], _053560_, _038256_);
  and g_128670_(out[451], _038256_, _038258_);
  and g_128671_(_021111_, _038256_, _038259_);
  and g_128672_(out[453], _038259_, _038260_);
  or g_128673_(out[454], _038260_, _038261_);
  and g_128674_(out[455], _038261_, _038262_);
  and g_128675_(out[456], _038262_, _038263_);
  or g_128676_(out[457], _038263_, _038264_);
  and g_128677_(out[458], _038264_, _038265_);
  xor g_128678_(out[459], _038265_, _038266_);
  xor g_128679_(_004795_, _038265_, _038267_);
  or g_128680_(out[433], out[432], _038269_);
  or g_128681_(out[432], _053386_, _038270_);
  and g_128682_(out[435], _038270_, _038271_);
  and g_128683_(_020958_, _038270_, _038272_);
  and g_128684_(out[437], _038272_, _038273_);
  or g_128685_(out[438], _038273_, _038274_);
  and g_128686_(out[439], _038274_, _038275_);
  and g_128687_(out[440], _038275_, _038276_);
  or g_128688_(out[441], _038276_, _038277_);
  and g_128689_(out[442], _038277_, _038278_);
  xor g_128690_(out[443], _038278_, _038280_);
  xor g_128691_(_004762_, _038278_, _038281_);
  or g_128692_(out[417], out[416], _038282_);
  or g_128693_(out[416], _053270_, _038283_);
  and g_128694_(out[419], _038283_, _038284_);
  and g_128695_(_020797_, _038283_, _038285_);
  and g_128696_(out[421], _038285_, _038286_);
  or g_128697_(out[422], _038286_, _038287_);
  and g_128698_(out[423], _038287_, _038288_);
  and g_128699_(out[424], _038288_, _038289_);
  or g_128700_(out[425], _038289_, _038291_);
  and g_128701_(out[426], _038291_, _038292_);
  xor g_128702_(out[427], _038292_, _038293_);
  xor g_128703_(_004729_, _038292_, _038294_);
  or g_128704_(out[401], out[400], _038295_);
  or g_128705_(out[400], _053009_, _038296_);
  and g_128706_(out[403], _038296_, _038297_);
  and g_128707_(_020576_, _038296_, _038298_);
  and g_128708_(out[405], _038298_, _038299_);
  or g_128709_(out[406], _038299_, _038300_);
  and g_128710_(out[407], _038300_, _038302_);
  and g_128711_(out[408], _038302_, _038303_);
  or g_128712_(out[409], _038303_, _038304_);
  and g_128713_(out[410], _038304_, _038305_);
  xor g_128714_(out[411], _038305_, _038306_);
  xor g_128715_(_004696_, _038305_, _038307_);
  or g_128716_(out[385], out[384], _038308_);
  or g_128717_(out[384], _052921_, _038309_);
  and g_128718_(out[387], _038309_, _038310_);
  and g_128719_(_020352_, _038309_, _038311_);
  and g_128720_(out[389], _038311_, _038313_);
  or g_128721_(out[390], _038313_, _038314_);
  and g_128722_(out[391], _038314_, _038315_);
  and g_128723_(out[392], _038315_, _038316_);
  or g_128724_(out[393], _038316_, _038317_);
  and g_128725_(out[394], _038317_, _038318_);
  xor g_128726_(out[395], _038318_, _038319_);
  xor g_128727_(_004663_, _038318_, _038320_);
  or g_128728_(out[369], out[368], _038321_);
  or g_128729_(out[368], _052741_, _038322_);
  and g_128730_(out[371], _038322_, _038324_);
  and g_128731_(_020134_, _038322_, _038325_);
  and g_128732_(out[373], _038325_, _038326_);
  or g_128733_(out[374], _038326_, _038327_);
  and g_128734_(out[375], _038327_, _038328_);
  and g_128735_(out[376], _038328_, _038329_);
  or g_128736_(out[377], _038329_, _038330_);
  and g_128737_(out[378], _038330_, _038331_);
  xor g_128738_(out[379], _038331_, _038332_);
  xor g_128739_(_004630_, _038331_, _038333_);
  or g_128740_(out[353], out[352], _038335_);
  or g_128741_(out[352], _052547_, _038336_);
  and g_128742_(out[355], _038336_, _038337_);
  and g_128743_(_019962_, _038336_, _038338_);
  and g_128744_(out[357], _038338_, _038339_);
  or g_128745_(out[358], _038339_, _038340_);
  and g_128746_(out[359], _038340_, _038341_);
  and g_128747_(out[360], _038341_, _038342_);
  or g_128748_(out[361], _038342_, _038343_);
  and g_128749_(out[362], _038343_, _038344_);
  xor g_128750_(out[363], _038344_, _038346_);
  xor g_128751_(_004597_, _038344_, _038347_);
  xor g_128752_(out[362], _038343_, _038348_);
  xor g_128753_(_004619_, _038343_, _038349_);
  or g_128754_(out[337], out[336], _038350_);
  or g_128755_(out[336], _052353_, _038351_);
  and g_128756_(out[339], _038351_, _038352_);
  and g_128757_(_019791_, _038351_, _038353_);
  and g_128758_(out[341], _038353_, _038354_);
  or g_128759_(out[342], _038354_, _038355_);
  and g_128760_(out[343], _038355_, _038357_);
  and g_128761_(out[344], _038357_, _038358_);
  or g_128762_(out[345], _038358_, _038359_);
  and g_128763_(out[346], _038359_, _038360_);
  xor g_128764_(out[346], _038359_, _038361_);
  not g_128765_(_038361_, _038362_);
  xor g_128766_(out[345], _038358_, _038363_);
  xor g_128767_(_053533_, _038358_, _038364_);
  or g_128768_(out[321], out[320], _038365_);
  or g_128769_(out[320], _052166_, _038366_);
  and g_128770_(out[323], _038366_, _038368_);
  and g_128771_(_019605_, _038366_, _038369_);
  and g_128772_(out[325], _038369_, _038370_);
  or g_128773_(out[326], _038370_, _038371_);
  and g_128774_(out[327], _038371_, _038372_);
  and g_128775_(out[328], _038372_, _038373_);
  or g_128776_(out[329], _038373_, _038374_);
  xor g_128777_(out[329], _038373_, _038375_);
  xor g_128778_(_053434_, _038373_, _038376_);
  xor g_128779_(out[326], _038370_, _038377_);
  xor g_128780_(_053379_, _038370_, _038379_);
  or g_128781_(out[177], out[176], _038380_);
  or g_128782_(out[176], _042679_, _038381_);
  and g_128783_(out[179], _038381_, _038382_);
  and g_128784_(_017755_, _038381_, _038383_);
  and g_128785_(out[181], _038383_, _038384_);
  or g_128786_(out[182], _038384_, _038385_);
  xor g_128787_(out[182], _038384_, _038386_);
  xor g_128788_(_003772_, _038384_, _038387_);
  or g_128789_(out[81], out[80], _038388_);
  or g_128790_(out[80], _026575_, _038390_);
  and g_128791_(out[83], _038390_, _038391_);
  and g_128792_(_016381_, _038390_, _038392_);
  and g_128793_(out[85], _038392_, _038393_);
  or g_128794_(out[86], _038393_, _038394_);
  and g_128795_(out[87], _038394_, _038395_);
  and g_128796_(out[88], _038395_, _038396_);
  or g_128797_(out[89], _038396_, _038397_);
  and g_128798_(out[90], _038397_, _038398_);
  xor g_128799_(out[90], _038397_, _038399_);
  not g_128800_(_038399_, _038401_);
  or g_128801_(out[65], out[64], _038402_);
  or g_128802_(out[64], _026608_, _038403_);
  and g_128803_(out[67], _038403_, _038404_);
  and g_128804_(_016164_, _038403_, _038405_);
  and g_128805_(out[69], _038405_, _038406_);
  or g_128806_(out[70], _038406_, _038407_);
  and g_128807_(out[71], _038407_, _038408_);
  and g_128808_(out[72], _038408_, _038409_);
  or g_128809_(out[73], _038409_, _038410_);
  and g_128810_(out[74], _038410_, _038412_);
  xor g_128811_(_002826_, _038412_, _038413_);
  not g_128812_(_038413_, _038414_);
  xor g_128813_(out[66], _038402_, _038415_);
  xor g_128814_(_002903_, _038402_, _038416_);
  or g_128815_(out[49], out[48], _038417_);
  or g_128816_(out[48], _010823_, _038418_);
  xor g_128817_(out[50], _038417_, _038419_);
  xor g_128818_(_002771_, _038417_, _038420_);
  and g_128819_(out[51], _038418_, _038421_);
  and g_128820_(_015987_, _038418_, _038423_);
  and g_128821_(out[53], _038423_, _038424_);
  or g_128822_(out[54], _038424_, _038425_);
  and g_128823_(out[55], _038425_, _038426_);
  and g_128824_(out[56], _038426_, _038427_);
  or g_128825_(out[57], _038427_, _038428_);
  and g_128826_(out[58], _038428_, _038429_);
  xor g_128827_(out[58], _038428_, _038430_);
  not g_128828_(_038430_, _038431_);
  or g_128829_(out[33], out[32], _038432_);
  or g_128830_(out[32], _007831_, _038434_);
  and g_128831_(out[35], _038434_, _038435_);
  and g_128832_(_015708_, _038434_, _038436_);
  and g_128833_(out[37], _038436_, _038437_);
  or g_128834_(out[38], _038437_, _038438_);
  and g_128835_(out[39], _038438_, _038439_);
  and g_128836_(out[40], _038439_, _038440_);
  or g_128837_(out[41], _038440_, _038441_);
  and g_128838_(out[42], _038441_, _038442_);
  xor g_128839_(out[42], _038441_, _038443_);
  not g_128840_(_038443_, _038445_);
  or g_128841_(out[1], out[0], _038446_);
  not g_128842_(_038446_, _038447_);
  or g_128843_(out[2], _038446_, _038448_);
  and g_128844_(out[3], _038448_, _038449_);
  and g_128845_(_015556_, _038448_, _038450_);
  and g_128846_(_015628_, _038448_, _038451_);
  or g_128847_(out[6], _038451_, _038452_);
  and g_128848_(out[7], _038452_, _038453_);
  and g_128849_(out[8], _038453_, _038454_);
  or g_128850_(out[9], _038454_, _038456_);
  and g_128851_(out[10], _038456_, _038457_);
  xor g_128852_(out[10], _038456_, _038458_);
  xor g_128853_(_002419_, _038456_, _038459_);
  xor g_128854_(out[9], _038454_, _038460_);
  xor g_128855_(_002408_, _038454_, _038461_);
  or g_128856_(out[17], out[16], _038462_);
  or g_128857_(out[16], _005818_, _038463_);
  and g_128858_(out[19], _038463_, _038464_);
  and g_128859_(_015567_, _038463_, _038465_);
  and g_128860_(_015632_, _038463_, _038467_);
  or g_128861_(out[22], _038467_, _038468_);
  and g_128862_(out[23], _038468_, _038469_);
  and g_128863_(out[24], _038469_, _038470_);
  or g_128864_(out[25], _038470_, _038471_);
  xor g_128865_(out[25], _038470_, _038472_);
  xor g_128866_(_002540_, _038470_, _038473_);
  and g_128867_(_038460_, _038473_, _038474_);
  or g_128868_(_038461_, _038472_, _038475_);
  and g_128869_(out[26], _038471_, _038476_);
  xor g_128870_(out[26], _038471_, _038478_);
  xor g_128871_(_002551_, _038471_, _038479_);
  and g_128872_(_038459_, _038478_, _038480_);
  or g_128873_(_038458_, _038479_, _038481_);
  and g_128874_(_038475_, _038481_, _038482_);
  or g_128875_(_038474_, _038480_, _038483_);
  and g_128876_(_038461_, _038472_, _038484_);
  or g_128877_(_038460_, _038473_, _038485_);
  xor g_128878_(out[24], _038469_, _038486_);
  xor g_128879_(_002529_, _038469_, _038487_);
  xor g_128880_(out[8], _038453_, _038489_);
  xor g_128881_(_002397_, _038453_, _038490_);
  and g_128882_(_038487_, _038489_, _038491_);
  or g_128883_(_038486_, _038490_, _038492_);
  and g_128884_(_038485_, _038492_, _038493_);
  or g_128885_(_038484_, _038491_, _038494_);
  xor g_128886_(out[7], _038452_, _038495_);
  xor g_128887_(_002309_, _038452_, _038496_);
  xor g_128888_(out[23], _038468_, _038497_);
  xor g_128889_(_002441_, _038468_, _038498_);
  and g_128890_(_038496_, _038497_, _038500_);
  or g_128891_(_038495_, _038498_, _038501_);
  and g_128892_(_038486_, _038490_, _038502_);
  or g_128893_(_038487_, _038489_, _038503_);
  and g_128894_(_038501_, _038503_, _038504_);
  or g_128895_(_038500_, _038502_, _038505_);
  and g_128896_(_038495_, _038498_, _038506_);
  or g_128897_(_038496_, _038497_, _038507_);
  xor g_128898_(out[4], _038449_, _038508_);
  xor g_128899_(_002342_, _038449_, _038509_);
  xor g_128900_(out[20], _038464_, _038511_);
  xor g_128901_(_002474_, _038464_, _038512_);
  and g_128902_(_038508_, _038512_, _038513_);
  or g_128903_(_038509_, _038511_, _038514_);
  xor g_128904_(out[6], _038451_, _038515_);
  xor g_128905_(_002320_, _038451_, _038516_);
  xor g_128906_(out[22], _038467_, _038517_);
  xor g_128907_(_002452_, _038467_, _038518_);
  and g_128908_(_038516_, _038517_, _038519_);
  or g_128909_(_038515_, _038518_, _038520_);
  xor g_128910_(out[21], _038465_, _038522_);
  xor g_128911_(_002463_, _038465_, _038523_);
  xor g_128912_(out[5], _038450_, _038524_);
  xor g_128913_(_002331_, _038450_, _038525_);
  and g_128914_(_038523_, _038524_, _038526_);
  or g_128915_(_038522_, _038525_, _038527_);
  and g_128916_(_038520_, _038527_, _038528_);
  or g_128917_(_038519_, _038526_, _038529_);
  and g_128918_(_038514_, _038528_, _038530_);
  or g_128919_(_038513_, _038529_, _038531_);
  and g_128920_(_038515_, _038518_, _038533_);
  or g_128921_(_038516_, _038517_, _038534_);
  and g_128922_(_038522_, _038525_, _038535_);
  or g_128923_(_038523_, _038524_, _038536_);
  and g_128924_(_038534_, _038536_, _038537_);
  or g_128925_(_038533_, _038535_, _038538_);
  and g_128926_(_038509_, _038511_, _038539_);
  or g_128927_(_038508_, _038512_, _038540_);
  and g_128928_(_006313_, _038540_, _038541_);
  or g_128929_(_006324_, _038539_, _038542_);
  and g_128930_(_038537_, _038541_, _038544_);
  or g_128931_(_038538_, _038542_, _038545_);
  and g_128932_(_038530_, _038544_, _038546_);
  or g_128933_(_038531_, _038545_, _038547_);
  and g_128934_(_038520_, _038538_, _038548_);
  or g_128935_(_038519_, _038537_, _038549_);
  and g_128936_(out[1], out[17], _038550_);
  not g_128937_(_038550_, _038551_);
  and g_128938_(_006038_, _038550_, _038552_);
  or g_128939_(_006027_, _038551_, _038553_);
  and g_128940_(_002485_, out[16], _038555_);
  or g_128941_(out[17], _002496_, _038556_);
  and g_128942_(_038446_, _038556_, _038557_);
  or g_128943_(_038447_, _038555_, _038558_);
  and g_128944_(_038553_, _038557_, _038559_);
  or g_128945_(_038552_, _038558_, _038560_);
  xor g_128946_(out[2], _038446_, _038561_);
  xor g_128947_(_002375_, _038446_, _038562_);
  xor g_128948_(out[18], _038462_, _038563_);
  xor g_128949_(_002507_, _038462_, _038564_);
  and g_128950_(_038561_, _038564_, _038566_);
  or g_128951_(_038562_, _038563_, _038567_);
  and g_128952_(_038560_, _038567_, _038568_);
  or g_128953_(_038559_, _038566_, _038569_);
  xor g_128954_(out[19], _038463_, _038570_);
  xor g_128955_(_002518_, _038463_, _038571_);
  xor g_128956_(out[3], _038448_, _038572_);
  xor g_128957_(_002386_, _038448_, _038573_);
  and g_128958_(_038571_, _038572_, _038574_);
  or g_128959_(_038570_, _038573_, _038575_);
  and g_128960_(_038562_, _038563_, _038577_);
  or g_128961_(_038561_, _038564_, _038578_);
  and g_128962_(_038575_, _038578_, _038579_);
  or g_128963_(_038574_, _038577_, _038580_);
  and g_128964_(_038569_, _038579_, _038581_);
  or g_128965_(_038568_, _038580_, _038582_);
  and g_128966_(_038570_, _038573_, _038583_);
  or g_128967_(_038571_, _038572_, _038584_);
  and g_128968_(_038540_, _038584_, _038585_);
  or g_128969_(_038539_, _038583_, _038586_);
  and g_128970_(_038582_, _038585_, _038588_);
  or g_128971_(_038581_, _038586_, _038589_);
  and g_128972_(_038530_, _038589_, _038590_);
  or g_128973_(_038531_, _038588_, _038591_);
  and g_128974_(_038549_, _038591_, _038592_);
  or g_128975_(_038548_, _038590_, _038593_);
  and g_128976_(_038547_, _038592_, _038594_);
  or g_128977_(_038546_, _038593_, _038595_);
  and g_128978_(_038507_, _038595_, _038596_);
  or g_128979_(_038506_, _038594_, _038597_);
  and g_128980_(_038504_, _038597_, _038599_);
  or g_128981_(_038505_, _038596_, _038600_);
  and g_128982_(_038493_, _038600_, _038601_);
  or g_128983_(_038494_, _038599_, _038602_);
  and g_128984_(_038482_, _038602_, _038603_);
  or g_128985_(_038483_, _038601_, _038604_);
  and g_128986_(_038458_, _038479_, _038605_);
  or g_128987_(_038459_, _038478_, _038606_);
  xor g_128988_(out[11], _038457_, _038607_);
  xor g_128989_(_002298_, _038457_, _038608_);
  xor g_128990_(out[27], _038476_, _038610_);
  xor g_128991_(_002430_, _038476_, _038611_);
  and g_128992_(_038607_, _038611_, _038612_);
  or g_128993_(_038608_, _038610_, _038613_);
  and g_128994_(_038606_, _038613_, _038614_);
  or g_128995_(_038605_, _038612_, _038615_);
  and g_128996_(_038604_, _038614_, _038616_);
  or g_128997_(_038603_, _038615_, _038617_);
  and g_128998_(_038608_, _038610_, _038618_);
  or g_128999_(_038607_, _038611_, _038619_);
  and g_129000_(_038617_, _038619_, _038621_);
  or g_129001_(_038616_, _038618_, _038622_);
  or g_129002_(_038458_, _038621_, _038623_);
  or g_129003_(_038478_, _038622_, _038624_);
  and g_129004_(_038623_, _038624_, _038625_);
  not g_129005_(_038625_, _038626_);
  and g_129006_(_038443_, _038626_, _038627_);
  or g_129007_(_038445_, _038625_, _038628_);
  and g_129008_(_038607_, _038610_, _038629_);
  or g_129009_(_038608_, _038611_, _038630_);
  xor g_129010_(out[43], _038442_, _038632_);
  xor g_129011_(_002562_, _038442_, _038633_);
  and g_129012_(_038630_, _038632_, _038634_);
  or g_129013_(_038629_, _038633_, _038635_);
  and g_129014_(_038628_, _038635_, _038636_);
  or g_129015_(_038627_, _038634_, _038637_);
  and g_129016_(_038629_, _038633_, _038638_);
  or g_129017_(_038630_, _038632_, _038639_);
  and g_129018_(_038637_, _038639_, _038640_);
  or g_129019_(_038636_, _038638_, _038641_);
  and g_129020_(_038460_, _038622_, _038643_);
  or g_129021_(_038461_, _038621_, _038644_);
  and g_129022_(_038472_, _038621_, _038645_);
  or g_129023_(_038473_, _038622_, _038646_);
  and g_129024_(_038644_, _038646_, _038647_);
  or g_129025_(_038643_, _038645_, _038648_);
  xor g_129026_(out[41], _038440_, _038649_);
  xor g_129027_(_002672_, _038440_, _038650_);
  and g_129028_(_038648_, _038650_, _038651_);
  or g_129029_(_038647_, _038649_, _038652_);
  xor g_129030_(out[40], _038439_, _038654_);
  not g_129031_(_038654_, _038655_);
  and g_129032_(_038490_, _038622_, _038656_);
  or g_129033_(_038489_, _038621_, _038657_);
  and g_129034_(_038487_, _038621_, _038658_);
  or g_129035_(_038486_, _038622_, _038659_);
  and g_129036_(_038657_, _038659_, _038660_);
  or g_129037_(_038656_, _038658_, _038661_);
  and g_129038_(_038654_, _038661_, _038662_);
  or g_129039_(_038655_, _038660_, _038663_);
  and g_129040_(_038652_, _038663_, _038665_);
  or g_129041_(_038651_, _038662_, _038666_);
  xor g_129042_(out[39], _038438_, _038667_);
  xor g_129043_(_002573_, _038438_, _038668_);
  and g_129044_(_038496_, _038622_, _038669_);
  or g_129045_(_038495_, _038621_, _038670_);
  and g_129046_(_038498_, _038621_, _038671_);
  or g_129047_(_038497_, _038622_, _038672_);
  and g_129048_(_038670_, _038672_, _038673_);
  or g_129049_(_038669_, _038671_, _038674_);
  and g_129050_(_038667_, _038674_, _038676_);
  or g_129051_(_038668_, _038673_, _038677_);
  xor g_129052_(_002617_, out[32], _038678_);
  not g_129053_(_038678_, _038679_);
  xor g_129054_(out[17], out[16], _038680_);
  xor g_129055_(_002485_, out[16], _038681_);
  and g_129056_(_038621_, _038681_, _038682_);
  or g_129057_(_038622_, _038680_, _038683_);
  xor g_129058_(out[1], out[0], _038684_);
  xor g_129059_(_002353_, out[0], _038685_);
  and g_129060_(_038622_, _038685_, _038687_);
  or g_129061_(_038621_, _038684_, _038688_);
  and g_129062_(_038683_, _038688_, _038689_);
  or g_129063_(_038682_, _038687_, _038690_);
  and g_129064_(_038679_, _038690_, _038691_);
  or g_129065_(_038678_, _038689_, _038692_);
  and g_129066_(out[16], _038621_, _038693_);
  or g_129067_(_002496_, _038622_, _038694_);
  and g_129068_(out[0], _038622_, _038695_);
  or g_129069_(_002364_, _038621_, _038696_);
  and g_129070_(_038694_, _038696_, _038698_);
  or g_129071_(_038693_, _038695_, _038699_);
  and g_129072_(out[32], _038698_, _038700_);
  or g_129073_(_002628_, _038699_, _038701_);
  and g_129074_(_038692_, _038701_, _038702_);
  or g_129075_(_038691_, _038700_, _038703_);
  xor g_129076_(out[34], _038432_, _038704_);
  xor g_129077_(_002639_, _038432_, _038705_);
  and g_129078_(_038563_, _038621_, _038706_);
  or g_129079_(_038564_, _038622_, _038707_);
  and g_129080_(_038561_, _038622_, _038709_);
  or g_129081_(_038562_, _038621_, _038710_);
  and g_129082_(_038707_, _038710_, _038711_);
  or g_129083_(_038706_, _038709_, _038712_);
  and g_129084_(_038705_, _038712_, _038713_);
  or g_129085_(_038704_, _038711_, _038714_);
  and g_129086_(out[33], _038689_, _038715_);
  or g_129087_(_002617_, _038690_, _038716_);
  and g_129088_(_038714_, _038716_, _038717_);
  or g_129089_(_038713_, _038715_, _038718_);
  and g_129090_(_038703_, _038717_, _038720_);
  or g_129091_(_038702_, _038718_, _038721_);
  xor g_129092_(out[35], _038434_, _038722_);
  xor g_129093_(_002650_, _038434_, _038723_);
  and g_129094_(_038573_, _038622_, _038724_);
  or g_129095_(_038572_, _038621_, _038725_);
  and g_129096_(_038571_, _038621_, _038726_);
  or g_129097_(_038570_, _038622_, _038727_);
  and g_129098_(_038725_, _038727_, _038728_);
  or g_129099_(_038724_, _038726_, _038729_);
  and g_129100_(_038723_, _038728_, _038731_);
  or g_129101_(_038722_, _038729_, _038732_);
  and g_129102_(_038704_, _038711_, _038733_);
  or g_129103_(_038705_, _038712_, _038734_);
  and g_129104_(_038732_, _038734_, _038735_);
  or g_129105_(_038731_, _038733_, _038736_);
  and g_129106_(_038721_, _038735_, _038737_);
  or g_129107_(_038720_, _038736_, _038738_);
  and g_129108_(_038722_, _038729_, _038739_);
  or g_129109_(_038723_, _038728_, _038740_);
  xor g_129110_(out[36], _038435_, _038742_);
  xor g_129111_(_002606_, _038435_, _038743_);
  and g_129112_(_038512_, _038621_, _038744_);
  or g_129113_(_038511_, _038622_, _038745_);
  and g_129114_(_038509_, _038622_, _038746_);
  or g_129115_(_038508_, _038621_, _038747_);
  and g_129116_(_038745_, _038747_, _038748_);
  or g_129117_(_038744_, _038746_, _038749_);
  and g_129118_(_038742_, _038749_, _038750_);
  or g_129119_(_038743_, _038748_, _038751_);
  and g_129120_(_038740_, _038751_, _038753_);
  or g_129121_(_038739_, _038750_, _038754_);
  and g_129122_(_038738_, _038753_, _038755_);
  or g_129123_(_038737_, _038754_, _038756_);
  and g_129124_(_038523_, _038621_, _038757_);
  or g_129125_(_038522_, _038622_, _038758_);
  and g_129126_(_038525_, _038622_, _038759_);
  or g_129127_(_038524_, _038621_, _038760_);
  and g_129128_(_038758_, _038760_, _038761_);
  or g_129129_(_038757_, _038759_, _038762_);
  xor g_129130_(out[37], _038436_, _038764_);
  xor g_129131_(_002595_, _038436_, _038765_);
  and g_129132_(_038761_, _038765_, _038766_);
  or g_129133_(_038762_, _038764_, _038767_);
  and g_129134_(_038743_, _038748_, _038768_);
  or g_129135_(_038742_, _038749_, _038769_);
  and g_129136_(_038767_, _038769_, _038770_);
  or g_129137_(_038766_, _038768_, _038771_);
  and g_129138_(_038756_, _038770_, _038772_);
  or g_129139_(_038755_, _038771_, _038773_);
  xor g_129140_(out[38], _038437_, _038775_);
  xor g_129141_(_002584_, _038437_, _038776_);
  and g_129142_(_038515_, _038622_, _038777_);
  or g_129143_(_038516_, _038621_, _038778_);
  and g_129144_(_038517_, _038621_, _038779_);
  or g_129145_(_038518_, _038622_, _038780_);
  and g_129146_(_038778_, _038780_, _038781_);
  or g_129147_(_038777_, _038779_, _038782_);
  and g_129148_(_038776_, _038782_, _038783_);
  or g_129149_(_038775_, _038781_, _038784_);
  and g_129150_(_038762_, _038764_, _038786_);
  or g_129151_(_038761_, _038765_, _038787_);
  and g_129152_(_038784_, _038787_, _038788_);
  or g_129153_(_038783_, _038786_, _038789_);
  and g_129154_(_038773_, _038788_, _038790_);
  or g_129155_(_038772_, _038789_, _038791_);
  and g_129156_(_038668_, _038673_, _038792_);
  or g_129157_(_038667_, _038674_, _038793_);
  and g_129158_(_038775_, _038781_, _038794_);
  or g_129159_(_038776_, _038782_, _038795_);
  and g_129160_(_038793_, _038795_, _038797_);
  or g_129161_(_038792_, _038794_, _038798_);
  and g_129162_(_038791_, _038797_, _038799_);
  or g_129163_(_038790_, _038798_, _038800_);
  and g_129164_(_038677_, _038800_, _038801_);
  or g_129165_(_038676_, _038799_, _038802_);
  and g_129166_(_038647_, _038649_, _038803_);
  or g_129167_(_038648_, _038650_, _038804_);
  and g_129168_(_038445_, _038625_, _038805_);
  or g_129169_(_038443_, _038626_, _038806_);
  and g_129170_(_038639_, _038806_, _038808_);
  or g_129171_(_038638_, _038805_, _038809_);
  and g_129172_(_038636_, _038808_, _038810_);
  or g_129173_(_038637_, _038809_, _038811_);
  and g_129174_(_038666_, _038810_, _038812_);
  or g_129175_(_038665_, _038811_, _038813_);
  and g_129176_(_038804_, _038812_, _038814_);
  or g_129177_(_038803_, _038813_, _038815_);
  xor g_129178_(_038655_, _038660_, _038816_);
  xor g_129179_(_038654_, _038660_, _038817_);
  and g_129180_(_038804_, _038816_, _038819_);
  or g_129181_(_038803_, _038817_, _038820_);
  and g_129182_(_038810_, _038819_, _038821_);
  or g_129183_(_038811_, _038820_, _038822_);
  and g_129184_(_038652_, _038821_, _038823_);
  or g_129185_(_038651_, _038822_, _038824_);
  and g_129186_(_038802_, _038823_, _038825_);
  or g_129187_(_038801_, _038824_, _038826_);
  and g_129188_(_038641_, _038826_, _038827_);
  or g_129189_(_038640_, _038825_, _038828_);
  and g_129190_(_038815_, _038827_, _038830_);
  or g_129191_(_038814_, _038828_, _038831_);
  or g_129192_(_038443_, _038831_, _038832_);
  or g_129193_(_038625_, _038830_, _038833_);
  and g_129194_(_038832_, _038833_, _038834_);
  not g_129195_(_038834_, _038835_);
  and g_129196_(_038431_, _038834_, _038836_);
  or g_129197_(_038430_, _038835_, _038837_);
  and g_129198_(_038629_, _038632_, _038838_);
  not g_129199_(_038838_, _038839_);
  xor g_129200_(out[59], _038429_, _038841_);
  not g_129201_(_038841_, _038842_);
  and g_129202_(_038838_, _038842_, _038843_);
  or g_129203_(_038839_, _038841_, _038844_);
  and g_129204_(_038837_, _038844_, _038845_);
  or g_129205_(_038836_, _038843_, _038846_);
  and g_129206_(_038430_, _038835_, _038847_);
  or g_129207_(_038431_, _038834_, _038848_);
  and g_129208_(_038839_, _038841_, _038849_);
  or g_129209_(_038838_, _038842_, _038850_);
  xor g_129210_(out[57], _038427_, _038852_);
  xor g_129211_(_002804_, _038427_, _038853_);
  and g_129212_(_038649_, _038830_, _038854_);
  or g_129213_(_038650_, _038831_, _038855_);
  and g_129214_(_038648_, _038831_, _038856_);
  or g_129215_(_038647_, _038830_, _038857_);
  and g_129216_(_038855_, _038857_, _038858_);
  or g_129217_(_038854_, _038856_, _038859_);
  and g_129218_(_038853_, _038859_, _038860_);
  or g_129219_(_038852_, _038858_, _038861_);
  and g_129220_(_038850_, _038861_, _038863_);
  or g_129221_(_038849_, _038860_, _038864_);
  and g_129222_(_038848_, _038863_, _038865_);
  or g_129223_(_038847_, _038864_, _038866_);
  and g_129224_(_038845_, _038865_, _038867_);
  or g_129225_(_038846_, _038866_, _038868_);
  and g_129226_(_038852_, _038858_, _038869_);
  or g_129227_(_038853_, _038859_, _038870_);
  xor g_129228_(out[56], _038426_, _038871_);
  xor g_129229_(_002793_, _038426_, _038872_);
  or g_129230_(_038654_, _038831_, _038874_);
  not g_129231_(_038874_, _038875_);
  and g_129232_(_038661_, _038831_, _038876_);
  or g_129233_(_038660_, _038830_, _038877_);
  and g_129234_(_038874_, _038877_, _038878_);
  or g_129235_(_038875_, _038876_, _038879_);
  and g_129236_(_038872_, _038878_, _038880_);
  or g_129237_(_038871_, _038879_, _038881_);
  and g_129238_(_038870_, _038881_, _038882_);
  or g_129239_(_038869_, _038880_, _038883_);
  and g_129240_(_038871_, _038879_, _038885_);
  or g_129241_(_038872_, _038878_, _038886_);
  and g_129242_(_038882_, _038886_, _038887_);
  or g_129243_(_038883_, _038885_, _038888_);
  and g_129244_(_038867_, _038887_, _038889_);
  or g_129245_(_038868_, _038888_, _038890_);
  and g_129246_(_038704_, _038830_, _038891_);
  or g_129247_(_038705_, _038831_, _038892_);
  and g_129248_(_038712_, _038831_, _038893_);
  or g_129249_(_038711_, _038830_, _038894_);
  and g_129250_(_038892_, _038894_, _038896_);
  or g_129251_(_038891_, _038893_, _038897_);
  and g_129252_(_038419_, _038896_, _038898_);
  or g_129253_(_038420_, _038897_, _038899_);
  xor g_129254_(out[51], _038418_, _038900_);
  xor g_129255_(_002782_, _038418_, _038901_);
  and g_129256_(_038723_, _038830_, _038902_);
  or g_129257_(_038722_, _038831_, _038903_);
  and g_129258_(_038729_, _038831_, _038904_);
  or g_129259_(_038728_, _038830_, _038905_);
  and g_129260_(_038903_, _038905_, _038907_);
  or g_129261_(_038902_, _038904_, _038908_);
  and g_129262_(_038901_, _038907_, _038909_);
  or g_129263_(_038900_, _038908_, _038910_);
  and g_129264_(_038899_, _038910_, _038911_);
  or g_129265_(_038898_, _038909_, _038912_);
  xor g_129266_(out[49], out[48], _038913_);
  not g_129267_(_038913_, _038914_);
  or g_129268_(_038678_, _038831_, _038915_);
  or g_129269_(_038690_, _038830_, _038916_);
  and g_129270_(_038915_, _038916_, _038918_);
  and g_129271_(_038913_, _038918_, _038919_);
  not g_129272_(_038919_, _038920_);
  and g_129273_(out[32], _038830_, _038921_);
  or g_129274_(_002628_, _038831_, _038922_);
  and g_129275_(_038699_, _038831_, _038923_);
  or g_129276_(_038698_, _038830_, _038924_);
  and g_129277_(_038922_, _038924_, _038925_);
  or g_129278_(_038921_, _038923_, _038926_);
  and g_129279_(_002760_, _038926_, _038927_);
  or g_129280_(out[48], _038925_, _038929_);
  xor g_129281_(_038913_, _038918_, _038930_);
  xor g_129282_(_038914_, _038918_, _038931_);
  and g_129283_(_038929_, _038930_, _038932_);
  or g_129284_(_038927_, _038931_, _038933_);
  and g_129285_(_038920_, _038933_, _038934_);
  or g_129286_(_038919_, _038932_, _038935_);
  and g_129287_(_038420_, _038897_, _038936_);
  or g_129288_(_038419_, _038896_, _038937_);
  and g_129289_(_038935_, _038937_, _038938_);
  or g_129290_(_038934_, _038936_, _038940_);
  and g_129291_(_038911_, _038940_, _038941_);
  or g_129292_(_038912_, _038938_, _038942_);
  and g_129293_(_038900_, _038908_, _038943_);
  or g_129294_(_038901_, _038907_, _038944_);
  xor g_129295_(out[54], _038424_, _038945_);
  xor g_129296_(_002716_, _038424_, _038946_);
  and g_129297_(_038775_, _038830_, _038947_);
  or g_129298_(_038776_, _038831_, _038948_);
  and g_129299_(_038782_, _038831_, _038949_);
  or g_129300_(_038781_, _038830_, _038951_);
  and g_129301_(_038948_, _038951_, _038952_);
  or g_129302_(_038947_, _038949_, _038953_);
  and g_129303_(_038945_, _038952_, _038954_);
  or g_129304_(_038946_, _038953_, _038955_);
  xor g_129305_(out[55], _038425_, _038956_);
  xor g_129306_(_002705_, _038425_, _038957_);
  and g_129307_(_038668_, _038830_, _038958_);
  or g_129308_(_038667_, _038831_, _038959_);
  and g_129309_(_038674_, _038831_, _038960_);
  or g_129310_(_038673_, _038830_, _038962_);
  and g_129311_(_038959_, _038962_, _038963_);
  or g_129312_(_038958_, _038960_, _038964_);
  and g_129313_(_038957_, _038963_, _038965_);
  or g_129314_(_038956_, _038964_, _038966_);
  and g_129315_(_038955_, _038966_, _038967_);
  or g_129316_(_038954_, _038965_, _038968_);
  and g_129317_(_038956_, _038964_, _038969_);
  or g_129318_(_038957_, _038963_, _038970_);
  and g_129319_(_038946_, _038953_, _038971_);
  or g_129320_(_038945_, _038952_, _038973_);
  and g_129321_(_038970_, _038973_, _038974_);
  or g_129322_(_038969_, _038971_, _038975_);
  and g_129323_(_038967_, _038974_, _038976_);
  or g_129324_(_038968_, _038975_, _038977_);
  and g_129325_(_038762_, _038831_, _038978_);
  or g_129326_(_038761_, _038830_, _038979_);
  and g_129327_(_038765_, _038830_, _038980_);
  or g_129328_(_038764_, _038831_, _038981_);
  and g_129329_(_038979_, _038981_, _038982_);
  or g_129330_(_038978_, _038980_, _038984_);
  xor g_129331_(out[53], _038423_, _038985_);
  xor g_129332_(_002727_, _038423_, _038986_);
  and g_129333_(_038982_, _038986_, _038987_);
  or g_129334_(_038984_, _038985_, _038988_);
  xor g_129335_(out[52], _038421_, _038989_);
  xor g_129336_(_002738_, _038421_, _038990_);
  and g_129337_(_038749_, _038831_, _038991_);
  or g_129338_(_038748_, _038830_, _038992_);
  and g_129339_(_038743_, _038830_, _038993_);
  or g_129340_(_038742_, _038831_, _038995_);
  and g_129341_(_038992_, _038995_, _038996_);
  or g_129342_(_038991_, _038993_, _038997_);
  and g_129343_(_038990_, _038996_, _038998_);
  or g_129344_(_038989_, _038997_, _038999_);
  and g_129345_(_038988_, _038999_, _039000_);
  or g_129346_(_038987_, _038998_, _039001_);
  and g_129347_(_038989_, _038997_, _039002_);
  or g_129348_(_038990_, _038996_, _039003_);
  and g_129349_(_038984_, _038985_, _039004_);
  or g_129350_(_038982_, _038986_, _039006_);
  and g_129351_(_039003_, _039006_, _039007_);
  or g_129352_(_039002_, _039004_, _039008_);
  and g_129353_(_039000_, _039007_, _039009_);
  or g_129354_(_039001_, _039008_, _039010_);
  and g_129355_(_038976_, _039009_, _039011_);
  or g_129356_(_038977_, _039010_, _039012_);
  and g_129357_(_038944_, _039011_, _039013_);
  or g_129358_(_038943_, _039012_, _039014_);
  and g_129359_(_038942_, _039013_, _039015_);
  or g_129360_(_038941_, _039014_, _039017_);
  and g_129361_(_038968_, _038970_, _039018_);
  or g_129362_(_038967_, _038969_, _039019_);
  and g_129363_(_039001_, _039006_, _039020_);
  or g_129364_(_039000_, _039004_, _039021_);
  and g_129365_(_038976_, _039020_, _039022_);
  or g_129366_(_038977_, _039021_, _039023_);
  and g_129367_(_039019_, _039023_, _039024_);
  or g_129368_(_039018_, _039022_, _039025_);
  and g_129369_(_039017_, _039024_, _039026_);
  or g_129370_(_039015_, _039025_, _039028_);
  and g_129371_(_038889_, _039028_, _039029_);
  or g_129372_(_038890_, _039026_, _039030_);
  and g_129373_(_038867_, _038883_, _039031_);
  or g_129374_(_038868_, _038882_, _039032_);
  and g_129375_(_038846_, _038850_, _039033_);
  or g_129376_(_038845_, _038849_, _039034_);
  and g_129377_(_039032_, _039034_, _039035_);
  or g_129378_(_039031_, _039033_, _039036_);
  and g_129379_(_039030_, _039035_, _039037_);
  or g_129380_(_039029_, _039036_, _039039_);
  and g_129381_(out[48], _038925_, _039040_);
  or g_129382_(_002760_, _038926_, _039041_);
  and g_129383_(_038937_, _038944_, _039042_);
  or g_129384_(_038936_, _038943_, _039043_);
  and g_129385_(_039041_, _039042_, _039044_);
  or g_129386_(_039040_, _039043_, _039045_);
  and g_129387_(_038911_, _039044_, _039046_);
  or g_129388_(_038912_, _039045_, _039047_);
  and g_129389_(_038932_, _039046_, _039048_);
  or g_129390_(_038933_, _039047_, _039050_);
  and g_129391_(_038889_, _039048_, _039051_);
  or g_129392_(_038890_, _039050_, _039052_);
  and g_129393_(_039011_, _039051_, _039053_);
  or g_129394_(_039012_, _039052_, _039054_);
  and g_129395_(_039039_, _039054_, _039055_);
  or g_129396_(_039037_, _039053_, _039056_);
  and g_129397_(_038419_, _039055_, _039057_);
  not g_129398_(_039057_, _039058_);
  or g_129399_(_038896_, _039055_, _039059_);
  not g_129400_(_039059_, _039061_);
  and g_129401_(_039058_, _039059_, _039062_);
  or g_129402_(_039057_, _039061_, _039063_);
  and g_129403_(_038415_, _039062_, _039064_);
  or g_129404_(_038416_, _039063_, _039065_);
  xor g_129405_(_002914_, _038403_, _039066_);
  or g_129406_(_038900_, _039056_, _039067_);
  or g_129407_(_038907_, _039055_, _039068_);
  and g_129408_(_039067_, _039068_, _039069_);
  and g_129409_(_039066_, _039069_, _039070_);
  not g_129410_(_039070_, _039072_);
  and g_129411_(_039065_, _039072_, _039073_);
  or g_129412_(_039064_, _039070_, _039074_);
  xor g_129413_(out[65], out[64], _039075_);
  not g_129414_(_039075_, _039076_);
  and g_129415_(_038913_, _039055_, _039077_);
  not g_129416_(_039077_, _039078_);
  or g_129417_(_038918_, _039055_, _039079_);
  not g_129418_(_039079_, _039080_);
  and g_129419_(_039078_, _039079_, _039081_);
  or g_129420_(_039077_, _039080_, _039083_);
  and g_129421_(_039075_, _039081_, _039084_);
  or g_129422_(_039076_, _039083_, _039085_);
  and g_129423_(out[48], _039055_, _039086_);
  not g_129424_(_039086_, _039087_);
  or g_129425_(_038925_, _039055_, _039088_);
  not g_129426_(_039088_, _039089_);
  and g_129427_(_039087_, _039088_, _039090_);
  or g_129428_(_039086_, _039089_, _039091_);
  and g_129429_(_002892_, _039091_, _039092_);
  or g_129430_(out[64], _039090_, _039094_);
  xor g_129431_(_039075_, _039081_, _039095_);
  xor g_129432_(_039076_, _039081_, _039096_);
  and g_129433_(_039094_, _039095_, _039097_);
  or g_129434_(_039092_, _039096_, _039098_);
  and g_129435_(_039085_, _039098_, _039099_);
  or g_129436_(_039084_, _039097_, _039100_);
  and g_129437_(_038416_, _039063_, _039101_);
  or g_129438_(_038415_, _039062_, _039102_);
  and g_129439_(_039100_, _039102_, _039103_);
  or g_129440_(_039099_, _039101_, _039105_);
  and g_129441_(_039073_, _039105_, _039106_);
  or g_129442_(_039074_, _039103_, _039107_);
  xor g_129443_(out[71], _038407_, _039108_);
  xor g_129444_(_002837_, _038407_, _039109_);
  and g_129445_(_038957_, _039055_, _039110_);
  or g_129446_(_038956_, _039056_, _039111_);
  and g_129447_(_038964_, _039056_, _039112_);
  or g_129448_(_038963_, _039055_, _039113_);
  and g_129449_(_039111_, _039113_, _039114_);
  or g_129450_(_039110_, _039112_, _039116_);
  and g_129451_(_039109_, _039114_, _039117_);
  not g_129452_(_039117_, _039118_);
  xor g_129453_(out[70], _038406_, _039119_);
  not g_129454_(_039119_, _039120_);
  and g_129455_(_038945_, _039055_, _039121_);
  or g_129456_(_038946_, _039056_, _039122_);
  and g_129457_(_038953_, _039056_, _039123_);
  or g_129458_(_038952_, _039055_, _039124_);
  and g_129459_(_039122_, _039124_, _039125_);
  or g_129460_(_039121_, _039123_, _039127_);
  and g_129461_(_039119_, _039125_, _039128_);
  not g_129462_(_039128_, _039129_);
  and g_129463_(_039118_, _039129_, _039130_);
  or g_129464_(_039117_, _039128_, _039131_);
  xor g_129465_(out[69], _038405_, _039132_);
  xor g_129466_(_002859_, _038405_, _039133_);
  or g_129467_(_038982_, _039055_, _039134_);
  not g_129468_(_039134_, _039135_);
  and g_129469_(_038986_, _039055_, _039136_);
  not g_129470_(_039136_, _039138_);
  and g_129471_(_039134_, _039138_, _039139_);
  or g_129472_(_039135_, _039136_, _039140_);
  and g_129473_(_039132_, _039140_, _039141_);
  or g_129474_(_039133_, _039139_, _039142_);
  and g_129475_(_039120_, _039127_, _039143_);
  or g_129476_(_039119_, _039125_, _039144_);
  and g_129477_(_039108_, _039116_, _039145_);
  or g_129478_(_039109_, _039114_, _039146_);
  and g_129479_(_039144_, _039146_, _039147_);
  or g_129480_(_039143_, _039145_, _039149_);
  and g_129481_(_039142_, _039147_, _039150_);
  or g_129482_(_039141_, _039149_, _039151_);
  and g_129483_(_039130_, _039150_, _039152_);
  or g_129484_(_039131_, _039151_, _039153_);
  xor g_129485_(out[74], _038410_, _039154_);
  xor g_129486_(_002947_, _038410_, _039155_);
  or g_129487_(_038430_, _039056_, _039156_);
  or g_129488_(_038834_, _039055_, _039157_);
  and g_129489_(_039156_, _039157_, _039158_);
  and g_129490_(_039155_, _039158_, _039160_);
  or g_129491_(_038841_, _039056_, _039161_);
  or g_129492_(_038838_, _039055_, _039162_);
  and g_129493_(_039161_, _039162_, _039163_);
  or g_129494_(_038413_, _039163_, _039164_);
  and g_129495_(_038413_, _039163_, _039165_);
  xor g_129496_(_039155_, _039158_, _039166_);
  xor g_129497_(_039154_, _039158_, _039167_);
  xor g_129498_(_038413_, _039163_, _039168_);
  xor g_129499_(_038414_, _039163_, _039169_);
  and g_129500_(_039166_, _039168_, _039171_);
  or g_129501_(_039167_, _039169_, _039172_);
  xor g_129502_(out[72], _038408_, _039173_);
  xor g_129503_(_002925_, _038408_, _039174_);
  and g_129504_(_038872_, _039055_, _039175_);
  or g_129505_(_038871_, _039056_, _039176_);
  and g_129506_(_038879_, _039056_, _039177_);
  or g_129507_(_038878_, _039055_, _039178_);
  and g_129508_(_039176_, _039178_, _039179_);
  or g_129509_(_039175_, _039177_, _039180_);
  and g_129510_(_039174_, _039179_, _039182_);
  or g_129511_(_039173_, _039180_, _039183_);
  xor g_129512_(out[73], _038409_, _039184_);
  not g_129513_(_039184_, _039185_);
  and g_129514_(_038852_, _039055_, _039186_);
  or g_129515_(_038853_, _039056_, _039187_);
  and g_129516_(_038859_, _039056_, _039188_);
  or g_129517_(_038858_, _039055_, _039189_);
  and g_129518_(_039187_, _039189_, _039190_);
  or g_129519_(_039186_, _039188_, _039191_);
  and g_129520_(_039184_, _039190_, _039193_);
  or g_129521_(_039185_, _039191_, _039194_);
  and g_129522_(_039183_, _039194_, _039195_);
  or g_129523_(_039182_, _039193_, _039196_);
  and g_129524_(_039185_, _039191_, _039197_);
  or g_129525_(_039184_, _039190_, _039198_);
  and g_129526_(_039173_, _039180_, _039199_);
  or g_129527_(_039174_, _039179_, _039200_);
  and g_129528_(_039198_, _039200_, _039201_);
  or g_129529_(_039197_, _039199_, _039202_);
  and g_129530_(_039195_, _039201_, _039204_);
  or g_129531_(_039196_, _039202_, _039205_);
  and g_129532_(_039171_, _039204_, _039206_);
  or g_129533_(_039172_, _039205_, _039207_);
  and g_129534_(_039152_, _039206_, _039208_);
  or g_129535_(_039153_, _039207_, _039209_);
  and g_129536_(_039133_, _039139_, _039210_);
  not g_129537_(_039210_, _039211_);
  xor g_129538_(out[68], _038404_, _039212_);
  xor g_129539_(_002870_, _038404_, _039213_);
  or g_129540_(_038989_, _039056_, _039215_);
  or g_129541_(_038996_, _039055_, _039216_);
  and g_129542_(_039215_, _039216_, _039217_);
  not g_129543_(_039217_, _039218_);
  and g_129544_(_039213_, _039217_, _039219_);
  or g_129545_(_039212_, _039218_, _039220_);
  and g_129546_(_039211_, _039220_, _039221_);
  or g_129547_(_039210_, _039219_, _039222_);
  or g_129548_(_039066_, _039069_, _039223_);
  or g_129549_(_039213_, _039217_, _039224_);
  and g_129550_(_039223_, _039224_, _039226_);
  not g_129551_(_039226_, _039227_);
  and g_129552_(_039221_, _039226_, _039228_);
  or g_129553_(_039222_, _039227_, _039229_);
  and g_129554_(_039208_, _039228_, _039230_);
  or g_129555_(_039209_, _039229_, _039231_);
  and g_129556_(_039107_, _039230_, _039232_);
  or g_129557_(_039106_, _039231_, _039233_);
  and g_129558_(_039208_, _039222_, _039234_);
  or g_129559_(_039209_, _039221_, _039235_);
  and g_129560_(_039171_, _039196_, _039237_);
  or g_129561_(_039172_, _039195_, _039238_);
  and g_129562_(_039198_, _039237_, _039239_);
  or g_129563_(_039197_, _039238_, _039240_);
  and g_129564_(_039160_, _039164_, _039241_);
  or g_129565_(_039165_, _039241_, _039242_);
  not g_129566_(_039242_, _039243_);
  and g_129567_(_039240_, _039243_, _039244_);
  or g_129568_(_039239_, _039242_, _039245_);
  and g_129569_(_039131_, _039146_, _039246_);
  not g_129570_(_039246_, _039248_);
  and g_129571_(_039206_, _039246_, _039249_);
  or g_129572_(_039207_, _039248_, _039250_);
  and g_129573_(_039244_, _039250_, _039251_);
  or g_129574_(_039245_, _039249_, _039252_);
  and g_129575_(_039235_, _039251_, _039253_);
  or g_129576_(_039234_, _039252_, _039254_);
  and g_129577_(_039233_, _039253_, _039255_);
  or g_129578_(_039232_, _039254_, _039256_);
  and g_129579_(out[64], _039090_, _039257_);
  or g_129580_(_039101_, _039257_, _039259_);
  or g_129581_(_039074_, _039259_, _039260_);
  not g_129582_(_039260_, _039261_);
  and g_129583_(_039097_, _039261_, _039262_);
  and g_129584_(_039230_, _039262_, _039263_);
  not g_129585_(_039263_, _039264_);
  and g_129586_(_039256_, _039264_, _039265_);
  or g_129587_(_039255_, _039263_, _039266_);
  and g_129588_(_038413_, _039265_, _039267_);
  not g_129589_(_039267_, _039268_);
  or g_129590_(_039163_, _039265_, _039270_);
  not g_129591_(_039270_, _039271_);
  and g_129592_(_039268_, _039270_, _039272_);
  or g_129593_(_039267_, _039271_, _039273_);
  xor g_129594_(out[91], _038398_, _039274_);
  xor g_129595_(_002958_, _038398_, _039275_);
  and g_129596_(_039273_, _039274_, _039276_);
  or g_129597_(_039273_, _039274_, _039277_);
  and g_129598_(_039155_, _039265_, _039278_);
  not g_129599_(_039278_, _039279_);
  or g_129600_(_039158_, _039265_, _039281_);
  not g_129601_(_039281_, _039282_);
  and g_129602_(_039279_, _039281_, _039283_);
  or g_129603_(_039278_, _039282_, _039284_);
  and g_129604_(_038399_, _039284_, _039285_);
  and g_129605_(_039277_, _039285_, _039286_);
  or g_129606_(_039276_, _039286_, _039287_);
  not g_129607_(_039287_, _039288_);
  xor g_129608_(out[89], _038396_, _039289_);
  xor g_129609_(_003068_, _038396_, _039290_);
  and g_129610_(_039184_, _039265_, _039292_);
  not g_129611_(_039292_, _039293_);
  or g_129612_(_039190_, _039265_, _039294_);
  not g_129613_(_039294_, _039295_);
  and g_129614_(_039293_, _039294_, _039296_);
  or g_129615_(_039292_, _039295_, _039297_);
  and g_129616_(_039290_, _039297_, _039298_);
  or g_129617_(_039289_, _039296_, _039299_);
  xor g_129618_(out[88], _038395_, _039300_);
  xor g_129619_(_003057_, _038395_, _039301_);
  and g_129620_(_039174_, _039265_, _039303_);
  not g_129621_(_039303_, _039304_);
  or g_129622_(_039179_, _039265_, _039305_);
  not g_129623_(_039305_, _039306_);
  and g_129624_(_039304_, _039305_, _039307_);
  or g_129625_(_039303_, _039306_, _039308_);
  and g_129626_(_039300_, _039308_, _039309_);
  or g_129627_(_039301_, _039307_, _039310_);
  and g_129628_(_039299_, _039310_, _039311_);
  or g_129629_(_039298_, _039309_, _039312_);
  and g_129630_(out[64], _039265_, _039314_);
  or g_129631_(_002892_, _039266_, _039315_);
  and g_129632_(_039091_, _039266_, _039316_);
  or g_129633_(_039090_, _039265_, _039317_);
  and g_129634_(_039315_, _039317_, _039318_);
  or g_129635_(_039314_, _039316_, _039319_);
  and g_129636_(out[80], _039318_, _039320_);
  or g_129637_(_003024_, _039319_, _039321_);
  and g_129638_(_039075_, _039265_, _039322_);
  or g_129639_(_039076_, _039266_, _039323_);
  and g_129640_(_039083_, _039266_, _039325_);
  or g_129641_(_039081_, _039265_, _039326_);
  and g_129642_(_039323_, _039326_, _039327_);
  or g_129643_(_039322_, _039325_, _039328_);
  and g_129644_(out[81], _039328_, _039329_);
  or g_129645_(_003013_, _039327_, _039330_);
  xor g_129646_(out[81], out[80], _039331_);
  xor g_129647_(_003013_, out[80], _039332_);
  and g_129648_(_039320_, _039330_, _039333_);
  or g_129649_(_039321_, _039329_, _039334_);
  xor g_129650_(out[82], _038388_, _039336_);
  xor g_129651_(_003035_, _038388_, _039337_);
  and g_129652_(_038415_, _039265_, _039338_);
  or g_129653_(_038416_, _039266_, _039339_);
  and g_129654_(_039063_, _039266_, _039340_);
  or g_129655_(_039062_, _039265_, _039341_);
  and g_129656_(_039339_, _039341_, _039342_);
  or g_129657_(_039338_, _039340_, _039343_);
  and g_129658_(_039336_, _039342_, _039344_);
  or g_129659_(_039337_, _039343_, _039345_);
  and g_129660_(_039327_, _039331_, _039347_);
  or g_129661_(_039328_, _039332_, _039348_);
  and g_129662_(_039345_, _039348_, _039349_);
  or g_129663_(_039344_, _039347_, _039350_);
  and g_129664_(_039334_, _039349_, _039351_);
  or g_129665_(_039333_, _039350_, _039352_);
  and g_129666_(_039066_, _039265_, _039353_);
  not g_129667_(_039353_, _039354_);
  or g_129668_(_039069_, _039265_, _039355_);
  not g_129669_(_039355_, _039356_);
  and g_129670_(_039354_, _039355_, _039358_);
  or g_129671_(_039353_, _039356_, _039359_);
  xor g_129672_(out[83], _038390_, _039360_);
  xor g_129673_(_003046_, _038390_, _039361_);
  and g_129674_(_039359_, _039360_, _039362_);
  or g_129675_(_039358_, _039361_, _039363_);
  and g_129676_(_039337_, _039343_, _039364_);
  or g_129677_(_039336_, _039342_, _039365_);
  and g_129678_(_039363_, _039365_, _039366_);
  or g_129679_(_039362_, _039364_, _039367_);
  and g_129680_(_039352_, _039366_, _039369_);
  or g_129681_(_039351_, _039367_, _039370_);
  xor g_129682_(out[84], _038391_, _039371_);
  xor g_129683_(_003002_, _038391_, _039372_);
  and g_129684_(_039213_, _039265_, _039373_);
  not g_129685_(_039373_, _039374_);
  or g_129686_(_039217_, _039265_, _039375_);
  not g_129687_(_039375_, _039376_);
  and g_129688_(_039374_, _039375_, _039377_);
  or g_129689_(_039373_, _039376_, _039378_);
  and g_129690_(_039372_, _039377_, _039380_);
  or g_129691_(_039371_, _039378_, _039381_);
  and g_129692_(_039358_, _039361_, _039382_);
  or g_129693_(_039359_, _039360_, _039383_);
  and g_129694_(_039381_, _039383_, _039384_);
  or g_129695_(_039380_, _039382_, _039385_);
  and g_129696_(_039370_, _039384_, _039386_);
  or g_129697_(_039369_, _039385_, _039387_);
  xor g_129698_(out[85], _038392_, _039388_);
  xor g_129699_(_002991_, _038392_, _039389_);
  and g_129700_(_039133_, _039265_, _039391_);
  not g_129701_(_039391_, _039392_);
  or g_129702_(_039139_, _039265_, _039393_);
  not g_129703_(_039393_, _039394_);
  and g_129704_(_039392_, _039393_, _039395_);
  or g_129705_(_039391_, _039394_, _039396_);
  and g_129706_(_039388_, _039396_, _039397_);
  or g_129707_(_039389_, _039395_, _039398_);
  and g_129708_(_039371_, _039378_, _039399_);
  or g_129709_(_039372_, _039377_, _039400_);
  and g_129710_(_039398_, _039400_, _039402_);
  or g_129711_(_039397_, _039399_, _039403_);
  and g_129712_(_039387_, _039402_, _039404_);
  or g_129713_(_039386_, _039403_, _039405_);
  xor g_129714_(out[86], _038393_, _039406_);
  xor g_129715_(_002980_, _038393_, _039407_);
  and g_129716_(_039119_, _039265_, _039408_);
  not g_129717_(_039408_, _039409_);
  or g_129718_(_039125_, _039265_, _039410_);
  not g_129719_(_039410_, _039411_);
  and g_129720_(_039409_, _039410_, _039413_);
  or g_129721_(_039408_, _039411_, _039414_);
  and g_129722_(_039406_, _039413_, _039415_);
  or g_129723_(_039407_, _039414_, _039416_);
  and g_129724_(_039389_, _039395_, _039417_);
  or g_129725_(_039388_, _039396_, _039418_);
  and g_129726_(_039416_, _039418_, _039419_);
  or g_129727_(_039415_, _039417_, _039420_);
  and g_129728_(_039405_, _039419_, _039421_);
  or g_129729_(_039404_, _039420_, _039422_);
  xor g_129730_(out[87], _038394_, _039424_);
  xor g_129731_(_002969_, _038394_, _039425_);
  and g_129732_(_039109_, _039265_, _039426_);
  not g_129733_(_039426_, _039427_);
  or g_129734_(_039114_, _039265_, _039428_);
  not g_129735_(_039428_, _039429_);
  and g_129736_(_039427_, _039428_, _039430_);
  or g_129737_(_039426_, _039429_, _039431_);
  and g_129738_(_039424_, _039431_, _039432_);
  or g_129739_(_039425_, _039430_, _039433_);
  and g_129740_(_039407_, _039414_, _039435_);
  or g_129741_(_039406_, _039413_, _039436_);
  and g_129742_(_039433_, _039436_, _039437_);
  or g_129743_(_039432_, _039435_, _039438_);
  and g_129744_(_039422_, _039437_, _039439_);
  or g_129745_(_039421_, _039438_, _039440_);
  and g_129746_(_039301_, _039307_, _039441_);
  or g_129747_(_039300_, _039308_, _039442_);
  and g_129748_(_039425_, _039430_, _039443_);
  or g_129749_(_039424_, _039431_, _039444_);
  and g_129750_(_039442_, _039444_, _039446_);
  or g_129751_(_039441_, _039443_, _039447_);
  and g_129752_(_039289_, _039296_, _039448_);
  or g_129753_(_039290_, _039297_, _039449_);
  xor g_129754_(_038401_, _039283_, _039450_);
  xor g_129755_(_038399_, _039283_, _039451_);
  xor g_129756_(_039273_, _039274_, _039452_);
  xor g_129757_(_039272_, _039274_, _039453_);
  and g_129758_(_039450_, _039452_, _039454_);
  or g_129759_(_039451_, _039453_, _039455_);
  and g_129760_(_039312_, _039454_, _039457_);
  or g_129761_(_039311_, _039455_, _039458_);
  and g_129762_(_039449_, _039457_, _039459_);
  or g_129763_(_039448_, _039458_, _039460_);
  and g_129764_(_039288_, _039460_, _039461_);
  or g_129765_(_039287_, _039459_, _039462_);
  and g_129766_(_039311_, _039449_, _039463_);
  or g_129767_(_039312_, _039448_, _039464_);
  and g_129768_(_039446_, _039463_, _039465_);
  or g_129769_(_039447_, _039464_, _039466_);
  and g_129770_(_039440_, _039465_, _039468_);
  or g_129771_(_039439_, _039466_, _039469_);
  and g_129772_(_039454_, _039468_, _039470_);
  or g_129773_(_039455_, _039469_, _039471_);
  and g_129774_(_039461_, _039471_, _039472_);
  or g_129775_(_039462_, _039470_, _039473_);
  and g_129776_(_038401_, _039472_, _039474_);
  or g_129777_(_038399_, _039473_, _039475_);
  and g_129778_(_039284_, _039473_, _039476_);
  or g_129779_(_039283_, _039472_, _039477_);
  and g_129780_(_039475_, _039477_, _039479_);
  or g_129781_(_039474_, _039476_, _039480_);
  or g_129782_(out[97], out[96], _039481_);
  or g_129783_(out[96], _031195_, _039482_);
  and g_129784_(out[99], _039482_, _039483_);
  xor g_129785_(out[99], _039482_, _039484_);
  xor g_129786_(_003178_, _039482_, _039485_);
  and g_129787_(_039361_, _039472_, _039486_);
  or g_129788_(_039360_, _039473_, _039487_);
  and g_129789_(_039359_, _039473_, _039488_);
  or g_129790_(_039358_, _039472_, _039490_);
  and g_129791_(_039487_, _039490_, _039491_);
  or g_129792_(_039486_, _039488_, _039492_);
  and g_129793_(_039484_, _039492_, _039493_);
  or g_129794_(_039485_, _039491_, _039494_);
  and g_129795_(_039485_, _039491_, _039495_);
  or g_129796_(_039484_, _039492_, _039496_);
  xor g_129797_(out[98], _039481_, _039497_);
  xor g_129798_(_003167_, _039481_, _039498_);
  and g_129799_(_039336_, _039472_, _039499_);
  or g_129800_(_039337_, _039473_, _039501_);
  and g_129801_(_039343_, _039473_, _039502_);
  or g_129802_(_039342_, _039472_, _039503_);
  and g_129803_(_039501_, _039503_, _039504_);
  or g_129804_(_039499_, _039502_, _039505_);
  and g_129805_(_039497_, _039504_, _039506_);
  or g_129806_(_039498_, _039505_, _039507_);
  and g_129807_(_039496_, _039507_, _039508_);
  or g_129808_(_039495_, _039506_, _039509_);
  and g_129809_(_039494_, _039509_, _039510_);
  or g_129810_(_039493_, _039508_, _039512_);
  xor g_129811_(out[97], out[96], _039513_);
  not g_129812_(_039513_, _039514_);
  and g_129813_(_039331_, _039472_, _039515_);
  or g_129814_(_039332_, _039473_, _039516_);
  and g_129815_(_039328_, _039473_, _039517_);
  or g_129816_(_039327_, _039472_, _039518_);
  and g_129817_(_039516_, _039518_, _039519_);
  or g_129818_(_039515_, _039517_, _039520_);
  and g_129819_(_039513_, _039519_, _039521_);
  or g_129820_(_039514_, _039520_, _039523_);
  and g_129821_(out[80], _039472_, _039524_);
  or g_129822_(_003024_, _039473_, _039525_);
  and g_129823_(_039319_, _039473_, _039526_);
  or g_129824_(_039318_, _039472_, _039527_);
  and g_129825_(_039525_, _039527_, _039528_);
  or g_129826_(_039524_, _039526_, _039529_);
  and g_129827_(_003156_, _039529_, _039530_);
  or g_129828_(out[96], _039528_, _039531_);
  xor g_129829_(_039513_, _039519_, _039532_);
  xor g_129830_(_039514_, _039519_, _039534_);
  and g_129831_(_039531_, _039532_, _039535_);
  or g_129832_(_039530_, _039534_, _039536_);
  and g_129833_(_039523_, _039536_, _039537_);
  or g_129834_(_039521_, _039535_, _039538_);
  and g_129835_(_039498_, _039505_, _039539_);
  or g_129836_(_039497_, _039504_, _039540_);
  and g_129837_(_039494_, _039540_, _039541_);
  or g_129838_(_039493_, _039539_, _039542_);
  and g_129839_(_039538_, _039541_, _039543_);
  or g_129840_(_039537_, _039542_, _039545_);
  and g_129841_(_039512_, _039545_, _039546_);
  or g_129842_(_039510_, _039543_, _039547_);
  and g_129843_(_039272_, _039274_, _039548_);
  or g_129844_(_039273_, _039275_, _039549_);
  and g_129845_(_016602_, _039482_, _039550_);
  and g_129846_(out[101], _039550_, _039551_);
  or g_129847_(out[102], _039551_, _039552_);
  and g_129848_(out[103], _039552_, _039553_);
  and g_129849_(out[104], _039553_, _039554_);
  or g_129850_(out[105], _039554_, _039556_);
  and g_129851_(out[106], _039556_, _039557_);
  xor g_129852_(out[107], _039557_, _039558_);
  xor g_129853_(_003090_, _039557_, _039559_);
  and g_129854_(_039548_, _039559_, _039560_);
  or g_129855_(_039549_, _039558_, _039561_);
  xor g_129856_(out[106], _039556_, _039562_);
  xor g_129857_(_003211_, _039556_, _039563_);
  and g_129858_(_039479_, _039563_, _039564_);
  or g_129859_(_039480_, _039562_, _039565_);
  and g_129860_(_039561_, _039565_, _039567_);
  or g_129861_(_039560_, _039564_, _039568_);
  and g_129862_(_039480_, _039562_, _039569_);
  or g_129863_(_039479_, _039563_, _039570_);
  and g_129864_(_039549_, _039558_, _039571_);
  or g_129865_(_039548_, _039559_, _039572_);
  xor g_129866_(out[105], _039554_, _039573_);
  xor g_129867_(_003200_, _039554_, _039574_);
  and g_129868_(_039289_, _039472_, _039575_);
  or g_129869_(_039290_, _039473_, _039576_);
  and g_129870_(_039297_, _039473_, _039578_);
  or g_129871_(_039296_, _039472_, _039579_);
  and g_129872_(_039576_, _039579_, _039580_);
  or g_129873_(_039575_, _039578_, _039581_);
  and g_129874_(_039574_, _039581_, _039582_);
  or g_129875_(_039573_, _039580_, _039583_);
  and g_129876_(_039570_, _039572_, _039584_);
  or g_129877_(_039569_, _039571_, _039585_);
  and g_129878_(_039567_, _039584_, _039586_);
  or g_129879_(_039568_, _039585_, _039587_);
  and g_129880_(_039583_, _039586_, _039589_);
  or g_129881_(_039582_, _039587_, _039590_);
  xor g_129882_(out[104], _039553_, _039591_);
  xor g_129883_(_003189_, _039553_, _039592_);
  and g_129884_(_039301_, _039472_, _039593_);
  or g_129885_(_039300_, _039473_, _039594_);
  and g_129886_(_039308_, _039473_, _039595_);
  or g_129887_(_039307_, _039472_, _039596_);
  and g_129888_(_039594_, _039596_, _039597_);
  or g_129889_(_039593_, _039595_, _039598_);
  and g_129890_(_039591_, _039598_, _039600_);
  or g_129891_(_039592_, _039597_, _039601_);
  and g_129892_(_039573_, _039580_, _039602_);
  or g_129893_(_039574_, _039581_, _039603_);
  and g_129894_(_039592_, _039597_, _039604_);
  or g_129895_(_039591_, _039598_, _039605_);
  and g_129896_(_039603_, _039605_, _039606_);
  or g_129897_(_039602_, _039604_, _039607_);
  and g_129898_(_039601_, _039606_, _039608_);
  or g_129899_(_039600_, _039607_, _039609_);
  and g_129900_(_039589_, _039608_, _039611_);
  or g_129901_(_039590_, _039609_, _039612_);
  xor g_129902_(out[102], _039551_, _039613_);
  xor g_129903_(_003112_, _039551_, _039614_);
  and g_129904_(_039406_, _039472_, _039615_);
  or g_129905_(_039407_, _039473_, _039616_);
  and g_129906_(_039414_, _039473_, _039617_);
  or g_129907_(_039413_, _039472_, _039618_);
  and g_129908_(_039616_, _039618_, _039619_);
  or g_129909_(_039615_, _039617_, _039620_);
  and g_129910_(_039613_, _039619_, _039622_);
  or g_129911_(_039614_, _039620_, _039623_);
  xor g_129912_(out[103], _039552_, _039624_);
  xor g_129913_(_003101_, _039552_, _039625_);
  and g_129914_(_039425_, _039472_, _039626_);
  or g_129915_(_039424_, _039473_, _039627_);
  and g_129916_(_039431_, _039473_, _039628_);
  or g_129917_(_039430_, _039472_, _039629_);
  and g_129918_(_039627_, _039629_, _039630_);
  or g_129919_(_039626_, _039628_, _039631_);
  and g_129920_(_039625_, _039630_, _039633_);
  or g_129921_(_039624_, _039631_, _039634_);
  and g_129922_(_039623_, _039634_, _039635_);
  or g_129923_(_039622_, _039633_, _039636_);
  and g_129924_(_039624_, _039631_, _039637_);
  or g_129925_(_039625_, _039630_, _039638_);
  and g_129926_(_039614_, _039620_, _039639_);
  or g_129927_(_039613_, _039619_, _039640_);
  and g_129928_(_039638_, _039640_, _039641_);
  or g_129929_(_039637_, _039639_, _039642_);
  and g_129930_(_039635_, _039641_, _039644_);
  or g_129931_(_039636_, _039642_, _039645_);
  xor g_129932_(out[101], _039550_, _039646_);
  xor g_129933_(_003123_, _039550_, _039647_);
  and g_129934_(_039389_, _039472_, _039648_);
  or g_129935_(_039388_, _039473_, _039649_);
  and g_129936_(_039396_, _039473_, _039650_);
  or g_129937_(_039395_, _039472_, _039651_);
  and g_129938_(_039649_, _039651_, _039652_);
  or g_129939_(_039648_, _039650_, _039653_);
  and g_129940_(_039647_, _039652_, _039655_);
  or g_129941_(_039646_, _039653_, _039656_);
  xor g_129942_(out[100], _039483_, _039657_);
  xor g_129943_(_003134_, _039483_, _039658_);
  and g_129944_(_039378_, _039473_, _039659_);
  or g_129945_(_039377_, _039472_, _039660_);
  and g_129946_(_039372_, _039472_, _039661_);
  or g_129947_(_039371_, _039473_, _039662_);
  and g_129948_(_039660_, _039662_, _039663_);
  or g_129949_(_039659_, _039661_, _039664_);
  and g_129950_(_039658_, _039663_, _039666_);
  or g_129951_(_039657_, _039664_, _039667_);
  and g_129952_(_039656_, _039667_, _039668_);
  or g_129953_(_039655_, _039666_, _039669_);
  and g_129954_(_039657_, _039664_, _039670_);
  or g_129955_(_039658_, _039663_, _039671_);
  and g_129956_(_039646_, _039653_, _039672_);
  or g_129957_(_039647_, _039652_, _039673_);
  and g_129958_(_039671_, _039673_, _039674_);
  or g_129959_(_039670_, _039672_, _039675_);
  and g_129960_(_039668_, _039674_, _039677_);
  or g_129961_(_039669_, _039675_, _039678_);
  and g_129962_(_039644_, _039677_, _039679_);
  or g_129963_(_039645_, _039678_, _039680_);
  and g_129964_(_039611_, _039679_, _039681_);
  or g_129965_(_039612_, _039680_, _039682_);
  and g_129966_(_039547_, _039681_, _039683_);
  or g_129967_(_039546_, _039682_, _039684_);
  and g_129968_(_039636_, _039638_, _039685_);
  or g_129969_(_039635_, _039637_, _039686_);
  and g_129970_(_039669_, _039673_, _039688_);
  or g_129971_(_039668_, _039672_, _039689_);
  and g_129972_(_039641_, _039688_, _039690_);
  or g_129973_(_039642_, _039689_, _039691_);
  and g_129974_(_039686_, _039691_, _039692_);
  or g_129975_(_039685_, _039690_, _039693_);
  and g_129976_(_039611_, _039693_, _039694_);
  or g_129977_(_039612_, _039692_, _039695_);
  and g_129978_(_039589_, _039607_, _039696_);
  or g_129979_(_039590_, _039606_, _039697_);
  and g_129980_(_039568_, _039572_, _039699_);
  or g_129981_(_039567_, _039571_, _039700_);
  and g_129982_(_039697_, _039700_, _039701_);
  or g_129983_(_039696_, _039699_, _039702_);
  and g_129984_(_039695_, _039701_, _039703_);
  or g_129985_(_039694_, _039702_, _039704_);
  and g_129986_(_039684_, _039703_, _039705_);
  or g_129987_(_039683_, _039704_, _039706_);
  and g_129988_(out[96], _039528_, _039707_);
  or g_129989_(_003156_, _039529_, _039708_);
  and g_129990_(_039508_, _039708_, _039710_);
  or g_129991_(_039509_, _039707_, _039711_);
  and g_129992_(_039541_, _039710_, _039712_);
  or g_129993_(_039542_, _039711_, _039713_);
  and g_129994_(_039535_, _039712_, _039714_);
  or g_129995_(_039536_, _039713_, _039715_);
  and g_129996_(_039681_, _039714_, _039716_);
  or g_129997_(_039682_, _039715_, _039717_);
  and g_129998_(_039706_, _039717_, _039718_);
  or g_129999_(_039705_, _039716_, _039719_);
  and g_130000_(_039480_, _039719_, _039721_);
  or g_130001_(_039479_, _039718_, _039722_);
  and g_130002_(_039563_, _039718_, _039723_);
  or g_130003_(_039562_, _039719_, _039724_);
  and g_130004_(_039722_, _039724_, _039725_);
  or g_130005_(_039721_, _039723_, _039726_);
  or g_130006_(out[113], out[112], _039727_);
  or g_130007_(out[112], _034110_, _039728_);
  and g_130008_(out[115], _039728_, _039729_);
  and g_130009_(_016847_, _039728_, _039730_);
  and g_130010_(out[117], _039730_, _039732_);
  or g_130011_(out[118], _039732_, _039733_);
  and g_130012_(out[119], _039733_, _039734_);
  xor g_130013_(out[119], _039733_, _039735_);
  xor g_130014_(_003233_, _039733_, _039736_);
  and g_130015_(_039631_, _039719_, _039737_);
  or g_130016_(_039630_, _039718_, _039738_);
  and g_130017_(_039625_, _039718_, _039739_);
  or g_130018_(_039624_, _039719_, _039740_);
  and g_130019_(_039738_, _039740_, _039741_);
  or g_130020_(_039737_, _039739_, _039743_);
  and g_130021_(_039735_, _039743_, _039744_);
  or g_130022_(_039736_, _039741_, _039745_);
  xor g_130023_(out[118], _039732_, _039746_);
  xor g_130024_(_003244_, _039732_, _039747_);
  and g_130025_(_039620_, _039719_, _039748_);
  or g_130026_(_039619_, _039718_, _039749_);
  and g_130027_(_039613_, _039718_, _039750_);
  or g_130028_(_039614_, _039719_, _039751_);
  and g_130029_(_039749_, _039751_, _039752_);
  or g_130030_(_039748_, _039750_, _039754_);
  and g_130031_(_039747_, _039754_, _039755_);
  or g_130032_(_039746_, _039752_, _039756_);
  xor g_130033_(out[117], _039730_, _039757_);
  xor g_130034_(_003255_, _039730_, _039758_);
  and g_130035_(_039653_, _039719_, _039759_);
  or g_130036_(_039652_, _039718_, _039760_);
  and g_130037_(_039647_, _039718_, _039761_);
  or g_130038_(_039646_, _039719_, _039762_);
  and g_130039_(_039760_, _039762_, _039763_);
  or g_130040_(_039759_, _039761_, _039765_);
  and g_130041_(_039758_, _039763_, _039766_);
  or g_130042_(_039757_, _039765_, _039767_);
  and g_130043_(out[96], _039718_, _039768_);
  or g_130044_(_003156_, _039719_, _039769_);
  and g_130045_(_039529_, _039719_, _039770_);
  or g_130046_(_039528_, _039718_, _039771_);
  and g_130047_(_039769_, _039771_, _039772_);
  or g_130048_(_039768_, _039770_, _039773_);
  and g_130049_(out[112], _039772_, _039774_);
  or g_130050_(_003288_, _039773_, _039776_);
  and g_130051_(_039520_, _039719_, _039777_);
  or g_130052_(_039519_, _039718_, _039778_);
  and g_130053_(_039513_, _039718_, _039779_);
  or g_130054_(_039514_, _039719_, _039780_);
  and g_130055_(_039778_, _039780_, _039781_);
  or g_130056_(_039777_, _039779_, _039782_);
  and g_130057_(out[113], _039782_, _039783_);
  or g_130058_(_003277_, _039781_, _039784_);
  xor g_130059_(out[113], out[112], _039785_);
  xor g_130060_(_003277_, out[112], _039787_);
  and g_130061_(_039774_, _039784_, _039788_);
  or g_130062_(_039776_, _039783_, _039789_);
  xor g_130063_(out[114], _039727_, _039790_);
  xor g_130064_(_003299_, _039727_, _039791_);
  and g_130065_(_039505_, _039719_, _039792_);
  or g_130066_(_039504_, _039718_, _039793_);
  and g_130067_(_039497_, _039718_, _039794_);
  or g_130068_(_039498_, _039719_, _039795_);
  and g_130069_(_039793_, _039795_, _039796_);
  or g_130070_(_039792_, _039794_, _039798_);
  and g_130071_(_039790_, _039796_, _039799_);
  or g_130072_(_039791_, _039798_, _039800_);
  and g_130073_(_039781_, _039785_, _039801_);
  or g_130074_(_039782_, _039787_, _039802_);
  and g_130075_(_039800_, _039802_, _039803_);
  or g_130076_(_039799_, _039801_, _039804_);
  and g_130077_(_039789_, _039803_, _039805_);
  or g_130078_(_039788_, _039804_, _039806_);
  xor g_130079_(out[115], _039728_, _039807_);
  xor g_130080_(_003310_, _039728_, _039809_);
  and g_130081_(_039485_, _039718_, _039810_);
  or g_130082_(_039484_, _039719_, _039811_);
  and g_130083_(_039492_, _039719_, _039812_);
  or g_130084_(_039491_, _039718_, _039813_);
  and g_130085_(_039811_, _039813_, _039814_);
  or g_130086_(_039810_, _039812_, _039815_);
  and g_130087_(_039807_, _039815_, _039816_);
  or g_130088_(_039809_, _039814_, _039817_);
  and g_130089_(_039791_, _039798_, _039818_);
  or g_130090_(_039790_, _039796_, _039820_);
  and g_130091_(_039817_, _039820_, _039821_);
  or g_130092_(_039816_, _039818_, _039822_);
  and g_130093_(_039806_, _039821_, _039823_);
  or g_130094_(_039805_, _039822_, _039824_);
  and g_130095_(_039809_, _039814_, _039825_);
  or g_130096_(_039807_, _039815_, _039826_);
  xor g_130097_(out[116], _039729_, _039827_);
  xor g_130098_(_003266_, _039729_, _039828_);
  and g_130099_(_039664_, _039719_, _039829_);
  or g_130100_(_039663_, _039718_, _039831_);
  and g_130101_(_039658_, _039718_, _039832_);
  or g_130102_(_039657_, _039719_, _039833_);
  and g_130103_(_039831_, _039833_, _039834_);
  or g_130104_(_039829_, _039832_, _039835_);
  and g_130105_(_039828_, _039834_, _039836_);
  or g_130106_(_039827_, _039835_, _039837_);
  and g_130107_(_039826_, _039837_, _039838_);
  or g_130108_(_039825_, _039836_, _039839_);
  and g_130109_(_039824_, _039838_, _039840_);
  or g_130110_(_039823_, _039839_, _039842_);
  and g_130111_(_039757_, _039765_, _039843_);
  or g_130112_(_039758_, _039763_, _039844_);
  and g_130113_(_039827_, _039835_, _039845_);
  or g_130114_(_039828_, _039834_, _039846_);
  and g_130115_(_039844_, _039846_, _039847_);
  or g_130116_(_039843_, _039845_, _039848_);
  and g_130117_(_039842_, _039847_, _039849_);
  or g_130118_(_039840_, _039848_, _039850_);
  and g_130119_(_039767_, _039850_, _039851_);
  or g_130120_(_039766_, _039849_, _039853_);
  and g_130121_(_039756_, _039853_, _039854_);
  or g_130122_(_039755_, _039851_, _039855_);
  and g_130123_(_039736_, _039741_, _039856_);
  or g_130124_(_039735_, _039743_, _039857_);
  and g_130125_(_039746_, _039752_, _039858_);
  or g_130126_(_039747_, _039754_, _039859_);
  and g_130127_(_039857_, _039859_, _039860_);
  or g_130128_(_039856_, _039858_, _039861_);
  and g_130129_(_039855_, _039860_, _039862_);
  or g_130130_(_039854_, _039861_, _039864_);
  and g_130131_(_039745_, _039864_, _039865_);
  or g_130132_(_039744_, _039862_, _039866_);
  and g_130133_(out[120], _039734_, _039867_);
  or g_130134_(out[121], _039867_, _039868_);
  and g_130135_(out[122], _039868_, _039869_);
  xor g_130136_(out[122], _039868_, _039870_);
  not g_130137_(_039870_, _039871_);
  and g_130138_(_039726_, _039870_, _039872_);
  or g_130139_(_039725_, _039871_, _039873_);
  and g_130140_(_039559_, _039718_, _039875_);
  or g_130141_(_039558_, _039719_, _039876_);
  and g_130142_(_039549_, _039719_, _039877_);
  or g_130143_(_039548_, _039718_, _039878_);
  and g_130144_(_039876_, _039878_, _039879_);
  or g_130145_(_039875_, _039877_, _039880_);
  xor g_130146_(out[123], _039869_, _039881_);
  xor g_130147_(_003222_, _039869_, _039882_);
  and g_130148_(_039880_, _039881_, _039883_);
  or g_130149_(_039879_, _039882_, _039884_);
  or g_130150_(_039872_, _039883_, _039886_);
  and g_130151_(_039725_, _039871_, _039887_);
  and g_130152_(_039879_, _039882_, _039888_);
  or g_130153_(_039880_, _039881_, _039889_);
  or g_130154_(_039887_, _039888_, _039890_);
  xor g_130155_(_039726_, _039870_, _039891_);
  and g_130156_(_039884_, _039889_, _039892_);
  and g_130157_(_039891_, _039892_, _039893_);
  or g_130158_(_039886_, _039890_, _039894_);
  xor g_130159_(out[120], _039734_, _039895_);
  xor g_130160_(_003321_, _039734_, _039897_);
  and g_130161_(_039598_, _039719_, _039898_);
  or g_130162_(_039597_, _039718_, _039899_);
  and g_130163_(_039592_, _039718_, _039900_);
  or g_130164_(_039591_, _039719_, _039901_);
  and g_130165_(_039899_, _039901_, _039902_);
  or g_130166_(_039898_, _039900_, _039903_);
  and g_130167_(_039895_, _039903_, _039904_);
  or g_130168_(_039897_, _039902_, _039905_);
  xor g_130169_(out[121], _039867_, _039906_);
  xor g_130170_(_003332_, _039867_, _039908_);
  and g_130171_(_039581_, _039719_, _039909_);
  or g_130172_(_039580_, _039718_, _039910_);
  and g_130173_(_039573_, _039718_, _039911_);
  or g_130174_(_039574_, _039719_, _039912_);
  and g_130175_(_039910_, _039912_, _039913_);
  or g_130176_(_039909_, _039911_, _039914_);
  and g_130177_(_039908_, _039914_, _039915_);
  or g_130178_(_039906_, _039913_, _039916_);
  and g_130179_(_039905_, _039916_, _039917_);
  or g_130180_(_039904_, _039915_, _039919_);
  and g_130181_(_039897_, _039902_, _039920_);
  or g_130182_(_039895_, _039903_, _039921_);
  and g_130183_(_039906_, _039913_, _039922_);
  or g_130184_(_039908_, _039914_, _039923_);
  and g_130185_(_039921_, _039923_, _039924_);
  or g_130186_(_039920_, _039922_, _039925_);
  and g_130187_(_039917_, _039924_, _039926_);
  or g_130188_(_039919_, _039925_, _039927_);
  and g_130189_(_039893_, _039926_, _039928_);
  or g_130190_(_039894_, _039927_, _039930_);
  and g_130191_(_039866_, _039928_, _039931_);
  or g_130192_(_039865_, _039930_, _039932_);
  and g_130193_(_039919_, _039923_, _039933_);
  or g_130194_(_039917_, _039922_, _039934_);
  and g_130195_(_039893_, _039933_, _039935_);
  or g_130196_(_039894_, _039934_, _039936_);
  and g_130197_(_039872_, _039889_, _039937_);
  or g_130198_(_039873_, _039888_, _039938_);
  and g_130199_(_039884_, _039938_, _039939_);
  or g_130200_(_039883_, _039937_, _039941_);
  and g_130201_(_039936_, _039939_, _039942_);
  or g_130202_(_039935_, _039941_, _039943_);
  and g_130203_(_039932_, _039942_, _039944_);
  or g_130204_(_039931_, _039943_, _039945_);
  and g_130205_(_039726_, _039945_, _039946_);
  or g_130206_(_039725_, _039944_, _039947_);
  and g_130207_(_039871_, _039944_, _039948_);
  or g_130208_(_039870_, _039945_, _039949_);
  and g_130209_(_039947_, _039949_, _039950_);
  or g_130210_(_039946_, _039948_, _039952_);
  or g_130211_(out[129], out[128], _039953_);
  or g_130212_(out[128], _036178_, _039954_);
  and g_130213_(out[131], _039954_, _039955_);
  xor g_130214_(out[131], _039954_, _039956_);
  xor g_130215_(_003442_, _039954_, _039957_);
  and g_130216_(_039809_, _039944_, _039958_);
  or g_130217_(_039807_, _039945_, _039959_);
  and g_130218_(_039815_, _039945_, _039960_);
  or g_130219_(_039814_, _039944_, _039961_);
  and g_130220_(_039959_, _039961_, _039963_);
  or g_130221_(_039958_, _039960_, _039964_);
  and g_130222_(_039956_, _039964_, _039965_);
  or g_130223_(_039957_, _039963_, _039966_);
  and g_130224_(_039957_, _039963_, _039967_);
  or g_130225_(_039956_, _039964_, _039968_);
  xor g_130226_(out[130], _039953_, _039969_);
  xor g_130227_(_003431_, _039953_, _039970_);
  and g_130228_(_039790_, _039944_, _039971_);
  or g_130229_(_039791_, _039945_, _039972_);
  and g_130230_(_039798_, _039945_, _039974_);
  or g_130231_(_039796_, _039944_, _039975_);
  and g_130232_(_039972_, _039975_, _039976_);
  or g_130233_(_039971_, _039974_, _039977_);
  and g_130234_(_039969_, _039976_, _039978_);
  or g_130235_(_039970_, _039977_, _039979_);
  and g_130236_(_039968_, _039979_, _039980_);
  or g_130237_(_039967_, _039978_, _039981_);
  and g_130238_(_039966_, _039981_, _039982_);
  or g_130239_(_039965_, _039980_, _039983_);
  xor g_130240_(out[129], out[128], _039985_);
  not g_130241_(_039985_, _039986_);
  and g_130242_(_039785_, _039944_, _039987_);
  or g_130243_(_039787_, _039945_, _039988_);
  and g_130244_(_039782_, _039945_, _039989_);
  or g_130245_(_039781_, _039944_, _039990_);
  and g_130246_(_039988_, _039990_, _039991_);
  or g_130247_(_039987_, _039989_, _039992_);
  and g_130248_(_039985_, _039991_, _039993_);
  or g_130249_(_039986_, _039992_, _039994_);
  and g_130250_(out[112], _039944_, _039996_);
  or g_130251_(_003288_, _039945_, _039997_);
  and g_130252_(_039773_, _039945_, _039998_);
  or g_130253_(_039772_, _039944_, _039999_);
  and g_130254_(_039997_, _039999_, _040000_);
  or g_130255_(_039996_, _039998_, _040001_);
  and g_130256_(_003420_, _040001_, _040002_);
  or g_130257_(out[128], _040000_, _040003_);
  xor g_130258_(_039985_, _039991_, _040004_);
  xor g_130259_(_039986_, _039991_, _040005_);
  and g_130260_(_040003_, _040004_, _040007_);
  or g_130261_(_040002_, _040005_, _040008_);
  and g_130262_(_039994_, _040008_, _040009_);
  or g_130263_(_039993_, _040007_, _040010_);
  and g_130264_(_039970_, _039977_, _040011_);
  or g_130265_(_039969_, _039976_, _040012_);
  and g_130266_(_039966_, _040012_, _040013_);
  or g_130267_(_039965_, _040011_, _040014_);
  and g_130268_(_040010_, _040013_, _040015_);
  or g_130269_(_040009_, _040014_, _040016_);
  and g_130270_(_039983_, _040016_, _040018_);
  or g_130271_(_039982_, _040015_, _040019_);
  and g_130272_(_017084_, _039954_, _040020_);
  and g_130273_(out[133], _040020_, _040021_);
  or g_130274_(out[134], _040021_, _040022_);
  and g_130275_(out[135], _040022_, _040023_);
  and g_130276_(out[136], _040023_, _040024_);
  or g_130277_(out[137], _040024_, _040025_);
  and g_130278_(out[138], _040025_, _040026_);
  xor g_130279_(out[138], _040025_, _040027_);
  xor g_130280_(_003475_, _040025_, _040029_);
  and g_130281_(_039952_, _040027_, _040030_);
  or g_130282_(_039950_, _040029_, _040031_);
  and g_130283_(_039879_, _039881_, _040032_);
  or g_130284_(_039880_, _039882_, _040033_);
  xor g_130285_(out[139], _040026_, _040034_);
  xor g_130286_(_003354_, _040026_, _040035_);
  and g_130287_(_040033_, _040034_, _040036_);
  or g_130288_(_040032_, _040035_, _040037_);
  and g_130289_(_040031_, _040037_, _040038_);
  or g_130290_(_040030_, _040036_, _040040_);
  xor g_130291_(out[136], _040023_, _040041_);
  xor g_130292_(_003453_, _040023_, _040042_);
  and g_130293_(_039903_, _039945_, _040043_);
  or g_130294_(_039902_, _039944_, _040044_);
  and g_130295_(_039897_, _039944_, _040045_);
  or g_130296_(_039895_, _039945_, _040046_);
  and g_130297_(_040044_, _040046_, _040047_);
  or g_130298_(_040043_, _040045_, _040048_);
  and g_130299_(_040041_, _040048_, _040049_);
  or g_130300_(_040042_, _040047_, _040051_);
  xor g_130301_(out[137], _040024_, _040052_);
  xor g_130302_(_003464_, _040024_, _040053_);
  and g_130303_(_039914_, _039945_, _040054_);
  or g_130304_(_039913_, _039944_, _040055_);
  and g_130305_(_039906_, _039944_, _040056_);
  or g_130306_(_039908_, _039945_, _040057_);
  and g_130307_(_040055_, _040057_, _040058_);
  or g_130308_(_040054_, _040056_, _040059_);
  and g_130309_(_040053_, _040059_, _040060_);
  or g_130310_(_040052_, _040058_, _040062_);
  and g_130311_(_040051_, _040062_, _040063_);
  or g_130312_(_040049_, _040060_, _040064_);
  and g_130313_(_039950_, _040029_, _040065_);
  or g_130314_(_039952_, _040027_, _040066_);
  and g_130315_(_040032_, _040035_, _040067_);
  or g_130316_(_040033_, _040034_, _040068_);
  and g_130317_(_040066_, _040068_, _040069_);
  or g_130318_(_040065_, _040067_, _040070_);
  and g_130319_(_040042_, _040047_, _040071_);
  or g_130320_(_040041_, _040048_, _040073_);
  and g_130321_(_040052_, _040058_, _040074_);
  or g_130322_(_040053_, _040059_, _040075_);
  and g_130323_(_040073_, _040075_, _040076_);
  or g_130324_(_040071_, _040074_, _040077_);
  and g_130325_(_040038_, _040069_, _040078_);
  or g_130326_(_040040_, _040070_, _040079_);
  and g_130327_(_040063_, _040076_, _040080_);
  or g_130328_(_040064_, _040077_, _040081_);
  and g_130329_(_040078_, _040080_, _040082_);
  or g_130330_(_040079_, _040081_, _040084_);
  xor g_130331_(out[134], _040021_, _040085_);
  xor g_130332_(_003376_, _040021_, _040086_);
  and g_130333_(_039754_, _039945_, _040087_);
  or g_130334_(_039752_, _039944_, _040088_);
  and g_130335_(_039746_, _039944_, _040089_);
  or g_130336_(_039747_, _039945_, _040090_);
  and g_130337_(_040088_, _040090_, _040091_);
  or g_130338_(_040087_, _040089_, _040092_);
  and g_130339_(_040085_, _040091_, _040093_);
  or g_130340_(_040086_, _040092_, _040095_);
  xor g_130341_(out[135], _040022_, _040096_);
  xor g_130342_(_003365_, _040022_, _040097_);
  and g_130343_(_039743_, _039945_, _040098_);
  or g_130344_(_039741_, _039944_, _040099_);
  and g_130345_(_039736_, _039944_, _040100_);
  or g_130346_(_039735_, _039945_, _040101_);
  and g_130347_(_040099_, _040101_, _040102_);
  or g_130348_(_040098_, _040100_, _040103_);
  and g_130349_(_040097_, _040102_, _040104_);
  or g_130350_(_040096_, _040103_, _040106_);
  and g_130351_(_040095_, _040106_, _040107_);
  or g_130352_(_040093_, _040104_, _040108_);
  xor g_130353_(out[132], _039955_, _040109_);
  xor g_130354_(_003398_, _039955_, _040110_);
  and g_130355_(_039835_, _039945_, _040111_);
  or g_130356_(_039834_, _039944_, _040112_);
  and g_130357_(_039828_, _039944_, _040113_);
  or g_130358_(_039827_, _039945_, _040114_);
  and g_130359_(_040112_, _040114_, _040115_);
  or g_130360_(_040111_, _040113_, _040117_);
  and g_130361_(_040109_, _040117_, _040118_);
  or g_130362_(_040110_, _040115_, _040119_);
  xor g_130363_(out[133], _040020_, _040120_);
  xor g_130364_(_003387_, _040020_, _040121_);
  and g_130365_(_039765_, _039945_, _040122_);
  or g_130366_(_039763_, _039944_, _040123_);
  and g_130367_(_039758_, _039944_, _040124_);
  or g_130368_(_039757_, _039945_, _040125_);
  and g_130369_(_040123_, _040125_, _040126_);
  or g_130370_(_040122_, _040124_, _040128_);
  and g_130371_(_040120_, _040128_, _040129_);
  or g_130372_(_040121_, _040126_, _040130_);
  and g_130373_(_040096_, _040103_, _040131_);
  or g_130374_(_040097_, _040102_, _040132_);
  and g_130375_(_040110_, _040115_, _040133_);
  or g_130376_(_040109_, _040117_, _040134_);
  and g_130377_(_040121_, _040126_, _040135_);
  or g_130378_(_040120_, _040128_, _040136_);
  and g_130379_(_040134_, _040136_, _040137_);
  or g_130380_(_040133_, _040135_, _040139_);
  and g_130381_(_040119_, _040137_, _040140_);
  or g_130382_(_040118_, _040139_, _040141_);
  xor g_130383_(_040085_, _040091_, _040142_);
  xor g_130384_(_040086_, _040091_, _040143_);
  xor g_130385_(_040097_, _040102_, _040144_);
  xor g_130386_(_040096_, _040102_, _040145_);
  and g_130387_(_040142_, _040144_, _040146_);
  or g_130388_(_040143_, _040145_, _040147_);
  and g_130389_(_040130_, _040146_, _040148_);
  or g_130390_(_040129_, _040147_, _040150_);
  and g_130391_(_040140_, _040148_, _040151_);
  or g_130392_(_040141_, _040150_, _040152_);
  and g_130393_(_040082_, _040151_, _040153_);
  or g_130394_(_040084_, _040152_, _040154_);
  and g_130395_(_040019_, _040153_, _040155_);
  or g_130396_(_040018_, _040154_, _040156_);
  and g_130397_(_040108_, _040132_, _040157_);
  or g_130398_(_040107_, _040131_, _040158_);
  and g_130399_(_040139_, _040146_, _040159_);
  or g_130400_(_040137_, _040147_, _040161_);
  and g_130401_(_040130_, _040159_, _040162_);
  or g_130402_(_040129_, _040161_, _040163_);
  and g_130403_(_040158_, _040163_, _040164_);
  or g_130404_(_040157_, _040162_, _040165_);
  and g_130405_(_040082_, _040165_, _040166_);
  or g_130406_(_040084_, _040164_, _040167_);
  and g_130407_(_040031_, _040062_, _040168_);
  or g_130408_(_040030_, _040060_, _040169_);
  and g_130409_(_040077_, _040168_, _040170_);
  or g_130410_(_040076_, _040169_, _040172_);
  and g_130411_(_040069_, _040172_, _040173_);
  or g_130412_(_040070_, _040170_, _040174_);
  and g_130413_(_040037_, _040174_, _040175_);
  or g_130414_(_040036_, _040173_, _040176_);
  and g_130415_(_040167_, _040176_, _040177_);
  or g_130416_(_040166_, _040175_, _040178_);
  and g_130417_(_040156_, _040177_, _040179_);
  or g_130418_(_040155_, _040178_, _040180_);
  and g_130419_(out[128], _040000_, _040181_);
  or g_130420_(_003420_, _040001_, _040183_);
  and g_130421_(_039980_, _040013_, _040184_);
  or g_130422_(_039981_, _040014_, _040185_);
  and g_130423_(_040183_, _040184_, _040186_);
  or g_130424_(_040181_, _040185_, _040187_);
  and g_130425_(_040007_, _040186_, _040188_);
  or g_130426_(_040008_, _040187_, _040189_);
  and g_130427_(_040153_, _040188_, _040190_);
  or g_130428_(_040154_, _040189_, _040191_);
  and g_130429_(_040180_, _040191_, _040192_);
  or g_130430_(_040179_, _040190_, _040194_);
  and g_130431_(_039952_, _040194_, _040195_);
  or g_130432_(_039950_, _040192_, _040196_);
  and g_130433_(_040029_, _040192_, _040197_);
  or g_130434_(_040027_, _040194_, _040198_);
  and g_130435_(_040196_, _040198_, _040199_);
  or g_130436_(_040195_, _040197_, _040200_);
  or g_130437_(out[145], out[144], _040201_);
  or g_130438_(out[144], _038455_, _040202_);
  and g_130439_(out[147], _040202_, _040203_);
  and g_130440_(_017316_, _040202_, _040205_);
  and g_130441_(out[149], _040205_, _040206_);
  or g_130442_(out[150], _040206_, _040207_);
  and g_130443_(out[151], _040207_, _040208_);
  xor g_130444_(out[151], _040207_, _040209_);
  xor g_130445_(_003497_, _040207_, _040210_);
  and g_130446_(_040103_, _040194_, _040211_);
  or g_130447_(_040102_, _040192_, _040212_);
  and g_130448_(_040097_, _040192_, _040213_);
  or g_130449_(_040096_, _040194_, _040214_);
  and g_130450_(_040212_, _040214_, _040216_);
  or g_130451_(_040211_, _040213_, _040217_);
  and g_130452_(_040209_, _040217_, _040218_);
  or g_130453_(_040210_, _040216_, _040219_);
  xor g_130454_(out[150], _040206_, _040220_);
  xor g_130455_(_003508_, _040206_, _040221_);
  and g_130456_(_040092_, _040194_, _040222_);
  or g_130457_(_040091_, _040192_, _040223_);
  and g_130458_(_040085_, _040192_, _040224_);
  or g_130459_(_040086_, _040194_, _040225_);
  and g_130460_(_040223_, _040225_, _040227_);
  or g_130461_(_040222_, _040224_, _040228_);
  and g_130462_(_040221_, _040228_, _040229_);
  or g_130463_(_040220_, _040227_, _040230_);
  xor g_130464_(out[149], _040205_, _040231_);
  xor g_130465_(_003519_, _040205_, _040232_);
  and g_130466_(_040128_, _040194_, _040233_);
  or g_130467_(_040126_, _040192_, _040234_);
  and g_130468_(_040121_, _040192_, _040235_);
  or g_130469_(_040120_, _040194_, _040236_);
  and g_130470_(_040234_, _040236_, _040238_);
  or g_130471_(_040233_, _040235_, _040239_);
  and g_130472_(_040232_, _040238_, _040240_);
  or g_130473_(_040231_, _040239_, _040241_);
  and g_130474_(out[128], _040192_, _040242_);
  or g_130475_(_003420_, _040194_, _040243_);
  and g_130476_(_040001_, _040194_, _040244_);
  or g_130477_(_040000_, _040192_, _040245_);
  and g_130478_(_040243_, _040245_, _040246_);
  or g_130479_(_040242_, _040244_, _040247_);
  and g_130480_(out[144], _040246_, _040249_);
  or g_130481_(_003552_, _040247_, _040250_);
  and g_130482_(_039992_, _040194_, _040251_);
  or g_130483_(_039991_, _040192_, _040252_);
  and g_130484_(_039985_, _040192_, _040253_);
  or g_130485_(_039986_, _040194_, _040254_);
  and g_130486_(_040252_, _040254_, _040255_);
  or g_130487_(_040251_, _040253_, _040256_);
  and g_130488_(out[145], _040256_, _040257_);
  or g_130489_(_003541_, _040255_, _040258_);
  xor g_130490_(out[145], out[144], _040260_);
  xor g_130491_(_003541_, out[144], _040261_);
  and g_130492_(_040249_, _040258_, _040262_);
  or g_130493_(_040250_, _040257_, _040263_);
  xor g_130494_(out[146], _040201_, _040264_);
  xor g_130495_(_003563_, _040201_, _040265_);
  and g_130496_(_039969_, _040192_, _040266_);
  or g_130497_(_039970_, _040194_, _040267_);
  and g_130498_(_039977_, _040194_, _040268_);
  or g_130499_(_039976_, _040192_, _040269_);
  and g_130500_(_040267_, _040269_, _040271_);
  or g_130501_(_040266_, _040268_, _040272_);
  and g_130502_(_040264_, _040271_, _040273_);
  or g_130503_(_040265_, _040272_, _040274_);
  and g_130504_(_040255_, _040260_, _040275_);
  or g_130505_(_040256_, _040261_, _040276_);
  and g_130506_(_040274_, _040276_, _040277_);
  or g_130507_(_040273_, _040275_, _040278_);
  and g_130508_(_040263_, _040277_, _040279_);
  or g_130509_(_040262_, _040278_, _040280_);
  xor g_130510_(out[147], _040202_, _040282_);
  xor g_130511_(_003574_, _040202_, _040283_);
  and g_130512_(_039957_, _040192_, _040284_);
  or g_130513_(_039956_, _040194_, _040285_);
  and g_130514_(_039964_, _040194_, _040286_);
  or g_130515_(_039963_, _040192_, _040287_);
  and g_130516_(_040285_, _040287_, _040288_);
  or g_130517_(_040284_, _040286_, _040289_);
  and g_130518_(_040282_, _040289_, _040290_);
  or g_130519_(_040283_, _040288_, _040291_);
  and g_130520_(_040265_, _040272_, _040293_);
  or g_130521_(_040264_, _040271_, _040294_);
  and g_130522_(_040291_, _040294_, _040295_);
  or g_130523_(_040290_, _040293_, _040296_);
  and g_130524_(_040280_, _040295_, _040297_);
  or g_130525_(_040279_, _040296_, _040298_);
  xor g_130526_(out[148], _040203_, _040299_);
  xor g_130527_(_003530_, _040203_, _040300_);
  and g_130528_(_040117_, _040194_, _040301_);
  or g_130529_(_040115_, _040192_, _040302_);
  and g_130530_(_040110_, _040192_, _040304_);
  or g_130531_(_040109_, _040194_, _040305_);
  and g_130532_(_040302_, _040305_, _040306_);
  or g_130533_(_040301_, _040304_, _040307_);
  and g_130534_(_040300_, _040306_, _040308_);
  or g_130535_(_040299_, _040307_, _040309_);
  and g_130536_(_040283_, _040288_, _040310_);
  or g_130537_(_040282_, _040289_, _040311_);
  and g_130538_(_040309_, _040311_, _040312_);
  or g_130539_(_040308_, _040310_, _040313_);
  and g_130540_(_040298_, _040312_, _040315_);
  or g_130541_(_040297_, _040313_, _040316_);
  and g_130542_(_040231_, _040239_, _040317_);
  or g_130543_(_040232_, _040238_, _040318_);
  and g_130544_(_040299_, _040307_, _040319_);
  or g_130545_(_040300_, _040306_, _040320_);
  and g_130546_(_040318_, _040320_, _040321_);
  or g_130547_(_040317_, _040319_, _040322_);
  and g_130548_(_040316_, _040321_, _040323_);
  or g_130549_(_040315_, _040322_, _040324_);
  and g_130550_(_040241_, _040324_, _040326_);
  or g_130551_(_040240_, _040323_, _040327_);
  and g_130552_(_040230_, _040327_, _040328_);
  or g_130553_(_040229_, _040326_, _040329_);
  and g_130554_(_040210_, _040216_, _040330_);
  or g_130555_(_040209_, _040217_, _040331_);
  and g_130556_(_040220_, _040227_, _040332_);
  or g_130557_(_040221_, _040228_, _040333_);
  and g_130558_(_040331_, _040333_, _040334_);
  or g_130559_(_040330_, _040332_, _040335_);
  and g_130560_(_040329_, _040334_, _040337_);
  or g_130561_(_040328_, _040335_, _040338_);
  and g_130562_(_040219_, _040338_, _040339_);
  or g_130563_(_040218_, _040337_, _040340_);
  and g_130564_(out[152], _040208_, _040341_);
  or g_130565_(out[153], _040341_, _040342_);
  and g_130566_(out[154], _040342_, _040343_);
  xor g_130567_(out[154], _040342_, _040344_);
  not g_130568_(_040344_, _040345_);
  and g_130569_(_040200_, _040344_, _040346_);
  or g_130570_(_040199_, _040345_, _040348_);
  xor g_130571_(out[155], _040343_, _040349_);
  xor g_130572_(_003486_, _040343_, _040350_);
  or g_130573_(_040034_, _040194_, _040351_);
  or g_130574_(_040032_, _040192_, _040352_);
  and g_130575_(_040351_, _040352_, _040353_);
  and g_130576_(_040032_, _040194_, _040354_);
  or g_130577_(_040033_, _040192_, _040355_);
  and g_130578_(_040034_, _040192_, _040356_);
  or g_130579_(_040035_, _040194_, _040357_);
  and g_130580_(_040355_, _040357_, _040359_);
  or g_130581_(_040354_, _040356_, _040360_);
  and g_130582_(_040349_, _040359_, _040361_);
  or g_130583_(_040350_, _040360_, _040362_);
  or g_130584_(_040346_, _040361_, _040363_);
  and g_130585_(_040199_, _040345_, _040364_);
  and g_130586_(_040350_, _040353_, _040365_);
  or g_130587_(_040364_, _040365_, _040366_);
  xor g_130588_(_040200_, _040344_, _040367_);
  or g_130589_(_040349_, _040359_, _040368_);
  and g_130590_(_040362_, _040368_, _040370_);
  and g_130591_(_040367_, _040370_, _040371_);
  or g_130592_(_040363_, _040366_, _040372_);
  xor g_130593_(out[153], _040341_, _040373_);
  xor g_130594_(_003596_, _040341_, _040374_);
  and g_130595_(_040059_, _040194_, _040375_);
  or g_130596_(_040058_, _040192_, _040376_);
  and g_130597_(_040052_, _040192_, _040377_);
  or g_130598_(_040053_, _040194_, _040378_);
  and g_130599_(_040376_, _040378_, _040379_);
  or g_130600_(_040375_, _040377_, _040381_);
  and g_130601_(_040374_, _040381_, _040382_);
  or g_130602_(_040373_, _040379_, _040383_);
  xor g_130603_(out[152], _040208_, _040384_);
  xor g_130604_(_003585_, _040208_, _040385_);
  and g_130605_(_040048_, _040194_, _040386_);
  or g_130606_(_040047_, _040192_, _040387_);
  and g_130607_(_040042_, _040192_, _040388_);
  or g_130608_(_040041_, _040194_, _040389_);
  and g_130609_(_040387_, _040389_, _040390_);
  or g_130610_(_040386_, _040388_, _040392_);
  and g_130611_(_040384_, _040392_, _040393_);
  or g_130612_(_040385_, _040390_, _040394_);
  and g_130613_(_040383_, _040394_, _040395_);
  or g_130614_(_040382_, _040393_, _040396_);
  and g_130615_(_040373_, _040379_, _040397_);
  or g_130616_(_040374_, _040381_, _040398_);
  and g_130617_(_040385_, _040390_, _040399_);
  or g_130618_(_040384_, _040392_, _040400_);
  and g_130619_(_040398_, _040400_, _040401_);
  or g_130620_(_040397_, _040399_, _040403_);
  and g_130621_(_040395_, _040401_, _040404_);
  or g_130622_(_040396_, _040403_, _040405_);
  and g_130623_(_040371_, _040404_, _040406_);
  or g_130624_(_040372_, _040405_, _040407_);
  and g_130625_(_040340_, _040406_, _040408_);
  or g_130626_(_040339_, _040407_, _040409_);
  and g_130627_(_040396_, _040398_, _040410_);
  or g_130628_(_040395_, _040397_, _040411_);
  and g_130629_(_040371_, _040410_, _040412_);
  or g_130630_(_040372_, _040411_, _040414_);
  and g_130631_(_040346_, _040368_, _040415_);
  or g_130632_(_040348_, _040365_, _040416_);
  and g_130633_(_040362_, _040416_, _040417_);
  or g_130634_(_040361_, _040415_, _040418_);
  and g_130635_(_040414_, _040417_, _040419_);
  or g_130636_(_040412_, _040418_, _040420_);
  and g_130637_(_040409_, _040419_, _040421_);
  or g_130638_(_040408_, _040420_, _040422_);
  and g_130639_(_040200_, _040422_, _040423_);
  not g_130640_(_040423_, _040425_);
  or g_130641_(_040344_, _040422_, _040426_);
  not g_130642_(_040426_, _040427_);
  and g_130643_(_040425_, _040426_, _040428_);
  or g_130644_(_040423_, _040427_, _040429_);
  or g_130645_(out[161], out[160], _040430_);
  or g_130646_(out[160], _040556_, _040431_);
  and g_130647_(out[163], _040431_, _040432_);
  and g_130648_(_017527_, _040431_, _040433_);
  and g_130649_(out[165], _040433_, _040434_);
  or g_130650_(out[166], _040434_, _040436_);
  and g_130651_(out[167], _040436_, _040437_);
  and g_130652_(out[168], _040437_, _040438_);
  or g_130653_(out[169], _040438_, _040439_);
  and g_130654_(out[170], _040439_, _040440_);
  xor g_130655_(out[171], _040440_, _040441_);
  xor g_130656_(_003618_, _040440_, _040442_);
  and g_130657_(_040349_, _040353_, _040443_);
  xor g_130658_(out[170], _040439_, _040444_);
  xor g_130659_(_003739_, _040439_, _040445_);
  and g_130660_(_040429_, _040444_, _040447_);
  or g_130661_(_040428_, _040445_, _040448_);
  and g_130662_(_040349_, _040360_, _040449_);
  or g_130663_(_040350_, _040359_, _040450_);
  and g_130664_(_040441_, _040450_, _040451_);
  or g_130665_(_040442_, _040449_, _040452_);
  and g_130666_(_040448_, _040452_, _040453_);
  or g_130667_(_040447_, _040451_, _040454_);
  and g_130668_(_040428_, _040445_, _040455_);
  or g_130669_(_040429_, _040444_, _040456_);
  xor g_130670_(out[169], _040438_, _040458_);
  xor g_130671_(_003728_, _040438_, _040459_);
  and g_130672_(_040381_, _040422_, _040460_);
  not g_130673_(_040460_, _040461_);
  or g_130674_(_040374_, _040422_, _040462_);
  not g_130675_(_040462_, _040463_);
  and g_130676_(_040461_, _040462_, _040464_);
  or g_130677_(_040460_, _040463_, _040465_);
  and g_130678_(_040458_, _040464_, _040466_);
  or g_130679_(_040459_, _040465_, _040467_);
  xor g_130680_(out[168], _040437_, _040469_);
  xor g_130681_(_003717_, _040437_, _040470_);
  and g_130682_(_040392_, _040422_, _040471_);
  not g_130683_(_040471_, _040472_);
  or g_130684_(_040384_, _040422_, _040473_);
  not g_130685_(_040473_, _040474_);
  and g_130686_(_040472_, _040473_, _040475_);
  or g_130687_(_040471_, _040474_, _040476_);
  and g_130688_(_040469_, _040476_, _040477_);
  or g_130689_(_040470_, _040475_, _040478_);
  and g_130690_(_040459_, _040465_, _040480_);
  or g_130691_(_040458_, _040464_, _040481_);
  and g_130692_(_040478_, _040481_, _040482_);
  or g_130693_(_040477_, _040480_, _040483_);
  and g_130694_(_040467_, _040483_, _040484_);
  or g_130695_(_040466_, _040482_, _040485_);
  xor g_130696_(out[162], _040430_, _040486_);
  xor g_130697_(_003695_, _040430_, _040487_);
  and g_130698_(_040272_, _040422_, _040488_);
  not g_130699_(_040488_, _040489_);
  or g_130700_(_040265_, _040422_, _040491_);
  not g_130701_(_040491_, _040492_);
  and g_130702_(_040489_, _040491_, _040493_);
  or g_130703_(_040488_, _040492_, _040494_);
  and g_130704_(_040486_, _040493_, _040495_);
  or g_130705_(_040487_, _040494_, _040496_);
  and g_130706_(_040260_, _040421_, _040497_);
  or g_130707_(_040261_, _040422_, _040498_);
  and g_130708_(_040256_, _040422_, _040499_);
  or g_130709_(_040255_, _040421_, _040500_);
  and g_130710_(_040498_, _040500_, _040502_);
  or g_130711_(_040497_, _040499_, _040503_);
  and g_130712_(out[161], _040503_, _040504_);
  not g_130713_(_040504_, _040505_);
  xor g_130714_(out[161], out[160], _040506_);
  xor g_130715_(_003673_, out[160], _040507_);
  and g_130716_(_040502_, _040506_, _040508_);
  or g_130717_(_040503_, _040507_, _040509_);
  and g_130718_(out[144], _040421_, _040510_);
  or g_130719_(_003552_, _040422_, _040511_);
  and g_130720_(_040247_, _040422_, _040513_);
  or g_130721_(_040246_, _040421_, _040514_);
  and g_130722_(_040511_, _040514_, _040515_);
  or g_130723_(_040510_, _040513_, _040516_);
  and g_130724_(out[160], _040515_, _040517_);
  or g_130725_(_003684_, _040516_, _040518_);
  and g_130726_(_040509_, _040518_, _040519_);
  or g_130727_(_040508_, _040517_, _040520_);
  and g_130728_(_040505_, _040520_, _040521_);
  or g_130729_(_040504_, _040519_, _040522_);
  and g_130730_(_040496_, _040522_, _040524_);
  or g_130731_(_040495_, _040521_, _040525_);
  and g_130732_(_040487_, _040494_, _040526_);
  or g_130733_(_040486_, _040493_, _040527_);
  xor g_130734_(out[163], _040431_, _040528_);
  xor g_130735_(_003706_, _040431_, _040529_);
  or g_130736_(_040282_, _040422_, _040530_);
  not g_130737_(_040530_, _040531_);
  and g_130738_(_040289_, _040422_, _040532_);
  not g_130739_(_040532_, _040533_);
  and g_130740_(_040530_, _040533_, _040535_);
  or g_130741_(_040531_, _040532_, _040536_);
  and g_130742_(_040528_, _040536_, _040537_);
  or g_130743_(_040529_, _040535_, _040538_);
  and g_130744_(_040527_, _040538_, _040539_);
  or g_130745_(_040526_, _040537_, _040540_);
  and g_130746_(_040525_, _040539_, _040541_);
  or g_130747_(_040524_, _040540_, _040542_);
  xor g_130748_(out[164], _040432_, _040543_);
  xor g_130749_(_003662_, _040432_, _040544_);
  or g_130750_(_040299_, _040422_, _040546_);
  not g_130751_(_040546_, _040547_);
  and g_130752_(_040307_, _040422_, _040548_);
  not g_130753_(_040548_, _040549_);
  and g_130754_(_040546_, _040549_, _040550_);
  or g_130755_(_040547_, _040548_, _040551_);
  and g_130756_(_040544_, _040550_, _040552_);
  or g_130757_(_040543_, _040551_, _040553_);
  and g_130758_(_040529_, _040535_, _040554_);
  or g_130759_(_040528_, _040536_, _040555_);
  and g_130760_(_040553_, _040555_, _040557_);
  or g_130761_(_040552_, _040554_, _040558_);
  and g_130762_(_040542_, _040557_, _040559_);
  or g_130763_(_040541_, _040558_, _040560_);
  xor g_130764_(out[165], _040433_, _040561_);
  xor g_130765_(_003651_, _040433_, _040562_);
  and g_130766_(_040239_, _040422_, _040563_);
  not g_130767_(_040563_, _040564_);
  or g_130768_(_040231_, _040422_, _040565_);
  not g_130769_(_040565_, _040566_);
  and g_130770_(_040564_, _040565_, _040568_);
  or g_130771_(_040563_, _040566_, _040569_);
  and g_130772_(_040561_, _040569_, _040570_);
  or g_130773_(_040562_, _040568_, _040571_);
  and g_130774_(_040543_, _040551_, _040572_);
  or g_130775_(_040544_, _040550_, _040573_);
  and g_130776_(_040571_, _040573_, _040574_);
  or g_130777_(_040570_, _040572_, _040575_);
  and g_130778_(_040560_, _040574_, _040576_);
  or g_130779_(_040559_, _040575_, _040577_);
  xor g_130780_(out[166], _040434_, _040579_);
  xor g_130781_(_003640_, _040434_, _040580_);
  and g_130782_(_040228_, _040422_, _040581_);
  not g_130783_(_040581_, _040582_);
  or g_130784_(_040221_, _040422_, _040583_);
  not g_130785_(_040583_, _040584_);
  and g_130786_(_040582_, _040583_, _040585_);
  or g_130787_(_040581_, _040584_, _040586_);
  and g_130788_(_040579_, _040585_, _040587_);
  or g_130789_(_040580_, _040586_, _040588_);
  and g_130790_(_040562_, _040568_, _040590_);
  or g_130791_(_040561_, _040569_, _040591_);
  and g_130792_(_040588_, _040591_, _040592_);
  or g_130793_(_040587_, _040590_, _040593_);
  and g_130794_(_040577_, _040592_, _040594_);
  or g_130795_(_040576_, _040593_, _040595_);
  xor g_130796_(out[167], _040436_, _040596_);
  xor g_130797_(_003629_, _040436_, _040597_);
  and g_130798_(_040217_, _040422_, _040598_);
  not g_130799_(_040598_, _040599_);
  or g_130800_(_040209_, _040422_, _040601_);
  not g_130801_(_040601_, _040602_);
  and g_130802_(_040599_, _040601_, _040603_);
  or g_130803_(_040598_, _040602_, _040604_);
  and g_130804_(_040596_, _040604_, _040605_);
  or g_130805_(_040597_, _040603_, _040606_);
  and g_130806_(_040580_, _040586_, _040607_);
  or g_130807_(_040579_, _040585_, _040608_);
  and g_130808_(_040606_, _040608_, _040609_);
  or g_130809_(_040605_, _040607_, _040610_);
  and g_130810_(_040595_, _040609_, _040612_);
  or g_130811_(_040594_, _040610_, _040613_);
  and g_130812_(_040467_, _040481_, _040614_);
  or g_130813_(_040466_, _040480_, _040615_);
  and g_130814_(_040597_, _040603_, _040616_);
  or g_130815_(_040596_, _040604_, _040617_);
  and g_130816_(_040470_, _040475_, _040618_);
  or g_130817_(_040469_, _040476_, _040619_);
  and g_130818_(_040442_, _040449_, _040620_);
  or g_130819_(_040441_, _040450_, _040621_);
  and g_130820_(_040454_, _040621_, _040623_);
  or g_130821_(_040453_, _040620_, _040624_);
  and g_130822_(_040617_, _040619_, _040625_);
  or g_130823_(_040616_, _040618_, _040626_);
  and g_130824_(_040614_, _040625_, _040627_);
  or g_130825_(_040615_, _040626_, _040628_);
  and g_130826_(_040456_, _040621_, _040629_);
  or g_130827_(_040455_, _040620_, _040630_);
  and g_130828_(_040453_, _040629_, _040631_);
  or g_130829_(_040454_, _040630_, _040632_);
  and g_130830_(_040627_, _040631_, _040634_);
  or g_130831_(_040628_, _040632_, _040635_);
  and g_130832_(_040478_, _040634_, _040636_);
  or g_130833_(_040477_, _040635_, _040637_);
  and g_130834_(_040613_, _040636_, _040638_);
  or g_130835_(_040612_, _040637_, _040639_);
  and g_130836_(_040484_, _040629_, _040640_);
  or g_130837_(_040485_, _040630_, _040641_);
  and g_130838_(_040639_, _040641_, _040642_);
  or g_130839_(_040638_, _040640_, _040643_);
  or g_130840_(_040623_, _040643_, _040645_);
  and g_130841_(_040624_, _040642_, _040646_);
  and g_130842_(_040429_, _040645_, _040647_);
  not g_130843_(_040647_, _040648_);
  or g_130844_(_040444_, _040645_, _040649_);
  not g_130845_(_040649_, _040650_);
  and g_130846_(_040648_, _040649_, _040651_);
  or g_130847_(_040647_, _040650_, _040652_);
  and g_130848_(out[183], _038385_, _040653_);
  and g_130849_(out[184], _040653_, _040654_);
  or g_130850_(out[185], _040654_, _040656_);
  and g_130851_(out[186], _040656_, _040657_);
  xor g_130852_(out[186], _040656_, _040658_);
  not g_130853_(_040658_, _040659_);
  and g_130854_(_040652_, _040658_, _040660_);
  or g_130855_(_040651_, _040659_, _040661_);
  xor g_130856_(out[187], _040657_, _040662_);
  xor g_130857_(_003750_, _040657_, _040663_);
  and g_130858_(_040441_, _040443_, _040664_);
  or g_130859_(_040442_, _040450_, _040665_);
  and g_130860_(_040662_, _040665_, _040667_);
  or g_130861_(_040663_, _040664_, _040668_);
  and g_130862_(_040661_, _040668_, _040669_);
  xor g_130863_(out[184], _040653_, _040670_);
  and g_130864_(_040476_, _040645_, _040671_);
  not g_130865_(_040671_, _040672_);
  or g_130866_(_040469_, _040645_, _040673_);
  not g_130867_(_040673_, _040674_);
  and g_130868_(_040672_, _040673_, _040675_);
  or g_130869_(_040671_, _040674_, _040676_);
  and g_130870_(_040670_, _040676_, _040678_);
  not g_130871_(_040678_, _040679_);
  xor g_130872_(_003860_, _040654_, _040680_);
  and g_130873_(_040465_, _040645_, _040681_);
  not g_130874_(_040681_, _040682_);
  and g_130875_(_040458_, _040646_, _040683_);
  or g_130876_(_040459_, _040645_, _040684_);
  and g_130877_(_040682_, _040684_, _040685_);
  or g_130878_(_040681_, _040683_, _040686_);
  and g_130879_(_040680_, _040686_, _040687_);
  not g_130880_(_040687_, _040689_);
  or g_130881_(_040678_, _040687_, _040690_);
  xor g_130882_(out[178], _038380_, _040691_);
  xor g_130883_(_003827_, _038380_, _040692_);
  and g_130884_(_040486_, _040646_, _040693_);
  or g_130885_(_040487_, _040645_, _040694_);
  and g_130886_(_040494_, _040645_, _040695_);
  or g_130887_(_040493_, _040646_, _040696_);
  and g_130888_(_040694_, _040696_, _040697_);
  or g_130889_(_040693_, _040695_, _040698_);
  and g_130890_(_040691_, _040697_, _040700_);
  or g_130891_(_040692_, _040698_, _040701_);
  and g_130892_(_040506_, _040646_, _040702_);
  or g_130893_(_040507_, _040645_, _040703_);
  and g_130894_(_040503_, _040645_, _040704_);
  or g_130895_(_040502_, _040646_, _040705_);
  and g_130896_(_040703_, _040705_, _040706_);
  or g_130897_(_040702_, _040704_, _040707_);
  and g_130898_(out[177], _040707_, _040708_);
  not g_130899_(_040708_, _040709_);
  xor g_130900_(out[177], out[176], _040711_);
  xor g_130901_(_003805_, out[176], _040712_);
  and g_130902_(_040706_, _040711_, _040713_);
  or g_130903_(_040707_, _040712_, _040714_);
  and g_130904_(_040516_, _040645_, _040715_);
  or g_130905_(_040515_, _040646_, _040716_);
  and g_130906_(out[160], _040646_, _040717_);
  or g_130907_(_003684_, _040645_, _040718_);
  and g_130908_(_040716_, _040718_, _040719_);
  or g_130909_(_040715_, _040717_, _040720_);
  and g_130910_(out[176], _040719_, _040722_);
  or g_130911_(_003816_, _040720_, _040723_);
  and g_130912_(_040714_, _040723_, _040724_);
  or g_130913_(_040713_, _040722_, _040725_);
  and g_130914_(_040709_, _040725_, _040726_);
  or g_130915_(_040708_, _040724_, _040727_);
  and g_130916_(_040701_, _040727_, _040728_);
  or g_130917_(_040700_, _040726_, _040729_);
  and g_130918_(_040692_, _040698_, _040730_);
  or g_130919_(_040691_, _040697_, _040731_);
  xor g_130920_(out[179], _038381_, _040733_);
  xor g_130921_(_003838_, _038381_, _040734_);
  and g_130922_(_040529_, _040646_, _040735_);
  or g_130923_(_040528_, _040645_, _040736_);
  and g_130924_(_040536_, _040645_, _040737_);
  or g_130925_(_040535_, _040646_, _040738_);
  and g_130926_(_040736_, _040738_, _040739_);
  or g_130927_(_040735_, _040737_, _040740_);
  and g_130928_(_040733_, _040740_, _040741_);
  or g_130929_(_040734_, _040739_, _040742_);
  and g_130930_(_040731_, _040742_, _040744_);
  or g_130931_(_040730_, _040741_, _040745_);
  and g_130932_(_040729_, _040744_, _040746_);
  or g_130933_(_040728_, _040745_, _040747_);
  xor g_130934_(out[180], _038382_, _040748_);
  xor g_130935_(_003794_, _038382_, _040749_);
  or g_130936_(_040543_, _040645_, _040750_);
  not g_130937_(_040750_, _040751_);
  and g_130938_(_040551_, _040645_, _040752_);
  not g_130939_(_040752_, _040753_);
  and g_130940_(_040750_, _040753_, _040755_);
  or g_130941_(_040751_, _040752_, _040756_);
  and g_130942_(_040749_, _040755_, _040757_);
  or g_130943_(_040748_, _040756_, _040758_);
  and g_130944_(_040734_, _040739_, _040759_);
  or g_130945_(_040733_, _040740_, _040760_);
  and g_130946_(_040758_, _040760_, _040761_);
  or g_130947_(_040757_, _040759_, _040762_);
  and g_130948_(_040747_, _040761_, _040763_);
  or g_130949_(_040746_, _040762_, _040764_);
  xor g_130950_(out[181], _038383_, _040766_);
  xor g_130951_(_003783_, _038383_, _040767_);
  or g_130952_(_040561_, _040645_, _040768_);
  not g_130953_(_040768_, _040769_);
  and g_130954_(_040569_, _040645_, _040770_);
  not g_130955_(_040770_, _040771_);
  and g_130956_(_040768_, _040771_, _040772_);
  or g_130957_(_040769_, _040770_, _040773_);
  and g_130958_(_040766_, _040773_, _040774_);
  or g_130959_(_040767_, _040772_, _040775_);
  and g_130960_(_040748_, _040756_, _040777_);
  or g_130961_(_040749_, _040755_, _040778_);
  and g_130962_(_040775_, _040778_, _040779_);
  or g_130963_(_040774_, _040777_, _040780_);
  and g_130964_(_040764_, _040779_, _040781_);
  or g_130965_(_040763_, _040780_, _040782_);
  and g_130966_(_040586_, _040645_, _040783_);
  not g_130967_(_040783_, _040784_);
  and g_130968_(_040579_, _040646_, _040785_);
  or g_130969_(_040580_, _040645_, _040786_);
  and g_130970_(_040784_, _040786_, _040788_);
  or g_130971_(_040783_, _040785_, _040789_);
  and g_130972_(_038386_, _040788_, _040790_);
  or g_130973_(_038387_, _040789_, _040791_);
  and g_130974_(_040767_, _040772_, _040792_);
  or g_130975_(_040766_, _040773_, _040793_);
  and g_130976_(_040791_, _040793_, _040794_);
  or g_130977_(_040790_, _040792_, _040795_);
  and g_130978_(_040782_, _040794_, _040796_);
  or g_130979_(_040781_, _040795_, _040797_);
  xor g_130980_(out[183], _038385_, _040799_);
  not g_130981_(_040799_, _040800_);
  and g_130982_(_040604_, _040645_, _040801_);
  not g_130983_(_040801_, _040802_);
  or g_130984_(_040596_, _040645_, _040803_);
  not g_130985_(_040803_, _040804_);
  and g_130986_(_040802_, _040803_, _040805_);
  or g_130987_(_040801_, _040804_, _040806_);
  and g_130988_(_040799_, _040806_, _040807_);
  or g_130989_(_040800_, _040805_, _040808_);
  and g_130990_(_038387_, _040789_, _040810_);
  or g_130991_(_038386_, _040788_, _040811_);
  and g_130992_(_040808_, _040811_, _040812_);
  or g_130993_(_040807_, _040810_, _040813_);
  and g_130994_(_040797_, _040812_, _040814_);
  or g_130995_(_040796_, _040813_, _040815_);
  or g_130996_(_040670_, _040676_, _040816_);
  or g_130997_(_040799_, _040806_, _040817_);
  or g_130998_(_040652_, _040658_, _040818_);
  or g_130999_(_040680_, _040686_, _040819_);
  or g_131000_(_040662_, _040665_, _040821_);
  and g_131001_(_040818_, _040821_, _040822_);
  and g_131002_(_040669_, _040822_, _040823_);
  and g_131003_(_040690_, _040819_, _040824_);
  and g_131004_(_040816_, _040819_, _040825_);
  and g_131005_(_040689_, _040817_, _040826_);
  and g_131006_(_040825_, _040826_, _040827_);
  and g_131007_(_040823_, _040827_, _040828_);
  not g_131008_(_040828_, _040829_);
  and g_131009_(_040679_, _040828_, _040830_);
  or g_131010_(_040678_, _040829_, _040832_);
  and g_131011_(_040815_, _040830_, _040833_);
  or g_131012_(_040814_, _040832_, _040834_);
  and g_131013_(_040823_, _040824_, _040835_);
  and g_131014_(_040660_, _040821_, _040836_);
  or g_131015_(_040835_, _040836_, _040837_);
  or g_131016_(_040667_, _040837_, _040838_);
  not g_131017_(_040838_, _040839_);
  and g_131018_(_040834_, _040839_, _040840_);
  or g_131019_(_040833_, _040838_, _040841_);
  or g_131020_(_038387_, _040841_, _040843_);
  not g_131021_(_040843_, _040844_);
  and g_131022_(_040789_, _040841_, _040845_);
  not g_131023_(_040845_, _040846_);
  and g_131024_(_040843_, _040846_, _040847_);
  or g_131025_(_040844_, _040845_, _040848_);
  or g_131026_(out[193], out[192], _040849_);
  or g_131027_(out[192], _044516_, _040850_);
  and g_131028_(out[195], _040850_, _040851_);
  and g_131029_(_017968_, _040850_, _040852_);
  and g_131030_(out[197], _040852_, _040854_);
  or g_131031_(out[198], _040854_, _040855_);
  and g_131032_(out[199], _040855_, _040856_);
  and g_131033_(out[200], _040856_, _040857_);
  or g_131034_(out[201], _040857_, _040858_);
  not g_131035_(_040858_, _040859_);
  and g_131036_(out[202], _040858_, _040860_);
  xor g_131037_(out[202], _040858_, _040861_);
  xor g_131038_(out[202], _040859_, _040862_);
  and g_131039_(_040659_, _040840_, _040863_);
  or g_131040_(_040658_, _040841_, _040865_);
  and g_131041_(_040652_, _040841_, _040866_);
  or g_131042_(_040651_, _040840_, _040867_);
  and g_131043_(_040865_, _040867_, _040868_);
  or g_131044_(_040863_, _040866_, _040869_);
  and g_131045_(_040862_, _040868_, _040870_);
  or g_131046_(_040861_, _040869_, _040871_);
  xor g_131047_(out[203], _040860_, _040872_);
  xor g_131048_(_003882_, _040860_, _040873_);
  and g_131049_(_040662_, _040664_, _040874_);
  and g_131050_(_040873_, _040874_, _040876_);
  or g_131051_(_040663_, _040665_, _040877_);
  or g_131052_(_040872_, _040877_, _040878_);
  and g_131053_(_040871_, _040878_, _040879_);
  or g_131054_(_040870_, _040876_, _040880_);
  and g_131055_(_040872_, _040877_, _040881_);
  or g_131056_(_040873_, _040874_, _040882_);
  and g_131057_(_040861_, _040869_, _040883_);
  or g_131058_(_040862_, _040868_, _040884_);
  and g_131059_(_040882_, _040884_, _040885_);
  or g_131060_(_040881_, _040883_, _040887_);
  and g_131061_(out[201], _040857_, _040888_);
  xor g_131062_(out[201], _040857_, _040889_);
  or g_131063_(_040859_, _040888_, _040890_);
  or g_131064_(_040680_, _040841_, _040891_);
  not g_131065_(_040891_, _040892_);
  and g_131066_(_040686_, _040841_, _040893_);
  or g_131067_(_040685_, _040840_, _040894_);
  and g_131068_(_040891_, _040894_, _040895_);
  or g_131069_(_040892_, _040893_, _040896_);
  and g_131070_(_040890_, _040896_, _040898_);
  or g_131071_(_040889_, _040895_, _040899_);
  and g_131072_(_040885_, _040899_, _040900_);
  and g_131073_(_040879_, _040900_, _040901_);
  or g_131074_(_040670_, _040841_, _040902_);
  not g_131075_(_040902_, _040903_);
  and g_131076_(_040676_, _040841_, _040904_);
  or g_131077_(_040675_, _040840_, _040905_);
  and g_131078_(_040902_, _040905_, _040906_);
  or g_131079_(_040903_, _040904_, _040907_);
  xor g_131080_(out[200], _040856_, _040909_);
  xor g_131081_(_003981_, _040856_, _040910_);
  and g_131082_(_040907_, _040909_, _040911_);
  not g_131083_(_040911_, _040912_);
  and g_131084_(_040889_, _040895_, _040913_);
  or g_131085_(_040890_, _040896_, _040914_);
  and g_131086_(_040906_, _040910_, _040915_);
  or g_131087_(_040907_, _040909_, _040916_);
  and g_131088_(_040914_, _040916_, _040917_);
  or g_131089_(_040913_, _040915_, _040918_);
  and g_131090_(_040912_, _040917_, _040920_);
  or g_131091_(_040880_, _040887_, _040921_);
  or g_131092_(_040898_, _040918_, _040922_);
  or g_131093_(_040911_, _040922_, _040923_);
  and g_131094_(_040901_, _040920_, _040924_);
  or g_131095_(_040921_, _040923_, _040925_);
  xor g_131096_(out[199], _040855_, _040926_);
  xor g_131097_(_003893_, _040855_, _040927_);
  or g_131098_(_040799_, _040841_, _040928_);
  not g_131099_(_040928_, _040929_);
  and g_131100_(_040806_, _040841_, _040931_);
  not g_131101_(_040931_, _040932_);
  and g_131102_(_040928_, _040932_, _040933_);
  or g_131103_(_040929_, _040931_, _040934_);
  and g_131104_(_040926_, _040934_, _040935_);
  or g_131105_(_040927_, _040933_, _040936_);
  xor g_131106_(out[198], _040854_, _040937_);
  xor g_131107_(_003904_, _040854_, _040938_);
  and g_131108_(_040848_, _040938_, _040939_);
  or g_131109_(_040847_, _040937_, _040940_);
  and g_131110_(_040936_, _040940_, _040942_);
  or g_131111_(_040935_, _040939_, _040943_);
  and g_131112_(_040847_, _040937_, _040944_);
  or g_131113_(_040848_, _040938_, _040945_);
  and g_131114_(_040927_, _040933_, _040946_);
  or g_131115_(_040926_, _040934_, _040947_);
  and g_131116_(_040945_, _040947_, _040948_);
  or g_131117_(_040944_, _040946_, _040949_);
  and g_131118_(_040942_, _040948_, _040950_);
  or g_131119_(_040943_, _040949_, _040951_);
  xor g_131120_(out[197], _040852_, _040953_);
  xor g_131121_(_003915_, _040852_, _040954_);
  and g_131122_(_040773_, _040841_, _040955_);
  or g_131123_(_040772_, _040840_, _040956_);
  and g_131124_(_040767_, _040840_, _040957_);
  or g_131125_(_040766_, _040841_, _040958_);
  and g_131126_(_040956_, _040958_, _040959_);
  or g_131127_(_040955_, _040957_, _040960_);
  and g_131128_(_040954_, _040959_, _040961_);
  or g_131129_(_040953_, _040960_, _040962_);
  xor g_131130_(out[196], _040851_, _040964_);
  xor g_131131_(_003926_, _040851_, _040965_);
  and g_131132_(_040749_, _040840_, _040966_);
  or g_131133_(_040748_, _040841_, _040967_);
  and g_131134_(_040756_, _040841_, _040968_);
  or g_131135_(_040755_, _040840_, _040969_);
  and g_131136_(_040967_, _040969_, _040970_);
  or g_131137_(_040966_, _040968_, _040971_);
  and g_131138_(_040965_, _040970_, _040972_);
  or g_131139_(_040964_, _040971_, _040973_);
  and g_131140_(_040962_, _040973_, _040975_);
  or g_131141_(_040961_, _040972_, _040976_);
  and g_131142_(_040964_, _040971_, _040977_);
  or g_131143_(_040965_, _040970_, _040978_);
  and g_131144_(_040953_, _040960_, _040979_);
  or g_131145_(_040954_, _040959_, _040980_);
  and g_131146_(_040978_, _040980_, _040981_);
  or g_131147_(_040977_, _040979_, _040982_);
  and g_131148_(_040975_, _040981_, _040983_);
  or g_131149_(_040976_, _040982_, _040984_);
  and g_131150_(_040950_, _040983_, _040986_);
  or g_131151_(_040951_, _040984_, _040987_);
  and g_131152_(_040924_, _040986_, _040988_);
  or g_131153_(_040925_, _040987_, _040989_);
  xor g_131154_(out[195], _040850_, _040990_);
  xor g_131155_(_003970_, _040850_, _040991_);
  or g_131156_(_040733_, _040841_, _040992_);
  not g_131157_(_040992_, _040993_);
  and g_131158_(_040740_, _040841_, _040994_);
  not g_131159_(_040994_, _040995_);
  and g_131160_(_040992_, _040995_, _040997_);
  or g_131161_(_040993_, _040994_, _040998_);
  and g_131162_(_040990_, _040998_, _040999_);
  or g_131163_(_040991_, _040997_, _041000_);
  xor g_131164_(out[194], _040849_, _041001_);
  not g_131165_(_041001_, _041002_);
  or g_131166_(_040692_, _040841_, _041003_);
  not g_131167_(_041003_, _041004_);
  and g_131168_(_040698_, _040841_, _041005_);
  not g_131169_(_041005_, _041006_);
  and g_131170_(_041003_, _041006_, _041008_);
  or g_131171_(_041004_, _041005_, _041009_);
  and g_131172_(_041001_, _041008_, _041010_);
  or g_131173_(_041002_, _041009_, _041011_);
  and g_131174_(_040991_, _040997_, _041012_);
  or g_131175_(_040990_, _040998_, _041013_);
  and g_131176_(_041011_, _041013_, _041014_);
  or g_131177_(_041010_, _041012_, _041015_);
  and g_131178_(_041000_, _041015_, _041016_);
  or g_131179_(_040999_, _041014_, _041017_);
  xor g_131180_(out[193], out[192], _041019_);
  not g_131181_(_041019_, _041020_);
  or g_131182_(_040712_, _040841_, _041021_);
  not g_131183_(_041021_, _041022_);
  and g_131184_(_040707_, _040841_, _041023_);
  not g_131185_(_041023_, _041024_);
  and g_131186_(_041021_, _041024_, _041025_);
  or g_131187_(_041022_, _041023_, _041026_);
  and g_131188_(_041019_, _041025_, _041027_);
  or g_131189_(_041020_, _041026_, _041028_);
  or g_131190_(_003816_, _040841_, _041030_);
  not g_131191_(_041030_, _041031_);
  and g_131192_(_040720_, _040841_, _041032_);
  not g_131193_(_041032_, _041033_);
  and g_131194_(_041030_, _041033_, _041034_);
  or g_131195_(_041031_, _041032_, _041035_);
  and g_131196_(_003948_, _041035_, _041036_);
  or g_131197_(out[192], _041034_, _041037_);
  xor g_131198_(_041019_, _041025_, _041038_);
  xor g_131199_(_041020_, _041025_, _041039_);
  and g_131200_(_041037_, _041038_, _041041_);
  or g_131201_(_041036_, _041039_, _041042_);
  and g_131202_(_041028_, _041042_, _041043_);
  or g_131203_(_041027_, _041041_, _041044_);
  xor g_131204_(_041001_, _041008_, _041045_);
  xor g_131205_(_041002_, _041008_, _041046_);
  and g_131206_(_041000_, _041013_, _041047_);
  or g_131207_(_040999_, _041012_, _041048_);
  and g_131208_(_041045_, _041047_, _041049_);
  or g_131209_(_041046_, _041048_, _041050_);
  and g_131210_(_041044_, _041049_, _041052_);
  or g_131211_(_041043_, _041050_, _041053_);
  and g_131212_(_041017_, _041053_, _041054_);
  or g_131213_(_041016_, _041052_, _041055_);
  and g_131214_(_040988_, _041055_, _041056_);
  or g_131215_(_040989_, _041054_, _041057_);
  and g_131216_(_040936_, _040949_, _041058_);
  or g_131217_(_040935_, _040948_, _041059_);
  and g_131218_(_040976_, _040980_, _041060_);
  or g_131219_(_040975_, _040979_, _041061_);
  and g_131220_(_040942_, _041060_, _041063_);
  or g_131221_(_040943_, _041061_, _041064_);
  and g_131222_(_041059_, _041064_, _041065_);
  or g_131223_(_041058_, _041063_, _041066_);
  and g_131224_(_040924_, _041066_, _041067_);
  or g_131225_(_040925_, _041065_, _041068_);
  or g_131226_(_040879_, _040881_, _041069_);
  not g_131227_(_041069_, _041070_);
  or g_131228_(_040917_, _040921_, _041071_);
  and g_131229_(_040901_, _040918_, _041072_);
  or g_131230_(_040898_, _041071_, _041074_);
  and g_131231_(_041069_, _041074_, _041075_);
  or g_131232_(_041070_, _041072_, _041076_);
  and g_131233_(_041068_, _041075_, _041077_);
  or g_131234_(_041067_, _041076_, _041078_);
  and g_131235_(_041057_, _041077_, _041079_);
  or g_131236_(_041056_, _041078_, _041080_);
  and g_131237_(out[192], _041034_, _041081_);
  or g_131238_(_003948_, _041035_, _041082_);
  and g_131239_(_040988_, _041082_, _041083_);
  or g_131240_(_040989_, _041081_, _041085_);
  and g_131241_(_041041_, _041049_, _041086_);
  or g_131242_(_041042_, _041050_, _041087_);
  and g_131243_(_041083_, _041086_, _041088_);
  or g_131244_(_041085_, _041087_, _041089_);
  and g_131245_(_041080_, _041089_, _041090_);
  or g_131246_(_041079_, _041088_, _041091_);
  or g_131247_(_040847_, _041090_, _041092_);
  not g_131248_(_041092_, _041093_);
  and g_131249_(_040937_, _041090_, _041094_);
  not g_131250_(_041094_, _041096_);
  and g_131251_(_041092_, _041096_, _041097_);
  or g_131252_(_041093_, _041094_, _041098_);
  or g_131253_(_040933_, _041090_, _041099_);
  not g_131254_(_041099_, _041100_);
  and g_131255_(_040927_, _041090_, _041101_);
  or g_131256_(_040926_, _041091_, _041102_);
  and g_131257_(_041099_, _041102_, _041103_);
  or g_131258_(_041100_, _041101_, _041104_);
  or g_131259_(out[209], out[208], _041105_);
  or g_131260_(out[208], _046870_, _041107_);
  and g_131261_(out[211], _041107_, _041108_);
  and g_131262_(_018164_, _041107_, _041109_);
  and g_131263_(out[213], _041109_, _041110_);
  or g_131264_(out[214], _041110_, _041111_);
  and g_131265_(out[215], _041111_, _041112_);
  xor g_131266_(out[215], _041111_, _041113_);
  xor g_131267_(_004003_, _041111_, _041114_);
  and g_131268_(_041104_, _041113_, _041115_);
  or g_131269_(_041103_, _041114_, _041116_);
  xor g_131270_(out[214], _041110_, _041118_);
  xor g_131271_(_004014_, _041110_, _041119_);
  and g_131272_(_041098_, _041119_, _041120_);
  or g_131273_(_041097_, _041118_, _041121_);
  xor g_131274_(out[213], _041109_, _041122_);
  xor g_131275_(_004025_, _041109_, _041123_);
  and g_131276_(_040954_, _041090_, _041124_);
  or g_131277_(_040953_, _041091_, _041125_);
  or g_131278_(_040959_, _041090_, _041126_);
  not g_131279_(_041126_, _041127_);
  and g_131280_(_041125_, _041126_, _041129_);
  or g_131281_(_041124_, _041127_, _041130_);
  and g_131282_(_041123_, _041129_, _041131_);
  or g_131283_(_041122_, _041130_, _041132_);
  xor g_131284_(out[210], _041105_, _041133_);
  xor g_131285_(_004069_, _041105_, _041134_);
  or g_131286_(_041008_, _041090_, _041135_);
  not g_131287_(_041135_, _041136_);
  and g_131288_(_041001_, _041090_, _041137_);
  not g_131289_(_041137_, _041138_);
  and g_131290_(_041135_, _041138_, _041140_);
  or g_131291_(_041136_, _041137_, _041141_);
  and g_131292_(_041133_, _041140_, _041142_);
  or g_131293_(_041134_, _041141_, _041143_);
  and g_131294_(_041026_, _041091_, _041144_);
  or g_131295_(_041025_, _041090_, _041145_);
  and g_131296_(_041019_, _041090_, _041146_);
  or g_131297_(_041020_, _041091_, _041147_);
  and g_131298_(_041145_, _041147_, _041148_);
  or g_131299_(_041144_, _041146_, _041149_);
  and g_131300_(out[209], _041149_, _041151_);
  not g_131301_(_041151_, _041152_);
  xor g_131302_(out[209], out[208], _041153_);
  xor g_131303_(_004047_, out[208], _041154_);
  and g_131304_(_041148_, _041153_, _041155_);
  or g_131305_(_041149_, _041154_, _041156_);
  and g_131306_(out[192], _041090_, _041157_);
  or g_131307_(_003948_, _041091_, _041158_);
  and g_131308_(_041035_, _041091_, _041159_);
  or g_131309_(_041034_, _041090_, _041160_);
  and g_131310_(_041158_, _041160_, _041162_);
  or g_131311_(_041157_, _041159_, _041163_);
  and g_131312_(out[208], _041162_, _041164_);
  or g_131313_(_004058_, _041163_, _041165_);
  and g_131314_(_041156_, _041165_, _041166_);
  or g_131315_(_041155_, _041164_, _041167_);
  and g_131316_(_041152_, _041167_, _041168_);
  or g_131317_(_041151_, _041166_, _041169_);
  and g_131318_(_041143_, _041169_, _041170_);
  or g_131319_(_041142_, _041168_, _041171_);
  and g_131320_(_041134_, _041141_, _041173_);
  or g_131321_(_041133_, _041140_, _041174_);
  xor g_131322_(out[211], _041107_, _041175_);
  xor g_131323_(_004080_, _041107_, _041176_);
  and g_131324_(_040991_, _041090_, _041177_);
  or g_131325_(_040990_, _041091_, _041178_);
  or g_131326_(_040997_, _041090_, _041179_);
  not g_131327_(_041179_, _041180_);
  and g_131328_(_041178_, _041179_, _041181_);
  or g_131329_(_041177_, _041180_, _041182_);
  and g_131330_(_041175_, _041182_, _041184_);
  or g_131331_(_041176_, _041181_, _041185_);
  and g_131332_(_041174_, _041185_, _041186_);
  or g_131333_(_041173_, _041184_, _041187_);
  and g_131334_(_041171_, _041186_, _041188_);
  or g_131335_(_041170_, _041187_, _041189_);
  xor g_131336_(out[212], _041108_, _041190_);
  xor g_131337_(_004036_, _041108_, _041191_);
  or g_131338_(_040970_, _041090_, _041192_);
  not g_131339_(_041192_, _041193_);
  and g_131340_(_040965_, _041090_, _041195_);
  or g_131341_(_040964_, _041091_, _041196_);
  and g_131342_(_041192_, _041196_, _041197_);
  or g_131343_(_041193_, _041195_, _041198_);
  and g_131344_(_041191_, _041197_, _041199_);
  or g_131345_(_041190_, _041198_, _041200_);
  and g_131346_(_041176_, _041181_, _041201_);
  or g_131347_(_041175_, _041182_, _041202_);
  and g_131348_(_041200_, _041202_, _041203_);
  or g_131349_(_041199_, _041201_, _041204_);
  and g_131350_(_041189_, _041203_, _041206_);
  or g_131351_(_041188_, _041204_, _041207_);
  and g_131352_(_041122_, _041130_, _041208_);
  or g_131353_(_041123_, _041129_, _041209_);
  and g_131354_(_041190_, _041198_, _041210_);
  or g_131355_(_041191_, _041197_, _041211_);
  and g_131356_(_041209_, _041211_, _041212_);
  or g_131357_(_041208_, _041210_, _041213_);
  and g_131358_(_041207_, _041212_, _041214_);
  or g_131359_(_041206_, _041213_, _041215_);
  and g_131360_(_041132_, _041215_, _041217_);
  or g_131361_(_041131_, _041214_, _041218_);
  and g_131362_(_041121_, _041218_, _041219_);
  or g_131363_(_041120_, _041217_, _041220_);
  and g_131364_(_041103_, _041114_, _041221_);
  or g_131365_(_041104_, _041113_, _041222_);
  and g_131366_(_041097_, _041118_, _041223_);
  or g_131367_(_041098_, _041119_, _041224_);
  and g_131368_(_041222_, _041224_, _041225_);
  or g_131369_(_041221_, _041223_, _041226_);
  and g_131370_(_041220_, _041225_, _041228_);
  or g_131371_(_041219_, _041226_, _041229_);
  and g_131372_(_041116_, _041229_, _041230_);
  or g_131373_(_041115_, _041228_, _041231_);
  and g_131374_(out[216], _041112_, _041232_);
  or g_131375_(out[217], _041232_, _041233_);
  and g_131376_(out[218], _041233_, _041234_);
  xor g_131377_(out[218], _041233_, _041235_);
  xor g_131378_(_004113_, _041233_, _041236_);
  and g_131379_(_040869_, _041091_, _041237_);
  and g_131380_(_040862_, _041090_, _041239_);
  or g_131381_(_041237_, _041239_, _041240_);
  and g_131382_(_041235_, _041240_, _041241_);
  xor g_131383_(out[219], _041234_, _041242_);
  xor g_131384_(_003992_, _041234_, _041243_);
  and g_131385_(_040873_, _041090_, _041244_);
  or g_131386_(_040872_, _041091_, _041245_);
  or g_131387_(_040874_, _041090_, _041246_);
  not g_131388_(_041246_, _041247_);
  and g_131389_(_041245_, _041246_, _041248_);
  or g_131390_(_041244_, _041247_, _041250_);
  or g_131391_(_040877_, _041090_, _041251_);
  not g_131392_(_041251_, _041252_);
  and g_131393_(_040872_, _041090_, _041253_);
  not g_131394_(_041253_, _041254_);
  and g_131395_(_041251_, _041254_, _041255_);
  or g_131396_(_041252_, _041253_, _041256_);
  and g_131397_(_041242_, _041255_, _041257_);
  or g_131398_(_041242_, _041250_, _041258_);
  xor g_131399_(_041235_, _041240_, _041259_);
  xor g_131400_(_041236_, _041240_, _041261_);
  xor g_131401_(_041243_, _041248_, _041262_);
  xor g_131402_(_041242_, _041248_, _041263_);
  and g_131403_(_041259_, _041262_, _041264_);
  or g_131404_(_041261_, _041263_, _041265_);
  and g_131405_(_040907_, _041091_, _041266_);
  and g_131406_(_040910_, _041090_, _041267_);
  or g_131407_(_041266_, _041267_, _041268_);
  xor g_131408_(out[216], _041112_, _041269_);
  xor g_131409_(_004091_, _041112_, _041270_);
  xor g_131410_(out[217], _041232_, _041272_);
  not g_131411_(_041272_, _041273_);
  and g_131412_(_040896_, _041091_, _041274_);
  and g_131413_(_040889_, _041090_, _041275_);
  or g_131414_(_041274_, _041275_, _041276_);
  or g_131415_(_041273_, _041276_, _041277_);
  and g_131416_(_041268_, _041269_, _041278_);
  and g_131417_(_041273_, _041276_, _041279_);
  or g_131418_(_041278_, _041279_, _041280_);
  xor g_131419_(_041268_, _041269_, _041281_);
  xor g_131420_(_041268_, _041270_, _041283_);
  xor g_131421_(_041273_, _041276_, _041284_);
  xor g_131422_(_041272_, _041276_, _041285_);
  and g_131423_(_041264_, _041284_, _041286_);
  or g_131424_(_041265_, _041285_, _041287_);
  and g_131425_(_041281_, _041286_, _041288_);
  or g_131426_(_041283_, _041287_, _041289_);
  and g_131427_(_041231_, _041288_, _041290_);
  or g_131428_(_041230_, _041289_, _041291_);
  and g_131429_(_041264_, _041280_, _041292_);
  and g_131430_(_041277_, _041292_, _041294_);
  and g_131431_(_041241_, _041258_, _041295_);
  or g_131432_(_041257_, _041295_, _041296_);
  or g_131433_(_041294_, _041296_, _041297_);
  not g_131434_(_041297_, _041298_);
  and g_131435_(_041291_, _041298_, _041299_);
  or g_131436_(_041290_, _041297_, _041300_);
  and g_131437_(_041098_, _041300_, _041301_);
  not g_131438_(_041301_, _041302_);
  or g_131439_(_041119_, _041300_, _041303_);
  not g_131440_(_041303_, _041305_);
  and g_131441_(_041302_, _041303_, _041306_);
  or g_131442_(_041301_, _041305_, _041307_);
  and g_131443_(_041104_, _041300_, _041308_);
  not g_131444_(_041308_, _041309_);
  or g_131445_(_041113_, _041300_, _041310_);
  not g_131446_(_041310_, _041311_);
  and g_131447_(_041309_, _041310_, _041312_);
  or g_131448_(_041308_, _041311_, _041313_);
  or g_131449_(out[225], out[224], _041314_);
  or g_131450_(out[224], _047805_, _041316_);
  and g_131451_(out[227], _041316_, _041317_);
  and g_131452_(_018335_, _041316_, _041318_);
  and g_131453_(out[229], _041318_, _041319_);
  or g_131454_(out[230], _041319_, _041320_);
  and g_131455_(out[231], _041320_, _041321_);
  xor g_131456_(out[231], _041320_, _041322_);
  not g_131457_(_041322_, _041323_);
  and g_131458_(_041313_, _041322_, _041324_);
  or g_131459_(_041312_, _041323_, _041325_);
  xor g_131460_(out[230], _041319_, _041327_);
  xor g_131461_(_004146_, _041319_, _041328_);
  and g_131462_(_041306_, _041327_, _041329_);
  or g_131463_(_041307_, _041328_, _041330_);
  xor g_131464_(out[229], _041318_, _041331_);
  not g_131465_(_041331_, _041332_);
  or g_131466_(_041122_, _041300_, _041333_);
  not g_131467_(_041333_, _041334_);
  and g_131468_(_041130_, _041300_, _041335_);
  not g_131469_(_041335_, _041336_);
  and g_131470_(_041333_, _041336_, _041338_);
  or g_131471_(_041334_, _041335_, _041339_);
  and g_131472_(_041332_, _041338_, _041340_);
  or g_131473_(_041331_, _041339_, _041341_);
  xor g_131474_(out[228], _041317_, _041342_);
  not g_131475_(_041342_, _041343_);
  or g_131476_(_041190_, _041300_, _041344_);
  not g_131477_(_041344_, _041345_);
  and g_131478_(_041198_, _041300_, _041346_);
  not g_131479_(_041346_, _041347_);
  and g_131480_(_041344_, _041347_, _041349_);
  or g_131481_(_041345_, _041346_, _041350_);
  and g_131482_(_041342_, _041350_, _041351_);
  or g_131483_(_041343_, _041349_, _041352_);
  xor g_131484_(out[226], _041314_, _041353_);
  xor g_131485_(_004201_, _041314_, _041354_);
  and g_131486_(_041133_, _041299_, _041355_);
  and g_131487_(_041141_, _041300_, _041356_);
  or g_131488_(_041355_, _041356_, _041357_);
  not g_131489_(_041357_, _041358_);
  and g_131490_(_041353_, _041358_, _041360_);
  or g_131491_(_041354_, _041357_, _041361_);
  and g_131492_(_041153_, _041299_, _041362_);
  or g_131493_(_041154_, _041300_, _041363_);
  and g_131494_(_041149_, _041300_, _041364_);
  or g_131495_(_041148_, _041299_, _041365_);
  and g_131496_(_041363_, _041365_, _041366_);
  or g_131497_(_041362_, _041364_, _041367_);
  and g_131498_(out[225], _041367_, _041368_);
  not g_131499_(_041368_, _041369_);
  xor g_131500_(out[225], out[224], _041371_);
  xor g_131501_(_004179_, out[224], _041372_);
  and g_131502_(_041366_, _041371_, _041373_);
  or g_131503_(_041367_, _041372_, _041374_);
  and g_131504_(out[208], _041299_, _041375_);
  or g_131505_(_004058_, _041300_, _041376_);
  and g_131506_(_041163_, _041300_, _041377_);
  or g_131507_(_041162_, _041299_, _041378_);
  and g_131508_(_041376_, _041378_, _041379_);
  or g_131509_(_041375_, _041377_, _041380_);
  and g_131510_(out[224], _041379_, _041382_);
  or g_131511_(_004190_, _041380_, _041383_);
  and g_131512_(_041374_, _041383_, _041384_);
  or g_131513_(_041373_, _041382_, _041385_);
  and g_131514_(_041369_, _041385_, _041386_);
  or g_131515_(_041368_, _041384_, _041387_);
  and g_131516_(_041361_, _041387_, _041388_);
  or g_131517_(_041360_, _041386_, _041389_);
  and g_131518_(_041354_, _041357_, _041390_);
  or g_131519_(_041353_, _041358_, _041391_);
  xor g_131520_(out[227], _041316_, _041393_);
  xor g_131521_(_004212_, _041316_, _041394_);
  or g_131522_(_041175_, _041300_, _041395_);
  not g_131523_(_041395_, _041396_);
  and g_131524_(_041182_, _041300_, _041397_);
  not g_131525_(_041397_, _041398_);
  and g_131526_(_041395_, _041398_, _041399_);
  or g_131527_(_041396_, _041397_, _041400_);
  and g_131528_(_041393_, _041400_, _041401_);
  or g_131529_(_041394_, _041399_, _041402_);
  and g_131530_(_041391_, _041402_, _041404_);
  or g_131531_(_041390_, _041401_, _041405_);
  and g_131532_(_041389_, _041404_, _041406_);
  or g_131533_(_041388_, _041405_, _041407_);
  or g_131534_(_041342_, _041350_, _041408_);
  or g_131535_(_041393_, _041400_, _041409_);
  and g_131536_(_041408_, _041409_, _041410_);
  not g_131537_(_041410_, _041411_);
  and g_131538_(_041407_, _041410_, _041412_);
  or g_131539_(_041406_, _041411_, _041413_);
  and g_131540_(_041352_, _041413_, _041415_);
  or g_131541_(_041351_, _041412_, _041416_);
  and g_131542_(_041341_, _041416_, _041417_);
  or g_131543_(_041340_, _041415_, _041418_);
  and g_131544_(_041307_, _041328_, _041419_);
  or g_131545_(_041306_, _041327_, _041420_);
  and g_131546_(_041331_, _041339_, _041421_);
  or g_131547_(_041332_, _041338_, _041422_);
  and g_131548_(_041420_, _041422_, _041423_);
  or g_131549_(_041419_, _041421_, _041424_);
  and g_131550_(_041418_, _041423_, _041426_);
  or g_131551_(_041417_, _041424_, _041427_);
  and g_131552_(_041330_, _041427_, _041428_);
  or g_131553_(_041329_, _041426_, _041429_);
  and g_131554_(_041325_, _041429_, _041430_);
  or g_131555_(_041324_, _041428_, _041431_);
  and g_131556_(out[232], _041321_, _041432_);
  or g_131557_(out[233], _041432_, _041433_);
  xor g_131558_(out[233], _041432_, _041434_);
  not g_131559_(_041434_, _041435_);
  and g_131560_(_041276_, _041300_, _041437_);
  not g_131561_(_041437_, _041438_);
  or g_131562_(_041273_, _041300_, _041439_);
  not g_131563_(_041439_, _041440_);
  and g_131564_(_041438_, _041439_, _041441_);
  or g_131565_(_041437_, _041440_, _041442_);
  and g_131566_(_041434_, _041441_, _041443_);
  or g_131567_(_041435_, _041442_, _041444_);
  and g_131568_(_041435_, _041442_, _041445_);
  or g_131569_(_041434_, _041441_, _041446_);
  xor g_131570_(out[232], _041321_, _041448_);
  not g_131571_(_041448_, _041449_);
  and g_131572_(_041268_, _041300_, _041450_);
  not g_131573_(_041450_, _041451_);
  or g_131574_(_041269_, _041300_, _041452_);
  not g_131575_(_041452_, _041453_);
  and g_131576_(_041451_, _041452_, _041454_);
  or g_131577_(_041450_, _041453_, _041455_);
  and g_131578_(_041448_, _041455_, _041456_);
  or g_131579_(_041449_, _041454_, _041457_);
  and g_131580_(_041446_, _041457_, _041459_);
  or g_131581_(_041445_, _041456_, _041460_);
  and g_131582_(_041444_, _041459_, _041461_);
  or g_131583_(_041443_, _041460_, _041462_);
  and g_131584_(out[234], _041433_, _041463_);
  xor g_131585_(out[234], _041433_, _041464_);
  not g_131586_(_041464_, _041465_);
  and g_131587_(_041240_, _041300_, _041466_);
  not g_131588_(_041466_, _041467_);
  or g_131589_(_041235_, _041300_, _041468_);
  not g_131590_(_041468_, _041470_);
  and g_131591_(_041467_, _041468_, _041471_);
  or g_131592_(_041466_, _041470_, _041472_);
  and g_131593_(_041465_, _041471_, _041473_);
  or g_131594_(_041464_, _041472_, _041474_);
  xor g_131595_(out[235], _041463_, _041475_);
  xor g_131596_(_004124_, _041463_, _041476_);
  and g_131597_(_041242_, _041248_, _041477_);
  or g_131598_(_041243_, _041250_, _041478_);
  and g_131599_(_041476_, _041477_, _041479_);
  or g_131600_(_041475_, _041478_, _041481_);
  and g_131601_(_041474_, _041481_, _041482_);
  or g_131602_(_041473_, _041479_, _041483_);
  and g_131603_(_041464_, _041472_, _041484_);
  or g_131604_(_041465_, _041471_, _041485_);
  and g_131605_(_041242_, _041256_, _041486_);
  or g_131606_(_041243_, _041255_, _041487_);
  and g_131607_(_041475_, _041487_, _041488_);
  or g_131608_(_041476_, _041477_, _041489_);
  and g_131609_(_041485_, _041489_, _041490_);
  or g_131610_(_041484_, _041488_, _041492_);
  and g_131611_(_041449_, _041454_, _041493_);
  or g_131612_(_041448_, _041455_, _041494_);
  and g_131613_(_041312_, _041323_, _041495_);
  or g_131614_(_041313_, _041322_, _041496_);
  and g_131615_(_041494_, _041496_, _041497_);
  or g_131616_(_041493_, _041495_, _041498_);
  and g_131617_(_041490_, _041497_, _041499_);
  or g_131618_(_041492_, _041498_, _041500_);
  and g_131619_(_041482_, _041499_, _041501_);
  or g_131620_(_041483_, _041500_, _041503_);
  and g_131621_(_041461_, _041501_, _041504_);
  or g_131622_(_041462_, _041503_, _041505_);
  and g_131623_(_041431_, _041504_, _041506_);
  or g_131624_(_041430_, _041505_, _041507_);
  and g_131625_(_041481_, _041492_, _041508_);
  or g_131626_(_041479_, _041490_, _041509_);
  and g_131627_(_041444_, _041482_, _041510_);
  or g_131628_(_041443_, _041483_, _041511_);
  and g_131629_(_041460_, _041510_, _041512_);
  or g_131630_(_041459_, _041511_, _041514_);
  and g_131631_(_041509_, _041514_, _041515_);
  or g_131632_(_041508_, _041512_, _041516_);
  and g_131633_(_041507_, _041515_, _041517_);
  or g_131634_(_041506_, _041516_, _041518_);
  and g_131635_(_041307_, _041518_, _041519_);
  not g_131636_(_041519_, _041520_);
  or g_131637_(_041328_, _041518_, _041521_);
  not g_131638_(_041521_, _041522_);
  and g_131639_(_041520_, _041521_, _041523_);
  or g_131640_(_041519_, _041522_, _041525_);
  or g_131641_(out[241], out[240], _041526_);
  or g_131642_(out[240], _050467_, _041527_);
  and g_131643_(out[243], _041527_, _041528_);
  and g_131644_(_018517_, _041527_, _041529_);
  and g_131645_(out[245], _041529_, _041530_);
  or g_131646_(out[246], _041530_, _041531_);
  and g_131647_(out[247], _041531_, _041532_);
  and g_131648_(out[248], _041532_, _041533_);
  or g_131649_(out[249], _041533_, _041534_);
  and g_131650_(out[250], _041534_, _041536_);
  xor g_131651_(out[250], _041534_, _041537_);
  not g_131652_(_041537_, _041538_);
  and g_131653_(_041472_, _041518_, _041539_);
  not g_131654_(_041539_, _041540_);
  or g_131655_(_041464_, _041518_, _041541_);
  not g_131656_(_041541_, _041542_);
  and g_131657_(_041540_, _041541_, _041543_);
  or g_131658_(_041539_, _041542_, _041544_);
  and g_131659_(_041537_, _041544_, _041545_);
  xor g_131660_(out[251], _041536_, _041547_);
  xor g_131661_(_004245_, _041536_, _041548_);
  and g_131662_(_041475_, _041477_, _041549_);
  and g_131663_(_041475_, _041486_, _041550_);
  or g_131664_(_041476_, _041487_, _041551_);
  and g_131665_(_041547_, _041551_, _041552_);
  xor g_131666_(_041538_, _041543_, _041553_);
  xor g_131667_(_041537_, _041543_, _041554_);
  or g_131668_(_041547_, _041551_, _041555_);
  xor g_131669_(_041548_, _041550_, _041556_);
  xor g_131670_(_041547_, _041550_, _041558_);
  and g_131671_(_041553_, _041556_, _041559_);
  or g_131672_(_041554_, _041558_, _041560_);
  xor g_131673_(out[249], _041533_, _041561_);
  xor g_131674_(_004344_, _041533_, _041562_);
  and g_131675_(_041442_, _041518_, _041563_);
  not g_131676_(_041563_, _041564_);
  or g_131677_(_041435_, _041518_, _041565_);
  not g_131678_(_041565_, _041566_);
  and g_131679_(_041564_, _041565_, _041567_);
  or g_131680_(_041563_, _041566_, _041569_);
  and g_131681_(_041561_, _041567_, _041570_);
  or g_131682_(_041562_, _041569_, _041571_);
  and g_131683_(_041455_, _041518_, _041572_);
  not g_131684_(_041572_, _041573_);
  or g_131685_(_041448_, _041518_, _041574_);
  not g_131686_(_041574_, _041575_);
  and g_131687_(_041573_, _041574_, _041576_);
  or g_131688_(_041572_, _041575_, _041577_);
  xor g_131689_(out[248], _041532_, _041578_);
  xor g_131690_(_004333_, _041532_, _041580_);
  and g_131691_(_041577_, _041578_, _041581_);
  or g_131692_(_041576_, _041580_, _041582_);
  and g_131693_(_041562_, _041569_, _041583_);
  or g_131694_(_041561_, _041567_, _041584_);
  or g_131695_(_041581_, _041583_, _041585_);
  and g_131696_(_041571_, _041585_, _041586_);
  xor g_131697_(out[242], _041526_, _041587_);
  xor g_131698_(_004311_, _041526_, _041588_);
  or g_131699_(_041354_, _041518_, _041589_);
  not g_131700_(_041589_, _041591_);
  and g_131701_(_041357_, _041518_, _041592_);
  not g_131702_(_041592_, _041593_);
  and g_131703_(_041589_, _041593_, _041594_);
  or g_131704_(_041591_, _041592_, _041595_);
  and g_131705_(_041587_, _041594_, _041596_);
  or g_131706_(_041588_, _041595_, _041597_);
  and g_131707_(_041371_, _041517_, _041598_);
  or g_131708_(_041372_, _041518_, _041599_);
  and g_131709_(_041367_, _041518_, _041600_);
  or g_131710_(_041366_, _041517_, _041602_);
  and g_131711_(_041599_, _041602_, _041603_);
  or g_131712_(_041598_, _041600_, _041604_);
  and g_131713_(out[241], _041604_, _041605_);
  not g_131714_(_041605_, _041606_);
  xor g_131715_(_053038_, out[240], _041607_);
  not g_131716_(_041607_, _041608_);
  and g_131717_(_041603_, _041608_, _041609_);
  or g_131718_(_041604_, _041607_, _041610_);
  and g_131719_(out[224], _041517_, _041611_);
  or g_131720_(_004190_, _041518_, _041613_);
  and g_131721_(_041380_, _041518_, _041614_);
  or g_131722_(_041379_, _041517_, _041615_);
  and g_131723_(_041613_, _041615_, _041616_);
  or g_131724_(_041611_, _041614_, _041617_);
  and g_131725_(out[240], _041616_, _041618_);
  or g_131726_(_004300_, _041617_, _041619_);
  and g_131727_(_041610_, _041619_, _041620_);
  or g_131728_(_041609_, _041618_, _041621_);
  and g_131729_(_041606_, _041621_, _041622_);
  or g_131730_(_041605_, _041620_, _041624_);
  and g_131731_(_041597_, _041624_, _041625_);
  or g_131732_(_041596_, _041622_, _041626_);
  and g_131733_(_041588_, _041595_, _041627_);
  or g_131734_(_041587_, _041594_, _041628_);
  xor g_131735_(out[243], _041527_, _041629_);
  xor g_131736_(_004322_, _041527_, _041630_);
  or g_131737_(_041393_, _041518_, _041631_);
  not g_131738_(_041631_, _041632_);
  and g_131739_(_041400_, _041518_, _041633_);
  not g_131740_(_041633_, _041635_);
  and g_131741_(_041631_, _041635_, _041636_);
  or g_131742_(_041632_, _041633_, _041637_);
  and g_131743_(_041629_, _041637_, _041638_);
  or g_131744_(_041630_, _041636_, _041639_);
  and g_131745_(_041628_, _041639_, _041640_);
  or g_131746_(_041627_, _041638_, _041641_);
  and g_131747_(_041626_, _041640_, _041642_);
  or g_131748_(_041625_, _041641_, _041643_);
  xor g_131749_(out[244], _041528_, _041644_);
  xor g_131750_(_004289_, _041528_, _041646_);
  or g_131751_(_041342_, _041518_, _041647_);
  not g_131752_(_041647_, _041648_);
  and g_131753_(_041350_, _041518_, _041649_);
  not g_131754_(_041649_, _041650_);
  and g_131755_(_041647_, _041650_, _041651_);
  or g_131756_(_041648_, _041649_, _041652_);
  and g_131757_(_041646_, _041651_, _041653_);
  or g_131758_(_041644_, _041652_, _041654_);
  and g_131759_(_041630_, _041636_, _041655_);
  or g_131760_(_041629_, _041637_, _041657_);
  and g_131761_(_041654_, _041657_, _041658_);
  or g_131762_(_041653_, _041655_, _041659_);
  and g_131763_(_041643_, _041658_, _041660_);
  or g_131764_(_041642_, _041659_, _041661_);
  xor g_131765_(out[245], _041529_, _041662_);
  xor g_131766_(_004278_, _041529_, _041663_);
  or g_131767_(_041331_, _041518_, _041664_);
  not g_131768_(_041664_, _041665_);
  and g_131769_(_041339_, _041518_, _041666_);
  not g_131770_(_041666_, _041668_);
  and g_131771_(_041664_, _041668_, _041669_);
  or g_131772_(_041665_, _041666_, _041670_);
  and g_131773_(_041662_, _041670_, _041671_);
  or g_131774_(_041663_, _041669_, _041672_);
  and g_131775_(_041644_, _041652_, _041673_);
  or g_131776_(_041646_, _041651_, _041674_);
  and g_131777_(_041672_, _041674_, _041675_);
  or g_131778_(_041671_, _041673_, _041676_);
  and g_131779_(_041661_, _041675_, _041677_);
  or g_131780_(_041660_, _041676_, _041679_);
  xor g_131781_(out[246], _041530_, _041680_);
  xor g_131782_(_004267_, _041530_, _041681_);
  and g_131783_(_041523_, _041680_, _041682_);
  or g_131784_(_041525_, _041681_, _041683_);
  and g_131785_(_041663_, _041669_, _041684_);
  or g_131786_(_041662_, _041670_, _041685_);
  and g_131787_(_041683_, _041685_, _041686_);
  or g_131788_(_041682_, _041684_, _041687_);
  and g_131789_(_041679_, _041686_, _041688_);
  or g_131790_(_041677_, _041687_, _041690_);
  xor g_131791_(out[247], _041531_, _041691_);
  xor g_131792_(_004256_, _041531_, _041692_);
  and g_131793_(_041313_, _041518_, _041693_);
  not g_131794_(_041693_, _041694_);
  or g_131795_(_041322_, _041518_, _041695_);
  not g_131796_(_041695_, _041696_);
  and g_131797_(_041694_, _041695_, _041697_);
  or g_131798_(_041693_, _041696_, _041698_);
  and g_131799_(_041691_, _041698_, _041699_);
  or g_131800_(_041692_, _041697_, _041701_);
  and g_131801_(_041525_, _041681_, _041702_);
  or g_131802_(_041523_, _041680_, _041703_);
  and g_131803_(_041701_, _041703_, _041704_);
  or g_131804_(_041699_, _041702_, _041705_);
  and g_131805_(_041690_, _041704_, _041706_);
  or g_131806_(_041688_, _041705_, _041707_);
  and g_131807_(_041576_, _041580_, _041708_);
  or g_131808_(_041577_, _041578_, _041709_);
  and g_131809_(_041692_, _041697_, _041710_);
  or g_131810_(_041691_, _041698_, _041712_);
  and g_131811_(_041571_, _041709_, _041713_);
  or g_131812_(_041570_, _041708_, _041714_);
  and g_131813_(_041584_, _041712_, _041715_);
  or g_131814_(_041583_, _041710_, _041716_);
  and g_131815_(_041713_, _041715_, _041717_);
  or g_131816_(_041714_, _041716_, _041718_);
  and g_131817_(_041559_, _041717_, _041719_);
  or g_131818_(_041560_, _041718_, _041720_);
  and g_131819_(_041707_, _041719_, _041721_);
  or g_131820_(_041706_, _041720_, _041723_);
  and g_131821_(_041582_, _041721_, _041724_);
  or g_131822_(_041581_, _041723_, _041725_);
  and g_131823_(_041559_, _041586_, _041726_);
  and g_131824_(_041545_, _041555_, _041727_);
  or g_131825_(_041726_, _041727_, _041728_);
  or g_131826_(_041552_, _041728_, _041729_);
  not g_131827_(_041729_, _041730_);
  and g_131828_(_041725_, _041730_, _041731_);
  or g_131829_(_041724_, _041729_, _041732_);
  and g_131830_(_041525_, _041732_, _041734_);
  or g_131831_(_041523_, _041731_, _041735_);
  and g_131832_(_041680_, _041731_, _041736_);
  or g_131833_(_041681_, _041732_, _041737_);
  and g_131834_(_041735_, _041737_, _041738_);
  or g_131835_(_041734_, _041736_, _041739_);
  or g_131836_(out[257], out[256], _041740_);
  or g_131837_(out[256], _051425_, _041741_);
  and g_131838_(out[259], _041741_, _041742_);
  and g_131839_(_018749_, _041741_, _041743_);
  and g_131840_(out[261], _041743_, _041745_);
  or g_131841_(out[262], _041745_, _041746_);
  and g_131842_(out[263], _041746_, _041747_);
  and g_131843_(out[264], _041747_, _041748_);
  xor g_131844_(out[264], _041747_, _041749_);
  xor g_131845_(_004399_, _041747_, _041750_);
  and g_131846_(_041577_, _041732_, _041751_);
  or g_131847_(_041576_, _041731_, _041752_);
  and g_131848_(_041580_, _041731_, _041753_);
  or g_131849_(_041578_, _041732_, _041754_);
  and g_131850_(_041752_, _041754_, _041756_);
  or g_131851_(_041751_, _041753_, _041757_);
  and g_131852_(_041750_, _041756_, _041758_);
  or g_131853_(_041749_, _041757_, _041759_);
  or g_131854_(out[265], _041748_, _041760_);
  xor g_131855_(out[265], _041748_, _041761_);
  xor g_131856_(_004410_, _041748_, _041762_);
  and g_131857_(_041569_, _041732_, _041763_);
  or g_131858_(_041567_, _041731_, _041764_);
  and g_131859_(_041561_, _041731_, _041765_);
  or g_131860_(_041562_, _041732_, _041767_);
  and g_131861_(_041764_, _041767_, _041768_);
  or g_131862_(_041763_, _041765_, _041769_);
  and g_131863_(_041761_, _041768_, _041770_);
  or g_131864_(_041762_, _041769_, _041771_);
  and g_131865_(_041759_, _041771_, _041772_);
  or g_131866_(_041758_, _041770_, _041773_);
  and g_131867_(out[266], _041760_, _041774_);
  xor g_131868_(out[267], _041774_, _041775_);
  xor g_131869_(_004366_, _041774_, _041776_);
  and g_131870_(_041547_, _041549_, _041778_);
  or g_131871_(_041548_, _041551_, _041779_);
  and g_131872_(_041775_, _041779_, _041780_);
  or g_131873_(_041776_, _041778_, _041781_);
  and g_131874_(_041749_, _041757_, _041782_);
  or g_131875_(_041750_, _041756_, _041783_);
  and g_131876_(_041781_, _041783_, _041784_);
  or g_131877_(_041780_, _041782_, _041785_);
  and g_131878_(_041772_, _041784_, _041786_);
  or g_131879_(_041773_, _041785_, _041787_);
  xor g_131880_(out[266], _041760_, _041789_);
  xor g_131881_(_004421_, _041760_, _041790_);
  and g_131882_(_041544_, _041732_, _041791_);
  or g_131883_(_041543_, _041731_, _041792_);
  and g_131884_(_041538_, _041731_, _041793_);
  or g_131885_(_041537_, _041732_, _041794_);
  and g_131886_(_041792_, _041794_, _041795_);
  or g_131887_(_041791_, _041793_, _041796_);
  and g_131888_(_041790_, _041795_, _041797_);
  or g_131889_(_041789_, _041796_, _041798_);
  and g_131890_(_041776_, _041778_, _041800_);
  or g_131891_(_041775_, _041779_, _041801_);
  and g_131892_(_041798_, _041801_, _041802_);
  or g_131893_(_041797_, _041800_, _041803_);
  and g_131894_(_041789_, _041796_, _041804_);
  or g_131895_(_041790_, _041795_, _041805_);
  and g_131896_(_041762_, _041769_, _041806_);
  or g_131897_(_041761_, _041768_, _041807_);
  and g_131898_(_041805_, _041807_, _041808_);
  or g_131899_(_041804_, _041806_, _041809_);
  and g_131900_(_041802_, _041808_, _041811_);
  or g_131901_(_041803_, _041809_, _041812_);
  and g_131902_(_041786_, _041811_, _041813_);
  or g_131903_(_041787_, _041812_, _041814_);
  and g_131904_(_041698_, _041732_, _041815_);
  or g_131905_(_041697_, _041731_, _041816_);
  and g_131906_(_041692_, _041731_, _041817_);
  or g_131907_(_041691_, _041732_, _041818_);
  and g_131908_(_041816_, _041818_, _041819_);
  or g_131909_(_041815_, _041817_, _041820_);
  xor g_131910_(out[263], _041746_, _041822_);
  not g_131911_(_041822_, _041823_);
  and g_131912_(_041819_, _041823_, _041824_);
  or g_131913_(_041820_, _041822_, _041825_);
  xor g_131914_(out[262], _041745_, _041826_);
  not g_131915_(_041826_, _041827_);
  and g_131916_(_041738_, _041826_, _041828_);
  or g_131917_(_041739_, _041827_, _041829_);
  and g_131918_(_041825_, _041829_, _041830_);
  or g_131919_(_041824_, _041828_, _041831_);
  and g_131920_(_041820_, _041822_, _041833_);
  or g_131921_(_041819_, _041823_, _041834_);
  and g_131922_(_041739_, _041827_, _041835_);
  or g_131923_(_041738_, _041826_, _041836_);
  and g_131924_(_041834_, _041836_, _041837_);
  or g_131925_(_041833_, _041835_, _041838_);
  and g_131926_(_041830_, _041837_, _041839_);
  or g_131927_(_041831_, _041838_, _041840_);
  xor g_131928_(out[261], _041743_, _041841_);
  xor g_131929_(_052972_, _041743_, _041842_);
  and g_131930_(_041663_, _041731_, _041844_);
  or g_131931_(_041662_, _041732_, _041845_);
  and g_131932_(_041670_, _041732_, _041846_);
  or g_131933_(_041669_, _041731_, _041847_);
  and g_131934_(_041845_, _041847_, _041848_);
  or g_131935_(_041844_, _041846_, _041849_);
  and g_131936_(_041842_, _041848_, _041850_);
  or g_131937_(_041841_, _041849_, _041851_);
  xor g_131938_(out[260], _041742_, _041852_);
  xor g_131939_(_052994_, _041742_, _041853_);
  and g_131940_(_041646_, _041731_, _041855_);
  or g_131941_(_041644_, _041732_, _041856_);
  and g_131942_(_041652_, _041732_, _041857_);
  or g_131943_(_041651_, _041731_, _041858_);
  and g_131944_(_041856_, _041858_, _041859_);
  or g_131945_(_041855_, _041857_, _041860_);
  and g_131946_(_041853_, _041859_, _041861_);
  or g_131947_(_041852_, _041860_, _041862_);
  and g_131948_(_041851_, _041862_, _041863_);
  or g_131949_(_041850_, _041861_, _041864_);
  and g_131950_(_041852_, _041860_, _041866_);
  or g_131951_(_041853_, _041859_, _041867_);
  and g_131952_(_041841_, _041849_, _041868_);
  or g_131953_(_041842_, _041848_, _041869_);
  and g_131954_(_041867_, _041869_, _041870_);
  or g_131955_(_041866_, _041868_, _041871_);
  and g_131956_(_041863_, _041870_, _041872_);
  or g_131957_(_041864_, _041871_, _041873_);
  and g_131958_(_041839_, _041872_, _041874_);
  or g_131959_(_041840_, _041873_, _041875_);
  and g_131960_(_041813_, _041874_, _041877_);
  or g_131961_(_041814_, _041875_, _041878_);
  xor g_131962_(out[258], _041740_, _041879_);
  not g_131963_(_041879_, _041880_);
  and g_131964_(_041587_, _041731_, _041881_);
  or g_131965_(_041588_, _041732_, _041882_);
  and g_131966_(_041595_, _041732_, _041883_);
  or g_131967_(_041594_, _041731_, _041884_);
  and g_131968_(_041882_, _041884_, _041885_);
  or g_131969_(_041881_, _041883_, _041886_);
  and g_131970_(_041879_, _041885_, _041888_);
  or g_131971_(_041880_, _041886_, _041889_);
  xor g_131972_(out[259], _041741_, _041890_);
  xor g_131973_(_053005_, _041741_, _041891_);
  and g_131974_(_041630_, _041731_, _041892_);
  or g_131975_(_041629_, _041732_, _041893_);
  and g_131976_(_041637_, _041732_, _041894_);
  or g_131977_(_041636_, _041731_, _041895_);
  and g_131978_(_041893_, _041895_, _041896_);
  or g_131979_(_041892_, _041894_, _041897_);
  and g_131980_(_041891_, _041896_, _041899_);
  or g_131981_(_041890_, _041897_, _041900_);
  and g_131982_(_041890_, _041897_, _041901_);
  or g_131983_(_041891_, _041896_, _041902_);
  xor g_131984_(_041879_, _041885_, _041903_);
  xor g_131985_(_041880_, _041885_, _041904_);
  and g_131986_(_041900_, _041902_, _041905_);
  or g_131987_(_041899_, _041901_, _041906_);
  and g_131988_(_041903_, _041905_, _041907_);
  or g_131989_(_041904_, _041906_, _041908_);
  xor g_131990_(out[257], out[256], _041910_);
  not g_131991_(_041910_, _041911_);
  or g_131992_(_041607_, _041732_, _041912_);
  or g_131993_(_041603_, _041731_, _041913_);
  and g_131994_(_041912_, _041913_, _041914_);
  not g_131995_(_041914_, _041915_);
  and g_131996_(_041910_, _041914_, _041916_);
  not g_131997_(_041916_, _041917_);
  and g_131998_(out[240], _041731_, _041918_);
  or g_131999_(_004300_, _041732_, _041919_);
  and g_132000_(_041617_, _041732_, _041921_);
  or g_132001_(_041616_, _041731_, _041922_);
  and g_132002_(_041919_, _041922_, _041923_);
  or g_132003_(_041918_, _041921_, _041924_);
  and g_132004_(_004388_, _041924_, _041925_);
  or g_132005_(out[256], _041923_, _041926_);
  xor g_132006_(_041910_, _041914_, _041927_);
  xor g_132007_(_041911_, _041914_, _041928_);
  and g_132008_(_041926_, _041927_, _041929_);
  or g_132009_(_041925_, _041928_, _041930_);
  and g_132010_(_041917_, _041930_, _041932_);
  or g_132011_(_041916_, _041929_, _041933_);
  and g_132012_(_041907_, _041933_, _041934_);
  or g_132013_(_041908_, _041932_, _041935_);
  and g_132014_(_041888_, _041902_, _041936_);
  or g_132015_(_041889_, _041901_, _041937_);
  and g_132016_(_041900_, _041937_, _041938_);
  or g_132017_(_041899_, _041936_, _041939_);
  and g_132018_(_041935_, _041938_, _041940_);
  or g_132019_(_041934_, _041939_, _041941_);
  and g_132020_(_041877_, _041941_, _041943_);
  or g_132021_(_041878_, _041940_, _041944_);
  and g_132022_(_041831_, _041834_, _041945_);
  or g_132023_(_041830_, _041833_, _041946_);
  and g_132024_(_041864_, _041869_, _041947_);
  or g_132025_(_041863_, _041868_, _041948_);
  and g_132026_(_041839_, _041947_, _041949_);
  or g_132027_(_041840_, _041948_, _041950_);
  and g_132028_(_041946_, _041950_, _041951_);
  or g_132029_(_041945_, _041949_, _041952_);
  and g_132030_(_041813_, _041952_, _041954_);
  or g_132031_(_041814_, _041951_, _041955_);
  and g_132032_(_041773_, _041808_, _041956_);
  or g_132033_(_041772_, _041809_, _041957_);
  and g_132034_(_041802_, _041957_, _041958_);
  or g_132035_(_041803_, _041956_, _041959_);
  and g_132036_(_041781_, _041959_, _041960_);
  or g_132037_(_041780_, _041958_, _041961_);
  and g_132038_(_041955_, _041961_, _041962_);
  or g_132039_(_041954_, _041960_, _041963_);
  and g_132040_(_041944_, _041962_, _041965_);
  or g_132041_(_041943_, _041963_, _041966_);
  and g_132042_(out[256], _041923_, _041967_);
  or g_132043_(_004388_, _041924_, _041968_);
  and g_132044_(_041907_, _041968_, _041969_);
  or g_132045_(_041908_, _041967_, _041970_);
  and g_132046_(_041929_, _041969_, _041971_);
  or g_132047_(_041930_, _041970_, _041972_);
  and g_132048_(_041877_, _041971_, _041973_);
  or g_132049_(_041878_, _041972_, _041974_);
  and g_132050_(_041966_, _041974_, _041976_);
  or g_132051_(_041965_, _041973_, _041977_);
  and g_132052_(_041739_, _041977_, _041978_);
  or g_132053_(_041738_, _041976_, _041979_);
  and g_132054_(_041826_, _041976_, _041980_);
  not g_132055_(_041980_, _041981_);
  and g_132056_(_041979_, _041981_, _041982_);
  or g_132057_(_041978_, _041980_, _041983_);
  or g_132058_(out[273], out[272], _041984_);
  or g_132059_(out[272], _051640_, _041985_);
  and g_132060_(out[275], _041985_, _041987_);
  and g_132061_(_018960_, _041985_, _041988_);
  and g_132062_(out[277], _041988_, _041989_);
  or g_132063_(out[278], _041989_, _041990_);
  and g_132064_(out[279], _041990_, _041991_);
  and g_132065_(out[280], _041991_, _041992_);
  xor g_132066_(out[280], _041991_, _041993_);
  xor g_132067_(_053060_, _041991_, _041994_);
  and g_132068_(_041757_, _041977_, _041995_);
  or g_132069_(_041756_, _041976_, _041996_);
  and g_132070_(_041750_, _041976_, _041998_);
  or g_132071_(_041749_, _041977_, _041999_);
  and g_132072_(_041996_, _041999_, _042000_);
  or g_132073_(_041995_, _041998_, _042001_);
  and g_132074_(_041993_, _042001_, _042002_);
  not g_132075_(_042002_, _042003_);
  or g_132076_(out[281], _041992_, _042004_);
  xor g_132077_(_053137_, _041992_, _042005_);
  and g_132078_(_041769_, _041977_, _042006_);
  and g_132079_(_041761_, _041976_, _042007_);
  or g_132080_(_042006_, _042007_, _042009_);
  and g_132081_(_042005_, _042009_, _042010_);
  not g_132082_(_042010_, _042011_);
  or g_132083_(_042002_, _042010_, _042012_);
  and g_132084_(_041820_, _041977_, _042013_);
  or g_132085_(_041819_, _041976_, _042014_);
  and g_132086_(_041823_, _041976_, _042015_);
  or g_132087_(_041822_, _041977_, _042016_);
  and g_132088_(_042014_, _042016_, _042017_);
  or g_132089_(_042013_, _042015_, _042018_);
  xor g_132090_(out[279], _041990_, _042020_);
  xor g_132091_(_053049_, _041990_, _042021_);
  and g_132092_(_042018_, _042020_, _042022_);
  or g_132093_(_042017_, _042021_, _042023_);
  xor g_132094_(out[273], out[272], _042024_);
  xor g_132095_(_053126_, out[272], _042025_);
  and g_132096_(_041915_, _041977_, _042026_);
  or g_132097_(_041914_, _041976_, _042027_);
  and g_132098_(_041910_, _041976_, _042028_);
  or g_132099_(_041911_, _041977_, _042029_);
  and g_132100_(_042027_, _042029_, _042031_);
  or g_132101_(_042026_, _042028_, _042032_);
  and g_132102_(_042024_, _042031_, _042033_);
  or g_132103_(_042025_, _042032_, _042034_);
  and g_132104_(out[256], _041976_, _042035_);
  or g_132105_(_004388_, _041977_, _042036_);
  and g_132106_(_041924_, _041977_, _042037_);
  or g_132107_(_041923_, _041976_, _042038_);
  and g_132108_(_042036_, _042038_, _042039_);
  or g_132109_(_042035_, _042037_, _042040_);
  and g_132110_(out[272], _042039_, _042042_);
  or g_132111_(_004443_, _042040_, _042043_);
  and g_132112_(_042034_, _042043_, _042044_);
  or g_132113_(_042033_, _042042_, _042045_);
  xor g_132114_(out[274], _041984_, _042046_);
  xor g_132115_(_053115_, _041984_, _042047_);
  and g_132116_(_041879_, _041976_, _042048_);
  or g_132117_(_041880_, _041977_, _042049_);
  and g_132118_(_041886_, _041977_, _042050_);
  or g_132119_(_041885_, _041976_, _042051_);
  and g_132120_(_042049_, _042051_, _042053_);
  or g_132121_(_042048_, _042050_, _042054_);
  and g_132122_(_042047_, _042054_, _042055_);
  or g_132123_(_042046_, _042053_, _042056_);
  and g_132124_(out[273], _042032_, _042057_);
  or g_132125_(_053126_, _042031_, _042058_);
  and g_132126_(_042056_, _042058_, _042059_);
  or g_132127_(_042055_, _042057_, _042060_);
  and g_132128_(_042045_, _042059_, _042061_);
  or g_132129_(_042044_, _042060_, _042062_);
  and g_132130_(_042046_, _042053_, _042064_);
  or g_132131_(_042047_, _042054_, _042065_);
  xor g_132132_(out[275], _041985_, _042066_);
  xor g_132133_(_053093_, _041985_, _042067_);
  and g_132134_(_041891_, _041976_, _042068_);
  or g_132135_(_041890_, _041977_, _042069_);
  and g_132136_(_041897_, _041977_, _042070_);
  or g_132137_(_041896_, _041976_, _042071_);
  and g_132138_(_042069_, _042071_, _042072_);
  or g_132139_(_042068_, _042070_, _042073_);
  and g_132140_(_042067_, _042072_, _042075_);
  or g_132141_(_042066_, _042073_, _042076_);
  and g_132142_(_042065_, _042076_, _042077_);
  or g_132143_(_042064_, _042075_, _042078_);
  and g_132144_(_042062_, _042077_, _042079_);
  or g_132145_(_042061_, _042078_, _042080_);
  and g_132146_(_042066_, _042073_, _042081_);
  or g_132147_(_042067_, _042072_, _042082_);
  xor g_132148_(out[276], _041987_, _042083_);
  xor g_132149_(_053104_, _041987_, _042084_);
  and g_132150_(_041853_, _041976_, _042086_);
  or g_132151_(_041852_, _041977_, _042087_);
  and g_132152_(_041860_, _041977_, _042088_);
  or g_132153_(_041859_, _041976_, _042089_);
  and g_132154_(_042087_, _042089_, _042090_);
  or g_132155_(_042086_, _042088_, _042091_);
  and g_132156_(_042083_, _042091_, _042092_);
  or g_132157_(_042084_, _042090_, _042093_);
  and g_132158_(_042082_, _042093_, _042094_);
  or g_132159_(_042081_, _042092_, _042095_);
  and g_132160_(_042080_, _042094_, _042097_);
  or g_132161_(_042079_, _042095_, _042098_);
  xor g_132162_(out[277], _041988_, _042099_);
  xor g_132163_(_053071_, _041988_, _042100_);
  and g_132164_(_041842_, _041976_, _042101_);
  or g_132165_(_041841_, _041977_, _042102_);
  and g_132166_(_041849_, _041977_, _042103_);
  or g_132167_(_041848_, _041976_, _042104_);
  and g_132168_(_042102_, _042104_, _042105_);
  or g_132169_(_042101_, _042103_, _042106_);
  and g_132170_(_042100_, _042105_, _042108_);
  or g_132171_(_042099_, _042106_, _042109_);
  and g_132172_(_042084_, _042090_, _042110_);
  or g_132173_(_042083_, _042091_, _042111_);
  and g_132174_(_042109_, _042111_, _042112_);
  or g_132175_(_042108_, _042110_, _042113_);
  and g_132176_(_042098_, _042112_, _042114_);
  or g_132177_(_042097_, _042113_, _042115_);
  xor g_132178_(out[278], _041989_, _042116_);
  xor g_132179_(_053082_, _041989_, _042117_);
  and g_132180_(_041983_, _042117_, _042119_);
  or g_132181_(_041982_, _042116_, _042120_);
  and g_132182_(_042099_, _042106_, _042121_);
  or g_132183_(_042100_, _042105_, _042122_);
  and g_132184_(_042120_, _042122_, _042123_);
  or g_132185_(_042119_, _042121_, _042124_);
  and g_132186_(_042115_, _042123_, _042125_);
  or g_132187_(_042114_, _042124_, _042126_);
  and g_132188_(_042017_, _042021_, _042127_);
  or g_132189_(_042018_, _042020_, _042128_);
  and g_132190_(_041982_, _042116_, _042130_);
  or g_132191_(_041983_, _042117_, _042131_);
  and g_132192_(_042128_, _042131_, _042132_);
  or g_132193_(_042127_, _042130_, _042133_);
  and g_132194_(_042126_, _042132_, _042134_);
  or g_132195_(_042125_, _042133_, _042135_);
  and g_132196_(_042023_, _042135_, _042136_);
  or g_132197_(_042022_, _042134_, _042137_);
  and g_132198_(_041994_, _042000_, _042138_);
  or g_132199_(_041993_, _042001_, _042139_);
  and g_132200_(_041796_, _041977_, _042141_);
  and g_132201_(_041790_, _041976_, _042142_);
  or g_132202_(_042141_, _042142_, _042143_);
  and g_132203_(out[282], _042004_, _042144_);
  xor g_132204_(out[282], _042004_, _042145_);
  and g_132205_(_042143_, _042145_, _042146_);
  xor g_132206_(out[283], _042144_, _042147_);
  not g_132207_(_042147_, _042148_);
  or g_132208_(_041775_, _041977_, _042149_);
  or g_132209_(_041778_, _041976_, _042150_);
  and g_132210_(_042149_, _042150_, _042152_);
  not g_132211_(_042152_, _042153_);
  or g_132212_(_041779_, _041976_, _042154_);
  or g_132213_(_041776_, _041977_, _042155_);
  and g_132214_(_042154_, _042155_, _042156_);
  not g_132215_(_042156_, _042157_);
  and g_132216_(_042147_, _042156_, _042158_);
  or g_132217_(_042005_, _042009_, _042159_);
  not g_132218_(_042159_, _042160_);
  xor g_132219_(_042143_, _042145_, _042161_);
  or g_132220_(_042147_, _042156_, _042163_);
  xor g_132221_(_042147_, _042156_, _042164_);
  and g_132222_(_042161_, _042164_, _042165_);
  not g_132223_(_042165_, _042166_);
  and g_132224_(_042012_, _042165_, _042167_);
  and g_132225_(_042003_, _042159_, _042168_);
  or g_132226_(_042002_, _042160_, _042169_);
  and g_132227_(_042011_, _042139_, _042170_);
  or g_132228_(_042010_, _042138_, _042171_);
  and g_132229_(_042165_, _042170_, _042172_);
  or g_132230_(_042166_, _042171_, _042174_);
  and g_132231_(_042168_, _042172_, _042175_);
  or g_132232_(_042169_, _042174_, _042176_);
  and g_132233_(_042137_, _042175_, _042177_);
  or g_132234_(_042136_, _042176_, _042178_);
  and g_132235_(_042146_, _042163_, _042179_);
  and g_132236_(_042159_, _042167_, _042180_);
  or g_132237_(_042158_, _042180_, _042181_);
  or g_132238_(_042179_, _042181_, _042182_);
  not g_132239_(_042182_, _042183_);
  and g_132240_(_042178_, _042183_, _042185_);
  or g_132241_(_042177_, _042182_, _042186_);
  and g_132242_(_041983_, _042186_, _042187_);
  not g_132243_(_042187_, _042188_);
  or g_132244_(_042117_, _042186_, _042189_);
  not g_132245_(_042189_, _042190_);
  and g_132246_(_042188_, _042189_, _042191_);
  or g_132247_(_042187_, _042190_, _042192_);
  or g_132248_(out[289], out[288], _042193_);
  or g_132249_(out[288], _051815_, _042194_);
  and g_132250_(out[291], _042194_, _042196_);
  and g_132251_(_019199_, _042194_, _042197_);
  and g_132252_(out[293], _042197_, _042198_);
  or g_132253_(out[294], _042198_, _042199_);
  and g_132254_(out[295], _042199_, _042200_);
  and g_132255_(out[296], _042200_, _042201_);
  or g_132256_(out[297], _042201_, _042202_);
  and g_132257_(out[298], _042202_, _042203_);
  xor g_132258_(out[299], _042203_, _042204_);
  xor g_132259_(_004465_, _042203_, _042205_);
  and g_132260_(_042147_, _042152_, _042207_);
  or g_132261_(_042148_, _042153_, _042208_);
  and g_132262_(_042205_, _042207_, _042209_);
  or g_132263_(_042204_, _042208_, _042210_);
  and g_132264_(_042143_, _042186_, _042211_);
  not g_132265_(_042211_, _042212_);
  or g_132266_(_042145_, _042186_, _042213_);
  not g_132267_(_042213_, _042214_);
  and g_132268_(_042212_, _042213_, _042215_);
  or g_132269_(_042211_, _042214_, _042216_);
  xor g_132270_(out[298], _042202_, _042218_);
  xor g_132271_(_004487_, _042202_, _042219_);
  and g_132272_(_042216_, _042218_, _042220_);
  or g_132273_(_042215_, _042219_, _042221_);
  and g_132274_(_042147_, _042157_, _042222_);
  and g_132275_(_042204_, _042208_, _042223_);
  or g_132276_(_042205_, _042207_, _042224_);
  and g_132277_(_042221_, _042224_, _042225_);
  or g_132278_(_042220_, _042223_, _042226_);
  and g_132279_(_042210_, _042226_, _042227_);
  or g_132280_(_042209_, _042225_, _042229_);
  and g_132281_(_042215_, _042219_, _042230_);
  or g_132282_(_042216_, _042218_, _042231_);
  and g_132283_(_042210_, _042231_, _042232_);
  or g_132284_(_042209_, _042230_, _042233_);
  and g_132285_(_042225_, _042232_, _042234_);
  or g_132286_(_042226_, _042233_, _042235_);
  xor g_132287_(out[290], _042193_, _042236_);
  xor g_132288_(_053214_, _042193_, _042237_);
  and g_132289_(_042054_, _042186_, _042238_);
  not g_132290_(_042238_, _042240_);
  or g_132291_(_042047_, _042186_, _042241_);
  not g_132292_(_042241_, _042242_);
  and g_132293_(_042240_, _042241_, _042243_);
  or g_132294_(_042238_, _042242_, _042244_);
  and g_132295_(_042236_, _042243_, _042245_);
  or g_132296_(_042237_, _042244_, _042246_);
  and g_132297_(_042024_, _042185_, _042247_);
  or g_132298_(_042025_, _042186_, _042248_);
  and g_132299_(_042032_, _042186_, _042249_);
  or g_132300_(_042031_, _042185_, _042251_);
  and g_132301_(_042248_, _042251_, _042252_);
  or g_132302_(_042247_, _042249_, _042253_);
  and g_132303_(out[289], _042253_, _042254_);
  not g_132304_(_042254_, _042255_);
  xor g_132305_(out[289], out[288], _042256_);
  xor g_132306_(_053225_, out[288], _042257_);
  and g_132307_(_042252_, _042256_, _042258_);
  or g_132308_(_042253_, _042257_, _042259_);
  and g_132309_(out[272], _042185_, _042260_);
  or g_132310_(_004443_, _042186_, _042262_);
  and g_132311_(_042040_, _042186_, _042263_);
  or g_132312_(_042039_, _042185_, _042264_);
  and g_132313_(_042262_, _042264_, _042265_);
  or g_132314_(_042260_, _042263_, _042266_);
  and g_132315_(out[288], _042265_, _042267_);
  or g_132316_(_004476_, _042266_, _042268_);
  and g_132317_(_042259_, _042268_, _042269_);
  or g_132318_(_042258_, _042267_, _042270_);
  and g_132319_(_042255_, _042270_, _042271_);
  or g_132320_(_042254_, _042269_, _042273_);
  and g_132321_(_042246_, _042273_, _042274_);
  or g_132322_(_042245_, _042271_, _042275_);
  and g_132323_(_042237_, _042244_, _042276_);
  or g_132324_(_042236_, _042243_, _042277_);
  xor g_132325_(out[291], _042194_, _042278_);
  xor g_132326_(_053192_, _042194_, _042279_);
  and g_132327_(_042073_, _042186_, _042280_);
  not g_132328_(_042280_, _042281_);
  or g_132329_(_042066_, _042186_, _042282_);
  not g_132330_(_042282_, _042284_);
  and g_132331_(_042281_, _042282_, _042285_);
  or g_132332_(_042280_, _042284_, _042286_);
  and g_132333_(_042278_, _042286_, _042287_);
  or g_132334_(_042279_, _042285_, _042288_);
  and g_132335_(_042277_, _042288_, _042289_);
  or g_132336_(_042276_, _042287_, _042290_);
  and g_132337_(_042275_, _042289_, _042291_);
  or g_132338_(_042274_, _042290_, _042292_);
  xor g_132339_(out[292], _042196_, _042293_);
  xor g_132340_(_053203_, _042196_, _042295_);
  and g_132341_(_042091_, _042186_, _042296_);
  not g_132342_(_042296_, _042297_);
  or g_132343_(_042083_, _042186_, _042298_);
  not g_132344_(_042298_, _042299_);
  and g_132345_(_042297_, _042298_, _042300_);
  or g_132346_(_042296_, _042299_, _042301_);
  and g_132347_(_042295_, _042300_, _042302_);
  or g_132348_(_042293_, _042301_, _042303_);
  and g_132349_(_042279_, _042285_, _042304_);
  or g_132350_(_042278_, _042286_, _042306_);
  and g_132351_(_042303_, _042306_, _042307_);
  or g_132352_(_042302_, _042304_, _042308_);
  and g_132353_(_042292_, _042307_, _042309_);
  or g_132354_(_042291_, _042308_, _042310_);
  xor g_132355_(out[293], _042197_, _042311_);
  xor g_132356_(_053170_, _042197_, _042312_);
  or g_132357_(_042099_, _042186_, _042313_);
  not g_132358_(_042313_, _042314_);
  and g_132359_(_042106_, _042186_, _042315_);
  not g_132360_(_042315_, _042317_);
  and g_132361_(_042313_, _042317_, _042318_);
  or g_132362_(_042314_, _042315_, _042319_);
  and g_132363_(_042311_, _042319_, _042320_);
  or g_132364_(_042312_, _042318_, _042321_);
  and g_132365_(_042293_, _042301_, _042322_);
  or g_132366_(_042295_, _042300_, _042323_);
  and g_132367_(_042321_, _042323_, _042324_);
  or g_132368_(_042320_, _042322_, _042325_);
  and g_132369_(_042310_, _042324_, _042326_);
  or g_132370_(_042309_, _042325_, _042328_);
  xor g_132371_(out[294], _042198_, _042329_);
  xor g_132372_(_053181_, _042198_, _042330_);
  and g_132373_(_042191_, _042329_, _042331_);
  or g_132374_(_042192_, _042330_, _042332_);
  and g_132375_(_042312_, _042318_, _042333_);
  or g_132376_(_042311_, _042319_, _042334_);
  and g_132377_(_042332_, _042334_, _042335_);
  or g_132378_(_042331_, _042333_, _042336_);
  and g_132379_(_042328_, _042335_, _042337_);
  or g_132380_(_042326_, _042336_, _042339_);
  and g_132381_(_042018_, _042186_, _042340_);
  not g_132382_(_042340_, _042341_);
  or g_132383_(_042020_, _042186_, _042342_);
  not g_132384_(_042342_, _042343_);
  and g_132385_(_042341_, _042342_, _042344_);
  or g_132386_(_042340_, _042343_, _042345_);
  xor g_132387_(out[295], _042199_, _042346_);
  xor g_132388_(_053148_, _042199_, _042347_);
  and g_132389_(_042345_, _042346_, _042348_);
  or g_132390_(_042344_, _042347_, _042350_);
  and g_132391_(_042192_, _042330_, _042351_);
  or g_132392_(_042191_, _042329_, _042352_);
  and g_132393_(_042350_, _042352_, _042353_);
  or g_132394_(_042348_, _042351_, _042354_);
  and g_132395_(_042339_, _042353_, _042355_);
  or g_132396_(_042337_, _042354_, _042356_);
  xor g_132397_(out[297], _042201_, _042357_);
  xor g_132398_(_053236_, _042201_, _042358_);
  and g_132399_(_042009_, _042186_, _042359_);
  not g_132400_(_042359_, _042361_);
  or g_132401_(_042005_, _042186_, _042362_);
  not g_132402_(_042362_, _042363_);
  and g_132403_(_042361_, _042362_, _042364_);
  or g_132404_(_042359_, _042363_, _042365_);
  and g_132405_(_042357_, _042364_, _042366_);
  or g_132406_(_042358_, _042365_, _042367_);
  and g_132407_(_042358_, _042365_, _042368_);
  or g_132408_(_042357_, _042364_, _042369_);
  xor g_132409_(out[296], _042200_, _042370_);
  xor g_132410_(_053159_, _042200_, _042372_);
  and g_132411_(_042001_, _042186_, _042373_);
  not g_132412_(_042373_, _042374_);
  or g_132413_(_041993_, _042186_, _042375_);
  not g_132414_(_042375_, _042376_);
  and g_132415_(_042374_, _042375_, _042377_);
  or g_132416_(_042373_, _042376_, _042378_);
  and g_132417_(_042372_, _042377_, _042379_);
  or g_132418_(_042370_, _042378_, _042380_);
  and g_132419_(_042370_, _042378_, _042381_);
  or g_132420_(_042372_, _042377_, _042383_);
  and g_132421_(_042344_, _042347_, _042384_);
  or g_132422_(_042345_, _042346_, _042385_);
  and g_132423_(_042369_, _042383_, _042386_);
  or g_132424_(_042368_, _042381_, _042387_);
  and g_132425_(_042234_, _042387_, _042388_);
  or g_132426_(_042235_, _042386_, _042389_);
  and g_132427_(_042367_, _042388_, _042390_);
  or g_132428_(_042366_, _042389_, _042391_);
  and g_132429_(_042367_, _042380_, _042392_);
  or g_132430_(_042366_, _042379_, _042394_);
  and g_132431_(_042369_, _042385_, _042395_);
  or g_132432_(_042368_, _042384_, _042396_);
  and g_132433_(_042392_, _042395_, _042397_);
  or g_132434_(_042394_, _042396_, _042398_);
  and g_132435_(_042234_, _042397_, _042399_);
  or g_132436_(_042235_, _042398_, _042400_);
  and g_132437_(_042383_, _042399_, _042401_);
  or g_132438_(_042381_, _042400_, _042402_);
  and g_132439_(_042356_, _042401_, _042403_);
  or g_132440_(_042355_, _042402_, _042405_);
  and g_132441_(_042229_, _042405_, _042406_);
  or g_132442_(_042227_, _042403_, _042407_);
  and g_132443_(_042391_, _042406_, _042408_);
  or g_132444_(_042390_, _042407_, _042409_);
  and g_132445_(_042192_, _042409_, _042410_);
  or g_132446_(_042191_, _042408_, _042411_);
  and g_132447_(_042329_, _042408_, _042412_);
  or g_132448_(_042330_, _042409_, _042413_);
  and g_132449_(_042411_, _042413_, _042414_);
  or g_132450_(_042410_, _042412_, _042416_);
  or g_132451_(out[305], out[304], _042417_);
  or g_132452_(out[304], _051956_, _042418_);
  xor g_132453_(out[306], _042417_, _042419_);
  xor g_132454_(_053313_, _042417_, _042420_);
  and g_132455_(_042244_, _042409_, _042421_);
  or g_132456_(_042243_, _042408_, _042422_);
  and g_132457_(_042236_, _042408_, _042423_);
  or g_132458_(_042237_, _042409_, _042424_);
  and g_132459_(_042422_, _042424_, _042425_);
  or g_132460_(_042421_, _042423_, _042427_);
  and g_132461_(_042419_, _042425_, _042428_);
  or g_132462_(_042420_, _042427_, _042429_);
  and g_132463_(_042256_, _042408_, _042430_);
  or g_132464_(_042257_, _042409_, _042431_);
  and g_132465_(_042253_, _042409_, _042432_);
  or g_132466_(_042252_, _042408_, _042433_);
  and g_132467_(_042431_, _042433_, _042434_);
  or g_132468_(_042430_, _042432_, _042435_);
  and g_132469_(out[305], _042435_, _042436_);
  not g_132470_(_042436_, _042438_);
  xor g_132471_(out[305], out[304], _042439_);
  xor g_132472_(_053324_, out[304], _042440_);
  and g_132473_(_042434_, _042439_, _042441_);
  or g_132474_(_042435_, _042440_, _042442_);
  and g_132475_(out[288], _042408_, _042443_);
  or g_132476_(_004476_, _042409_, _042444_);
  and g_132477_(_042266_, _042409_, _042445_);
  or g_132478_(_042265_, _042408_, _042446_);
  and g_132479_(_042444_, _042446_, _042447_);
  or g_132480_(_042443_, _042445_, _042449_);
  and g_132481_(out[304], _042447_, _042450_);
  or g_132482_(_004509_, _042449_, _042451_);
  and g_132483_(_042442_, _042451_, _042452_);
  or g_132484_(_042441_, _042450_, _042453_);
  and g_132485_(_042438_, _042453_, _042454_);
  or g_132486_(_042436_, _042452_, _042455_);
  and g_132487_(_042429_, _042455_, _042456_);
  or g_132488_(_042428_, _042454_, _042457_);
  and g_132489_(_042420_, _042427_, _042458_);
  or g_132490_(_042419_, _042425_, _042460_);
  and g_132491_(out[307], _042418_, _042461_);
  xor g_132492_(out[307], _042418_, _042462_);
  xor g_132493_(_053302_, _042418_, _042463_);
  and g_132494_(_042279_, _042408_, _042464_);
  or g_132495_(_042278_, _042409_, _042465_);
  and g_132496_(_042286_, _042409_, _042466_);
  or g_132497_(_042285_, _042408_, _042467_);
  and g_132498_(_042465_, _042467_, _042468_);
  or g_132499_(_042464_, _042466_, _042469_);
  and g_132500_(_042462_, _042469_, _042471_);
  or g_132501_(_042463_, _042468_, _042472_);
  and g_132502_(_042460_, _042472_, _042473_);
  or g_132503_(_042458_, _042471_, _042474_);
  and g_132504_(_042457_, _042473_, _042475_);
  or g_132505_(_042456_, _042474_, _042476_);
  and g_132506_(_019371_, _042418_, _042477_);
  xor g_132507_(out[308], _042461_, _042478_);
  xor g_132508_(_053291_, _042461_, _042479_);
  and g_132509_(_042295_, _042408_, _042480_);
  or g_132510_(_042293_, _042409_, _042482_);
  and g_132511_(_042301_, _042409_, _042483_);
  or g_132512_(_042300_, _042408_, _042484_);
  and g_132513_(_042482_, _042484_, _042485_);
  or g_132514_(_042480_, _042483_, _042486_);
  and g_132515_(_042479_, _042485_, _042487_);
  or g_132516_(_042478_, _042486_, _042488_);
  and g_132517_(_042463_, _042468_, _042489_);
  or g_132518_(_042462_, _042469_, _042490_);
  and g_132519_(_042488_, _042490_, _042491_);
  or g_132520_(_042487_, _042489_, _042493_);
  and g_132521_(_042476_, _042491_, _042494_);
  or g_132522_(_042475_, _042493_, _042495_);
  and g_132523_(out[309], _042477_, _042496_);
  xor g_132524_(out[309], _042477_, _042497_);
  xor g_132525_(_053269_, _042477_, _042498_);
  and g_132526_(_042312_, _042408_, _042499_);
  or g_132527_(_042311_, _042409_, _042500_);
  and g_132528_(_042319_, _042409_, _042501_);
  or g_132529_(_042318_, _042408_, _042502_);
  and g_132530_(_042500_, _042502_, _042504_);
  or g_132531_(_042499_, _042501_, _042505_);
  and g_132532_(_042497_, _042505_, _042506_);
  or g_132533_(_042498_, _042504_, _042507_);
  and g_132534_(_042478_, _042486_, _042508_);
  or g_132535_(_042479_, _042485_, _042509_);
  and g_132536_(_042507_, _042509_, _042510_);
  or g_132537_(_042506_, _042508_, _042511_);
  and g_132538_(_042495_, _042510_, _042512_);
  or g_132539_(_042494_, _042511_, _042513_);
  or g_132540_(out[310], _042496_, _042515_);
  xor g_132541_(out[310], _042496_, _042516_);
  xor g_132542_(_053280_, _042496_, _042517_);
  and g_132543_(_042414_, _042516_, _042518_);
  or g_132544_(_042416_, _042517_, _042519_);
  and g_132545_(_042498_, _042504_, _042520_);
  or g_132546_(_042497_, _042505_, _042521_);
  and g_132547_(_042519_, _042521_, _042522_);
  or g_132548_(_042518_, _042520_, _042523_);
  and g_132549_(_042513_, _042522_, _042524_);
  or g_132550_(_042512_, _042523_, _042526_);
  and g_132551_(_042345_, _042409_, _042527_);
  or g_132552_(_042344_, _042408_, _042528_);
  and g_132553_(_042347_, _042408_, _042529_);
  or g_132554_(_042346_, _042409_, _042530_);
  and g_132555_(_042528_, _042530_, _042531_);
  or g_132556_(_042527_, _042529_, _042532_);
  and g_132557_(out[311], _042515_, _042533_);
  xor g_132558_(out[311], _042515_, _042534_);
  xor g_132559_(_053247_, _042515_, _042535_);
  and g_132560_(_042532_, _042534_, _042537_);
  or g_132561_(_042531_, _042535_, _042538_);
  and g_132562_(_042416_, _042517_, _042539_);
  or g_132563_(_042414_, _042516_, _042540_);
  and g_132564_(_042538_, _042540_, _042541_);
  or g_132565_(_042537_, _042539_, _042542_);
  and g_132566_(_042526_, _042541_, _042543_);
  or g_132567_(_042524_, _042542_, _042544_);
  and g_132568_(_042531_, _042535_, _042545_);
  or g_132569_(_042532_, _042534_, _042546_);
  and g_132570_(out[312], _042533_, _042548_);
  or g_132571_(out[313], _042548_, _042549_);
  and g_132572_(out[314], _042549_, _042550_);
  xor g_132573_(out[314], _042549_, _042551_);
  xor g_132574_(_004520_, _042549_, _042552_);
  and g_132575_(_042216_, _042409_, _042553_);
  or g_132576_(_042215_, _042408_, _042554_);
  and g_132577_(_042219_, _042408_, _042555_);
  or g_132578_(_042218_, _042409_, _042556_);
  and g_132579_(_042554_, _042556_, _042557_);
  or g_132580_(_042553_, _042555_, _042559_);
  and g_132581_(_042552_, _042557_, _042560_);
  or g_132582_(_042551_, _042559_, _042561_);
  xor g_132583_(out[312], _042533_, _042562_);
  xor g_132584_(_053258_, _042533_, _042563_);
  and g_132585_(_042378_, _042409_, _042564_);
  or g_132586_(_042377_, _042408_, _042565_);
  and g_132587_(_042372_, _042408_, _042566_);
  or g_132588_(_042370_, _042409_, _042567_);
  and g_132589_(_042565_, _042567_, _042568_);
  or g_132590_(_042564_, _042566_, _042570_);
  and g_132591_(_042563_, _042568_, _042571_);
  or g_132592_(_042562_, _042570_, _042572_);
  and g_132593_(_042561_, _042572_, _042573_);
  or g_132594_(_042560_, _042571_, _042574_);
  and g_132595_(_042546_, _042573_, _042575_);
  or g_132596_(_042545_, _042574_, _042576_);
  and g_132597_(_042551_, _042559_, _042577_);
  or g_132598_(_042552_, _042557_, _042578_);
  xor g_132599_(out[315], _042550_, _042579_);
  xor g_132600_(_004498_, _042550_, _042581_);
  and g_132601_(_042204_, _042207_, _042582_);
  or g_132602_(_042205_, _042208_, _042583_);
  and g_132603_(_042204_, _042222_, _042584_);
  and g_132604_(_042579_, _042583_, _042585_);
  or g_132605_(_042581_, _042582_, _042586_);
  and g_132606_(_042578_, _042586_, _042587_);
  or g_132607_(_042577_, _042585_, _042588_);
  xor g_132608_(out[313], _042548_, _042589_);
  xor g_132609_(_053335_, _042548_, _042590_);
  and g_132610_(_042365_, _042409_, _042592_);
  or g_132611_(_042364_, _042408_, _042593_);
  and g_132612_(_042357_, _042408_, _042594_);
  or g_132613_(_042358_, _042409_, _042595_);
  and g_132614_(_042593_, _042595_, _042596_);
  or g_132615_(_042592_, _042594_, _042597_);
  and g_132616_(_042590_, _042597_, _042598_);
  or g_132617_(_042589_, _042596_, _042599_);
  and g_132618_(_042581_, _042582_, _042600_);
  or g_132619_(_042579_, _042583_, _042601_);
  and g_132620_(_042599_, _042601_, _042603_);
  or g_132621_(_042598_, _042600_, _042604_);
  and g_132622_(_042589_, _042596_, _042605_);
  or g_132623_(_042590_, _042597_, _042606_);
  and g_132624_(_042562_, _042570_, _042607_);
  or g_132625_(_042563_, _042568_, _042608_);
  and g_132626_(_042606_, _042608_, _042609_);
  or g_132627_(_042605_, _042607_, _042610_);
  and g_132628_(_042603_, _042609_, _042611_);
  or g_132629_(_042604_, _042610_, _042612_);
  and g_132630_(_042587_, _042611_, _042614_);
  or g_132631_(_042588_, _042612_, _042615_);
  and g_132632_(_042575_, _042614_, _042616_);
  or g_132633_(_042576_, _042615_, _042617_);
  and g_132634_(_042544_, _042616_, _042618_);
  or g_132635_(_042543_, _042617_, _042619_);
  and g_132636_(_042599_, _042608_, _042620_);
  or g_132637_(_042598_, _042607_, _042621_);
  and g_132638_(_042561_, _042606_, _042622_);
  or g_132639_(_042560_, _042605_, _042623_);
  and g_132640_(_042621_, _042622_, _042625_);
  or g_132641_(_042620_, _042623_, _042626_);
  and g_132642_(_042587_, _042626_, _042627_);
  or g_132643_(_042588_, _042625_, _042628_);
  and g_132644_(_042601_, _042628_, _042629_);
  or g_132645_(_042600_, _042627_, _042630_);
  and g_132646_(_042619_, _042630_, _042631_);
  or g_132647_(_042618_, _042629_, _042632_);
  and g_132648_(_042416_, _042632_, _042633_);
  or g_132649_(_042414_, _042631_, _042634_);
  and g_132650_(_042516_, _042631_, _042636_);
  or g_132651_(_042517_, _042632_, _042637_);
  and g_132652_(_042634_, _042637_, _042638_);
  or g_132653_(_042633_, _042636_, _042639_);
  and g_132654_(_038377_, _042638_, _042640_);
  or g_132655_(_038379_, _042639_, _042641_);
  xor g_132656_(out[327], _038371_, _042642_);
  xor g_132657_(_053346_, _038371_, _042643_);
  and g_132658_(_042532_, _042632_, _042644_);
  or g_132659_(_042531_, _042631_, _042645_);
  and g_132660_(_042535_, _042631_, _042647_);
  or g_132661_(_042534_, _042632_, _042648_);
  and g_132662_(_042645_, _042648_, _042649_);
  or g_132663_(_042644_, _042647_, _042650_);
  and g_132664_(_042643_, _042649_, _042651_);
  or g_132665_(_042642_, _042650_, _042652_);
  and g_132666_(_042641_, _042652_, _042653_);
  or g_132667_(_042640_, _042651_, _042654_);
  and g_132668_(_038379_, _042639_, _042655_);
  or g_132669_(_038377_, _042638_, _042656_);
  and g_132670_(_042642_, _042650_, _042658_);
  or g_132671_(_042643_, _042649_, _042659_);
  xor g_132672_(out[325], _038369_, _042660_);
  xor g_132673_(_053368_, _038369_, _042661_);
  and g_132674_(_042505_, _042632_, _042662_);
  not g_132675_(_042662_, _042663_);
  or g_132676_(_042497_, _042632_, _042664_);
  not g_132677_(_042664_, _042665_);
  and g_132678_(_042663_, _042664_, _042666_);
  or g_132679_(_042662_, _042665_, _042667_);
  and g_132680_(_042660_, _042667_, _042669_);
  or g_132681_(_042661_, _042666_, _042670_);
  and g_132682_(_042656_, _042659_, _042671_);
  or g_132683_(_042655_, _042658_, _042672_);
  and g_132684_(_042653_, _042671_, _042673_);
  or g_132685_(_042654_, _042672_, _042674_);
  and g_132686_(_042670_, _042673_, _042675_);
  or g_132687_(_042669_, _042674_, _042676_);
  xor g_132688_(out[324], _038368_, _042677_);
  xor g_132689_(_053401_, _038368_, _042678_);
  and g_132690_(_042486_, _042632_, _042680_);
  not g_132691_(_042680_, _042681_);
  or g_132692_(_042478_, _042632_, _042682_);
  not g_132693_(_042682_, _042683_);
  and g_132694_(_042681_, _042682_, _042684_);
  or g_132695_(_042680_, _042683_, _042685_);
  and g_132696_(_042678_, _042684_, _042686_);
  or g_132697_(_042677_, _042685_, _042687_);
  and g_132698_(_042661_, _042666_, _042688_);
  or g_132699_(_042660_, _042667_, _042689_);
  and g_132700_(_042687_, _042689_, _042691_);
  or g_132701_(_042686_, _042688_, _042692_);
  and g_132702_(_042677_, _042685_, _042693_);
  or g_132703_(_042678_, _042684_, _042694_);
  and g_132704_(_042691_, _042694_, _042695_);
  or g_132705_(_042692_, _042693_, _042696_);
  and g_132706_(_042675_, _042695_, _042697_);
  or g_132707_(_042676_, _042696_, _042698_);
  xor g_132708_(out[323], _038366_, _042699_);
  xor g_132709_(_053390_, _038366_, _042700_);
  and g_132710_(_042469_, _042632_, _042702_);
  not g_132711_(_042702_, _042703_);
  or g_132712_(_042462_, _042632_, _042704_);
  not g_132713_(_042704_, _042705_);
  and g_132714_(_042703_, _042704_, _042706_);
  or g_132715_(_042702_, _042705_, _042707_);
  and g_132716_(_042699_, _042707_, _042708_);
  or g_132717_(_042700_, _042706_, _042709_);
  and g_132718_(_042700_, _042706_, _042710_);
  or g_132719_(_042699_, _042707_, _042711_);
  xor g_132720_(out[322], _038365_, _042713_);
  xor g_132721_(_053412_, _038365_, _042714_);
  and g_132722_(_042427_, _042632_, _042715_);
  not g_132723_(_042715_, _042716_);
  or g_132724_(_042420_, _042632_, _042717_);
  not g_132725_(_042717_, _042718_);
  and g_132726_(_042716_, _042717_, _042719_);
  or g_132727_(_042715_, _042718_, _042720_);
  and g_132728_(_042713_, _042719_, _042721_);
  or g_132729_(_042714_, _042720_, _042722_);
  and g_132730_(_042711_, _042722_, _042724_);
  or g_132731_(_042710_, _042721_, _042725_);
  and g_132732_(_042709_, _042725_, _042726_);
  or g_132733_(_042708_, _042724_, _042727_);
  and g_132734_(_042439_, _042631_, _042728_);
  and g_132735_(_042435_, _042632_, _042729_);
  or g_132736_(_042728_, _042729_, _042730_);
  not g_132737_(_042730_, _042731_);
  xor g_132738_(out[321], out[320], _042732_);
  xor g_132739_(_053423_, out[320], _042733_);
  or g_132740_(_042730_, _042733_, _042735_);
  not g_132741_(_042735_, _042736_);
  and g_132742_(out[304], _042631_, _042737_);
  or g_132743_(_004509_, _042632_, _042738_);
  and g_132744_(_042449_, _042632_, _042739_);
  or g_132745_(_042447_, _042631_, _042740_);
  and g_132746_(_042738_, _042740_, _042741_);
  or g_132747_(_042737_, _042739_, _042742_);
  and g_132748_(_004542_, _042742_, _042743_);
  or g_132749_(out[320], _042741_, _042744_);
  xor g_132750_(_042730_, _042733_, _042746_);
  xor g_132751_(_042730_, _042732_, _042747_);
  and g_132752_(_042744_, _042746_, _042748_);
  or g_132753_(_042743_, _042747_, _042749_);
  and g_132754_(_042735_, _042749_, _042750_);
  or g_132755_(_042736_, _042748_, _042751_);
  and g_132756_(_042714_, _042720_, _042752_);
  or g_132757_(_042713_, _042719_, _042753_);
  and g_132758_(_042709_, _042753_, _042754_);
  or g_132759_(_042708_, _042752_, _042755_);
  and g_132760_(_042751_, _042754_, _042757_);
  or g_132761_(_042750_, _042755_, _042758_);
  and g_132762_(_042727_, _042758_, _042759_);
  or g_132763_(_042726_, _042757_, _042760_);
  and g_132764_(_042697_, _042760_, _042761_);
  or g_132765_(_042698_, _042759_, _042762_);
  and g_132766_(_042675_, _042692_, _042763_);
  or g_132767_(_042676_, _042691_, _042764_);
  and g_132768_(_042654_, _042659_, _042765_);
  or g_132769_(_042653_, _042658_, _042766_);
  and g_132770_(_042764_, _042766_, _042768_);
  or g_132771_(_042763_, _042765_, _042769_);
  and g_132772_(_042762_, _042768_, _042770_);
  or g_132773_(_042761_, _042769_, _042771_);
  and g_132774_(out[330], _038374_, _042772_);
  xor g_132775_(out[330], _038374_, _042773_);
  not g_132776_(_042773_, _042774_);
  and g_132777_(_042559_, _042632_, _042775_);
  not g_132778_(_042775_, _042776_);
  or g_132779_(_042551_, _042632_, _042777_);
  not g_132780_(_042777_, _042779_);
  and g_132781_(_042776_, _042777_, _042780_);
  or g_132782_(_042775_, _042779_, _042781_);
  and g_132783_(_042774_, _042780_, _042782_);
  or g_132784_(_042773_, _042781_, _042783_);
  xor g_132785_(out[331], _042772_, _042784_);
  xor g_132786_(_004531_, _042772_, _042785_);
  and g_132787_(_042579_, _042582_, _042786_);
  or g_132788_(_042581_, _042583_, _042787_);
  and g_132789_(_042785_, _042786_, _042788_);
  or g_132790_(_042784_, _042787_, _042790_);
  and g_132791_(_042783_, _042790_, _042791_);
  or g_132792_(_042782_, _042788_, _042792_);
  and g_132793_(_042579_, _042584_, _042793_);
  and g_132794_(_042784_, _042787_, _042794_);
  or g_132795_(_042785_, _042786_, _042795_);
  and g_132796_(_042773_, _042781_, _042796_);
  or g_132797_(_042774_, _042780_, _042797_);
  and g_132798_(_042795_, _042797_, _042798_);
  or g_132799_(_042794_, _042796_, _042799_);
  and g_132800_(_042791_, _042798_, _042801_);
  or g_132801_(_042792_, _042799_, _042802_);
  xor g_132802_(out[328], _038372_, _042803_);
  xor g_132803_(_053357_, _038372_, _042804_);
  and g_132804_(_042570_, _042632_, _042805_);
  not g_132805_(_042805_, _042806_);
  or g_132806_(_042562_, _042632_, _042807_);
  not g_132807_(_042807_, _042808_);
  and g_132808_(_042806_, _042807_, _042809_);
  or g_132809_(_042805_, _042808_, _042810_);
  and g_132810_(_042804_, _042809_, _042812_);
  or g_132811_(_042803_, _042810_, _042813_);
  and g_132812_(_042597_, _042632_, _042814_);
  not g_132813_(_042814_, _042815_);
  or g_132814_(_042590_, _042632_, _042816_);
  not g_132815_(_042816_, _042817_);
  and g_132816_(_042815_, _042816_, _042818_);
  or g_132817_(_042814_, _042817_, _042819_);
  and g_132818_(_038376_, _042819_, _042820_);
  or g_132819_(_038375_, _042818_, _042821_);
  and g_132820_(_042813_, _042821_, _042823_);
  or g_132821_(_042812_, _042820_, _042824_);
  and g_132822_(_038375_, _042818_, _042825_);
  or g_132823_(_038376_, _042819_, _042826_);
  and g_132824_(_042803_, _042810_, _042827_);
  or g_132825_(_042804_, _042809_, _042828_);
  and g_132826_(_042826_, _042828_, _042829_);
  or g_132827_(_042825_, _042827_, _042830_);
  and g_132828_(_042823_, _042829_, _042831_);
  or g_132829_(_042824_, _042830_, _042832_);
  and g_132830_(_042801_, _042831_, _042834_);
  or g_132831_(_042802_, _042832_, _042835_);
  and g_132832_(_042771_, _042834_, _042836_);
  or g_132833_(_042770_, _042835_, _042837_);
  and g_132834_(_042792_, _042795_, _042838_);
  or g_132835_(_042791_, _042794_, _042839_);
  and g_132836_(_042813_, _042826_, _042840_);
  or g_132837_(_042812_, _042825_, _042841_);
  and g_132838_(_042821_, _042841_, _042842_);
  or g_132839_(_042820_, _042840_, _042843_);
  and g_132840_(_042801_, _042842_, _042845_);
  or g_132841_(_042802_, _042843_, _042846_);
  and g_132842_(_042839_, _042846_, _042847_);
  or g_132843_(_042838_, _042845_, _042848_);
  and g_132844_(_042837_, _042847_, _042849_);
  or g_132845_(_042836_, _042848_, _042850_);
  and g_132846_(out[320], _042741_, _042851_);
  or g_132847_(_004542_, _042742_, _042852_);
  and g_132848_(_042724_, _042852_, _042853_);
  or g_132849_(_042725_, _042851_, _042854_);
  and g_132850_(_042754_, _042853_, _042856_);
  or g_132851_(_042755_, _042854_, _042857_);
  and g_132852_(_042748_, _042856_, _042858_);
  or g_132853_(_042749_, _042857_, _042859_);
  and g_132854_(_042697_, _042834_, _042860_);
  or g_132855_(_042698_, _042835_, _042861_);
  and g_132856_(_042858_, _042860_, _042862_);
  or g_132857_(_042859_, _042861_, _042863_);
  and g_132858_(_042850_, _042863_, _042864_);
  or g_132859_(_042849_, _042862_, _042865_);
  and g_132860_(_038375_, _042864_, _042867_);
  or g_132861_(_038376_, _042865_, _042868_);
  and g_132862_(_042819_, _042865_, _042869_);
  or g_132863_(_042818_, _042864_, _042870_);
  and g_132864_(_042868_, _042870_, _042871_);
  or g_132865_(_042867_, _042869_, _042872_);
  and g_132866_(_038364_, _042872_, _042873_);
  or g_132867_(_038363_, _042871_, _042874_);
  xor g_132868_(out[344], _038357_, _042875_);
  xor g_132869_(_053456_, _038357_, _042876_);
  and g_132870_(_042804_, _042864_, _042878_);
  or g_132871_(_042803_, _042865_, _042879_);
  and g_132872_(_042810_, _042865_, _042880_);
  or g_132873_(_042809_, _042864_, _042881_);
  and g_132874_(_042879_, _042881_, _042882_);
  or g_132875_(_042878_, _042880_, _042883_);
  and g_132876_(_042875_, _042883_, _042884_);
  or g_132877_(_042876_, _042882_, _042885_);
  and g_132878_(_042874_, _042885_, _042886_);
  or g_132879_(_042873_, _042884_, _042887_);
  and g_132880_(out[320], _042864_, _042889_);
  or g_132881_(_004542_, _042865_, _042890_);
  and g_132882_(_042742_, _042865_, _042891_);
  or g_132883_(_042741_, _042864_, _042892_);
  and g_132884_(_042890_, _042892_, _042893_);
  or g_132885_(_042889_, _042891_, _042894_);
  and g_132886_(out[336], _042893_, _042895_);
  or g_132887_(_004575_, _042894_, _042896_);
  and g_132888_(_042730_, _042865_, _042897_);
  or g_132889_(_042731_, _042864_, _042898_);
  and g_132890_(_042732_, _042864_, _042900_);
  or g_132891_(_042733_, _042865_, _042901_);
  and g_132892_(_042898_, _042901_, _042902_);
  or g_132893_(_042897_, _042900_, _042903_);
  and g_132894_(out[337], _042903_, _042904_);
  or g_132895_(_053522_, _042902_, _042905_);
  xor g_132896_(out[337], out[336], _042906_);
  xor g_132897_(_053522_, out[336], _042907_);
  and g_132898_(_042895_, _042905_, _042908_);
  or g_132899_(_042896_, _042904_, _042909_);
  xor g_132900_(out[338], _038350_, _042911_);
  xor g_132901_(_053511_, _038350_, _042912_);
  and g_132902_(_042713_, _042864_, _042913_);
  or g_132903_(_042714_, _042865_, _042914_);
  and g_132904_(_042720_, _042865_, _042915_);
  or g_132905_(_042719_, _042864_, _042916_);
  and g_132906_(_042914_, _042916_, _042917_);
  or g_132907_(_042913_, _042915_, _042918_);
  and g_132908_(_042911_, _042917_, _042919_);
  or g_132909_(_042912_, _042918_, _042920_);
  and g_132910_(_042902_, _042906_, _042922_);
  or g_132911_(_042903_, _042907_, _042923_);
  and g_132912_(_042920_, _042923_, _042924_);
  or g_132913_(_042919_, _042922_, _042925_);
  and g_132914_(_042909_, _042924_, _042926_);
  or g_132915_(_042908_, _042925_, _042927_);
  xor g_132916_(out[339], _038351_, _042928_);
  xor g_132917_(_053489_, _038351_, _042929_);
  and g_132918_(_042700_, _042864_, _042930_);
  or g_132919_(_042699_, _042865_, _042931_);
  and g_132920_(_042707_, _042865_, _042933_);
  or g_132921_(_042706_, _042864_, _042934_);
  and g_132922_(_042931_, _042934_, _042935_);
  or g_132923_(_042930_, _042933_, _042936_);
  and g_132924_(_042928_, _042936_, _042937_);
  or g_132925_(_042929_, _042935_, _042938_);
  and g_132926_(_042912_, _042918_, _042939_);
  or g_132927_(_042911_, _042917_, _042940_);
  and g_132928_(_042938_, _042940_, _042941_);
  or g_132929_(_042937_, _042939_, _042942_);
  and g_132930_(_042927_, _042941_, _042944_);
  or g_132931_(_042926_, _042942_, _042945_);
  xor g_132932_(out[340], _038352_, _042946_);
  xor g_132933_(_053500_, _038352_, _042947_);
  and g_132934_(_042678_, _042864_, _042948_);
  or g_132935_(_042677_, _042865_, _042949_);
  and g_132936_(_042685_, _042865_, _042950_);
  or g_132937_(_042684_, _042864_, _042951_);
  and g_132938_(_042949_, _042951_, _042952_);
  or g_132939_(_042948_, _042950_, _042953_);
  and g_132940_(_042947_, _042952_, _042955_);
  or g_132941_(_042946_, _042953_, _042956_);
  and g_132942_(_042929_, _042935_, _042957_);
  or g_132943_(_042928_, _042936_, _042958_);
  and g_132944_(_042956_, _042958_, _042959_);
  or g_132945_(_042955_, _042957_, _042960_);
  and g_132946_(_042945_, _042959_, _042961_);
  or g_132947_(_042944_, _042960_, _042962_);
  xor g_132948_(out[341], _038353_, _042963_);
  xor g_132949_(_053467_, _038353_, _042964_);
  and g_132950_(_042661_, _042864_, _042966_);
  or g_132951_(_042660_, _042865_, _042967_);
  and g_132952_(_042667_, _042865_, _042968_);
  or g_132953_(_042666_, _042864_, _042969_);
  and g_132954_(_042967_, _042969_, _042970_);
  or g_132955_(_042966_, _042968_, _042971_);
  and g_132956_(_042963_, _042971_, _042972_);
  or g_132957_(_042964_, _042970_, _042973_);
  and g_132958_(_042946_, _042953_, _042974_);
  or g_132959_(_042947_, _042952_, _042975_);
  and g_132960_(_042973_, _042975_, _042977_);
  or g_132961_(_042972_, _042974_, _042978_);
  and g_132962_(_042962_, _042977_, _042979_);
  or g_132963_(_042961_, _042978_, _042980_);
  xor g_132964_(out[342], _038354_, _042981_);
  xor g_132965_(_053478_, _038354_, _042982_);
  and g_132966_(_038377_, _042864_, _042983_);
  or g_132967_(_038379_, _042865_, _042984_);
  and g_132968_(_042639_, _042865_, _042985_);
  or g_132969_(_042638_, _042864_, _042986_);
  and g_132970_(_042984_, _042986_, _042988_);
  or g_132971_(_042983_, _042985_, _042989_);
  and g_132972_(_042981_, _042988_, _042990_);
  or g_132973_(_042982_, _042989_, _042991_);
  and g_132974_(_042964_, _042970_, _042992_);
  or g_132975_(_042963_, _042971_, _042993_);
  and g_132976_(_042991_, _042993_, _042994_);
  or g_132977_(_042990_, _042992_, _042995_);
  and g_132978_(_042980_, _042994_, _042996_);
  or g_132979_(_042979_, _042995_, _042997_);
  xor g_132980_(out[343], _038355_, _042999_);
  xor g_132981_(_053445_, _038355_, _043000_);
  and g_132982_(_042643_, _042864_, _043001_);
  or g_132983_(_042642_, _042865_, _043002_);
  and g_132984_(_042650_, _042865_, _043003_);
  or g_132985_(_042649_, _042864_, _043004_);
  and g_132986_(_043002_, _043004_, _043005_);
  or g_132987_(_043001_, _043003_, _043006_);
  and g_132988_(_042999_, _043006_, _043007_);
  or g_132989_(_043000_, _043005_, _043008_);
  and g_132990_(_042982_, _042989_, _043010_);
  or g_132991_(_042981_, _042988_, _043011_);
  and g_132992_(_043008_, _043011_, _043012_);
  or g_132993_(_043007_, _043010_, _043013_);
  and g_132994_(_042997_, _043012_, _043014_);
  or g_132995_(_042996_, _043013_, _043015_);
  and g_132996_(_043000_, _043005_, _043016_);
  or g_132997_(_042999_, _043006_, _043017_);
  and g_132998_(_042876_, _042882_, _043018_);
  or g_132999_(_042875_, _042883_, _043019_);
  and g_133000_(_043017_, _043019_, _043021_);
  or g_133001_(_043016_, _043018_, _043022_);
  and g_133002_(_043015_, _043021_, _043023_);
  or g_133003_(_043014_, _043022_, _043024_);
  and g_133004_(_042886_, _043024_, _043025_);
  or g_133005_(_042887_, _043023_, _043026_);
  xor g_133006_(out[347], _038360_, _043027_);
  xor g_133007_(_004564_, _038360_, _043028_);
  and g_133008_(_042785_, _042864_, _043029_);
  or g_133009_(_042784_, _042865_, _043030_);
  and g_133010_(_042787_, _042865_, _043032_);
  or g_133011_(_042786_, _042864_, _043033_);
  and g_133012_(_043030_, _043033_, _043034_);
  or g_133013_(_043029_, _043032_, _043035_);
  and g_133014_(_042793_, _042865_, _043036_);
  not g_133015_(_043036_, _043037_);
  and g_133016_(_042784_, _042864_, _043038_);
  or g_133017_(_042785_, _042865_, _043039_);
  and g_133018_(_043037_, _043039_, _043040_);
  or g_133019_(_043036_, _043038_, _043041_);
  and g_133020_(_043027_, _043035_, _043043_);
  or g_133021_(_043028_, _043041_, _043044_);
  and g_133022_(_043028_, _043034_, _043045_);
  or g_133023_(_043027_, _043035_, _043046_);
  or g_133024_(_042773_, _042865_, _043047_);
  not g_133025_(_043047_, _043048_);
  and g_133026_(_042781_, _042865_, _043049_);
  or g_133027_(_042780_, _042864_, _043050_);
  and g_133028_(_043047_, _043050_, _043051_);
  or g_133029_(_043048_, _043049_, _043052_);
  and g_133030_(_038361_, _043052_, _043054_);
  or g_133031_(_038362_, _043051_, _043055_);
  and g_133032_(_038363_, _042871_, _043056_);
  or g_133033_(_038364_, _042872_, _043057_);
  and g_133034_(_043044_, _043057_, _043058_);
  or g_133035_(_043043_, _043056_, _043059_);
  xor g_133036_(_038362_, _043051_, _043060_);
  xor g_133037_(_038361_, _043051_, _043061_);
  and g_133038_(_043046_, _043060_, _043062_);
  or g_133039_(_043045_, _043061_, _043063_);
  and g_133040_(_043058_, _043062_, _043065_);
  or g_133041_(_043059_, _043063_, _043066_);
  and g_133042_(_043026_, _043065_, _043067_);
  or g_133043_(_043025_, _043066_, _043068_);
  and g_133044_(_043046_, _043054_, _043069_);
  or g_133045_(_043045_, _043055_, _043070_);
  and g_133046_(_043044_, _043070_, _043071_);
  or g_133047_(_043043_, _043069_, _043072_);
  and g_133048_(_043068_, _043071_, _043073_);
  or g_133049_(_043067_, _043072_, _043074_);
  or g_133050_(_038361_, _043074_, _043076_);
  not g_133051_(_043076_, _043077_);
  and g_133052_(_043052_, _043074_, _043078_);
  not g_133053_(_043078_, _043079_);
  and g_133054_(_043076_, _043079_, _043080_);
  or g_133055_(_043077_, _043078_, _043081_);
  and g_133056_(_038349_, _043080_, _043082_);
  or g_133057_(_038348_, _043081_, _043083_);
  and g_133058_(_043027_, _043034_, _043084_);
  or g_133059_(_043028_, _043035_, _043085_);
  and g_133060_(_043027_, _043041_, _043087_);
  or g_133061_(_043028_, _043040_, _043088_);
  and g_133062_(_038347_, _043087_, _043089_);
  or g_133063_(_038346_, _043088_, _043090_);
  and g_133064_(_043083_, _043090_, _043091_);
  or g_133065_(_043082_, _043089_, _043092_);
  and g_133066_(_038348_, _043081_, _043093_);
  or g_133067_(_038349_, _043080_, _043094_);
  and g_133068_(_038346_, _043085_, _043095_);
  or g_133069_(_038347_, _043087_, _043096_);
  xor g_133070_(out[361], _038342_, _043098_);
  xor g_133071_(_053632_, _038342_, _043099_);
  or g_133072_(_038364_, _043074_, _043100_);
  not g_133073_(_043100_, _043101_);
  and g_133074_(_042872_, _043074_, _043102_);
  not g_133075_(_043102_, _043103_);
  and g_133076_(_043100_, _043103_, _043104_);
  or g_133077_(_043101_, _043102_, _043105_);
  and g_133078_(_043099_, _043105_, _043106_);
  or g_133079_(_043098_, _043104_, _043107_);
  and g_133080_(_043096_, _043107_, _043109_);
  or g_133081_(_043095_, _043106_, _043110_);
  and g_133082_(_043094_, _043109_, _043111_);
  or g_133083_(_043093_, _043110_, _043112_);
  and g_133084_(_043091_, _043111_, _043113_);
  or g_133085_(_043092_, _043112_, _043114_);
  xor g_133086_(out[360], _038341_, _043115_);
  xor g_133087_(_053555_, _038341_, _043116_);
  or g_133088_(_042875_, _043074_, _043117_);
  not g_133089_(_043117_, _043118_);
  and g_133090_(_042883_, _043074_, _043120_);
  not g_133091_(_043120_, _043121_);
  and g_133092_(_043117_, _043121_, _043122_);
  or g_133093_(_043118_, _043120_, _043123_);
  and g_133094_(_043116_, _043122_, _043124_);
  or g_133095_(_043115_, _043123_, _043125_);
  and g_133096_(_043098_, _043104_, _043126_);
  or g_133097_(_043099_, _043105_, _043127_);
  and g_133098_(_043125_, _043127_, _043128_);
  or g_133099_(_043124_, _043126_, _043129_);
  and g_133100_(_043115_, _043123_, _043131_);
  or g_133101_(_043116_, _043122_, _043132_);
  and g_133102_(_043128_, _043132_, _043133_);
  or g_133103_(_043129_, _043131_, _043134_);
  and g_133104_(_043113_, _043133_, _043135_);
  or g_133105_(_043114_, _043134_, _043136_);
  xor g_133106_(out[354], _038335_, _043137_);
  xor g_133107_(_053610_, _038335_, _043138_);
  or g_133108_(_042912_, _043074_, _043139_);
  not g_133109_(_043139_, _043140_);
  and g_133110_(_042918_, _043074_, _043142_);
  not g_133111_(_043142_, _043143_);
  and g_133112_(_043139_, _043143_, _043144_);
  or g_133113_(_043140_, _043142_, _043145_);
  and g_133114_(_043137_, _043144_, _043146_);
  or g_133115_(_043138_, _043145_, _043147_);
  xor g_133116_(out[355], _038336_, _043148_);
  xor g_133117_(_053588_, _038336_, _043149_);
  and g_133118_(_042936_, _043074_, _043150_);
  not g_133119_(_043150_, _043151_);
  or g_133120_(_042928_, _043074_, _043153_);
  not g_133121_(_043153_, _043154_);
  and g_133122_(_043151_, _043153_, _043155_);
  or g_133123_(_043150_, _043154_, _043156_);
  and g_133124_(_043149_, _043155_, _043157_);
  or g_133125_(_043148_, _043156_, _043158_);
  and g_133126_(_043147_, _043158_, _043159_);
  or g_133127_(_043146_, _043157_, _043160_);
  and g_133128_(_043138_, _043145_, _043161_);
  or g_133129_(_043137_, _043144_, _043162_);
  xor g_133130_(out[353], out[352], _043164_);
  not g_133131_(_043164_, _043165_);
  or g_133132_(_042907_, _043074_, _043166_);
  not g_133133_(_043166_, _043167_);
  and g_133134_(_042903_, _043074_, _043168_);
  not g_133135_(_043168_, _043169_);
  and g_133136_(_043166_, _043169_, _043170_);
  or g_133137_(_043167_, _043168_, _043171_);
  and g_133138_(_043164_, _043170_, _043172_);
  or g_133139_(_043165_, _043171_, _043173_);
  or g_133140_(_004575_, _043074_, _043175_);
  not g_133141_(_043175_, _043176_);
  and g_133142_(_042894_, _043074_, _043177_);
  not g_133143_(_043177_, _043178_);
  and g_133144_(_043175_, _043178_, _043179_);
  or g_133145_(_043176_, _043177_, _043180_);
  and g_133146_(_004608_, _043180_, _043181_);
  or g_133147_(out[352], _043179_, _043182_);
  xor g_133148_(_043164_, _043170_, _043183_);
  xor g_133149_(_043165_, _043170_, _043184_);
  and g_133150_(_043182_, _043183_, _043186_);
  or g_133151_(_043181_, _043184_, _043187_);
  and g_133152_(_043173_, _043187_, _043188_);
  or g_133153_(_043172_, _043186_, _043189_);
  and g_133154_(_043162_, _043189_, _043190_);
  or g_133155_(_043161_, _043188_, _043191_);
  and g_133156_(_043159_, _043191_, _043192_);
  or g_133157_(_043160_, _043190_, _043193_);
  xor g_133158_(out[358], _038339_, _043194_);
  xor g_133159_(_053577_, _038339_, _043195_);
  and g_133160_(_042981_, _043073_, _043197_);
  or g_133161_(_042982_, _043074_, _043198_);
  and g_133162_(_042989_, _043074_, _043199_);
  or g_133163_(_042988_, _043073_, _043200_);
  and g_133164_(_043198_, _043200_, _043201_);
  or g_133165_(_043197_, _043199_, _043202_);
  and g_133166_(_043194_, _043201_, _043203_);
  or g_133167_(_043195_, _043202_, _043204_);
  xor g_133168_(out[359], _038340_, _043205_);
  xor g_133169_(_053544_, _038340_, _043206_);
  and g_133170_(_043000_, _043073_, _043208_);
  or g_133171_(_042999_, _043074_, _043209_);
  and g_133172_(_043006_, _043074_, _043210_);
  or g_133173_(_043005_, _043073_, _043211_);
  and g_133174_(_043209_, _043211_, _043212_);
  or g_133175_(_043208_, _043210_, _043213_);
  and g_133176_(_043206_, _043212_, _043214_);
  or g_133177_(_043205_, _043213_, _043215_);
  and g_133178_(_043204_, _043215_, _043216_);
  or g_133179_(_043203_, _043214_, _043217_);
  xor g_133180_(out[357], _038338_, _043219_);
  xor g_133181_(_053566_, _038338_, _043220_);
  or g_133182_(_042963_, _043074_, _043221_);
  not g_133183_(_043221_, _043222_);
  and g_133184_(_042971_, _043074_, _043223_);
  not g_133185_(_043223_, _043224_);
  and g_133186_(_043221_, _043224_, _043225_);
  or g_133187_(_043222_, _043223_, _043226_);
  and g_133188_(_043219_, _043226_, _043227_);
  or g_133189_(_043220_, _043225_, _043228_);
  and g_133190_(_043205_, _043213_, _043230_);
  or g_133191_(_043206_, _043212_, _043231_);
  and g_133192_(_043195_, _043202_, _043232_);
  or g_133193_(_043194_, _043201_, _043233_);
  and g_133194_(_043216_, _043233_, _043234_);
  or g_133195_(_043217_, _043232_, _043235_);
  and g_133196_(_043228_, _043231_, _043236_);
  or g_133197_(_043227_, _043230_, _043237_);
  and g_133198_(_043234_, _043236_, _043238_);
  or g_133199_(_043235_, _043237_, _043239_);
  xor g_133200_(out[356], _038337_, _043241_);
  xor g_133201_(_053599_, _038337_, _043242_);
  and g_133202_(_042953_, _043074_, _043243_);
  not g_133203_(_043243_, _043244_);
  or g_133204_(_042946_, _043074_, _043245_);
  not g_133205_(_043245_, _043246_);
  and g_133206_(_043244_, _043245_, _043247_);
  or g_133207_(_043243_, _043246_, _043248_);
  and g_133208_(_043242_, _043247_, _043249_);
  or g_133209_(_043241_, _043248_, _043250_);
  and g_133210_(_043220_, _043225_, _043252_);
  or g_133211_(_043219_, _043226_, _043253_);
  and g_133212_(_043250_, _043253_, _043254_);
  or g_133213_(_043249_, _043252_, _043255_);
  and g_133214_(_043241_, _043248_, _043256_);
  or g_133215_(_043242_, _043247_, _043257_);
  and g_133216_(_043254_, _043257_, _043258_);
  or g_133217_(_043255_, _043256_, _043259_);
  and g_133218_(_043238_, _043258_, _043260_);
  or g_133219_(_043239_, _043259_, _043261_);
  and g_133220_(_043148_, _043156_, _043263_);
  or g_133221_(_043149_, _043155_, _043264_);
  and g_133222_(_043260_, _043264_, _043265_);
  or g_133223_(_043261_, _043263_, _043266_);
  and g_133224_(_043193_, _043265_, _043267_);
  or g_133225_(_043192_, _043266_, _043268_);
  and g_133226_(_043217_, _043231_, _043269_);
  or g_133227_(_043216_, _043230_, _043270_);
  and g_133228_(_043238_, _043255_, _043271_);
  or g_133229_(_043239_, _043254_, _043272_);
  and g_133230_(_043270_, _043272_, _043274_);
  or g_133231_(_043269_, _043271_, _043275_);
  and g_133232_(_043268_, _043274_, _043276_);
  or g_133233_(_043267_, _043275_, _043277_);
  and g_133234_(_043135_, _043277_, _043278_);
  or g_133235_(_043136_, _043276_, _043279_);
  and g_133236_(_043113_, _043129_, _043280_);
  or g_133237_(_043114_, _043128_, _043281_);
  and g_133238_(_043092_, _043096_, _043282_);
  or g_133239_(_043091_, _043095_, _043283_);
  and g_133240_(_043281_, _043283_, _043285_);
  or g_133241_(_043280_, _043282_, _043286_);
  and g_133242_(_043279_, _043285_, _043287_);
  or g_133243_(_043278_, _043286_, _043288_);
  and g_133244_(out[352], _043179_, _043289_);
  and g_133245_(_043159_, _043162_, _043290_);
  or g_133246_(_043160_, _043161_, _043291_);
  or g_133247_(_043263_, _043289_, _043292_);
  not g_133248_(_043292_, _043293_);
  and g_133249_(_043290_, _043293_, _043294_);
  or g_133250_(_043291_, _043292_, _043296_);
  and g_133251_(_043186_, _043294_, _043297_);
  or g_133252_(_043187_, _043296_, _043298_);
  and g_133253_(_043135_, _043297_, _043299_);
  or g_133254_(_043136_, _043298_, _043300_);
  and g_133255_(_043260_, _043299_, _043301_);
  or g_133256_(_043261_, _043300_, _043302_);
  and g_133257_(_043288_, _043302_, _043303_);
  or g_133258_(_043287_, _043301_, _043304_);
  and g_133259_(_038347_, _043303_, _043305_);
  or g_133260_(_038346_, _043304_, _043307_);
  and g_133261_(_043085_, _043304_, _043308_);
  or g_133262_(_043084_, _043303_, _043309_);
  and g_133263_(_043307_, _043309_, _043310_);
  or g_133264_(_043305_, _043308_, _043311_);
  and g_133265_(_038332_, _043310_, _043312_);
  or g_133266_(_038333_, _043311_, _043313_);
  and g_133267_(_038319_, _043312_, _043314_);
  or g_133268_(_038320_, _043313_, _043315_);
  and g_133269_(_038306_, _043314_, _043316_);
  or g_133270_(_038307_, _043315_, _043318_);
  and g_133271_(_038293_, _043316_, _043319_);
  or g_133272_(_038294_, _043318_, _043320_);
  and g_133273_(_038280_, _043319_, _043321_);
  not g_133274_(_043321_, _043322_);
  and g_133275_(_038266_, _043321_, _043323_);
  not g_133276_(_043323_, _043324_);
  or g_133277_(out[945], out[944], _043325_);
  or g_133278_(out[944], _002904_, _043326_);
  and g_133279_(out[947], _043326_, _043327_);
  and g_133280_(_027322_, _043326_, _043329_);
  and g_133281_(out[949], _043329_, _043330_);
  or g_133282_(out[950], _043330_, _043331_);
  and g_133283_(out[951], _043331_, _043332_);
  and g_133284_(out[952], _043332_, _043333_);
  or g_133285_(out[953], _043333_, _043334_);
  and g_133286_(out[954], _043334_, _043335_);
  xor g_133287_(out[955], _043335_, _043336_);
  not g_133288_(_043336_, _043337_);
  xor g_133289_(out[950], _043330_, _043338_);
  not g_133290_(_043338_, _043340_);
  or g_133291_(out[865], out[864], _043341_);
  or g_133292_(out[864], _002016_, _043342_);
  and g_133293_(out[867], _043342_, _043343_);
  and g_133294_(_026347_, _043342_, _043344_);
  and g_133295_(out[869], _043344_, _043345_);
  or g_133296_(out[870], _043345_, _043346_);
  xor g_133297_(out[870], _043345_, _043347_);
  xor g_133298_(_001572_, _043345_, _043348_);
  and g_133299_(out[871], _043346_, _043349_);
  xor g_133300_(out[871], _043346_, _043351_);
  xor g_133301_(_001561_, _043346_, _043352_);
  or g_133302_(out[849], out[848], _043353_);
  or g_133303_(out[848], _001844_, _043354_);
  and g_133304_(out[851], _043354_, _043355_);
  and g_133305_(_026144_, _043354_, _043356_);
  and g_133306_(out[853], _043356_, _043357_);
  or g_133307_(out[854], _043357_, _043358_);
  and g_133308_(out[855], _043358_, _043359_);
  xor g_133309_(_001429_, _043358_, _043360_);
  not g_133310_(_043360_, _043362_);
  xor g_133311_(out[851], _043354_, _043363_);
  xor g_133312_(_001506_, _043354_, _043364_);
  or g_133313_(out[833], out[832], _043365_);
  or g_133314_(out[832], _001514_, _043366_);
  and g_133315_(out[835], _043366_, _043367_);
  xor g_133316_(out[835], _043366_, _043368_);
  xor g_133317_(_001374_, _043366_, _043369_);
  and g_133318_(_025997_, _043366_, _043370_);
  and g_133319_(out[837], _043370_, _043371_);
  or g_133320_(out[838], _043371_, _043373_);
  and g_133321_(out[839], _043373_, _043374_);
  xor g_133322_(out[839], _043373_, _043375_);
  not g_133323_(_043375_, _043376_);
  or g_133324_(out[817], out[816], _043377_);
  or g_133325_(out[816], _001338_, _043378_);
  and g_133326_(out[819], _043378_, _043379_);
  and g_133327_(_025751_, _043378_, _043380_);
  and g_133328_(out[821], _043380_, _043381_);
  or g_133329_(out[822], _043381_, _043382_);
  and g_133330_(out[823], _043382_, _043384_);
  xor g_133331_(out[823], _043382_, _043385_);
  not g_133332_(_043385_, _043386_);
  xor g_133333_(out[820], _043379_, _043387_);
  xor g_133334_(_001198_, _043379_, _043388_);
  or g_133335_(out[785], out[784], _043389_);
  or g_133336_(out[784], _001009_, _043390_);
  and g_133337_(out[787], _043390_, _043391_);
  and g_133338_(_025352_, _043390_, _043392_);
  xor g_133339_(out[788], _043391_, _043393_);
  xor g_133340_(_000934_, _043391_, _043395_);
  and g_133341_(out[789], _043392_, _043396_);
  or g_133342_(out[790], _043396_, _043397_);
  and g_133343_(out[791], _043397_, _043398_);
  and g_133344_(out[792], _043398_, _043399_);
  or g_133345_(out[793], _043399_, _043400_);
  and g_133346_(out[794], _043400_, _043401_);
  xor g_133347_(out[794], _043400_, _043402_);
  or g_133348_(out[737], out[736], _043403_);
  or g_133349_(out[736], _000361_, _043404_);
  and g_133350_(out[739], _043404_, _043406_);
  and g_133351_(_024779_, _043404_, _043407_);
  and g_133352_(out[741], _043407_, _043408_);
  or g_133353_(out[742], _043408_, _043409_);
  and g_133354_(out[743], _043409_, _043410_);
  and g_133355_(out[744], _043410_, _043411_);
  or g_133356_(out[745], _043411_, _043412_);
  and g_133357_(out[746], _043412_, _043413_);
  xor g_133358_(out[746], _043412_, _043414_);
  not g_133359_(_043414_, _043415_);
  xor g_133360_(out[743], _043409_, _043417_);
  xor g_133361_(_000505_, _043409_, _043418_);
  or g_133362_(out[657], out[656], _043419_);
  or g_133363_(out[656], _055437_, _043420_);
  and g_133364_(out[659], _043420_, _043421_);
  and g_133365_(_023710_, _043420_, _043422_);
  and g_133366_(out[661], _043422_, _043423_);
  or g_133367_(out[662], _043423_, _043424_);
  and g_133368_(out[663], _043424_, _043425_);
  xor g_133369_(out[663], _043424_, _043426_);
  xor g_133370_(_055810_, _043424_, _043428_);
  and g_133371_(out[664], _043425_, _043429_);
  or g_133372_(out[665], _043429_, _043430_);
  and g_133373_(out[666], _043430_, _043431_);
  xor g_133374_(out[666], _043430_, _043432_);
  xor g_133375_(_055920_, _043430_, _043433_);
  or g_133376_(out[513], out[512], _043434_);
  or g_133377_(out[512], _019073_, _043435_);
  and g_133378_(out[515], _043435_, _043436_);
  and g_133379_(_021667_, _043435_, _043437_);
  and g_133380_(out[517], _043437_, _043439_);
  or g_133381_(out[518], _043439_, _043440_);
  and g_133382_(out[519], _043440_, _043441_);
  and g_133383_(out[520], _043441_, _043442_);
  or g_133384_(out[521], _043442_, _043443_);
  and g_133385_(out[522], _043443_, _043444_);
  xor g_133386_(out[522], _043443_, _043445_);
  xor g_133387_(_054732_, _043443_, _043446_);
  and g_133388_(_054534_, _054545_, _043447_);
  or g_133389_(out[497], out[496], _043448_);
  or g_133390_(out[496], _016356_, _043450_);
  and g_133391_(out[499], _043450_, _043451_);
  and g_133392_(_021530_, _043450_, _043452_);
  and g_133393_(out[501], _043452_, _043453_);
  or g_133394_(out[502], _043453_, _043454_);
  and g_133395_(out[503], _043454_, _043455_);
  and g_133396_(out[504], _043455_, _043456_);
  or g_133397_(out[505], _043456_, _043457_);
  and g_133398_(out[506], _043457_, _043458_);
  xor g_133399_(out[506], _043457_, _043459_);
  xor g_133400_(_054600_, _043457_, _043461_);
  or g_133401_(out[480], _016389_, _043462_);
  and g_133402_(out[483], _043462_, _043463_);
  not g_133403_(_043463_, _043464_);
  and g_133404_(_021520_, _043462_, _043465_);
  and g_133405_(out[485], _043465_, _043466_);
  or g_133406_(out[486], _043466_, _043467_);
  and g_133407_(out[487], _043467_, _043468_);
  and g_133408_(out[488], _043468_, _043469_);
  or g_133409_(out[489], _043469_, _043470_);
  and g_133410_(out[490], _043470_, _043472_);
  xor g_133411_(out[491], _043472_, _043473_);
  xor g_133412_(_054358_, _043472_, _043474_);
  xor g_133413_(out[507], _043458_, _043475_);
  xor g_133414_(_054479_, _043458_, _043476_);
  and g_133415_(_043474_, _043475_, _043477_);
  or g_133416_(_043473_, _043476_, _043478_);
  xor g_133417_(out[488], _043468_, _043479_);
  xor g_133418_(_054446_, _043468_, _043480_);
  xor g_133419_(out[504], _043455_, _043481_);
  xor g_133420_(_054578_, _043455_, _043483_);
  and g_133421_(_043480_, _043481_, _043484_);
  or g_133422_(_043479_, _043483_, _043485_);
  and g_133423_(out[481], out[497], _043486_);
  not g_133424_(_043486_, _043487_);
  and g_133425_(_016851_, _043486_, _043488_);
  or g_133426_(_016840_, _043487_, _043489_);
  and g_133427_(out[480], _054413_, _043490_);
  or g_133428_(_054347_, out[481], _043491_);
  and g_133429_(_043448_, _043491_, _043492_);
  or g_133430_(_043447_, _043490_, _043494_);
  and g_133431_(_043489_, _043492_, _043495_);
  or g_133432_(_043488_, _043494_, _043496_);
  xor g_133433_(out[498], _043448_, _043497_);
  xor g_133434_(_054556_, _043448_, _043498_);
  or g_133435_(out[480], _016400_, _043499_);
  not g_133436_(_043499_, _043500_);
  and g_133437_(out[480], out[482], _043501_);
  not g_133438_(_043501_, _043502_);
  or g_133439_(_043500_, _043501_, _043503_);
  and g_133440_(_043499_, _043502_, _043505_);
  or g_133441_(out[480], _009411_, _043506_);
  not g_133442_(_043506_, _043507_);
  and g_133443_(_043464_, _043506_, _043508_);
  or g_133444_(_043463_, _043507_, _043509_);
  xor g_133445_(out[499], _043450_, _043510_);
  xor g_133446_(_054567_, _043450_, _043511_);
  and g_133447_(_043509_, _043510_, _043512_);
  or g_133448_(_043508_, _043511_, _043513_);
  and g_133449_(_043496_, _043498_, _043514_);
  or g_133450_(_043495_, _043497_, _043516_);
  and g_133451_(_043495_, _043497_, _043517_);
  or g_133452_(_043496_, _043498_, _043518_);
  and g_133453_(_043503_, _043516_, _043519_);
  or g_133454_(_043505_, _043514_, _043520_);
  and g_133455_(_043518_, _043520_, _043521_);
  or g_133456_(_043517_, _043519_, _043522_);
  and g_133457_(_043513_, _043522_, _043523_);
  or g_133458_(_043512_, _043521_, _043524_);
  xor g_133459_(out[484], _043463_, _043525_);
  xor g_133460_(_054402_, _043463_, _043527_);
  xor g_133461_(out[500], _043451_, _043528_);
  xor g_133462_(_054523_, _043451_, _043529_);
  and g_133463_(_043525_, _043529_, _043530_);
  or g_133464_(_043527_, _043528_, _043531_);
  and g_133465_(_043508_, _043511_, _043532_);
  or g_133466_(_043509_, _043510_, _043533_);
  and g_133467_(_043531_, _043533_, _043534_);
  or g_133468_(_043530_, _043532_, _043535_);
  and g_133469_(_043524_, _043534_, _043536_);
  or g_133470_(_043523_, _043535_, _043538_);
  and g_133471_(_043527_, _043528_, _043539_);
  or g_133472_(_043525_, _043529_, _043540_);
  xor g_133473_(out[485], _043465_, _043541_);
  xor g_133474_(_054391_, _043465_, _043542_);
  xor g_133475_(out[501], _043452_, _043543_);
  xor g_133476_(_054512_, _043452_, _043544_);
  and g_133477_(_043542_, _043543_, _043545_);
  or g_133478_(_043541_, _043544_, _043546_);
  and g_133479_(_043540_, _043546_, _043547_);
  or g_133480_(_043539_, _043545_, _043549_);
  and g_133481_(_043538_, _043547_, _043550_);
  or g_133482_(_043536_, _043549_, _043551_);
  xor g_133483_(out[486], _043466_, _043552_);
  xor g_133484_(_054380_, _043466_, _043553_);
  xor g_133485_(out[502], _043453_, _043554_);
  xor g_133486_(_054501_, _043453_, _043555_);
  and g_133487_(_043553_, _043554_, _043556_);
  or g_133488_(_043552_, _043555_, _043557_);
  and g_133489_(_043541_, _043544_, _043558_);
  or g_133490_(_043542_, _043543_, _043560_);
  and g_133491_(_043557_, _043560_, _043561_);
  or g_133492_(_043556_, _043558_, _043562_);
  and g_133493_(_043551_, _043561_, _043563_);
  or g_133494_(_043550_, _043562_, _043564_);
  xor g_133495_(out[487], _043467_, _043565_);
  xor g_133496_(_054369_, _043467_, _043566_);
  xor g_133497_(out[503], _043454_, _043567_);
  xor g_133498_(_054490_, _043454_, _043568_);
  and g_133499_(_043566_, _043567_, _043569_);
  or g_133500_(_043565_, _043568_, _043571_);
  and g_133501_(_043552_, _043555_, _043572_);
  or g_133502_(_043553_, _043554_, _043573_);
  and g_133503_(_043571_, _043573_, _043574_);
  or g_133504_(_043569_, _043572_, _043575_);
  and g_133505_(_043564_, _043574_, _043576_);
  or g_133506_(_043563_, _043575_, _043577_);
  and g_133507_(_043565_, _043568_, _043578_);
  or g_133508_(_043566_, _043567_, _043579_);
  xor g_133509_(out[489], _043469_, _043580_);
  xor g_133510_(_054457_, _043469_, _043582_);
  xor g_133511_(out[505], _043456_, _043583_);
  xor g_133512_(_054589_, _043456_, _043584_);
  and g_133513_(_043582_, _043583_, _043585_);
  or g_133514_(_043580_, _043584_, _043586_);
  and g_133515_(_043479_, _043483_, _043587_);
  or g_133516_(_043480_, _043481_, _043588_);
  and g_133517_(_043579_, _043588_, _043589_);
  or g_133518_(_043578_, _043587_, _043590_);
  and g_133519_(_043577_, _043589_, _043591_);
  or g_133520_(_043576_, _043590_, _043593_);
  and g_133521_(_043485_, _043593_, _043594_);
  or g_133522_(_043484_, _043591_, _043595_);
  and g_133523_(_043586_, _043595_, _043596_);
  or g_133524_(_043585_, _043594_, _043597_);
  and g_133525_(_043580_, _043584_, _043598_);
  or g_133526_(_043582_, _043583_, _043599_);
  xor g_133527_(out[490], _043470_, _043600_);
  xor g_133528_(_054468_, _043470_, _043601_);
  and g_133529_(_043459_, _043601_, _043602_);
  or g_133530_(_043461_, _043600_, _043604_);
  and g_133531_(_043599_, _043604_, _043605_);
  or g_133532_(_043598_, _043602_, _043606_);
  and g_133533_(_043597_, _043605_, _043607_);
  or g_133534_(_043596_, _043606_, _043608_);
  and g_133535_(_043461_, _043600_, _043609_);
  or g_133536_(_043459_, _043601_, _043610_);
  and g_133537_(_043473_, _043476_, _043611_);
  or g_133538_(_043474_, _043475_, _043612_);
  and g_133539_(_043610_, _043612_, _043613_);
  or g_133540_(_043609_, _043611_, _043615_);
  and g_133541_(_043608_, _043613_, _043616_);
  or g_133542_(_043607_, _043615_, _043617_);
  and g_133543_(_043478_, _043617_, _043618_);
  or g_133544_(_043477_, _043616_, _043619_);
  and g_133545_(_043461_, _043618_, _043620_);
  or g_133546_(_043459_, _043619_, _043621_);
  and g_133547_(_043601_, _043619_, _043622_);
  or g_133548_(_043600_, _043618_, _043623_);
  and g_133549_(_043621_, _043623_, _043624_);
  or g_133550_(_043620_, _043622_, _043626_);
  and g_133551_(_043445_, _043626_, _043627_);
  or g_133552_(_043446_, _043624_, _043628_);
  and g_133553_(_043473_, _043475_, _043629_);
  or g_133554_(_043474_, _043476_, _043630_);
  xor g_133555_(out[523], _043444_, _043631_);
  xor g_133556_(_054611_, _043444_, _043632_);
  and g_133557_(_043630_, _043631_, _043633_);
  or g_133558_(_043629_, _043632_, _043634_);
  and g_133559_(_043628_, _043634_, _043635_);
  or g_133560_(_043627_, _043633_, _043637_);
  and g_133561_(_043629_, _043632_, _043638_);
  or g_133562_(_043630_, _043631_, _043639_);
  and g_133563_(_043637_, _043639_, _043640_);
  or g_133564_(_043635_, _043638_, _043641_);
  xor g_133565_(out[521], _043442_, _043642_);
  xor g_133566_(_054721_, _043442_, _043643_);
  and g_133567_(_043583_, _043618_, _043644_);
  or g_133568_(_043584_, _043619_, _043645_);
  and g_133569_(_043580_, _043619_, _043646_);
  or g_133570_(_043582_, _043618_, _043648_);
  and g_133571_(_043645_, _043648_, _043649_);
  or g_133572_(_043644_, _043646_, _043650_);
  and g_133573_(_043643_, _043650_, _043651_);
  or g_133574_(_043642_, _043649_, _043652_);
  xor g_133575_(out[520], _043441_, _043653_);
  not g_133576_(_043653_, _043654_);
  and g_133577_(_043483_, _043618_, _043655_);
  or g_133578_(_043481_, _043619_, _043656_);
  and g_133579_(_043480_, _043619_, _043657_);
  or g_133580_(_043479_, _043618_, _043659_);
  and g_133581_(_043656_, _043659_, _043660_);
  or g_133582_(_043655_, _043657_, _043661_);
  and g_133583_(_043653_, _043661_, _043662_);
  or g_133584_(_043654_, _043660_, _043663_);
  xor g_133585_(out[514], _043434_, _043664_);
  xor g_133586_(_054688_, _043434_, _043665_);
  and g_133587_(_043505_, _043619_, _043666_);
  or g_133588_(_043503_, _043618_, _043667_);
  and g_133589_(_043497_, _043618_, _043668_);
  or g_133590_(_043498_, _043619_, _043670_);
  and g_133591_(_043667_, _043670_, _043671_);
  or g_133592_(_043666_, _043668_, _043672_);
  and g_133593_(_043664_, _043671_, _043673_);
  or g_133594_(_043665_, _043672_, _043674_);
  xor g_133595_(_054347_, out[481], _043675_);
  xor g_133596_(out[480], out[481], _043676_);
  and g_133597_(_043619_, _043676_, _043677_);
  or g_133598_(_043618_, _043675_, _043678_);
  xor g_133599_(out[497], out[496], _043679_);
  xor g_133600_(_054534_, out[496], _043681_);
  and g_133601_(_043618_, _043679_, _043682_);
  or g_133602_(_043619_, _043681_, _043683_);
  and g_133603_(_043678_, _043683_, _043684_);
  or g_133604_(_043677_, _043682_, _043685_);
  and g_133605_(out[513], _043685_, _043686_);
  not g_133606_(_043686_, _043687_);
  xor g_133607_(out[513], out[512], _043688_);
  xor g_133608_(_054666_, out[512], _043689_);
  and g_133609_(_043684_, _043688_, _043690_);
  or g_133610_(_043685_, _043689_, _043692_);
  and g_133611_(out[496], _043618_, _043693_);
  or g_133612_(_054545_, _043619_, _043694_);
  and g_133613_(out[480], _043619_, _043695_);
  or g_133614_(_054347_, _043618_, _043696_);
  and g_133615_(_043694_, _043696_, _043697_);
  or g_133616_(_043693_, _043695_, _043698_);
  and g_133617_(out[512], _043697_, _043699_);
  or g_133618_(_054677_, _043698_, _043700_);
  and g_133619_(_043692_, _043700_, _043701_);
  or g_133620_(_043690_, _043699_, _043703_);
  and g_133621_(_043687_, _043703_, _043704_);
  or g_133622_(_043686_, _043701_, _043705_);
  and g_133623_(_043674_, _043705_, _043706_);
  or g_133624_(_043673_, _043704_, _043707_);
  and g_133625_(_043665_, _043672_, _043708_);
  or g_133626_(_043664_, _043671_, _043709_);
  xor g_133627_(out[515], _043435_, _043710_);
  xor g_133628_(_054699_, _043435_, _043711_);
  and g_133629_(_043511_, _043618_, _043712_);
  or g_133630_(_043510_, _043619_, _043714_);
  and g_133631_(_043509_, _043619_, _043715_);
  or g_133632_(_043508_, _043618_, _043716_);
  and g_133633_(_043714_, _043716_, _043717_);
  or g_133634_(_043712_, _043715_, _043718_);
  and g_133635_(_043710_, _043718_, _043719_);
  or g_133636_(_043711_, _043717_, _043720_);
  and g_133637_(_043709_, _043720_, _043721_);
  or g_133638_(_043708_, _043719_, _043722_);
  and g_133639_(_043707_, _043721_, _043723_);
  or g_133640_(_043706_, _043722_, _043725_);
  xor g_133641_(out[516], _043436_, _043726_);
  xor g_133642_(_054655_, _043436_, _043727_);
  and g_133643_(_043527_, _043619_, _043728_);
  or g_133644_(_043525_, _043618_, _043729_);
  and g_133645_(_043529_, _043618_, _043730_);
  or g_133646_(_043528_, _043619_, _043731_);
  and g_133647_(_043729_, _043731_, _043732_);
  or g_133648_(_043728_, _043730_, _043733_);
  and g_133649_(_043727_, _043732_, _043734_);
  or g_133650_(_043726_, _043733_, _043736_);
  and g_133651_(_043711_, _043717_, _043737_);
  or g_133652_(_043710_, _043718_, _043738_);
  and g_133653_(_043736_, _043738_, _043739_);
  or g_133654_(_043734_, _043737_, _043740_);
  and g_133655_(_043725_, _043739_, _043741_);
  or g_133656_(_043723_, _043740_, _043742_);
  and g_133657_(_043726_, _043733_, _043743_);
  or g_133658_(_043727_, _043732_, _043744_);
  xor g_133659_(out[517], _043437_, _043745_);
  xor g_133660_(_054644_, _043437_, _043747_);
  and g_133661_(_043542_, _043619_, _043748_);
  or g_133662_(_043541_, _043618_, _043749_);
  and g_133663_(_043544_, _043618_, _043750_);
  or g_133664_(_043543_, _043619_, _043751_);
  and g_133665_(_043749_, _043751_, _043752_);
  or g_133666_(_043748_, _043750_, _043753_);
  and g_133667_(_043745_, _043753_, _043754_);
  or g_133668_(_043747_, _043752_, _043755_);
  and g_133669_(_043744_, _043755_, _043756_);
  or g_133670_(_043743_, _043754_, _043758_);
  and g_133671_(_043742_, _043756_, _043759_);
  or g_133672_(_043741_, _043758_, _043760_);
  xor g_133673_(out[518], _043439_, _043761_);
  xor g_133674_(_054633_, _043439_, _043762_);
  and g_133675_(_043554_, _043618_, _043763_);
  or g_133676_(_043555_, _043619_, _043764_);
  and g_133677_(_043552_, _043619_, _043765_);
  or g_133678_(_043553_, _043618_, _043766_);
  and g_133679_(_043764_, _043766_, _043767_);
  or g_133680_(_043763_, _043765_, _043769_);
  and g_133681_(_043761_, _043767_, _043770_);
  or g_133682_(_043762_, _043769_, _043771_);
  and g_133683_(_043747_, _043752_, _043772_);
  or g_133684_(_043745_, _043753_, _043773_);
  and g_133685_(_043771_, _043773_, _043774_);
  or g_133686_(_043770_, _043772_, _043775_);
  and g_133687_(_043760_, _043774_, _043776_);
  or g_133688_(_043759_, _043775_, _043777_);
  xor g_133689_(out[519], _043440_, _043778_);
  xor g_133690_(_054622_, _043440_, _043780_);
  and g_133691_(_043568_, _043618_, _043781_);
  or g_133692_(_043567_, _043619_, _043782_);
  and g_133693_(_043566_, _043619_, _043783_);
  or g_133694_(_043565_, _043618_, _043784_);
  and g_133695_(_043782_, _043784_, _043785_);
  or g_133696_(_043781_, _043783_, _043786_);
  and g_133697_(_043778_, _043786_, _043787_);
  or g_133698_(_043780_, _043785_, _043788_);
  and g_133699_(_043762_, _043769_, _043789_);
  or g_133700_(_043761_, _043767_, _043791_);
  and g_133701_(_043788_, _043791_, _043792_);
  or g_133702_(_043787_, _043789_, _043793_);
  and g_133703_(_043777_, _043792_, _043794_);
  or g_133704_(_043776_, _043793_, _043795_);
  and g_133705_(_043780_, _043785_, _043796_);
  or g_133706_(_043778_, _043786_, _043797_);
  and g_133707_(_043446_, _043624_, _043798_);
  or g_133708_(_043445_, _043626_, _043799_);
  and g_133709_(_043642_, _043649_, _043800_);
  or g_133710_(_043643_, _043650_, _043802_);
  and g_133711_(_043639_, _043799_, _043803_);
  or g_133712_(_043638_, _043798_, _043804_);
  and g_133713_(_043635_, _043803_, _043805_);
  or g_133714_(_043637_, _043804_, _043806_);
  and g_133715_(_043662_, _043802_, _043807_);
  or g_133716_(_043663_, _043800_, _043808_);
  and g_133717_(_043652_, _043808_, _043809_);
  or g_133718_(_043651_, _043807_, _043810_);
  and g_133719_(_043805_, _043810_, _043811_);
  or g_133720_(_043806_, _043809_, _043813_);
  xor g_133721_(_043654_, _043660_, _043814_);
  xor g_133722_(_043653_, _043660_, _043815_);
  and g_133723_(_043652_, _043797_, _043816_);
  or g_133724_(_043651_, _043796_, _043817_);
  and g_133725_(_043802_, _043816_, _043818_);
  or g_133726_(_043800_, _043817_, _043819_);
  and g_133727_(_043805_, _043818_, _043820_);
  or g_133728_(_043806_, _043819_, _043821_);
  and g_133729_(_043814_, _043820_, _043822_);
  or g_133730_(_043815_, _043821_, _043824_);
  and g_133731_(_043795_, _043822_, _043825_);
  or g_133732_(_043794_, _043824_, _043826_);
  or g_133733_(_043811_, _043825_, _043827_);
  and g_133734_(_043813_, _043826_, _043828_);
  and g_133735_(_043641_, _043828_, _043829_);
  or g_133736_(_043640_, _043827_, _043830_);
  and g_133737_(_043446_, _043829_, _043831_);
  or g_133738_(_043445_, _043830_, _043832_);
  and g_133739_(_043626_, _043830_, _043833_);
  or g_133740_(_043624_, _043829_, _043835_);
  and g_133741_(_043832_, _043835_, _043836_);
  or g_133742_(_043831_, _043833_, _043837_);
  and g_133743_(_043629_, _043631_, _043838_);
  or g_133744_(_043630_, _043632_, _043839_);
  or g_133745_(out[529], out[528], _043840_);
  or g_133746_(out[528], _020976_, _043841_);
  and g_133747_(out[531], _043841_, _043842_);
  and g_133748_(_021888_, _043841_, _043843_);
  and g_133749_(out[533], _043843_, _043844_);
  or g_133750_(out[534], _043844_, _043846_);
  and g_133751_(out[535], _043846_, _043847_);
  and g_133752_(out[536], _043847_, _043848_);
  or g_133753_(out[537], _043848_, _043849_);
  and g_133754_(out[538], _043849_, _043850_);
  xor g_133755_(out[539], _043850_, _043851_);
  xor g_133756_(_054743_, _043850_, _043852_);
  and g_133757_(_043838_, _043852_, _043853_);
  or g_133758_(_043839_, _043851_, _043854_);
  xor g_133759_(out[538], _043849_, _043855_);
  xor g_133760_(_054864_, _043849_, _043857_);
  and g_133761_(_043837_, _043855_, _043858_);
  or g_133762_(_043836_, _043857_, _043859_);
  and g_133763_(_043839_, _043851_, _043860_);
  or g_133764_(_043838_, _043852_, _043861_);
  and g_133765_(_043859_, _043861_, _043862_);
  or g_133766_(_043858_, _043860_, _043863_);
  and g_133767_(_043854_, _043863_, _043864_);
  or g_133768_(_043853_, _043862_, _043865_);
  and g_133769_(_043836_, _043857_, _043866_);
  or g_133770_(_043837_, _043855_, _043868_);
  and g_133771_(_043854_, _043868_, _043869_);
  or g_133772_(_043853_, _043866_, _043870_);
  and g_133773_(_043862_, _043869_, _043871_);
  or g_133774_(_043863_, _043870_, _043872_);
  and g_133775_(_043642_, _043829_, _043873_);
  or g_133776_(_043643_, _043830_, _043874_);
  and g_133777_(_043650_, _043830_, _043875_);
  or g_133778_(_043649_, _043829_, _043876_);
  and g_133779_(_043874_, _043876_, _043877_);
  or g_133780_(_043873_, _043875_, _043879_);
  xor g_133781_(out[537], _043848_, _043880_);
  xor g_133782_(_054853_, _043848_, _043881_);
  and g_133783_(_043877_, _043880_, _043882_);
  or g_133784_(_043879_, _043881_, _043883_);
  xor g_133785_(out[536], _043847_, _043884_);
  xor g_133786_(_054842_, _043847_, _043885_);
  or g_133787_(_043653_, _043830_, _043886_);
  not g_133788_(_043886_, _043887_);
  and g_133789_(_043661_, _043830_, _043888_);
  or g_133790_(_043660_, _043829_, _043890_);
  and g_133791_(_043886_, _043890_, _043891_);
  or g_133792_(_043887_, _043888_, _043892_);
  and g_133793_(_043884_, _043892_, _043893_);
  or g_133794_(_043885_, _043891_, _043894_);
  and g_133795_(_043879_, _043881_, _043895_);
  or g_133796_(_043877_, _043880_, _043896_);
  and g_133797_(_043894_, _043896_, _043897_);
  or g_133798_(_043893_, _043895_, _043898_);
  and g_133799_(_043883_, _043898_, _043899_);
  or g_133800_(_043882_, _043897_, _043901_);
  xor g_133801_(out[535], _043846_, _043902_);
  xor g_133802_(_054754_, _043846_, _043903_);
  and g_133803_(_043780_, _043829_, _043904_);
  or g_133804_(_043778_, _043830_, _043905_);
  and g_133805_(_043786_, _043830_, _043906_);
  or g_133806_(_043785_, _043829_, _043907_);
  and g_133807_(_043905_, _043907_, _043908_);
  or g_133808_(_043904_, _043906_, _043909_);
  and g_133809_(_043902_, _043909_, _043910_);
  or g_133810_(_043903_, _043908_, _043912_);
  xor g_133811_(out[534], _043844_, _043913_);
  xor g_133812_(_054765_, _043844_, _043914_);
  and g_133813_(_043761_, _043829_, _043915_);
  or g_133814_(_043762_, _043830_, _043916_);
  and g_133815_(_043769_, _043830_, _043917_);
  or g_133816_(_043767_, _043829_, _043918_);
  and g_133817_(_043916_, _043918_, _043919_);
  or g_133818_(_043915_, _043917_, _043920_);
  and g_133819_(_043913_, _043919_, _043921_);
  or g_133820_(_043914_, _043920_, _043923_);
  xor g_133821_(out[531], _043841_, _043924_);
  xor g_133822_(_054831_, _043841_, _043925_);
  and g_133823_(_043711_, _043829_, _043926_);
  or g_133824_(_043710_, _043830_, _043927_);
  and g_133825_(_043718_, _043830_, _043928_);
  or g_133826_(_043717_, _043829_, _043929_);
  and g_133827_(_043927_, _043929_, _043930_);
  or g_133828_(_043926_, _043928_, _043931_);
  and g_133829_(_043925_, _043930_, _043932_);
  or g_133830_(_043924_, _043931_, _043934_);
  xor g_133831_(out[530], _043840_, _043935_);
  xor g_133832_(_054820_, _043840_, _043936_);
  and g_133833_(_043664_, _043829_, _043937_);
  or g_133834_(_043665_, _043830_, _043938_);
  and g_133835_(_043672_, _043830_, _043939_);
  or g_133836_(_043671_, _043829_, _043940_);
  and g_133837_(_043938_, _043940_, _043941_);
  or g_133838_(_043937_, _043939_, _043942_);
  and g_133839_(_043936_, _043942_, _043943_);
  or g_133840_(_043935_, _043941_, _043945_);
  xor g_133841_(out[529], out[528], _043946_);
  xor g_133842_(_054798_, out[528], _043947_);
  and g_133843_(_043688_, _043829_, _043948_);
  or g_133844_(_043689_, _043830_, _043949_);
  and g_133845_(_043685_, _043830_, _043950_);
  or g_133846_(_043684_, _043829_, _043951_);
  and g_133847_(_043949_, _043951_, _043952_);
  or g_133848_(_043948_, _043950_, _043953_);
  and g_133849_(_043946_, _043952_, _043954_);
  or g_133850_(_043947_, _043953_, _043956_);
  and g_133851_(out[512], _043829_, _043957_);
  or g_133852_(_054677_, _043830_, _043958_);
  and g_133853_(_043698_, _043830_, _043959_);
  or g_133854_(_043697_, _043829_, _043960_);
  and g_133855_(_043958_, _043960_, _043961_);
  or g_133856_(_043957_, _043959_, _043962_);
  and g_133857_(out[528], _043961_, _043963_);
  or g_133858_(_054809_, _043962_, _043964_);
  and g_133859_(_043956_, _043964_, _043965_);
  or g_133860_(_043954_, _043963_, _043967_);
  and g_133861_(out[529], _043953_, _043968_);
  or g_133862_(_054798_, _043952_, _043969_);
  and g_133863_(_043935_, _043941_, _043970_);
  or g_133864_(_043936_, _043942_, _043971_);
  and g_133865_(_043945_, _043969_, _043972_);
  or g_133866_(_043943_, _043968_, _043973_);
  and g_133867_(_043967_, _043972_, _043974_);
  or g_133868_(_043965_, _043973_, _043975_);
  and g_133869_(_043934_, _043971_, _043976_);
  or g_133870_(_043932_, _043970_, _043978_);
  and g_133871_(_043975_, _043976_, _043979_);
  or g_133872_(_043974_, _043978_, _043980_);
  and g_133873_(_043924_, _043931_, _043981_);
  or g_133874_(_043925_, _043930_, _043982_);
  xor g_133875_(out[532], _043842_, _043983_);
  xor g_133876_(_054787_, _043842_, _043984_);
  and g_133877_(_043727_, _043829_, _043985_);
  or g_133878_(_043726_, _043830_, _043986_);
  and g_133879_(_043733_, _043830_, _043987_);
  or g_133880_(_043732_, _043829_, _043989_);
  and g_133881_(_043986_, _043989_, _043990_);
  or g_133882_(_043985_, _043987_, _043991_);
  and g_133883_(_043983_, _043991_, _043992_);
  or g_133884_(_043984_, _043990_, _043993_);
  and g_133885_(_043982_, _043993_, _043994_);
  or g_133886_(_043981_, _043992_, _043995_);
  and g_133887_(_043980_, _043994_, _043996_);
  or g_133888_(_043979_, _043995_, _043997_);
  xor g_133889_(out[533], _043843_, _043998_);
  xor g_133890_(_054776_, _043843_, _044000_);
  and g_133891_(_043747_, _043829_, _044001_);
  or g_133892_(_043745_, _043830_, _044002_);
  and g_133893_(_043753_, _043830_, _044003_);
  or g_133894_(_043752_, _043829_, _044004_);
  and g_133895_(_044002_, _044004_, _044005_);
  or g_133896_(_044001_, _044003_, _044006_);
  and g_133897_(_044000_, _044005_, _044007_);
  or g_133898_(_043998_, _044006_, _044008_);
  and g_133899_(_043984_, _043990_, _044009_);
  or g_133900_(_043983_, _043991_, _044011_);
  and g_133901_(_044008_, _044011_, _044012_);
  or g_133902_(_044007_, _044009_, _044013_);
  and g_133903_(_043997_, _044012_, _044014_);
  or g_133904_(_043996_, _044013_, _044015_);
  and g_133905_(_043914_, _043920_, _044016_);
  or g_133906_(_043913_, _043919_, _044017_);
  and g_133907_(_043998_, _044006_, _044018_);
  or g_133908_(_044000_, _044005_, _044019_);
  and g_133909_(_044017_, _044019_, _044020_);
  or g_133910_(_044016_, _044018_, _044022_);
  and g_133911_(_044015_, _044020_, _044023_);
  or g_133912_(_044014_, _044022_, _044024_);
  and g_133913_(_043923_, _044024_, _044025_);
  or g_133914_(_043921_, _044023_, _044026_);
  and g_133915_(_043912_, _044026_, _044027_);
  or g_133916_(_043910_, _044025_, _044028_);
  and g_133917_(_043885_, _043891_, _044029_);
  or g_133918_(_043884_, _043892_, _044030_);
  and g_133919_(_043903_, _043908_, _044031_);
  or g_133920_(_043902_, _043909_, _044033_);
  and g_133921_(_043883_, _043897_, _044034_);
  or g_133922_(_043882_, _043898_, _044035_);
  and g_133923_(_044030_, _044033_, _044036_);
  or g_133924_(_044029_, _044031_, _044037_);
  and g_133925_(_043871_, _044036_, _044038_);
  or g_133926_(_043872_, _044037_, _044039_);
  and g_133927_(_044034_, _044038_, _044040_);
  or g_133928_(_044035_, _044039_, _044041_);
  and g_133929_(_044028_, _044040_, _044042_);
  or g_133930_(_044027_, _044041_, _044044_);
  and g_133931_(_043871_, _043899_, _044045_);
  or g_133932_(_043872_, _043901_, _044046_);
  and g_133933_(_043865_, _044046_, _044047_);
  or g_133934_(_043864_, _044045_, _044048_);
  and g_133935_(_044044_, _044047_, _044049_);
  or g_133936_(_044042_, _044048_, _044050_);
  and g_133937_(_043837_, _044050_, _044051_);
  or g_133938_(_043836_, _044049_, _044052_);
  and g_133939_(_043857_, _044049_, _044053_);
  or g_133940_(_043855_, _044050_, _044055_);
  and g_133941_(_044052_, _044055_, _044056_);
  or g_133942_(_044051_, _044053_, _044057_);
  or g_133943_(out[545], out[544], _044058_);
  or g_133944_(out[544], _054003_, _044059_);
  and g_133945_(out[547], _044059_, _044060_);
  and g_133946_(_022114_, _044059_, _044061_);
  and g_133947_(out[549], _044061_, _044062_);
  or g_133948_(out[550], _044062_, _044063_);
  and g_133949_(out[551], _044063_, _044064_);
  xor g_133950_(out[551], _044063_, _044066_);
  xor g_133951_(_054886_, _044063_, _044067_);
  and g_133952_(_043909_, _044050_, _044068_);
  or g_133953_(_043908_, _044049_, _044069_);
  and g_133954_(_043903_, _044049_, _044070_);
  or g_133955_(_043902_, _044050_, _044071_);
  and g_133956_(_044069_, _044071_, _044072_);
  or g_133957_(_044068_, _044070_, _044073_);
  and g_133958_(_044066_, _044073_, _044074_);
  or g_133959_(_044067_, _044072_, _044075_);
  xor g_133960_(out[547], _044059_, _044077_);
  xor g_133961_(_054963_, _044059_, _044078_);
  and g_133962_(_043925_, _044049_, _044079_);
  or g_133963_(_043924_, _044050_, _044080_);
  and g_133964_(_043931_, _044050_, _044081_);
  or g_133965_(_043930_, _044049_, _044082_);
  and g_133966_(_044080_, _044082_, _044083_);
  or g_133967_(_044079_, _044081_, _044084_);
  and g_133968_(_044078_, _044083_, _044085_);
  or g_133969_(_044077_, _044084_, _044086_);
  xor g_133970_(out[546], _044058_, _044088_);
  xor g_133971_(_054952_, _044058_, _044089_);
  and g_133972_(_043942_, _044050_, _044090_);
  or g_133973_(_043941_, _044049_, _044091_);
  and g_133974_(_043935_, _044049_, _044092_);
  or g_133975_(_043936_, _044050_, _044093_);
  and g_133976_(_044091_, _044093_, _044094_);
  or g_133977_(_044090_, _044092_, _044095_);
  and g_133978_(_044089_, _044095_, _044096_);
  or g_133979_(_044088_, _044094_, _044097_);
  and g_133980_(_044088_, _044094_, _044099_);
  or g_133981_(_044089_, _044095_, _044100_);
  xor g_133982_(out[545], out[544], _044101_);
  xor g_133983_(_054930_, out[544], _044102_);
  and g_133984_(_043946_, _044049_, _044103_);
  or g_133985_(_043947_, _044050_, _044104_);
  and g_133986_(_043953_, _044050_, _044105_);
  or g_133987_(_043952_, _044049_, _044106_);
  and g_133988_(_044104_, _044106_, _044107_);
  or g_133989_(_044103_, _044105_, _044108_);
  and g_133990_(_044101_, _044107_, _044110_);
  or g_133991_(_044102_, _044108_, _044111_);
  and g_133992_(out[528], _044049_, _044112_);
  or g_133993_(_054809_, _044050_, _044113_);
  and g_133994_(_043962_, _044050_, _044114_);
  or g_133995_(_043961_, _044049_, _044115_);
  and g_133996_(_044113_, _044115_, _044116_);
  or g_133997_(_044112_, _044114_, _044117_);
  and g_133998_(out[544], _044116_, _044118_);
  or g_133999_(_054941_, _044117_, _044119_);
  and g_134000_(_044111_, _044119_, _044121_);
  or g_134001_(_044110_, _044118_, _044122_);
  and g_134002_(out[545], _044108_, _044123_);
  or g_134003_(_054930_, _044107_, _044124_);
  and g_134004_(_044097_, _044124_, _044125_);
  or g_134005_(_044096_, _044123_, _044126_);
  and g_134006_(_044122_, _044125_, _044127_);
  or g_134007_(_044121_, _044126_, _044128_);
  and g_134008_(_044086_, _044100_, _044129_);
  or g_134009_(_044085_, _044099_, _044130_);
  and g_134010_(_044128_, _044129_, _044132_);
  or g_134011_(_044127_, _044130_, _044133_);
  xor g_134012_(out[548], _044060_, _044134_);
  xor g_134013_(_054919_, _044060_, _044135_);
  and g_134014_(_043984_, _044049_, _044136_);
  or g_134015_(_043983_, _044050_, _044137_);
  and g_134016_(_043991_, _044050_, _044138_);
  or g_134017_(_043990_, _044049_, _044139_);
  and g_134018_(_044137_, _044139_, _044140_);
  or g_134019_(_044136_, _044138_, _044141_);
  and g_134020_(_044134_, _044141_, _044143_);
  or g_134021_(_044135_, _044140_, _044144_);
  and g_134022_(_044077_, _044084_, _044145_);
  or g_134023_(_044078_, _044083_, _044146_);
  and g_134024_(_044144_, _044146_, _044147_);
  or g_134025_(_044143_, _044145_, _044148_);
  and g_134026_(_044133_, _044147_, _044149_);
  or g_134027_(_044132_, _044148_, _044150_);
  xor g_134028_(out[549], _044061_, _044151_);
  xor g_134029_(_054908_, _044061_, _044152_);
  and g_134030_(_044000_, _044049_, _044154_);
  or g_134031_(_043998_, _044050_, _044155_);
  and g_134032_(_044006_, _044050_, _044156_);
  or g_134033_(_044005_, _044049_, _044157_);
  and g_134034_(_044155_, _044157_, _044158_);
  or g_134035_(_044154_, _044156_, _044159_);
  and g_134036_(_044152_, _044158_, _044160_);
  or g_134037_(_044151_, _044159_, _044161_);
  and g_134038_(_044135_, _044140_, _044162_);
  or g_134039_(_044134_, _044141_, _044163_);
  and g_134040_(_044161_, _044163_, _044165_);
  or g_134041_(_044160_, _044162_, _044166_);
  and g_134042_(_044150_, _044165_, _044167_);
  or g_134043_(_044149_, _044166_, _044168_);
  xor g_134044_(out[550], _044062_, _044169_);
  xor g_134045_(_054897_, _044062_, _044170_);
  and g_134046_(_043920_, _044050_, _044171_);
  or g_134047_(_043919_, _044049_, _044172_);
  and g_134048_(_043913_, _044049_, _044173_);
  or g_134049_(_043914_, _044050_, _044174_);
  and g_134050_(_044172_, _044174_, _044176_);
  or g_134051_(_044171_, _044173_, _044177_);
  and g_134052_(_044170_, _044177_, _044178_);
  or g_134053_(_044169_, _044176_, _044179_);
  and g_134054_(_044151_, _044159_, _044180_);
  or g_134055_(_044152_, _044158_, _044181_);
  and g_134056_(_044179_, _044181_, _044182_);
  or g_134057_(_044178_, _044180_, _044183_);
  and g_134058_(_044168_, _044182_, _044184_);
  or g_134059_(_044167_, _044183_, _044185_);
  and g_134060_(_044067_, _044072_, _044187_);
  or g_134061_(_044066_, _044073_, _044188_);
  and g_134062_(_044169_, _044176_, _044189_);
  or g_134063_(_044170_, _044177_, _044190_);
  and g_134064_(_044188_, _044190_, _044191_);
  or g_134065_(_044187_, _044189_, _044192_);
  and g_134066_(_044185_, _044191_, _044193_);
  or g_134067_(_044184_, _044192_, _044194_);
  and g_134068_(_044075_, _044194_, _044195_);
  or g_134069_(_044074_, _044193_, _044196_);
  and g_134070_(out[552], _044064_, _044198_);
  or g_134071_(out[553], _044198_, _044199_);
  and g_134072_(out[554], _044199_, _044200_);
  xor g_134073_(out[554], _044199_, _044201_);
  xor g_134074_(_054996_, _044199_, _044202_);
  and g_134075_(_044057_, _044201_, _044203_);
  or g_134076_(_044056_, _044202_, _044204_);
  and g_134077_(_043838_, _043851_, _044205_);
  or g_134078_(_043839_, _043852_, _044206_);
  xor g_134079_(out[555], _044200_, _044207_);
  xor g_134080_(_054875_, _044200_, _044209_);
  and g_134081_(_044206_, _044207_, _044210_);
  or g_134082_(_044205_, _044209_, _044211_);
  and g_134083_(_044204_, _044211_, _044212_);
  or g_134084_(_044203_, _044210_, _044213_);
  and g_134085_(_044205_, _044209_, _044214_);
  or g_134086_(_044206_, _044207_, _044215_);
  and g_134087_(_044056_, _044202_, _044216_);
  or g_134088_(_044057_, _044201_, _044217_);
  and g_134089_(_044215_, _044217_, _044218_);
  or g_134090_(_044214_, _044216_, _044220_);
  and g_134091_(_044212_, _044218_, _044221_);
  or g_134092_(_044213_, _044220_, _044222_);
  and g_134093_(_043879_, _044050_, _044223_);
  or g_134094_(_043877_, _044049_, _044224_);
  and g_134095_(_043880_, _044049_, _044225_);
  or g_134096_(_043881_, _044050_, _044226_);
  and g_134097_(_044224_, _044226_, _044227_);
  or g_134098_(_044223_, _044225_, _044228_);
  xor g_134099_(out[553], _044198_, _044229_);
  xor g_134100_(_054985_, _044198_, _044231_);
  and g_134101_(_044228_, _044231_, _044232_);
  or g_134102_(_044227_, _044229_, _044233_);
  xor g_134103_(out[552], _044064_, _044234_);
  xor g_134104_(_054974_, _044064_, _044235_);
  and g_134105_(_043892_, _044050_, _044236_);
  or g_134106_(_043891_, _044049_, _044237_);
  and g_134107_(_043885_, _044049_, _044238_);
  or g_134108_(_043884_, _044050_, _044239_);
  and g_134109_(_044237_, _044239_, _044240_);
  or g_134110_(_044236_, _044238_, _044242_);
  and g_134111_(_044234_, _044242_, _044243_);
  or g_134112_(_044235_, _044240_, _044244_);
  and g_134113_(_044233_, _044244_, _044245_);
  or g_134114_(_044232_, _044243_, _044246_);
  and g_134115_(_044227_, _044229_, _044247_);
  or g_134116_(_044228_, _044231_, _044248_);
  and g_134117_(_044235_, _044240_, _044249_);
  or g_134118_(_044234_, _044242_, _044250_);
  and g_134119_(_044248_, _044250_, _044251_);
  or g_134120_(_044247_, _044249_, _044253_);
  and g_134121_(_044245_, _044251_, _044254_);
  or g_134122_(_044246_, _044253_, _044255_);
  and g_134123_(_044221_, _044254_, _044256_);
  or g_134124_(_044222_, _044255_, _044257_);
  and g_134125_(_044196_, _044256_, _044258_);
  or g_134126_(_044195_, _044257_, _044259_);
  and g_134127_(_044213_, _044215_, _044260_);
  or g_134128_(_044212_, _044214_, _044261_);
  and g_134129_(_044246_, _044248_, _044262_);
  or g_134130_(_044245_, _044247_, _044264_);
  and g_134131_(_044221_, _044262_, _044265_);
  or g_134132_(_044222_, _044264_, _044266_);
  and g_134133_(_044261_, _044266_, _044267_);
  or g_134134_(_044260_, _044265_, _044268_);
  and g_134135_(_044259_, _044267_, _044269_);
  or g_134136_(_044258_, _044268_, _044270_);
  and g_134137_(_044057_, _044270_, _044271_);
  or g_134138_(_044056_, _044269_, _044272_);
  and g_134139_(_044202_, _044269_, _044273_);
  or g_134140_(_044201_, _044270_, _044275_);
  and g_134141_(_044272_, _044275_, _044276_);
  or g_134142_(_044271_, _044273_, _044277_);
  or g_134143_(out[561], out[560], _044278_);
  or g_134144_(out[560], _054260_, _044279_);
  and g_134145_(out[563], _044279_, _044280_);
  and g_134146_(_022344_, _044279_, _044281_);
  and g_134147_(out[565], _044281_, _044282_);
  or g_134148_(out[566], _044282_, _044283_);
  and g_134149_(out[567], _044283_, _044284_);
  xor g_134150_(out[567], _044283_, _044286_);
  xor g_134151_(_055018_, _044283_, _044287_);
  and g_134152_(_044073_, _044270_, _044288_);
  or g_134153_(_044072_, _044269_, _044289_);
  and g_134154_(_044067_, _044269_, _044290_);
  or g_134155_(_044066_, _044270_, _044291_);
  and g_134156_(_044289_, _044291_, _044292_);
  or g_134157_(_044288_, _044290_, _044293_);
  and g_134158_(_044286_, _044293_, _044294_);
  or g_134159_(_044287_, _044292_, _044295_);
  xor g_134160_(out[566], _044282_, _044297_);
  xor g_134161_(_055029_, _044282_, _044298_);
  and g_134162_(_044177_, _044270_, _044299_);
  or g_134163_(_044176_, _044269_, _044300_);
  and g_134164_(_044169_, _044269_, _044301_);
  or g_134165_(_044170_, _044270_, _044302_);
  and g_134166_(_044300_, _044302_, _044303_);
  or g_134167_(_044299_, _044301_, _044304_);
  and g_134168_(_044297_, _044303_, _044305_);
  or g_134169_(_044298_, _044304_, _044306_);
  xor g_134170_(out[561], out[560], _044308_);
  xor g_134171_(_055062_, out[560], _044309_);
  and g_134172_(_044101_, _044269_, _044310_);
  or g_134173_(_044102_, _044270_, _044311_);
  and g_134174_(_044108_, _044270_, _044312_);
  or g_134175_(_044107_, _044269_, _044313_);
  and g_134176_(_044311_, _044313_, _044314_);
  or g_134177_(_044310_, _044312_, _044315_);
  and g_134178_(_044308_, _044314_, _044316_);
  or g_134179_(_044309_, _044315_, _044317_);
  and g_134180_(out[544], _044269_, _044319_);
  or g_134181_(_054941_, _044270_, _044320_);
  and g_134182_(_044117_, _044270_, _044321_);
  or g_134183_(_044116_, _044269_, _044322_);
  and g_134184_(_044320_, _044322_, _044323_);
  or g_134185_(_044319_, _044321_, _044324_);
  and g_134186_(out[560], _044323_, _044325_);
  or g_134187_(_055073_, _044324_, _044326_);
  and g_134188_(_044317_, _044326_, _044327_);
  or g_134189_(_044316_, _044325_, _044328_);
  xor g_134190_(out[562], _044278_, _044330_);
  xor g_134191_(_055084_, _044278_, _044331_);
  and g_134192_(_044095_, _044270_, _044332_);
  or g_134193_(_044094_, _044269_, _044333_);
  and g_134194_(_044088_, _044269_, _044334_);
  or g_134195_(_044089_, _044270_, _044335_);
  and g_134196_(_044333_, _044335_, _044336_);
  or g_134197_(_044332_, _044334_, _044337_);
  and g_134198_(_044331_, _044337_, _044338_);
  or g_134199_(_044330_, _044336_, _044339_);
  and g_134200_(out[561], _044315_, _044341_);
  or g_134201_(_055062_, _044314_, _044342_);
  and g_134202_(_044339_, _044342_, _044343_);
  or g_134203_(_044338_, _044341_, _044344_);
  and g_134204_(_044328_, _044343_, _044345_);
  or g_134205_(_044327_, _044344_, _044346_);
  xor g_134206_(out[563], _044279_, _044347_);
  xor g_134207_(_055095_, _044279_, _044348_);
  and g_134208_(_044078_, _044269_, _044349_);
  or g_134209_(_044077_, _044270_, _044350_);
  and g_134210_(_044084_, _044270_, _044352_);
  or g_134211_(_044083_, _044269_, _044353_);
  and g_134212_(_044350_, _044353_, _044354_);
  or g_134213_(_044349_, _044352_, _044355_);
  and g_134214_(_044348_, _044354_, _044356_);
  or g_134215_(_044347_, _044355_, _044357_);
  and g_134216_(_044330_, _044336_, _044358_);
  or g_134217_(_044331_, _044337_, _044359_);
  and g_134218_(_044357_, _044359_, _044360_);
  or g_134219_(_044356_, _044358_, _044361_);
  and g_134220_(_044346_, _044360_, _044363_);
  or g_134221_(_044345_, _044361_, _044364_);
  xor g_134222_(out[564], _044280_, _044365_);
  xor g_134223_(_055051_, _044280_, _044366_);
  and g_134224_(_044135_, _044269_, _044367_);
  or g_134225_(_044134_, _044270_, _044368_);
  and g_134226_(_044141_, _044270_, _044369_);
  or g_134227_(_044140_, _044269_, _044370_);
  and g_134228_(_044368_, _044370_, _044371_);
  or g_134229_(_044367_, _044369_, _044372_);
  and g_134230_(_044365_, _044372_, _044374_);
  or g_134231_(_044366_, _044371_, _044375_);
  and g_134232_(_044347_, _044355_, _044376_);
  or g_134233_(_044348_, _044354_, _044377_);
  and g_134234_(_044375_, _044377_, _044378_);
  or g_134235_(_044374_, _044376_, _044379_);
  and g_134236_(_044364_, _044378_, _044380_);
  or g_134237_(_044363_, _044379_, _044381_);
  xor g_134238_(out[565], _044281_, _044382_);
  xor g_134239_(_055040_, _044281_, _044383_);
  and g_134240_(_044159_, _044270_, _044385_);
  or g_134241_(_044158_, _044269_, _044386_);
  and g_134242_(_044152_, _044269_, _044387_);
  or g_134243_(_044151_, _044270_, _044388_);
  and g_134244_(_044386_, _044388_, _044389_);
  or g_134245_(_044385_, _044387_, _044390_);
  and g_134246_(_044383_, _044389_, _044391_);
  or g_134247_(_044382_, _044390_, _044392_);
  and g_134248_(_044366_, _044371_, _044393_);
  or g_134249_(_044365_, _044372_, _044394_);
  and g_134250_(_044392_, _044394_, _044396_);
  or g_134251_(_044391_, _044393_, _044397_);
  and g_134252_(_044381_, _044396_, _044398_);
  or g_134253_(_044380_, _044397_, _044399_);
  and g_134254_(_044298_, _044304_, _044400_);
  or g_134255_(_044297_, _044303_, _044401_);
  and g_134256_(_044382_, _044390_, _044402_);
  or g_134257_(_044383_, _044389_, _044403_);
  and g_134258_(_044401_, _044403_, _044404_);
  or g_134259_(_044400_, _044402_, _044405_);
  and g_134260_(_044399_, _044404_, _044407_);
  or g_134261_(_044398_, _044405_, _044408_);
  and g_134262_(_044306_, _044408_, _044409_);
  or g_134263_(_044305_, _044407_, _044410_);
  and g_134264_(_044295_, _044410_, _044411_);
  or g_134265_(_044294_, _044409_, _044412_);
  and g_134266_(_044205_, _044207_, _044413_);
  or g_134267_(_044206_, _044209_, _044414_);
  and g_134268_(out[568], _044284_, _044415_);
  or g_134269_(out[569], _044415_, _044416_);
  and g_134270_(out[570], _044416_, _044418_);
  xor g_134271_(out[571], _044418_, _044419_);
  xor g_134272_(_055007_, _044418_, _044420_);
  and g_134273_(_044414_, _044419_, _044421_);
  or g_134274_(_044413_, _044420_, _044422_);
  xor g_134275_(out[570], _044416_, _044423_);
  xor g_134276_(_055128_, _044416_, _044424_);
  and g_134277_(_044277_, _044423_, _044425_);
  or g_134278_(_044276_, _044424_, _044426_);
  and g_134279_(_044422_, _044426_, _044427_);
  or g_134280_(_044421_, _044425_, _044429_);
  and g_134281_(_044276_, _044424_, _044430_);
  or g_134282_(_044277_, _044423_, _044431_);
  and g_134283_(_044413_, _044420_, _044432_);
  or g_134284_(_044414_, _044419_, _044433_);
  and g_134285_(_044431_, _044433_, _044434_);
  or g_134286_(_044430_, _044432_, _044435_);
  and g_134287_(_044427_, _044434_, _044436_);
  or g_134288_(_044429_, _044435_, _044437_);
  xor g_134289_(out[568], _044284_, _044438_);
  xor g_134290_(_055106_, _044284_, _044440_);
  and g_134291_(_044242_, _044270_, _044441_);
  or g_134292_(_044240_, _044269_, _044442_);
  and g_134293_(_044235_, _044269_, _044443_);
  or g_134294_(_044234_, _044270_, _044444_);
  and g_134295_(_044442_, _044444_, _044445_);
  or g_134296_(_044441_, _044443_, _044446_);
  and g_134297_(_044438_, _044446_, _044447_);
  or g_134298_(_044440_, _044445_, _044448_);
  xor g_134299_(out[569], _044415_, _044449_);
  xor g_134300_(_055117_, _044415_, _044451_);
  and g_134301_(_044228_, _044270_, _044452_);
  or g_134302_(_044227_, _044269_, _044453_);
  and g_134303_(_044229_, _044269_, _044454_);
  or g_134304_(_044231_, _044270_, _044455_);
  and g_134305_(_044453_, _044455_, _044456_);
  or g_134306_(_044452_, _044454_, _044457_);
  and g_134307_(_044451_, _044457_, _044458_);
  or g_134308_(_044449_, _044456_, _044459_);
  and g_134309_(_044448_, _044459_, _044460_);
  or g_134310_(_044447_, _044458_, _044462_);
  and g_134311_(_044449_, _044456_, _044463_);
  or g_134312_(_044451_, _044457_, _044464_);
  and g_134313_(_044440_, _044445_, _044465_);
  or g_134314_(_044438_, _044446_, _044466_);
  and g_134315_(_044464_, _044466_, _044467_);
  or g_134316_(_044463_, _044465_, _044468_);
  and g_134317_(_044287_, _044292_, _044469_);
  or g_134318_(_044286_, _044293_, _044470_);
  and g_134319_(_044467_, _044470_, _044471_);
  or g_134320_(_044468_, _044469_, _044473_);
  and g_134321_(_044460_, _044471_, _044474_);
  or g_134322_(_044462_, _044473_, _044475_);
  and g_134323_(_044436_, _044474_, _044476_);
  or g_134324_(_044437_, _044475_, _044477_);
  and g_134325_(_044412_, _044476_, _044478_);
  or g_134326_(_044411_, _044477_, _044479_);
  and g_134327_(_044462_, _044464_, _044480_);
  or g_134328_(_044460_, _044463_, _044481_);
  and g_134329_(_044436_, _044480_, _044482_);
  or g_134330_(_044437_, _044481_, _044484_);
  and g_134331_(_044429_, _044433_, _044485_);
  or g_134332_(_044427_, _044432_, _044486_);
  and g_134333_(_044484_, _044486_, _044487_);
  or g_134334_(_044482_, _044485_, _044488_);
  and g_134335_(_044479_, _044487_, _044489_);
  or g_134336_(_044478_, _044488_, _044490_);
  and g_134337_(_044277_, _044490_, _044491_);
  or g_134338_(_044276_, _044489_, _044492_);
  and g_134339_(_044424_, _044489_, _044493_);
  or g_134340_(_044423_, _044490_, _044495_);
  and g_134341_(_044492_, _044495_, _044496_);
  or g_134342_(_044491_, _044493_, _044497_);
  or g_134343_(out[577], out[576], _044498_);
  or g_134344_(out[576], _054570_, _044499_);
  and g_134345_(out[579], _044499_, _044500_);
  and g_134346_(_022564_, _044499_, _044501_);
  and g_134347_(out[581], _044501_, _044502_);
  or g_134348_(out[582], _044502_, _044503_);
  and g_134349_(out[583], _044503_, _044504_);
  xor g_134350_(out[583], _044503_, _044506_);
  xor g_134351_(_055150_, _044503_, _044507_);
  and g_134352_(_044293_, _044490_, _044508_);
  or g_134353_(_044292_, _044489_, _044509_);
  and g_134354_(_044287_, _044489_, _044510_);
  or g_134355_(_044286_, _044490_, _044511_);
  and g_134356_(_044509_, _044511_, _044512_);
  or g_134357_(_044508_, _044510_, _044513_);
  and g_134358_(_044506_, _044513_, _044514_);
  or g_134359_(_044507_, _044512_, _044515_);
  xor g_134360_(out[582], _044502_, _044517_);
  xor g_134361_(_055161_, _044502_, _044518_);
  and g_134362_(_044304_, _044490_, _044519_);
  or g_134363_(_044303_, _044489_, _044520_);
  and g_134364_(_044297_, _044489_, _044521_);
  or g_134365_(_044298_, _044490_, _044522_);
  and g_134366_(_044520_, _044522_, _044523_);
  or g_134367_(_044519_, _044521_, _044524_);
  and g_134368_(_044517_, _044523_, _044525_);
  or g_134369_(_044518_, _044524_, _044526_);
  xor g_134370_(out[577], out[576], _044528_);
  xor g_134371_(_055194_, out[576], _044529_);
  and g_134372_(_044308_, _044489_, _044530_);
  or g_134373_(_044309_, _044490_, _044531_);
  and g_134374_(_044315_, _044490_, _044532_);
  or g_134375_(_044314_, _044489_, _044533_);
  and g_134376_(_044531_, _044533_, _044534_);
  or g_134377_(_044530_, _044532_, _044535_);
  and g_134378_(_044528_, _044534_, _044536_);
  or g_134379_(_044529_, _044535_, _044537_);
  and g_134380_(out[560], _044489_, _044539_);
  or g_134381_(_055073_, _044490_, _044540_);
  and g_134382_(_044324_, _044490_, _044541_);
  or g_134383_(_044323_, _044489_, _044542_);
  and g_134384_(_044540_, _044542_, _044543_);
  or g_134385_(_044539_, _044541_, _044544_);
  and g_134386_(out[576], _044543_, _044545_);
  or g_134387_(_055205_, _044544_, _044546_);
  and g_134388_(_044537_, _044546_, _044547_);
  or g_134389_(_044536_, _044545_, _044548_);
  xor g_134390_(out[578], _044498_, _044550_);
  xor g_134391_(_055216_, _044498_, _044551_);
  and g_134392_(_044330_, _044489_, _044552_);
  or g_134393_(_044331_, _044490_, _044553_);
  and g_134394_(_044337_, _044490_, _044554_);
  or g_134395_(_044336_, _044489_, _044555_);
  and g_134396_(_044553_, _044555_, _044556_);
  or g_134397_(_044552_, _044554_, _044557_);
  and g_134398_(_044551_, _044557_, _044558_);
  or g_134399_(_044550_, _044556_, _044559_);
  and g_134400_(out[577], _044535_, _044561_);
  or g_134401_(_055194_, _044534_, _044562_);
  and g_134402_(_044559_, _044562_, _044563_);
  or g_134403_(_044558_, _044561_, _044564_);
  and g_134404_(_044548_, _044563_, _044565_);
  or g_134405_(_044547_, _044564_, _044566_);
  and g_134406_(_044550_, _044556_, _044567_);
  or g_134407_(_044551_, _044557_, _044568_);
  xor g_134408_(out[579], _044499_, _044569_);
  xor g_134409_(_055227_, _044499_, _044570_);
  and g_134410_(_044348_, _044489_, _044572_);
  or g_134411_(_044347_, _044490_, _044573_);
  and g_134412_(_044355_, _044490_, _044574_);
  or g_134413_(_044354_, _044489_, _044575_);
  and g_134414_(_044573_, _044575_, _044576_);
  or g_134415_(_044572_, _044574_, _044577_);
  and g_134416_(_044570_, _044576_, _044578_);
  or g_134417_(_044569_, _044577_, _044579_);
  and g_134418_(_044568_, _044579_, _044580_);
  or g_134419_(_044567_, _044578_, _044581_);
  and g_134420_(_044566_, _044580_, _044583_);
  or g_134421_(_044565_, _044581_, _044584_);
  and g_134422_(_044569_, _044577_, _044585_);
  or g_134423_(_044570_, _044576_, _044586_);
  xor g_134424_(out[580], _044500_, _044587_);
  xor g_134425_(_055183_, _044500_, _044588_);
  and g_134426_(_044372_, _044490_, _044589_);
  or g_134427_(_044371_, _044489_, _044590_);
  and g_134428_(_044366_, _044489_, _044591_);
  or g_134429_(_044365_, _044490_, _044592_);
  and g_134430_(_044590_, _044592_, _044594_);
  or g_134431_(_044589_, _044591_, _044595_);
  and g_134432_(_044587_, _044595_, _044596_);
  or g_134433_(_044588_, _044594_, _044597_);
  and g_134434_(_044586_, _044597_, _044598_);
  or g_134435_(_044585_, _044596_, _044599_);
  and g_134436_(_044584_, _044598_, _044600_);
  or g_134437_(_044583_, _044599_, _044601_);
  xor g_134438_(out[581], _044501_, _044602_);
  xor g_134439_(_055172_, _044501_, _044603_);
  and g_134440_(_044390_, _044490_, _044605_);
  or g_134441_(_044389_, _044489_, _044606_);
  and g_134442_(_044383_, _044489_, _044607_);
  or g_134443_(_044382_, _044490_, _044608_);
  and g_134444_(_044606_, _044608_, _044609_);
  or g_134445_(_044605_, _044607_, _044610_);
  and g_134446_(_044603_, _044609_, _044611_);
  or g_134447_(_044602_, _044610_, _044612_);
  and g_134448_(_044588_, _044594_, _044613_);
  or g_134449_(_044587_, _044595_, _044614_);
  and g_134450_(_044612_, _044614_, _044616_);
  or g_134451_(_044611_, _044613_, _044617_);
  and g_134452_(_044601_, _044616_, _044618_);
  or g_134453_(_044600_, _044617_, _044619_);
  and g_134454_(_044518_, _044524_, _044620_);
  or g_134455_(_044517_, _044523_, _044621_);
  and g_134456_(_044602_, _044610_, _044622_);
  or g_134457_(_044603_, _044609_, _044623_);
  and g_134458_(_044621_, _044623_, _044624_);
  or g_134459_(_044620_, _044622_, _044625_);
  and g_134460_(_044619_, _044624_, _044627_);
  or g_134461_(_044618_, _044625_, _044628_);
  and g_134462_(_044526_, _044628_, _044629_);
  or g_134463_(_044525_, _044627_, _044630_);
  and g_134464_(_044515_, _044630_, _044631_);
  or g_134465_(_044514_, _044629_, _044632_);
  and g_134466_(out[584], _044504_, _044633_);
  or g_134467_(out[585], _044633_, _044634_);
  and g_134468_(out[586], _044634_, _044635_);
  xor g_134469_(out[586], _044634_, _044636_);
  xor g_134470_(_055260_, _044634_, _044638_);
  and g_134471_(_044497_, _044636_, _044639_);
  or g_134472_(_044496_, _044638_, _044640_);
  and g_134473_(_044413_, _044419_, _044641_);
  or g_134474_(_044414_, _044420_, _044642_);
  xor g_134475_(out[587], _044635_, _044643_);
  xor g_134476_(_055139_, _044635_, _044644_);
  and g_134477_(_044642_, _044643_, _044645_);
  or g_134478_(_044641_, _044644_, _044646_);
  and g_134479_(_044640_, _044646_, _044647_);
  or g_134480_(_044639_, _044645_, _044649_);
  and g_134481_(_044496_, _044638_, _044650_);
  or g_134482_(_044497_, _044636_, _044651_);
  and g_134483_(_044641_, _044644_, _044652_);
  or g_134484_(_044642_, _044643_, _044653_);
  and g_134485_(_044651_, _044653_, _044654_);
  or g_134486_(_044650_, _044652_, _044655_);
  and g_134487_(_044647_, _044654_, _044656_);
  or g_134488_(_044649_, _044655_, _044657_);
  and g_134489_(_044457_, _044490_, _044658_);
  or g_134490_(_044456_, _044489_, _044660_);
  and g_134491_(_044449_, _044489_, _044661_);
  or g_134492_(_044451_, _044490_, _044662_);
  and g_134493_(_044660_, _044662_, _044663_);
  or g_134494_(_044658_, _044661_, _044664_);
  xor g_134495_(out[585], _044633_, _044665_);
  xor g_134496_(_055249_, _044633_, _044666_);
  and g_134497_(_044664_, _044666_, _044667_);
  or g_134498_(_044663_, _044665_, _044668_);
  xor g_134499_(out[584], _044504_, _044669_);
  xor g_134500_(_055238_, _044504_, _044671_);
  and g_134501_(_044446_, _044490_, _044672_);
  or g_134502_(_044445_, _044489_, _044673_);
  and g_134503_(_044440_, _044489_, _044674_);
  or g_134504_(_044438_, _044490_, _044675_);
  and g_134505_(_044673_, _044675_, _044676_);
  or g_134506_(_044672_, _044674_, _044677_);
  and g_134507_(_044669_, _044677_, _044678_);
  or g_134508_(_044671_, _044676_, _044679_);
  and g_134509_(_044668_, _044679_, _044680_);
  or g_134510_(_044667_, _044678_, _044682_);
  and g_134511_(_044671_, _044676_, _044683_);
  or g_134512_(_044669_, _044677_, _044684_);
  and g_134513_(_044663_, _044665_, _044685_);
  or g_134514_(_044664_, _044666_, _044686_);
  and g_134515_(_044507_, _044512_, _044687_);
  or g_134516_(_044506_, _044513_, _044688_);
  and g_134517_(_044686_, _044688_, _044689_);
  or g_134518_(_044685_, _044687_, _044690_);
  and g_134519_(_044684_, _044689_, _044691_);
  or g_134520_(_044683_, _044690_, _044693_);
  and g_134521_(_044680_, _044691_, _044694_);
  or g_134522_(_044682_, _044693_, _044695_);
  and g_134523_(_044656_, _044694_, _044696_);
  or g_134524_(_044657_, _044695_, _044697_);
  and g_134525_(_044632_, _044696_, _044698_);
  or g_134526_(_044631_, _044697_, _044699_);
  and g_134527_(_044682_, _044686_, _044700_);
  or g_134528_(_044680_, _044685_, _044701_);
  and g_134529_(_044656_, _044700_, _044702_);
  or g_134530_(_044657_, _044701_, _044704_);
  and g_134531_(_044649_, _044653_, _044705_);
  or g_134532_(_044647_, _044652_, _044706_);
  and g_134533_(_044704_, _044706_, _044707_);
  or g_134534_(_044702_, _044705_, _044708_);
  and g_134535_(_044699_, _044707_, _044709_);
  or g_134536_(_044698_, _044708_, _044710_);
  and g_134537_(_044497_, _044710_, _044711_);
  or g_134538_(_044496_, _044709_, _044712_);
  and g_134539_(_044638_, _044709_, _044713_);
  or g_134540_(_044636_, _044710_, _044715_);
  and g_134541_(_044712_, _044715_, _044716_);
  or g_134542_(_044711_, _044713_, _044717_);
  or g_134543_(out[593], out[592], _044718_);
  or g_134544_(out[592], _054791_, _044719_);
  and g_134545_(out[595], _044719_, _044720_);
  xor g_134546_(out[595], _044719_, _044721_);
  xor g_134547_(_055359_, _044719_, _044722_);
  and g_134548_(_044570_, _044709_, _044723_);
  or g_134549_(_044569_, _044710_, _044724_);
  and g_134550_(_044577_, _044710_, _044726_);
  or g_134551_(_044576_, _044709_, _044727_);
  and g_134552_(_044724_, _044727_, _044728_);
  or g_134553_(_044723_, _044726_, _044729_);
  and g_134554_(_044721_, _044729_, _044730_);
  or g_134555_(_044722_, _044728_, _044731_);
  and g_134556_(_044722_, _044728_, _044732_);
  or g_134557_(_044721_, _044729_, _044733_);
  xor g_134558_(out[594], _044718_, _044734_);
  xor g_134559_(_055348_, _044718_, _044735_);
  and g_134560_(_044557_, _044710_, _044737_);
  or g_134561_(_044556_, _044709_, _044738_);
  and g_134562_(_044550_, _044709_, _044739_);
  or g_134563_(_044551_, _044710_, _044740_);
  and g_134564_(_044738_, _044740_, _044741_);
  or g_134565_(_044737_, _044739_, _044742_);
  and g_134566_(_044734_, _044741_, _044743_);
  or g_134567_(_044735_, _044742_, _044744_);
  and g_134568_(_044733_, _044744_, _044745_);
  or g_134569_(_044732_, _044743_, _044746_);
  and g_134570_(_044731_, _044746_, _044748_);
  or g_134571_(_044730_, _044745_, _044749_);
  xor g_134572_(out[593], out[592], _044750_);
  not g_134573_(_044750_, _044751_);
  and g_134574_(_044528_, _044709_, _044752_);
  or g_134575_(_044529_, _044710_, _044753_);
  and g_134576_(_044535_, _044710_, _044754_);
  or g_134577_(_044534_, _044709_, _044755_);
  and g_134578_(_044753_, _044755_, _044756_);
  or g_134579_(_044752_, _044754_, _044757_);
  and g_134580_(_044750_, _044756_, _044759_);
  or g_134581_(_044751_, _044757_, _044760_);
  and g_134582_(out[576], _044709_, _044761_);
  or g_134583_(_055205_, _044710_, _044762_);
  and g_134584_(_044544_, _044710_, _044763_);
  or g_134585_(_044543_, _044709_, _044764_);
  and g_134586_(_044762_, _044764_, _044765_);
  or g_134587_(_044761_, _044763_, _044766_);
  and g_134588_(_055337_, _044766_, _044767_);
  or g_134589_(out[592], _044765_, _044768_);
  xor g_134590_(_044750_, _044756_, _044770_);
  xor g_134591_(_044751_, _044756_, _044771_);
  and g_134592_(_044768_, _044770_, _044772_);
  or g_134593_(_044767_, _044771_, _044773_);
  and g_134594_(_044760_, _044773_, _044774_);
  or g_134595_(_044759_, _044772_, _044775_);
  and g_134596_(_044735_, _044742_, _044776_);
  or g_134597_(_044734_, _044741_, _044777_);
  and g_134598_(_044731_, _044777_, _044778_);
  or g_134599_(_044730_, _044776_, _044779_);
  and g_134600_(_044775_, _044778_, _044781_);
  or g_134601_(_044774_, _044779_, _044782_);
  and g_134602_(_044749_, _044782_, _044783_);
  or g_134603_(_044748_, _044781_, _044784_);
  and g_134604_(_022798_, _044719_, _044785_);
  and g_134605_(out[597], _044785_, _044786_);
  or g_134606_(out[598], _044786_, _044787_);
  and g_134607_(out[599], _044787_, _044788_);
  and g_134608_(out[600], _044788_, _044789_);
  or g_134609_(out[601], _044789_, _044790_);
  and g_134610_(out[602], _044790_, _044792_);
  xor g_134611_(out[603], _044792_, _044793_);
  xor g_134612_(_055271_, _044792_, _044794_);
  and g_134613_(_044641_, _044643_, _044795_);
  or g_134614_(_044642_, _044644_, _044796_);
  and g_134615_(_044794_, _044795_, _044797_);
  or g_134616_(_044793_, _044796_, _044798_);
  xor g_134617_(out[602], _044790_, _044799_);
  xor g_134618_(_055392_, _044790_, _044800_);
  and g_134619_(_044716_, _044800_, _044801_);
  or g_134620_(_044717_, _044799_, _044803_);
  and g_134621_(_044798_, _044803_, _044804_);
  or g_134622_(_044797_, _044801_, _044805_);
  and g_134623_(_044717_, _044799_, _044806_);
  or g_134624_(_044716_, _044800_, _044807_);
  and g_134625_(_044793_, _044796_, _044808_);
  or g_134626_(_044794_, _044795_, _044809_);
  and g_134627_(_044807_, _044809_, _044810_);
  or g_134628_(_044806_, _044808_, _044811_);
  and g_134629_(_044804_, _044810_, _044812_);
  or g_134630_(_044805_, _044811_, _044814_);
  xor g_134631_(out[601], _044789_, _044815_);
  xor g_134632_(_055381_, _044789_, _044816_);
  and g_134633_(_044664_, _044710_, _044817_);
  or g_134634_(_044663_, _044709_, _044818_);
  and g_134635_(_044665_, _044709_, _044819_);
  or g_134636_(_044666_, _044710_, _044820_);
  and g_134637_(_044818_, _044820_, _044821_);
  or g_134638_(_044817_, _044819_, _044822_);
  and g_134639_(_044815_, _044821_, _044823_);
  or g_134640_(_044816_, _044822_, _044825_);
  xor g_134641_(out[600], _044788_, _044826_);
  xor g_134642_(_055370_, _044788_, _044827_);
  and g_134643_(_044677_, _044710_, _044828_);
  or g_134644_(_044676_, _044709_, _044829_);
  and g_134645_(_044671_, _044709_, _044830_);
  or g_134646_(_044669_, _044710_, _044831_);
  and g_134647_(_044829_, _044831_, _044832_);
  or g_134648_(_044828_, _044830_, _044833_);
  and g_134649_(_044827_, _044832_, _044834_);
  or g_134650_(_044826_, _044833_, _044836_);
  and g_134651_(_044825_, _044836_, _044837_);
  or g_134652_(_044823_, _044834_, _044838_);
  and g_134653_(_044826_, _044833_, _044839_);
  or g_134654_(_044827_, _044832_, _044840_);
  and g_134655_(_044816_, _044822_, _044841_);
  or g_134656_(_044815_, _044821_, _044842_);
  and g_134657_(_044840_, _044842_, _044843_);
  or g_134658_(_044839_, _044841_, _044844_);
  and g_134659_(_044837_, _044843_, _044845_);
  or g_134660_(_044838_, _044844_, _044847_);
  and g_134661_(_044812_, _044845_, _044848_);
  or g_134662_(_044814_, _044847_, _044849_);
  xor g_134663_(out[599], _044787_, _044850_);
  xor g_134664_(_055282_, _044787_, _044851_);
  and g_134665_(_044513_, _044710_, _044852_);
  or g_134666_(_044512_, _044709_, _044853_);
  and g_134667_(_044507_, _044709_, _044854_);
  or g_134668_(_044506_, _044710_, _044855_);
  and g_134669_(_044853_, _044855_, _044856_);
  or g_134670_(_044852_, _044854_, _044858_);
  and g_134671_(_044851_, _044856_, _044859_);
  or g_134672_(_044850_, _044858_, _044860_);
  xor g_134673_(out[598], _044786_, _044861_);
  xor g_134674_(_055293_, _044786_, _044862_);
  and g_134675_(_044524_, _044710_, _044863_);
  or g_134676_(_044523_, _044709_, _044864_);
  and g_134677_(_044517_, _044709_, _044865_);
  or g_134678_(_044518_, _044710_, _044866_);
  and g_134679_(_044864_, _044866_, _044867_);
  or g_134680_(_044863_, _044865_, _044869_);
  and g_134681_(_044861_, _044867_, _044870_);
  or g_134682_(_044862_, _044869_, _044871_);
  and g_134683_(_044860_, _044871_, _044872_);
  or g_134684_(_044859_, _044870_, _044873_);
  and g_134685_(_044862_, _044869_, _044874_);
  or g_134686_(_044861_, _044867_, _044875_);
  and g_134687_(_044850_, _044858_, _044876_);
  or g_134688_(_044851_, _044856_, _044877_);
  and g_134689_(_044875_, _044877_, _044878_);
  or g_134690_(_044874_, _044876_, _044880_);
  and g_134691_(_044872_, _044878_, _044881_);
  or g_134692_(_044873_, _044880_, _044882_);
  xor g_134693_(out[597], _044785_, _044883_);
  xor g_134694_(_055304_, _044785_, _044884_);
  and g_134695_(_044603_, _044709_, _044885_);
  or g_134696_(_044602_, _044710_, _044886_);
  and g_134697_(_044610_, _044710_, _044887_);
  or g_134698_(_044609_, _044709_, _044888_);
  and g_134699_(_044886_, _044888_, _044889_);
  or g_134700_(_044885_, _044887_, _044891_);
  and g_134701_(_044884_, _044889_, _044892_);
  or g_134702_(_044883_, _044891_, _044893_);
  xor g_134703_(out[596], _044720_, _044894_);
  xor g_134704_(_055315_, _044720_, _044895_);
  and g_134705_(_044588_, _044709_, _044896_);
  or g_134706_(_044587_, _044710_, _044897_);
  and g_134707_(_044595_, _044710_, _044898_);
  or g_134708_(_044594_, _044709_, _044899_);
  and g_134709_(_044897_, _044899_, _044900_);
  or g_134710_(_044896_, _044898_, _044902_);
  and g_134711_(_044895_, _044900_, _044903_);
  or g_134712_(_044894_, _044902_, _044904_);
  and g_134713_(_044893_, _044904_, _044905_);
  or g_134714_(_044892_, _044903_, _044906_);
  and g_134715_(_044894_, _044902_, _044907_);
  or g_134716_(_044895_, _044900_, _044908_);
  and g_134717_(_044883_, _044891_, _044909_);
  or g_134718_(_044884_, _044889_, _044910_);
  and g_134719_(_044908_, _044910_, _044911_);
  or g_134720_(_044907_, _044909_, _044913_);
  and g_134721_(_044905_, _044911_, _044914_);
  or g_134722_(_044906_, _044913_, _044915_);
  and g_134723_(_044881_, _044914_, _044916_);
  or g_134724_(_044882_, _044915_, _044917_);
  and g_134725_(_044848_, _044916_, _044918_);
  or g_134726_(_044849_, _044917_, _044919_);
  and g_134727_(_044784_, _044918_, _044920_);
  or g_134728_(_044783_, _044919_, _044921_);
  and g_134729_(_044873_, _044877_, _044922_);
  or g_134730_(_044872_, _044876_, _044924_);
  and g_134731_(_044906_, _044910_, _044925_);
  or g_134732_(_044905_, _044909_, _044926_);
  and g_134733_(_044881_, _044925_, _044927_);
  or g_134734_(_044882_, _044926_, _044928_);
  and g_134735_(_044924_, _044928_, _044929_);
  or g_134736_(_044922_, _044927_, _044930_);
  and g_134737_(_044848_, _044930_, _044931_);
  or g_134738_(_044849_, _044929_, _044932_);
  and g_134739_(_044838_, _044842_, _044933_);
  or g_134740_(_044837_, _044841_, _044935_);
  and g_134741_(_044812_, _044933_, _044936_);
  or g_134742_(_044814_, _044935_, _044937_);
  and g_134743_(_044805_, _044809_, _044938_);
  or g_134744_(_044804_, _044808_, _044939_);
  and g_134745_(_044937_, _044939_, _044940_);
  or g_134746_(_044936_, _044938_, _044941_);
  and g_134747_(_044932_, _044940_, _044942_);
  or g_134748_(_044931_, _044941_, _044943_);
  and g_134749_(_044921_, _044942_, _044944_);
  or g_134750_(_044920_, _044943_, _044946_);
  and g_134751_(out[592], _044765_, _044947_);
  or g_134752_(_055337_, _044766_, _044948_);
  and g_134753_(_044745_, _044778_, _044949_);
  or g_134754_(_044746_, _044779_, _044950_);
  and g_134755_(_044948_, _044949_, _044951_);
  or g_134756_(_044947_, _044950_, _044952_);
  and g_134757_(_044772_, _044951_, _044953_);
  or g_134758_(_044773_, _044952_, _044954_);
  and g_134759_(_044918_, _044953_, _044955_);
  or g_134760_(_044919_, _044954_, _044957_);
  and g_134761_(_044946_, _044957_, _044958_);
  or g_134762_(_044944_, _044955_, _044959_);
  and g_134763_(_044717_, _044959_, _044960_);
  or g_134764_(_044716_, _044958_, _044961_);
  and g_134765_(_044800_, _044958_, _044962_);
  or g_134766_(_044799_, _044959_, _044963_);
  and g_134767_(_044961_, _044963_, _044964_);
  or g_134768_(_044960_, _044962_, _044965_);
  or g_134769_(out[609], out[608], _044966_);
  or g_134770_(out[608], _054977_, _044968_);
  and g_134771_(out[611], _044968_, _044969_);
  and g_134772_(_023032_, _044968_, _044970_);
  and g_134773_(out[613], _044970_, _044971_);
  or g_134774_(out[614], _044971_, _044972_);
  xor g_134775_(out[614], _044971_, _044973_);
  xor g_134776_(_055425_, _044971_, _044974_);
  and g_134777_(_044869_, _044959_, _044975_);
  or g_134778_(_044867_, _044958_, _044976_);
  and g_134779_(_044861_, _044958_, _044977_);
  or g_134780_(_044862_, _044959_, _044979_);
  and g_134781_(_044976_, _044979_, _044980_);
  or g_134782_(_044975_, _044977_, _044981_);
  and g_134783_(_044973_, _044980_, _044982_);
  or g_134784_(_044974_, _044981_, _044983_);
  xor g_134785_(out[613], _044970_, _044984_);
  xor g_134786_(_055436_, _044970_, _044985_);
  and g_134787_(_044891_, _044959_, _044986_);
  or g_134788_(_044889_, _044958_, _044987_);
  and g_134789_(_044884_, _044958_, _044988_);
  or g_134790_(_044883_, _044959_, _044990_);
  and g_134791_(_044987_, _044990_, _044991_);
  or g_134792_(_044986_, _044988_, _044992_);
  and g_134793_(_044984_, _044992_, _044993_);
  or g_134794_(_044985_, _044991_, _044994_);
  xor g_134795_(_055458_, out[608], _044995_);
  not g_134796_(_044995_, _044996_);
  and g_134797_(_044757_, _044959_, _044997_);
  or g_134798_(_044756_, _044958_, _044998_);
  and g_134799_(_044750_, _044958_, _044999_);
  or g_134800_(_044751_, _044959_, _045001_);
  and g_134801_(_044998_, _045001_, _045002_);
  or g_134802_(_044997_, _044999_, _045003_);
  and g_134803_(_044996_, _045002_, _045004_);
  or g_134804_(_044995_, _045003_, _045005_);
  and g_134805_(out[592], _044958_, _045006_);
  or g_134806_(_055337_, _044959_, _045007_);
  and g_134807_(_044766_, _044959_, _045008_);
  or g_134808_(_044765_, _044958_, _045009_);
  and g_134809_(_045007_, _045009_, _045010_);
  or g_134810_(_045006_, _045008_, _045012_);
  and g_134811_(out[608], _045010_, _045013_);
  or g_134812_(_055469_, _045012_, _045014_);
  and g_134813_(_045005_, _045014_, _045015_);
  or g_134814_(_045004_, _045013_, _045016_);
  xor g_134815_(out[610], _044966_, _045017_);
  xor g_134816_(_055480_, _044966_, _045018_);
  and g_134817_(_044742_, _044959_, _045019_);
  or g_134818_(_044741_, _044958_, _045020_);
  and g_134819_(_044734_, _044958_, _045021_);
  or g_134820_(_044735_, _044959_, _045023_);
  and g_134821_(_045020_, _045023_, _045024_);
  or g_134822_(_045019_, _045021_, _045025_);
  and g_134823_(_045018_, _045025_, _045026_);
  or g_134824_(_045017_, _045024_, _045027_);
  and g_134825_(out[609], _045003_, _045028_);
  or g_134826_(_055458_, _045002_, _045029_);
  and g_134827_(_045027_, _045029_, _045030_);
  or g_134828_(_045026_, _045028_, _045031_);
  and g_134829_(_045016_, _045030_, _045032_);
  or g_134830_(_045015_, _045031_, _045034_);
  xor g_134831_(out[611], _044968_, _045035_);
  xor g_134832_(_055491_, _044968_, _045036_);
  and g_134833_(_044722_, _044958_, _045037_);
  or g_134834_(_044721_, _044959_, _045038_);
  and g_134835_(_044729_, _044959_, _045039_);
  or g_134836_(_044728_, _044958_, _045040_);
  and g_134837_(_045038_, _045040_, _045041_);
  or g_134838_(_045037_, _045039_, _045042_);
  and g_134839_(_045036_, _045041_, _045043_);
  or g_134840_(_045035_, _045042_, _045045_);
  and g_134841_(_045017_, _045024_, _045046_);
  or g_134842_(_045018_, _045025_, _045047_);
  and g_134843_(_045045_, _045047_, _045048_);
  or g_134844_(_045043_, _045046_, _045049_);
  and g_134845_(_045034_, _045048_, _045050_);
  or g_134846_(_045032_, _045049_, _045051_);
  xor g_134847_(out[612], _044969_, _045052_);
  xor g_134848_(_055447_, _044969_, _045053_);
  and g_134849_(_044902_, _044959_, _045054_);
  or g_134850_(_044900_, _044958_, _045056_);
  and g_134851_(_044895_, _044958_, _045057_);
  or g_134852_(_044894_, _044959_, _045058_);
  and g_134853_(_045056_, _045058_, _045059_);
  or g_134854_(_045054_, _045057_, _045060_);
  and g_134855_(_045052_, _045060_, _045061_);
  or g_134856_(_045053_, _045059_, _045062_);
  and g_134857_(_045035_, _045042_, _045063_);
  or g_134858_(_045036_, _045041_, _045064_);
  and g_134859_(_045062_, _045064_, _045065_);
  or g_134860_(_045061_, _045063_, _045067_);
  and g_134861_(_045051_, _045065_, _045068_);
  or g_134862_(_045050_, _045067_, _045069_);
  and g_134863_(_044985_, _044991_, _045070_);
  or g_134864_(_044984_, _044992_, _045071_);
  and g_134865_(_045053_, _045059_, _045072_);
  or g_134866_(_045052_, _045060_, _045073_);
  and g_134867_(_045071_, _045073_, _045074_);
  or g_134868_(_045070_, _045072_, _045075_);
  and g_134869_(_045069_, _045074_, _045076_);
  or g_134870_(_045068_, _045075_, _045078_);
  and g_134871_(_044994_, _045078_, _045079_);
  or g_134872_(_044993_, _045076_, _045080_);
  and g_134873_(_044983_, _045080_, _045081_);
  or g_134874_(_044982_, _045079_, _045082_);
  and g_134875_(out[615], _044972_, _045083_);
  xor g_134876_(out[615], _044972_, _045084_);
  xor g_134877_(_055414_, _044972_, _045085_);
  and g_134878_(_044858_, _044959_, _045086_);
  or g_134879_(_044856_, _044958_, _045087_);
  and g_134880_(_044851_, _044958_, _045089_);
  or g_134881_(_044850_, _044959_, _045090_);
  and g_134882_(_045087_, _045090_, _045091_);
  or g_134883_(_045086_, _045089_, _045092_);
  and g_134884_(_045084_, _045092_, _045093_);
  or g_134885_(_045085_, _045091_, _045094_);
  and g_134886_(_044974_, _044981_, _045095_);
  or g_134887_(_044973_, _044980_, _045096_);
  and g_134888_(_045094_, _045096_, _045097_);
  or g_134889_(_045093_, _045095_, _045098_);
  and g_134890_(_045082_, _045097_, _045100_);
  or g_134891_(_045081_, _045098_, _045101_);
  and g_134892_(out[616], _045083_, _045102_);
  or g_134893_(out[617], _045102_, _045103_);
  and g_134894_(out[618], _045103_, _045104_);
  xor g_134895_(out[618], _045103_, _045105_);
  xor g_134896_(_055524_, _045103_, _045106_);
  and g_134897_(_044965_, _045105_, _045107_);
  or g_134898_(_044964_, _045106_, _045108_);
  and g_134899_(_044794_, _044958_, _045109_);
  or g_134900_(_044793_, _044959_, _045111_);
  and g_134901_(_044796_, _044959_, _045112_);
  or g_134902_(_044795_, _044958_, _045113_);
  and g_134903_(_045111_, _045113_, _045114_);
  or g_134904_(_045109_, _045112_, _045115_);
  xor g_134905_(out[619], _045104_, _045116_);
  xor g_134906_(_055403_, _045104_, _045117_);
  and g_134907_(_045115_, _045116_, _045118_);
  or g_134908_(_045114_, _045117_, _045119_);
  and g_134909_(_045108_, _045119_, _045120_);
  or g_134910_(_045107_, _045118_, _045122_);
  and g_134911_(_045114_, _045117_, _045123_);
  or g_134912_(_045115_, _045116_, _045124_);
  and g_134913_(_044964_, _045106_, _045125_);
  or g_134914_(_044965_, _045105_, _045126_);
  and g_134915_(_045124_, _045126_, _045127_);
  or g_134916_(_045123_, _045125_, _045128_);
  and g_134917_(_045120_, _045127_, _045129_);
  or g_134918_(_045122_, _045128_, _045130_);
  and g_134919_(_044822_, _044959_, _045131_);
  or g_134920_(_044821_, _044958_, _045133_);
  and g_134921_(_044815_, _044958_, _045134_);
  or g_134922_(_044816_, _044959_, _045135_);
  and g_134923_(_045133_, _045135_, _045136_);
  or g_134924_(_045131_, _045134_, _045137_);
  xor g_134925_(out[617], _045102_, _045138_);
  not g_134926_(_045138_, _045139_);
  and g_134927_(_045137_, _045139_, _045140_);
  or g_134928_(_045136_, _045138_, _045141_);
  xor g_134929_(out[616], _045083_, _045142_);
  not g_134930_(_045142_, _045144_);
  and g_134931_(_044833_, _044959_, _045145_);
  or g_134932_(_044832_, _044958_, _045146_);
  and g_134933_(_044827_, _044958_, _045147_);
  or g_134934_(_044826_, _044959_, _045148_);
  and g_134935_(_045146_, _045148_, _045149_);
  or g_134936_(_045145_, _045147_, _045150_);
  and g_134937_(_045142_, _045150_, _045151_);
  or g_134938_(_045144_, _045149_, _045152_);
  and g_134939_(_045141_, _045152_, _045153_);
  or g_134940_(_045140_, _045151_, _045155_);
  and g_134941_(_045085_, _045091_, _045156_);
  or g_134942_(_045084_, _045092_, _045157_);
  and g_134943_(_045136_, _045138_, _045158_);
  or g_134944_(_045137_, _045139_, _045159_);
  and g_134945_(_045144_, _045149_, _045160_);
  or g_134946_(_045142_, _045150_, _045161_);
  and g_134947_(_045159_, _045161_, _045162_);
  or g_134948_(_045158_, _045160_, _045163_);
  and g_134949_(_045157_, _045162_, _045164_);
  or g_134950_(_045156_, _045163_, _045166_);
  and g_134951_(_045153_, _045164_, _045167_);
  or g_134952_(_045155_, _045166_, _045168_);
  and g_134953_(_045129_, _045167_, _045169_);
  or g_134954_(_045130_, _045168_, _045170_);
  and g_134955_(_045101_, _045169_, _045171_);
  or g_134956_(_045100_, _045170_, _045172_);
  and g_134957_(_045155_, _045159_, _045173_);
  or g_134958_(_045153_, _045158_, _045174_);
  and g_134959_(_045129_, _045173_, _045175_);
  or g_134960_(_045130_, _045174_, _045177_);
  and g_134961_(_045122_, _045124_, _045178_);
  or g_134962_(_045120_, _045123_, _045179_);
  and g_134963_(_045177_, _045179_, _045180_);
  or g_134964_(_045175_, _045178_, _045181_);
  and g_134965_(_045172_, _045180_, _045182_);
  or g_134966_(_045171_, _045181_, _045183_);
  and g_134967_(_044965_, _045183_, _045184_);
  or g_134968_(_044964_, _045182_, _045185_);
  and g_134969_(_045106_, _045182_, _045186_);
  or g_134970_(_045105_, _045183_, _045188_);
  and g_134971_(_045185_, _045188_, _045189_);
  or g_134972_(_045184_, _045186_, _045190_);
  and g_134973_(_045114_, _045116_, _045191_);
  or g_134974_(_045115_, _045117_, _045192_);
  or g_134975_(out[625], out[624], _045193_);
  or g_134976_(out[624], _055090_, _045194_);
  and g_134977_(out[627], _045194_, _045195_);
  and g_134978_(_023247_, _045194_, _045196_);
  and g_134979_(out[629], _045196_, _045197_);
  or g_134980_(out[630], _045197_, _045199_);
  and g_134981_(out[631], _045199_, _045200_);
  and g_134982_(out[632], _045200_, _045201_);
  or g_134983_(out[633], _045201_, _045202_);
  and g_134984_(out[634], _045202_, _045203_);
  xor g_134985_(out[635], _045203_, _045204_);
  xor g_134986_(_055535_, _045203_, _045205_);
  and g_134987_(_045192_, _045204_, _045206_);
  or g_134988_(_045191_, _045205_, _045207_);
  xor g_134989_(out[633], _045201_, _045208_);
  xor g_134990_(_055645_, _045201_, _045210_);
  and g_134991_(_045137_, _045183_, _045211_);
  or g_134992_(_045136_, _045182_, _045212_);
  and g_134993_(_045138_, _045182_, _045213_);
  or g_134994_(_045139_, _045183_, _045214_);
  and g_134995_(_045212_, _045214_, _045215_);
  or g_134996_(_045211_, _045213_, _045216_);
  and g_134997_(_045210_, _045216_, _045217_);
  or g_134998_(_045208_, _045215_, _045218_);
  and g_134999_(_045207_, _045218_, _045219_);
  or g_135000_(_045206_, _045217_, _045221_);
  xor g_135001_(out[634], _045202_, _045222_);
  xor g_135002_(_055656_, _045202_, _045223_);
  and g_135003_(_045190_, _045222_, _045224_);
  or g_135004_(_045189_, _045223_, _045225_);
  xor g_135005_(out[632], _045200_, _045226_);
  xor g_135006_(_055634_, _045200_, _045227_);
  and g_135007_(_045150_, _045183_, _045228_);
  or g_135008_(_045149_, _045182_, _045229_);
  and g_135009_(_045144_, _045182_, _045230_);
  or g_135010_(_045142_, _045183_, _045232_);
  and g_135011_(_045229_, _045232_, _045233_);
  or g_135012_(_045228_, _045230_, _045234_);
  and g_135013_(_045226_, _045234_, _045235_);
  or g_135014_(_045227_, _045233_, _045236_);
  and g_135015_(_045225_, _045236_, _045237_);
  or g_135016_(_045224_, _045235_, _045238_);
  and g_135017_(_045219_, _045237_, _045239_);
  or g_135018_(_045221_, _045238_, _045240_);
  and g_135019_(_045189_, _045223_, _045241_);
  or g_135020_(_045190_, _045222_, _045243_);
  and g_135021_(_045191_, _045205_, _045244_);
  or g_135022_(_045192_, _045204_, _045245_);
  and g_135023_(_045243_, _045245_, _045246_);
  or g_135024_(_045241_, _045244_, _045247_);
  and g_135025_(_045208_, _045215_, _045248_);
  or g_135026_(_045210_, _045216_, _045249_);
  and g_135027_(_045227_, _045233_, _045250_);
  or g_135028_(_045226_, _045234_, _045251_);
  and g_135029_(_045249_, _045251_, _045252_);
  or g_135030_(_045248_, _045250_, _045254_);
  and g_135031_(_045246_, _045252_, _045255_);
  or g_135032_(_045247_, _045254_, _045256_);
  and g_135033_(_045239_, _045255_, _045257_);
  or g_135034_(_045240_, _045256_, _045258_);
  xor g_135035_(out[630], _045197_, _045259_);
  xor g_135036_(_055557_, _045197_, _045260_);
  and g_135037_(_044981_, _045183_, _045261_);
  or g_135038_(_044980_, _045182_, _045262_);
  and g_135039_(_044973_, _045182_, _045263_);
  or g_135040_(_044974_, _045183_, _045265_);
  and g_135041_(_045262_, _045265_, _045266_);
  or g_135042_(_045261_, _045263_, _045267_);
  and g_135043_(_045260_, _045267_, _045268_);
  or g_135044_(_045259_, _045266_, _045269_);
  xor g_135045_(out[631], _045199_, _045270_);
  xor g_135046_(_055546_, _045199_, _045271_);
  and g_135047_(_045092_, _045183_, _045272_);
  or g_135048_(_045091_, _045182_, _045273_);
  and g_135049_(_045085_, _045182_, _045274_);
  or g_135050_(_045084_, _045183_, _045276_);
  and g_135051_(_045273_, _045276_, _045277_);
  or g_135052_(_045272_, _045274_, _045278_);
  and g_135053_(_045270_, _045278_, _045279_);
  or g_135054_(_045271_, _045277_, _045280_);
  xor g_135055_(out[629], _045196_, _045281_);
  xor g_135056_(_055568_, _045196_, _045282_);
  and g_135057_(_044985_, _045182_, _045283_);
  or g_135058_(_044984_, _045183_, _045284_);
  and g_135059_(_044992_, _045183_, _045285_);
  or g_135060_(_044991_, _045182_, _045287_);
  and g_135061_(_045284_, _045287_, _045288_);
  or g_135062_(_045283_, _045285_, _045289_);
  and g_135063_(_045281_, _045289_, _045290_);
  or g_135064_(_045282_, _045288_, _045291_);
  and g_135065_(_045282_, _045288_, _045292_);
  or g_135066_(_045281_, _045289_, _045293_);
  xor g_135067_(out[628], _045195_, _045294_);
  xor g_135068_(_055579_, _045195_, _045295_);
  and g_135069_(_045060_, _045183_, _045296_);
  or g_135070_(_045059_, _045182_, _045298_);
  and g_135071_(_045053_, _045182_, _045299_);
  or g_135072_(_045052_, _045183_, _045300_);
  and g_135073_(_045298_, _045300_, _045301_);
  or g_135074_(_045296_, _045299_, _045302_);
  and g_135075_(_045295_, _045301_, _045303_);
  or g_135076_(_045294_, _045302_, _045304_);
  and g_135077_(_045293_, _045304_, _045305_);
  or g_135078_(_045292_, _045303_, _045306_);
  and g_135079_(_045259_, _045266_, _045307_);
  or g_135080_(_045260_, _045267_, _045309_);
  and g_135081_(_045271_, _045277_, _045310_);
  or g_135082_(_045270_, _045278_, _045311_);
  and g_135083_(_045309_, _045311_, _045312_);
  or g_135084_(_045307_, _045310_, _045313_);
  and g_135085_(_045294_, _045302_, _045314_);
  or g_135086_(_045295_, _045301_, _045315_);
  and g_135087_(_045269_, _045280_, _045316_);
  or g_135088_(_045268_, _045279_, _045317_);
  and g_135089_(_045312_, _045316_, _045318_);
  or g_135090_(_045313_, _045317_, _045320_);
  and g_135091_(_045291_, _045315_, _045321_);
  or g_135092_(_045290_, _045314_, _045322_);
  and g_135093_(_045305_, _045321_, _045323_);
  or g_135094_(_045306_, _045322_, _045324_);
  and g_135095_(_045257_, _045323_, _045325_);
  or g_135096_(_045258_, _045324_, _045326_);
  and g_135097_(_045318_, _045325_, _045327_);
  or g_135098_(_045320_, _045326_, _045328_);
  xor g_135099_(out[626], _045193_, _045329_);
  not g_135100_(_045329_, _045331_);
  and g_135101_(_045025_, _045183_, _045332_);
  or g_135102_(_045024_, _045182_, _045333_);
  and g_135103_(_045017_, _045182_, _045334_);
  or g_135104_(_045018_, _045183_, _045335_);
  and g_135105_(_045333_, _045335_, _045336_);
  or g_135106_(_045332_, _045334_, _045337_);
  and g_135107_(_045329_, _045336_, _045338_);
  or g_135108_(_045331_, _045337_, _045339_);
  xor g_135109_(out[627], _045194_, _045340_);
  xor g_135110_(_055623_, _045194_, _045342_);
  and g_135111_(_045036_, _045182_, _045343_);
  or g_135112_(_045035_, _045183_, _045344_);
  and g_135113_(_045042_, _045183_, _045345_);
  or g_135114_(_045041_, _045182_, _045346_);
  and g_135115_(_045344_, _045346_, _045347_);
  or g_135116_(_045343_, _045345_, _045348_);
  and g_135117_(_045342_, _045347_, _045349_);
  or g_135118_(_045340_, _045348_, _045350_);
  and g_135119_(_045339_, _045350_, _045351_);
  or g_135120_(_045338_, _045349_, _045353_);
  and g_135121_(_045340_, _045348_, _045354_);
  or g_135122_(_045342_, _045347_, _045355_);
  and g_135123_(_045331_, _045337_, _045356_);
  or g_135124_(_045329_, _045336_, _045357_);
  and g_135125_(_045355_, _045357_, _045358_);
  or g_135126_(_045354_, _045356_, _045359_);
  and g_135127_(_045351_, _045358_, _045360_);
  or g_135128_(_045353_, _045359_, _045361_);
  xor g_135129_(out[625], out[624], _045362_);
  not g_135130_(_045362_, _045364_);
  or g_135131_(_044995_, _045183_, _045365_);
  or g_135132_(_045002_, _045182_, _045366_);
  and g_135133_(_045365_, _045366_, _045367_);
  not g_135134_(_045367_, _045368_);
  and g_135135_(_045362_, _045367_, _045369_);
  not g_135136_(_045369_, _045370_);
  and g_135137_(out[608], _045182_, _045371_);
  or g_135138_(_055469_, _045183_, _045372_);
  and g_135139_(_045012_, _045183_, _045373_);
  or g_135140_(_045010_, _045182_, _045375_);
  and g_135141_(_045372_, _045375_, _045376_);
  or g_135142_(_045371_, _045373_, _045377_);
  and g_135143_(_055601_, _045377_, _045378_);
  or g_135144_(out[624], _045376_, _045379_);
  xor g_135145_(_045362_, _045367_, _045380_);
  xor g_135146_(_045364_, _045367_, _045381_);
  and g_135147_(_045379_, _045380_, _045382_);
  or g_135148_(_045378_, _045381_, _045383_);
  and g_135149_(_045370_, _045383_, _045384_);
  or g_135150_(_045369_, _045382_, _045386_);
  and g_135151_(_045360_, _045386_, _045387_);
  or g_135152_(_045361_, _045384_, _045388_);
  and g_135153_(_045353_, _045355_, _045389_);
  or g_135154_(_045351_, _045354_, _045390_);
  and g_135155_(_045388_, _045390_, _045391_);
  or g_135156_(_045387_, _045389_, _045392_);
  and g_135157_(_045327_, _045392_, _045393_);
  or g_135158_(_045328_, _045391_, _045394_);
  and g_135159_(_045280_, _045313_, _045395_);
  or g_135160_(_045279_, _045312_, _045397_);
  and g_135161_(_045291_, _045306_, _045398_);
  or g_135162_(_045290_, _045305_, _045399_);
  and g_135163_(_045316_, _045398_, _045400_);
  or g_135164_(_045317_, _045399_, _045401_);
  and g_135165_(_045397_, _045401_, _045402_);
  or g_135166_(_045395_, _045400_, _045403_);
  and g_135167_(_045257_, _045403_, _045404_);
  or g_135168_(_045258_, _045402_, _045405_);
  and g_135169_(_045218_, _045225_, _045406_);
  or g_135170_(_045217_, _045224_, _045408_);
  and g_135171_(_045254_, _045406_, _045409_);
  or g_135172_(_045252_, _045408_, _045410_);
  and g_135173_(_045246_, _045410_, _045411_);
  or g_135174_(_045247_, _045409_, _045412_);
  and g_135175_(_045207_, _045412_, _045413_);
  or g_135176_(_045206_, _045411_, _045414_);
  and g_135177_(_045405_, _045414_, _045415_);
  or g_135178_(_045404_, _045413_, _045416_);
  and g_135179_(_045394_, _045415_, _045417_);
  or g_135180_(_045393_, _045416_, _045419_);
  and g_135181_(out[624], _045376_, _045420_);
  or g_135182_(_055601_, _045377_, _045421_);
  and g_135183_(_045360_, _045421_, _045422_);
  or g_135184_(_045361_, _045420_, _045423_);
  and g_135185_(_045382_, _045422_, _045424_);
  or g_135186_(_045383_, _045423_, _045425_);
  and g_135187_(_045327_, _045424_, _045426_);
  or g_135188_(_045328_, _045425_, _045427_);
  and g_135189_(_045419_, _045427_, _045428_);
  or g_135190_(_045417_, _045426_, _045430_);
  and g_135191_(_045190_, _045430_, _045431_);
  or g_135192_(_045189_, _045428_, _045432_);
  and g_135193_(_045223_, _045428_, _045433_);
  or g_135194_(_045222_, _045430_, _045434_);
  and g_135195_(_045432_, _045434_, _045435_);
  or g_135196_(_045431_, _045433_, _045436_);
  or g_135197_(out[641], out[640], _045437_);
  or g_135198_(out[640], _055356_, _045438_);
  and g_135199_(out[643], _045438_, _045439_);
  and g_135200_(_023479_, _045438_, _045441_);
  xor g_135201_(out[644], _045439_, _045442_);
  xor g_135202_(_055711_, _045439_, _045443_);
  and g_135203_(_045295_, _045428_, _045444_);
  or g_135204_(_045294_, _045430_, _045445_);
  and g_135205_(_045302_, _045430_, _045446_);
  or g_135206_(_045301_, _045428_, _045447_);
  and g_135207_(_045445_, _045447_, _045448_);
  or g_135208_(_045444_, _045446_, _045449_);
  and g_135209_(_045443_, _045448_, _045450_);
  or g_135210_(_045442_, _045449_, _045452_);
  xor g_135211_(out[643], _045438_, _045453_);
  xor g_135212_(_055755_, _045438_, _045454_);
  and g_135213_(_045342_, _045428_, _045455_);
  or g_135214_(_045340_, _045430_, _045456_);
  and g_135215_(_045348_, _045430_, _045457_);
  or g_135216_(_045347_, _045428_, _045458_);
  and g_135217_(_045456_, _045458_, _045459_);
  or g_135218_(_045455_, _045457_, _045460_);
  and g_135219_(_045453_, _045460_, _045461_);
  or g_135220_(_045454_, _045459_, _045463_);
  xor g_135221_(_055722_, out[640], _045464_);
  not g_135222_(_045464_, _045465_);
  and g_135223_(_045368_, _045430_, _045466_);
  or g_135224_(_045367_, _045428_, _045467_);
  and g_135225_(_045362_, _045428_, _045468_);
  or g_135226_(_045364_, _045430_, _045469_);
  and g_135227_(_045467_, _045469_, _045470_);
  or g_135228_(_045466_, _045468_, _045471_);
  and g_135229_(_045465_, _045470_, _045472_);
  or g_135230_(_045464_, _045471_, _045474_);
  and g_135231_(out[624], _045428_, _045475_);
  or g_135232_(_055601_, _045430_, _045476_);
  and g_135233_(_045377_, _045430_, _045477_);
  or g_135234_(_045376_, _045428_, _045478_);
  and g_135235_(_045476_, _045478_, _045479_);
  or g_135236_(_045475_, _045477_, _045480_);
  and g_135237_(out[640], _045479_, _045481_);
  or g_135238_(_055733_, _045480_, _045482_);
  and g_135239_(_045474_, _045482_, _045483_);
  or g_135240_(_045472_, _045481_, _045485_);
  xor g_135241_(out[642], _045437_, _045486_);
  not g_135242_(_045486_, _045487_);
  and g_135243_(_045329_, _045428_, _045488_);
  or g_135244_(_045331_, _045430_, _045489_);
  and g_135245_(_045337_, _045430_, _045490_);
  or g_135246_(_045336_, _045428_, _045491_);
  and g_135247_(_045489_, _045491_, _045492_);
  or g_135248_(_045488_, _045490_, _045493_);
  and g_135249_(_045487_, _045493_, _045494_);
  or g_135250_(_045486_, _045492_, _045496_);
  and g_135251_(out[641], _045471_, _045497_);
  or g_135252_(_055722_, _045470_, _045498_);
  and g_135253_(_045496_, _045498_, _045499_);
  or g_135254_(_045494_, _045497_, _045500_);
  and g_135255_(_045485_, _045499_, _045501_);
  or g_135256_(_045483_, _045500_, _045502_);
  and g_135257_(_045454_, _045459_, _045503_);
  or g_135258_(_045453_, _045460_, _045504_);
  and g_135259_(_045486_, _045492_, _045505_);
  or g_135260_(_045487_, _045493_, _045507_);
  and g_135261_(_045504_, _045507_, _045508_);
  or g_135262_(_045503_, _045505_, _045509_);
  and g_135263_(_045502_, _045508_, _045510_);
  or g_135264_(_045501_, _045509_, _045511_);
  and g_135265_(_045463_, _045511_, _045512_);
  or g_135266_(_045461_, _045510_, _045513_);
  and g_135267_(_045452_, _045513_, _045514_);
  or g_135268_(_045450_, _045512_, _045515_);
  and g_135269_(out[645], _045441_, _045516_);
  xor g_135270_(out[645], _045441_, _045518_);
  xor g_135271_(_055700_, _045441_, _045519_);
  and g_135272_(_045282_, _045428_, _045520_);
  or g_135273_(_045281_, _045430_, _045521_);
  and g_135274_(_045289_, _045430_, _045522_);
  or g_135275_(_045288_, _045428_, _045523_);
  and g_135276_(_045521_, _045523_, _045524_);
  or g_135277_(_045520_, _045522_, _045525_);
  and g_135278_(_045518_, _045525_, _045526_);
  or g_135279_(_045519_, _045524_, _045527_);
  and g_135280_(_045442_, _045449_, _045529_);
  or g_135281_(_045443_, _045448_, _045530_);
  and g_135282_(_045527_, _045530_, _045531_);
  or g_135283_(_045526_, _045529_, _045532_);
  and g_135284_(_045515_, _045531_, _045533_);
  or g_135285_(_045514_, _045532_, _045534_);
  or g_135286_(out[646], _045516_, _045535_);
  xor g_135287_(out[646], _045516_, _045536_);
  xor g_135288_(_055689_, _045516_, _045537_);
  and g_135289_(_045267_, _045430_, _045538_);
  or g_135290_(_045266_, _045428_, _045540_);
  and g_135291_(_045259_, _045428_, _045541_);
  or g_135292_(_045260_, _045430_, _045542_);
  and g_135293_(_045540_, _045542_, _045543_);
  or g_135294_(_045538_, _045541_, _045544_);
  and g_135295_(_045536_, _045543_, _045545_);
  or g_135296_(_045537_, _045544_, _045546_);
  and g_135297_(_045519_, _045524_, _045547_);
  or g_135298_(_045518_, _045525_, _045548_);
  and g_135299_(_045546_, _045548_, _045549_);
  or g_135300_(_045545_, _045547_, _045551_);
  and g_135301_(_045534_, _045549_, _045552_);
  or g_135302_(_045533_, _045551_, _045553_);
  and g_135303_(out[647], _045535_, _045554_);
  xor g_135304_(out[647], _045535_, _045555_);
  xor g_135305_(_055678_, _045535_, _045556_);
  and g_135306_(_045278_, _045430_, _045557_);
  or g_135307_(_045277_, _045428_, _045558_);
  and g_135308_(_045271_, _045428_, _045559_);
  or g_135309_(_045270_, _045430_, _045560_);
  and g_135310_(_045558_, _045560_, _045562_);
  or g_135311_(_045557_, _045559_, _045563_);
  and g_135312_(_045555_, _045563_, _045564_);
  or g_135313_(_045556_, _045562_, _045565_);
  and g_135314_(_045537_, _045544_, _045566_);
  or g_135315_(_045536_, _045543_, _045567_);
  and g_135316_(_045565_, _045567_, _045568_);
  or g_135317_(_045564_, _045566_, _045569_);
  and g_135318_(_045553_, _045568_, _045570_);
  or g_135319_(_045552_, _045569_, _045571_);
  and g_135320_(out[648], _045554_, _045573_);
  or g_135321_(out[649], _045573_, _045574_);
  and g_135322_(out[650], _045574_, _045575_);
  xor g_135323_(out[651], _045575_, _045576_);
  xor g_135324_(_055667_, _045575_, _045577_);
  and g_135325_(_045205_, _045428_, _045578_);
  or g_135326_(_045204_, _045430_, _045579_);
  and g_135327_(_045192_, _045430_, _045580_);
  or g_135328_(_045191_, _045428_, _045581_);
  and g_135329_(_045579_, _045581_, _045582_);
  or g_135330_(_045578_, _045580_, _045584_);
  and g_135331_(_045577_, _045582_, _045585_);
  or g_135332_(_045576_, _045584_, _045586_);
  xor g_135333_(out[650], _045574_, _045587_);
  xor g_135334_(_055788_, _045574_, _045588_);
  and g_135335_(_045435_, _045588_, _045589_);
  or g_135336_(_045436_, _045587_, _045590_);
  and g_135337_(_045556_, _045562_, _045591_);
  or g_135338_(_045555_, _045563_, _045592_);
  and g_135339_(_045436_, _045587_, _045593_);
  or g_135340_(_045435_, _045588_, _045595_);
  or g_135341_(_045192_, _045428_, _045596_);
  or g_135342_(_045205_, _045430_, _045597_);
  and g_135343_(_045596_, _045597_, _045598_);
  and g_135344_(_045576_, _045584_, _045599_);
  or g_135345_(_045577_, _045582_, _045600_);
  and g_135346_(_045595_, _045600_, _045601_);
  or g_135347_(_045593_, _045599_, _045602_);
  xor g_135348_(out[649], _045573_, _045603_);
  xor g_135349_(_055777_, _045573_, _045604_);
  and g_135350_(_045216_, _045430_, _045606_);
  or g_135351_(_045215_, _045428_, _045607_);
  and g_135352_(_045208_, _045428_, _045608_);
  or g_135353_(_045210_, _045430_, _045609_);
  and g_135354_(_045607_, _045609_, _045610_);
  or g_135355_(_045606_, _045608_, _045611_);
  and g_135356_(_045604_, _045611_, _045612_);
  or g_135357_(_045603_, _045610_, _045613_);
  xor g_135358_(out[648], _045554_, _045614_);
  not g_135359_(_045614_, _045615_);
  and g_135360_(_045234_, _045430_, _045617_);
  or g_135361_(_045233_, _045428_, _045618_);
  and g_135362_(_045227_, _045428_, _045619_);
  or g_135363_(_045226_, _045430_, _045620_);
  and g_135364_(_045618_, _045620_, _045621_);
  or g_135365_(_045617_, _045619_, _045622_);
  and g_135366_(_045603_, _045610_, _045623_);
  or g_135367_(_045604_, _045611_, _045624_);
  and g_135368_(_045614_, _045622_, _045625_);
  or g_135369_(_045615_, _045621_, _045626_);
  and g_135370_(_045590_, _045601_, _045628_);
  or g_135371_(_045589_, _045602_, _045629_);
  and g_135372_(_045586_, _045628_, _045630_);
  or g_135373_(_045585_, _045629_, _045631_);
  xor g_135374_(_045615_, _045621_, _045632_);
  xor g_135375_(_045614_, _045621_, _045633_);
  and g_135376_(_045613_, _045624_, _045634_);
  or g_135377_(_045612_, _045623_, _045635_);
  and g_135378_(_045592_, _045634_, _045636_);
  or g_135379_(_045591_, _045635_, _045637_);
  and g_135380_(_045632_, _045636_, _045639_);
  or g_135381_(_045633_, _045637_, _045640_);
  and g_135382_(_045630_, _045639_, _045641_);
  or g_135383_(_045631_, _045640_, _045642_);
  and g_135384_(_045571_, _045641_, _045643_);
  or g_135385_(_045570_, _045642_, _045644_);
  and g_135386_(_045613_, _045626_, _045645_);
  or g_135387_(_045612_, _045625_, _045646_);
  or g_135388_(_045623_, _045645_, _045647_);
  and g_135389_(_045624_, _045646_, _045648_);
  and g_135390_(_045590_, _045648_, _045650_);
  or g_135391_(_045589_, _045647_, _045651_);
  and g_135392_(_045601_, _045651_, _045652_);
  or g_135393_(_045602_, _045650_, _045653_);
  and g_135394_(_045586_, _045653_, _045654_);
  or g_135395_(_045585_, _045652_, _045655_);
  and g_135396_(_045644_, _045655_, _045656_);
  or g_135397_(_045643_, _045654_, _045657_);
  and g_135398_(_045436_, _045657_, _045658_);
  or g_135399_(_045435_, _045656_, _045659_);
  and g_135400_(_045588_, _045656_, _045661_);
  or g_135401_(_045587_, _045657_, _045662_);
  and g_135402_(_045659_, _045662_, _045663_);
  or g_135403_(_045658_, _045661_, _045664_);
  and g_135404_(_043433_, _045663_, _045665_);
  or g_135405_(_043432_, _045664_, _045666_);
  xor g_135406_(out[667], _043431_, _045667_);
  xor g_135407_(_055799_, _043431_, _045668_);
  and g_135408_(_045576_, _045582_, _045669_);
  or g_135409_(_045577_, _045584_, _045670_);
  and g_135410_(_045668_, _045669_, _045672_);
  or g_135411_(_045667_, _045670_, _045673_);
  or g_135412_(_045577_, _045598_, _045674_);
  and g_135413_(_045666_, _045673_, _045675_);
  or g_135414_(_045665_, _045672_, _045676_);
  and g_135415_(_045667_, _045670_, _045677_);
  or g_135416_(_045668_, _045669_, _045678_);
  and g_135417_(_043432_, _045664_, _045679_);
  or g_135418_(_043433_, _045663_, _045680_);
  and g_135419_(_045678_, _045680_, _045681_);
  or g_135420_(_045677_, _045679_, _045683_);
  and g_135421_(_045675_, _045681_, _045684_);
  or g_135422_(_045676_, _045683_, _045685_);
  xor g_135423_(out[664], _043425_, _045686_);
  xor g_135424_(_055898_, _043425_, _045687_);
  and g_135425_(_045622_, _045657_, _045688_);
  or g_135426_(_045621_, _045656_, _045689_);
  and g_135427_(_045615_, _045656_, _045690_);
  or g_135428_(_045614_, _045657_, _045691_);
  and g_135429_(_045689_, _045691_, _045692_);
  or g_135430_(_045688_, _045690_, _045694_);
  and g_135431_(_045687_, _045692_, _045695_);
  or g_135432_(_045686_, _045694_, _045696_);
  xor g_135433_(out[665], _043429_, _045697_);
  xor g_135434_(_055909_, _043429_, _045698_);
  and g_135435_(_045611_, _045657_, _045699_);
  or g_135436_(_045610_, _045656_, _045700_);
  and g_135437_(_045603_, _045656_, _045701_);
  or g_135438_(_045604_, _045657_, _045702_);
  and g_135439_(_045700_, _045702_, _045703_);
  or g_135440_(_045699_, _045701_, _045705_);
  and g_135441_(_045697_, _045703_, _045706_);
  or g_135442_(_045698_, _045705_, _045707_);
  and g_135443_(_045696_, _045707_, _045708_);
  or g_135444_(_045695_, _045706_, _045709_);
  and g_135445_(_045698_, _045705_, _045710_);
  or g_135446_(_045697_, _045703_, _045711_);
  and g_135447_(_045686_, _045694_, _045712_);
  or g_135448_(_045687_, _045692_, _045713_);
  and g_135449_(_045711_, _045713_, _045714_);
  or g_135450_(_045710_, _045712_, _045716_);
  and g_135451_(_045708_, _045714_, _045717_);
  or g_135452_(_045709_, _045716_, _045718_);
  and g_135453_(_045684_, _045717_, _045719_);
  or g_135454_(_045685_, _045718_, _045720_);
  xor g_135455_(out[660], _043421_, _045721_);
  xor g_135456_(_055843_, _043421_, _045722_);
  and g_135457_(_045443_, _045656_, _045723_);
  or g_135458_(_045442_, _045657_, _045724_);
  and g_135459_(_045449_, _045657_, _045725_);
  or g_135460_(_045448_, _045656_, _045727_);
  and g_135461_(_045724_, _045727_, _045728_);
  or g_135462_(_045723_, _045725_, _045729_);
  and g_135463_(_045722_, _045728_, _045730_);
  or g_135464_(_045721_, _045729_, _045731_);
  xor g_135465_(out[661], _043422_, _045732_);
  xor g_135466_(_055832_, _043422_, _045733_);
  and g_135467_(_045519_, _045656_, _045734_);
  or g_135468_(_045518_, _045657_, _045735_);
  and g_135469_(_045525_, _045657_, _045736_);
  or g_135470_(_045524_, _045656_, _045738_);
  and g_135471_(_045735_, _045738_, _045739_);
  or g_135472_(_045734_, _045736_, _045740_);
  and g_135473_(_045733_, _045739_, _045741_);
  or g_135474_(_045732_, _045740_, _045742_);
  and g_135475_(_045731_, _045742_, _045743_);
  or g_135476_(_045730_, _045741_, _045744_);
  xor g_135477_(out[662], _043423_, _045745_);
  not g_135478_(_045745_, _045746_);
  or g_135479_(_045543_, _045656_, _045747_);
  not g_135480_(_045747_, _045749_);
  and g_135481_(_045536_, _045656_, _045750_);
  not g_135482_(_045750_, _045751_);
  and g_135483_(_045747_, _045751_, _045752_);
  or g_135484_(_045749_, _045750_, _045753_);
  and g_135485_(_045745_, _045752_, _045754_);
  or g_135486_(_045746_, _045753_, _045755_);
  and g_135487_(_045563_, _045657_, _045756_);
  or g_135488_(_045562_, _045656_, _045757_);
  and g_135489_(_045556_, _045656_, _045758_);
  or g_135490_(_045555_, _045657_, _045760_);
  and g_135491_(_045757_, _045760_, _045761_);
  or g_135492_(_045756_, _045758_, _045762_);
  and g_135493_(_043426_, _045762_, _045763_);
  or g_135494_(_043428_, _045761_, _045764_);
  and g_135495_(_045732_, _045740_, _045765_);
  or g_135496_(_045733_, _045739_, _045766_);
  and g_135497_(_043428_, _045761_, _045767_);
  or g_135498_(_043426_, _045762_, _045768_);
  xor g_135499_(_045745_, _045752_, _045769_);
  xor g_135500_(_045746_, _045752_, _045771_);
  and g_135501_(_045764_, _045768_, _045772_);
  or g_135502_(_045763_, _045767_, _045773_);
  and g_135503_(_045769_, _045772_, _045774_);
  or g_135504_(_045771_, _045773_, _045775_);
  and g_135505_(_045766_, _045774_, _045776_);
  or g_135506_(_045765_, _045775_, _045777_);
  and g_135507_(_045744_, _045776_, _045778_);
  or g_135508_(_045743_, _045777_, _045779_);
  and g_135509_(_045754_, _045764_, _045780_);
  or g_135510_(_045755_, _045763_, _045782_);
  and g_135511_(_045768_, _045782_, _045783_);
  or g_135512_(_045767_, _045780_, _045784_);
  and g_135513_(_045779_, _045783_, _045785_);
  or g_135514_(_045778_, _045784_, _045786_);
  and g_135515_(_045719_, _045786_, _045787_);
  or g_135516_(_045720_, _045785_, _045788_);
  xor g_135517_(out[659], _043420_, _045789_);
  xor g_135518_(_055887_, _043420_, _045790_);
  and g_135519_(_045454_, _045656_, _045791_);
  not g_135520_(_045791_, _045793_);
  or g_135521_(_045459_, _045656_, _045794_);
  not g_135522_(_045794_, _045795_);
  and g_135523_(_045793_, _045794_, _045796_);
  or g_135524_(_045791_, _045795_, _045797_);
  and g_135525_(_045790_, _045796_, _045798_);
  or g_135526_(_045789_, _045797_, _045799_);
  xor g_135527_(out[658], _043419_, _045800_);
  xor g_135528_(_055876_, _043419_, _045801_);
  or g_135529_(_045492_, _045656_, _045802_);
  not g_135530_(_045802_, _045804_);
  and g_135531_(_045486_, _045656_, _045805_);
  not g_135532_(_045805_, _045806_);
  and g_135533_(_045802_, _045806_, _045807_);
  or g_135534_(_045804_, _045805_, _045808_);
  and g_135535_(_045800_, _045807_, _045809_);
  or g_135536_(_045801_, _045808_, _045810_);
  and g_135537_(_045799_, _045810_, _045811_);
  or g_135538_(_045798_, _045809_, _045812_);
  and g_135539_(_045789_, _045797_, _045813_);
  or g_135540_(_045790_, _045796_, _045815_);
  and g_135541_(_045812_, _045815_, _045816_);
  or g_135542_(_045811_, _045813_, _045817_);
  and g_135543_(_045801_, _045808_, _045818_);
  or g_135544_(_045800_, _045807_, _045819_);
  and g_135545_(_045815_, _045819_, _045820_);
  or g_135546_(_045813_, _045818_, _045821_);
  xor g_135547_(out[657], out[656], _045822_);
  not g_135548_(_045822_, _045823_);
  or g_135549_(_045464_, _045657_, _045824_);
  or g_135550_(_045470_, _045656_, _045826_);
  and g_135551_(_045824_, _045826_, _045827_);
  not g_135552_(_045827_, _045828_);
  and g_135553_(_045822_, _045827_, _045829_);
  not g_135554_(_045829_, _045830_);
  and g_135555_(out[640], _045656_, _045831_);
  or g_135556_(_055733_, _045657_, _045832_);
  and g_135557_(_045480_, _045657_, _045833_);
  or g_135558_(_045479_, _045656_, _045834_);
  and g_135559_(_045832_, _045834_, _045835_);
  or g_135560_(_045831_, _045833_, _045837_);
  and g_135561_(_055865_, _045837_, _045838_);
  or g_135562_(out[656], _045835_, _045839_);
  xor g_135563_(_045822_, _045827_, _045840_);
  xor g_135564_(_045823_, _045827_, _045841_);
  and g_135565_(_045839_, _045840_, _045842_);
  or g_135566_(_045838_, _045841_, _045843_);
  and g_135567_(_045830_, _045843_, _045844_);
  or g_135568_(_045829_, _045842_, _045845_);
  and g_135569_(_045820_, _045845_, _045846_);
  or g_135570_(_045821_, _045844_, _045848_);
  and g_135571_(_045817_, _045848_, _045849_);
  or g_135572_(_045816_, _045846_, _045850_);
  and g_135573_(_045721_, _045729_, _045851_);
  or g_135574_(_045722_, _045728_, _045852_);
  and g_135575_(_045766_, _045852_, _045853_);
  or g_135576_(_045765_, _045851_, _045854_);
  and g_135577_(_045743_, _045853_, _045855_);
  or g_135578_(_045744_, _045854_, _045856_);
  and g_135579_(_045774_, _045855_, _045857_);
  or g_135580_(_045775_, _045856_, _045859_);
  and g_135581_(_045719_, _045857_, _045860_);
  or g_135582_(_045720_, _045859_, _045861_);
  and g_135583_(_045850_, _045860_, _045862_);
  or g_135584_(_045849_, _045861_, _045863_);
  and g_135585_(_045676_, _045678_, _045864_);
  or g_135586_(_045675_, _045677_, _045865_);
  and g_135587_(_045709_, _045711_, _045866_);
  or g_135588_(_045708_, _045710_, _045867_);
  and g_135589_(_045684_, _045866_, _045868_);
  or g_135590_(_045685_, _045867_, _045870_);
  and g_135591_(_045865_, _045870_, _045871_);
  or g_135592_(_045864_, _045868_, _045872_);
  and g_135593_(_045863_, _045871_, _045873_);
  or g_135594_(_045862_, _045872_, _045874_);
  and g_135595_(_045788_, _045873_, _045875_);
  or g_135596_(_045787_, _045874_, _045876_);
  and g_135597_(out[656], _045835_, _045877_);
  or g_135598_(_055865_, _045837_, _045878_);
  and g_135599_(_045811_, _045878_, _045879_);
  or g_135600_(_045812_, _045877_, _045881_);
  and g_135601_(_045820_, _045879_, _045882_);
  or g_135602_(_045821_, _045881_, _045883_);
  and g_135603_(_045860_, _045882_, _045884_);
  or g_135604_(_045861_, _045883_, _045885_);
  and g_135605_(_045842_, _045884_, _045886_);
  or g_135606_(_045843_, _045885_, _045887_);
  and g_135607_(_045876_, _045887_, _045888_);
  or g_135608_(_045875_, _045886_, _045889_);
  and g_135609_(_043428_, _045888_, _045890_);
  not g_135610_(_045890_, _045892_);
  or g_135611_(_045761_, _045888_, _045893_);
  not g_135612_(_045893_, _045894_);
  and g_135613_(_045892_, _045893_, _045895_);
  or g_135614_(_045890_, _045894_, _045896_);
  or g_135615_(out[673], out[672], _045897_);
  or g_135616_(out[672], _055741_, _045898_);
  xor g_135617_(out[674], _045897_, _045899_);
  xor g_135618_(_000043_, _045897_, _045900_);
  and g_135619_(_045800_, _045888_, _045901_);
  not g_135620_(_045901_, _045903_);
  or g_135621_(_045807_, _045888_, _045904_);
  not g_135622_(_045904_, _045905_);
  and g_135623_(_045903_, _045904_, _045906_);
  or g_135624_(_045901_, _045905_, _045907_);
  and g_135625_(_045899_, _045906_, _045908_);
  or g_135626_(_045900_, _045907_, _045909_);
  and g_135627_(_045828_, _045889_, _045910_);
  or g_135628_(_045827_, _045888_, _045911_);
  and g_135629_(_045822_, _045888_, _045912_);
  or g_135630_(_045823_, _045889_, _045914_);
  and g_135631_(_045911_, _045914_, _045915_);
  or g_135632_(_045910_, _045912_, _045916_);
  and g_135633_(out[673], _045916_, _045917_);
  or g_135634_(_000021_, _045915_, _045918_);
  xor g_135635_(out[673], out[672], _045919_);
  xor g_135636_(_000021_, out[672], _045920_);
  and g_135637_(_045915_, _045919_, _045921_);
  or g_135638_(_045916_, _045920_, _045922_);
  and g_135639_(out[656], _045888_, _045923_);
  or g_135640_(_055865_, _045889_, _045925_);
  and g_135641_(_045837_, _045889_, _045926_);
  or g_135642_(_045835_, _045888_, _045927_);
  and g_135643_(_045925_, _045927_, _045928_);
  or g_135644_(_045923_, _045926_, _045929_);
  and g_135645_(out[672], _045928_, _045930_);
  or g_135646_(_000032_, _045929_, _045931_);
  and g_135647_(_045922_, _045931_, _045932_);
  or g_135648_(_045921_, _045930_, _045933_);
  and g_135649_(_045918_, _045933_, _045934_);
  or g_135650_(_045917_, _045932_, _045936_);
  and g_135651_(_045909_, _045936_, _045937_);
  or g_135652_(_045908_, _045934_, _045938_);
  and g_135653_(_045900_, _045907_, _045939_);
  or g_135654_(_045899_, _045906_, _045940_);
  and g_135655_(out[675], _045898_, _045941_);
  xor g_135656_(out[675], _045898_, _045942_);
  xor g_135657_(_000054_, _045898_, _045943_);
  and g_135658_(_045790_, _045888_, _045944_);
  not g_135659_(_045944_, _045945_);
  or g_135660_(_045796_, _045888_, _045947_);
  not g_135661_(_045947_, _045948_);
  and g_135662_(_045945_, _045947_, _045949_);
  or g_135663_(_045944_, _045948_, _045950_);
  and g_135664_(_045942_, _045950_, _045951_);
  or g_135665_(_045943_, _045949_, _045952_);
  and g_135666_(_045940_, _045952_, _045953_);
  or g_135667_(_045939_, _045951_, _045954_);
  and g_135668_(_045938_, _045953_, _045955_);
  or g_135669_(_045937_, _045954_, _045956_);
  and g_135670_(_023933_, _045898_, _045958_);
  xor g_135671_(out[676], _045941_, _045959_);
  xor g_135672_(_000010_, _045941_, _045960_);
  and g_135673_(_045722_, _045888_, _045961_);
  not g_135674_(_045961_, _045962_);
  or g_135675_(_045728_, _045888_, _045963_);
  not g_135676_(_045963_, _045964_);
  and g_135677_(_045962_, _045963_, _045965_);
  or g_135678_(_045961_, _045964_, _045966_);
  and g_135679_(_045960_, _045965_, _045967_);
  or g_135680_(_045959_, _045966_, _045969_);
  and g_135681_(_045943_, _045949_, _045970_);
  or g_135682_(_045942_, _045950_, _045971_);
  and g_135683_(_045969_, _045971_, _045972_);
  or g_135684_(_045967_, _045970_, _045973_);
  and g_135685_(_045956_, _045972_, _045974_);
  or g_135686_(_045955_, _045973_, _045975_);
  and g_135687_(out[677], _045958_, _045976_);
  xor g_135688_(out[677], _045958_, _045977_);
  xor g_135689_(_055964_, _045958_, _045978_);
  and g_135690_(_045733_, _045888_, _045980_);
  not g_135691_(_045980_, _045981_);
  or g_135692_(_045739_, _045888_, _045982_);
  not g_135693_(_045982_, _045983_);
  and g_135694_(_045981_, _045982_, _045984_);
  or g_135695_(_045980_, _045983_, _045985_);
  and g_135696_(_045977_, _045985_, _045986_);
  or g_135697_(_045978_, _045984_, _045987_);
  and g_135698_(_045959_, _045966_, _045988_);
  or g_135699_(_045960_, _045965_, _045989_);
  and g_135700_(_045987_, _045989_, _045991_);
  or g_135701_(_045986_, _045988_, _045992_);
  and g_135702_(_045975_, _045991_, _045993_);
  or g_135703_(_045974_, _045992_, _045994_);
  or g_135704_(out[678], _045976_, _045995_);
  xor g_135705_(out[678], _045976_, _045996_);
  xor g_135706_(_055953_, _045976_, _045997_);
  and g_135707_(_045745_, _045888_, _045998_);
  not g_135708_(_045998_, _045999_);
  or g_135709_(_045752_, _045888_, _046000_);
  not g_135710_(_046000_, _046002_);
  and g_135711_(_045999_, _046000_, _046003_);
  or g_135712_(_045998_, _046002_, _046004_);
  and g_135713_(_045996_, _046003_, _046005_);
  or g_135714_(_045997_, _046004_, _046006_);
  and g_135715_(_045978_, _045984_, _046007_);
  or g_135716_(_045977_, _045985_, _046008_);
  and g_135717_(_046006_, _046008_, _046009_);
  or g_135718_(_046005_, _046007_, _046010_);
  and g_135719_(_045994_, _046009_, _046011_);
  or g_135720_(_045993_, _046010_, _046013_);
  and g_135721_(out[679], _045995_, _046014_);
  xor g_135722_(out[679], _045995_, _046015_);
  xor g_135723_(_055942_, _045995_, _046016_);
  and g_135724_(_045896_, _046015_, _046017_);
  or g_135725_(_045895_, _046016_, _046018_);
  and g_135726_(_045997_, _046004_, _046019_);
  or g_135727_(_045996_, _046003_, _046020_);
  and g_135728_(_046018_, _046020_, _046021_);
  or g_135729_(_046017_, _046019_, _046022_);
  and g_135730_(_046013_, _046021_, _046024_);
  or g_135731_(_046011_, _046022_, _046025_);
  and g_135732_(out[680], _046014_, _046026_);
  or g_135733_(out[681], _046026_, _046027_);
  and g_135734_(out[682], _046027_, _046028_);
  xor g_135735_(out[682], _046027_, _046029_);
  and g_135736_(_043433_, _045888_, _046030_);
  not g_135737_(_046030_, _046031_);
  or g_135738_(_045663_, _045888_, _046032_);
  not g_135739_(_046032_, _046033_);
  and g_135740_(_046031_, _046032_, _046035_);
  or g_135741_(_046030_, _046033_, _046036_);
  and g_135742_(_046029_, _046036_, _046037_);
  xor g_135743_(out[683], _046028_, _046038_);
  xor g_135744_(_055931_, _046028_, _046039_);
  and g_135745_(_045668_, _045888_, _046040_);
  not g_135746_(_046040_, _046041_);
  or g_135747_(_045669_, _045888_, _046042_);
  not g_135748_(_046042_, _046043_);
  and g_135749_(_046041_, _046042_, _046044_);
  or g_135750_(_046040_, _046043_, _046046_);
  or g_135751_(_045674_, _045888_, _046047_);
  not g_135752_(_046047_, _046048_);
  and g_135753_(_045667_, _045888_, _046049_);
  not g_135754_(_046049_, _046050_);
  and g_135755_(_046047_, _046050_, _046051_);
  or g_135756_(_046048_, _046049_, _046052_);
  and g_135757_(_046038_, _046051_, _046053_);
  or g_135758_(_046038_, _046046_, _046054_);
  xor g_135759_(_046029_, _046036_, _046055_);
  xor g_135760_(_046029_, _046035_, _046057_);
  xor g_135761_(_046038_, _046051_, _046058_);
  xor g_135762_(_046039_, _046051_, _046059_);
  and g_135763_(_046055_, _046058_, _046060_);
  or g_135764_(_046057_, _046059_, _046061_);
  xor g_135765_(out[680], _046014_, _046062_);
  xor g_135766_(_000065_, _046014_, _046063_);
  and g_135767_(_045687_, _045888_, _046064_);
  not g_135768_(_046064_, _046065_);
  or g_135769_(_045692_, _045888_, _046066_);
  not g_135770_(_046066_, _046068_);
  and g_135771_(_046065_, _046066_, _046069_);
  or g_135772_(_046064_, _046068_, _046070_);
  and g_135773_(_046063_, _046069_, _046071_);
  or g_135774_(_046062_, _046070_, _046072_);
  xor g_135775_(out[681], _046026_, _046073_);
  xor g_135776_(_000076_, _046026_, _046074_);
  and g_135777_(_045697_, _045888_, _046075_);
  not g_135778_(_046075_, _046076_);
  or g_135779_(_045703_, _045888_, _046077_);
  not g_135780_(_046077_, _046079_);
  and g_135781_(_046076_, _046077_, _046080_);
  or g_135782_(_046075_, _046079_, _046081_);
  and g_135783_(_046074_, _046081_, _046082_);
  or g_135784_(_046073_, _046080_, _046083_);
  and g_135785_(_046073_, _046080_, _046084_);
  or g_135786_(_046074_, _046081_, _046085_);
  and g_135787_(_046062_, _046070_, _046086_);
  or g_135788_(_046063_, _046069_, _046087_);
  and g_135789_(_045895_, _046016_, _046088_);
  or g_135790_(_045896_, _046015_, _046090_);
  and g_135791_(_046072_, _046090_, _046091_);
  or g_135792_(_046071_, _046088_, _046092_);
  and g_135793_(_046083_, _046085_, _046093_);
  or g_135794_(_046082_, _046084_, _046094_);
  and g_135795_(_046091_, _046093_, _046095_);
  or g_135796_(_046092_, _046094_, _046096_);
  and g_135797_(_046060_, _046095_, _046097_);
  or g_135798_(_046061_, _046096_, _046098_);
  and g_135799_(_046087_, _046097_, _046099_);
  or g_135800_(_046086_, _046098_, _046101_);
  and g_135801_(_046025_, _046099_, _046102_);
  or g_135802_(_046024_, _046101_, _046103_);
  and g_135803_(_046083_, _046087_, _046104_);
  or g_135804_(_046082_, _046086_, _046105_);
  and g_135805_(_046060_, _046105_, _046106_);
  or g_135806_(_046061_, _046104_, _046107_);
  and g_135807_(_046085_, _046106_, _046108_);
  or g_135808_(_046084_, _046107_, _046109_);
  and g_135809_(_046037_, _046054_, _046110_);
  or g_135810_(_046053_, _046110_, _046112_);
  not g_135811_(_046112_, _046113_);
  and g_135812_(_046109_, _046113_, _046114_);
  or g_135813_(_046108_, _046112_, _046115_);
  and g_135814_(_046103_, _046114_, _046116_);
  or g_135815_(_046102_, _046115_, _046117_);
  and g_135816_(_045896_, _046117_, _046118_);
  not g_135817_(_046118_, _046119_);
  or g_135818_(_046015_, _046117_, _046120_);
  not g_135819_(_046120_, _046121_);
  and g_135820_(_046119_, _046120_, _046123_);
  or g_135821_(_046118_, _046121_, _046124_);
  or g_135822_(out[689], out[688], _046125_);
  or g_135823_(out[688], _055929_, _046126_);
  and g_135824_(out[691], _046126_, _046127_);
  and g_135825_(_024161_, _046126_, _046128_);
  and g_135826_(out[693], _046128_, _046129_);
  or g_135827_(out[694], _046129_, _046130_);
  and g_135828_(out[695], _046130_, _046131_);
  xor g_135829_(out[695], _046130_, _046132_);
  xor g_135830_(_000109_, _046130_, _046134_);
  and g_135831_(_046124_, _046132_, _046135_);
  or g_135832_(_046123_, _046134_, _046136_);
  xor g_135833_(out[694], _046129_, _046137_);
  xor g_135834_(_000120_, _046129_, _046138_);
  and g_135835_(_046004_, _046117_, _046139_);
  not g_135836_(_046139_, _046140_);
  or g_135837_(_045997_, _046117_, _046141_);
  not g_135838_(_046141_, _046142_);
  and g_135839_(_046140_, _046141_, _046143_);
  or g_135840_(_046139_, _046142_, _046145_);
  and g_135841_(_046137_, _046143_, _046146_);
  or g_135842_(_046138_, _046145_, _046147_);
  xor g_135843_(out[691], _046126_, _046148_);
  xor g_135844_(_000186_, _046126_, _046149_);
  or g_135845_(_045942_, _046117_, _046150_);
  not g_135846_(_046150_, _046151_);
  and g_135847_(_045950_, _046117_, _046152_);
  not g_135848_(_046152_, _046153_);
  and g_135849_(_046150_, _046153_, _046154_);
  or g_135850_(_046151_, _046152_, _046156_);
  and g_135851_(_046149_, _046154_, _046157_);
  or g_135852_(_046148_, _046156_, _046158_);
  xor g_135853_(out[690], _046125_, _046159_);
  xor g_135854_(_000175_, _046125_, _046160_);
  and g_135855_(_045899_, _046116_, _046161_);
  or g_135856_(_045900_, _046117_, _046162_);
  and g_135857_(_045907_, _046117_, _046163_);
  or g_135858_(_045906_, _046116_, _046164_);
  and g_135859_(_046162_, _046164_, _046165_);
  or g_135860_(_046161_, _046163_, _046167_);
  and g_135861_(_046160_, _046167_, _046168_);
  or g_135862_(_046159_, _046165_, _046169_);
  and g_135863_(out[672], _046116_, _046170_);
  or g_135864_(_000032_, _046117_, _046171_);
  and g_135865_(_045929_, _046117_, _046172_);
  or g_135866_(_045928_, _046116_, _046173_);
  and g_135867_(_046171_, _046173_, _046174_);
  or g_135868_(_046170_, _046172_, _046175_);
  and g_135869_(out[688], _046174_, _046176_);
  or g_135870_(_000164_, _046175_, _046178_);
  and g_135871_(_045919_, _046116_, _046179_);
  or g_135872_(_045920_, _046117_, _046180_);
  and g_135873_(_045916_, _046117_, _046181_);
  or g_135874_(_045915_, _046116_, _046182_);
  and g_135875_(_046180_, _046182_, _046183_);
  or g_135876_(_046179_, _046181_, _046184_);
  and g_135877_(out[689], _046184_, _046185_);
  or g_135878_(_000153_, _046183_, _046186_);
  xor g_135879_(out[689], out[688], _046187_);
  xor g_135880_(_000153_, out[688], _046189_);
  and g_135881_(_046176_, _046186_, _046190_);
  or g_135882_(_046178_, _046185_, _046191_);
  and g_135883_(_046159_, _046165_, _046192_);
  or g_135884_(_046160_, _046167_, _046193_);
  and g_135885_(_046183_, _046187_, _046194_);
  or g_135886_(_046184_, _046189_, _046195_);
  and g_135887_(_046193_, _046195_, _046196_);
  or g_135888_(_046192_, _046194_, _046197_);
  and g_135889_(_046191_, _046196_, _046198_);
  or g_135890_(_046190_, _046197_, _046200_);
  and g_135891_(_046169_, _046200_, _046201_);
  or g_135892_(_046168_, _046198_, _046202_);
  and g_135893_(_046158_, _046202_, _046203_);
  or g_135894_(_046157_, _046201_, _046204_);
  and g_135895_(_046148_, _046156_, _046205_);
  or g_135896_(_046149_, _046154_, _046206_);
  xor g_135897_(out[692], _046127_, _046207_);
  xor g_135898_(_000142_, _046127_, _046208_);
  or g_135899_(_045959_, _046117_, _046209_);
  not g_135900_(_046209_, _046211_);
  and g_135901_(_045966_, _046117_, _046212_);
  not g_135902_(_046212_, _046213_);
  and g_135903_(_046209_, _046213_, _046214_);
  or g_135904_(_046211_, _046212_, _046215_);
  and g_135905_(_046207_, _046215_, _046216_);
  or g_135906_(_046208_, _046214_, _046217_);
  and g_135907_(_046206_, _046217_, _046218_);
  or g_135908_(_046205_, _046216_, _046219_);
  and g_135909_(_046204_, _046218_, _046220_);
  or g_135910_(_046203_, _046219_, _046222_);
  xor g_135911_(out[693], _046128_, _046223_);
  xor g_135912_(_000131_, _046128_, _046224_);
  or g_135913_(_045977_, _046117_, _046225_);
  not g_135914_(_046225_, _046226_);
  and g_135915_(_045985_, _046117_, _046227_);
  not g_135916_(_046227_, _046228_);
  and g_135917_(_046225_, _046228_, _046229_);
  or g_135918_(_046226_, _046227_, _046230_);
  and g_135919_(_046224_, _046229_, _046231_);
  or g_135920_(_046223_, _046230_, _046233_);
  and g_135921_(_046208_, _046214_, _046234_);
  or g_135922_(_046207_, _046215_, _046235_);
  and g_135923_(_046233_, _046235_, _046236_);
  or g_135924_(_046231_, _046234_, _046237_);
  and g_135925_(_046222_, _046236_, _046238_);
  or g_135926_(_046220_, _046237_, _046239_);
  and g_135927_(_046138_, _046145_, _046240_);
  or g_135928_(_046137_, _046143_, _046241_);
  and g_135929_(_046223_, _046230_, _046242_);
  or g_135930_(_046224_, _046229_, _046244_);
  and g_135931_(_046241_, _046244_, _046245_);
  or g_135932_(_046240_, _046242_, _046246_);
  and g_135933_(_046239_, _046245_, _046247_);
  or g_135934_(_046238_, _046246_, _046248_);
  and g_135935_(_046147_, _046248_, _046249_);
  or g_135936_(_046146_, _046247_, _046250_);
  and g_135937_(_046136_, _046250_, _046251_);
  or g_135938_(_046135_, _046249_, _046252_);
  and g_135939_(out[696], _046131_, _046253_);
  or g_135940_(out[697], _046253_, _046255_);
  and g_135941_(out[698], _046255_, _046256_);
  xor g_135942_(out[698], _046255_, _046257_);
  xor g_135943_(_000219_, _046255_, _046258_);
  and g_135944_(_046036_, _046117_, _046259_);
  not g_135945_(_046259_, _046260_);
  or g_135946_(_046029_, _046117_, _046261_);
  not g_135947_(_046261_, _046262_);
  and g_135948_(_046260_, _046261_, _046263_);
  or g_135949_(_046259_, _046262_, _046264_);
  and g_135950_(_046257_, _046264_, _046266_);
  or g_135951_(_046258_, _046263_, _046267_);
  xor g_135952_(out[699], _046256_, _046268_);
  xor g_135953_(_000098_, _046256_, _046269_);
  and g_135954_(_046038_, _046044_, _046270_);
  or g_135955_(_046039_, _046046_, _046271_);
  and g_135956_(_046038_, _046052_, _046272_);
  or g_135957_(_046039_, _046051_, _046273_);
  and g_135958_(_046268_, _046273_, _046274_);
  or g_135959_(_046269_, _046272_, _046275_);
  and g_135960_(_046267_, _046275_, _046277_);
  or g_135961_(_046266_, _046274_, _046278_);
  and g_135962_(_046258_, _046263_, _046279_);
  or g_135963_(_046257_, _046264_, _046280_);
  and g_135964_(_046269_, _046270_, _046281_);
  or g_135965_(_046268_, _046271_, _046282_);
  and g_135966_(_046280_, _046282_, _046283_);
  or g_135967_(_046279_, _046281_, _046284_);
  and g_135968_(_046277_, _046283_, _046285_);
  or g_135969_(_046278_, _046284_, _046286_);
  xor g_135970_(out[696], _046131_, _046288_);
  xor g_135971_(_000197_, _046131_, _046289_);
  and g_135972_(_046070_, _046117_, _046290_);
  not g_135973_(_046290_, _046291_);
  or g_135974_(_046062_, _046117_, _046292_);
  not g_135975_(_046292_, _046293_);
  and g_135976_(_046291_, _046292_, _046294_);
  or g_135977_(_046290_, _046293_, _046295_);
  and g_135978_(_046288_, _046295_, _046296_);
  or g_135979_(_046289_, _046294_, _046297_);
  xor g_135980_(out[697], _046253_, _046299_);
  xor g_135981_(_000208_, _046253_, _046300_);
  and g_135982_(_046081_, _046117_, _046301_);
  not g_135983_(_046301_, _046302_);
  or g_135984_(_046074_, _046117_, _046303_);
  not g_135985_(_046303_, _046304_);
  and g_135986_(_046302_, _046303_, _046305_);
  or g_135987_(_046301_, _046304_, _046306_);
  and g_135988_(_046300_, _046306_, _046307_);
  or g_135989_(_046299_, _046305_, _046308_);
  and g_135990_(_046297_, _046308_, _046310_);
  or g_135991_(_046296_, _046307_, _046311_);
  and g_135992_(_046289_, _046294_, _046312_);
  or g_135993_(_046288_, _046295_, _046313_);
  and g_135994_(_046123_, _046134_, _046314_);
  or g_135995_(_046124_, _046132_, _046315_);
  and g_135996_(_046299_, _046305_, _046316_);
  or g_135997_(_046300_, _046306_, _046317_);
  and g_135998_(_046313_, _046317_, _046318_);
  or g_135999_(_046312_, _046316_, _046319_);
  and g_136000_(_046310_, _046318_, _046321_);
  or g_136001_(_046311_, _046319_, _046322_);
  and g_136002_(_046285_, _046321_, _046323_);
  or g_136003_(_046286_, _046322_, _046324_);
  and g_136004_(_046315_, _046323_, _046325_);
  or g_136005_(_046314_, _046324_, _046326_);
  and g_136006_(_046252_, _046325_, _046327_);
  or g_136007_(_046251_, _046326_, _046328_);
  and g_136008_(_046311_, _046317_, _046329_);
  or g_136009_(_046310_, _046316_, _046330_);
  and g_136010_(_046285_, _046329_, _046332_);
  or g_136011_(_046286_, _046330_, _046333_);
  and g_136012_(_046278_, _046282_, _046334_);
  or g_136013_(_046277_, _046281_, _046335_);
  and g_136014_(_046333_, _046335_, _046336_);
  or g_136015_(_046332_, _046334_, _046337_);
  and g_136016_(_046328_, _046336_, _046338_);
  or g_136017_(_046327_, _046337_, _046339_);
  and g_136018_(_046124_, _046339_, _046340_);
  or g_136019_(_046123_, _046338_, _046341_);
  and g_136020_(_046134_, _046338_, _046343_);
  or g_136021_(_046132_, _046339_, _046344_);
  and g_136022_(_046341_, _046344_, _046345_);
  or g_136023_(_046340_, _046343_, _046346_);
  or g_136024_(out[705], out[704], _046347_);
  or g_136025_(out[704], _000140_, _046348_);
  and g_136026_(out[707], _046348_, _046349_);
  and g_136027_(_024374_, _046348_, _046350_);
  and g_136028_(out[709], _046350_, _046351_);
  or g_136029_(out[710], _046351_, _046352_);
  and g_136030_(out[711], _046352_, _046354_);
  xor g_136031_(out[711], _046352_, _046355_);
  xor g_136032_(_000241_, _046352_, _046356_);
  and g_136033_(_046346_, _046355_, _046357_);
  or g_136034_(_046345_, _046356_, _046358_);
  xor g_136035_(out[710], _046351_, _046359_);
  xor g_136036_(_000252_, _046351_, _046360_);
  and g_136037_(_046145_, _046339_, _046361_);
  or g_136038_(_046143_, _046338_, _046362_);
  and g_136039_(_046137_, _046338_, _046363_);
  or g_136040_(_046138_, _046339_, _046365_);
  and g_136041_(_046362_, _046365_, _046366_);
  or g_136042_(_046361_, _046363_, _046367_);
  and g_136043_(_046359_, _046366_, _046368_);
  or g_136044_(_046360_, _046367_, _046369_);
  xor g_136045_(out[709], _046350_, _046370_);
  xor g_136046_(_000263_, _046350_, _046371_);
  and g_136047_(_046224_, _046338_, _046372_);
  or g_136048_(_046223_, _046339_, _046373_);
  and g_136049_(_046230_, _046339_, _046374_);
  or g_136050_(_046229_, _046338_, _046376_);
  and g_136051_(_046373_, _046376_, _046377_);
  or g_136052_(_046372_, _046374_, _046378_);
  and g_136053_(_046371_, _046377_, _046379_);
  or g_136054_(_046370_, _046378_, _046380_);
  xor g_136055_(out[708], _046349_, _046381_);
  xor g_136056_(_000274_, _046349_, _046382_);
  and g_136057_(_046215_, _046339_, _046383_);
  or g_136058_(_046214_, _046338_, _046384_);
  and g_136059_(_046208_, _046338_, _046385_);
  or g_136060_(_046207_, _046339_, _046387_);
  and g_136061_(_046384_, _046387_, _046388_);
  or g_136062_(_046383_, _046385_, _046389_);
  and g_136063_(_046381_, _046389_, _046390_);
  or g_136064_(_046382_, _046388_, _046391_);
  and g_136065_(out[688], _046338_, _046392_);
  or g_136066_(_000164_, _046339_, _046393_);
  and g_136067_(_046175_, _046339_, _046394_);
  or g_136068_(_046174_, _046338_, _046395_);
  and g_136069_(_046393_, _046395_, _046396_);
  or g_136070_(_046392_, _046394_, _046398_);
  and g_136071_(out[704], _046396_, _046399_);
  or g_136072_(_000296_, _046398_, _046400_);
  and g_136073_(_046187_, _046338_, _046401_);
  or g_136074_(_046189_, _046339_, _046402_);
  and g_136075_(_046184_, _046339_, _046403_);
  or g_136076_(_046183_, _046338_, _046404_);
  and g_136077_(_046402_, _046404_, _046405_);
  or g_136078_(_046401_, _046403_, _046406_);
  and g_136079_(out[705], _046406_, _046407_);
  or g_136080_(_000285_, _046405_, _046409_);
  xor g_136081_(out[705], out[704], _046410_);
  xor g_136082_(_000285_, out[704], _046411_);
  and g_136083_(_046399_, _046409_, _046412_);
  or g_136084_(_046400_, _046407_, _046413_);
  xor g_136085_(out[706], _046347_, _046414_);
  xor g_136086_(_000307_, _046347_, _046415_);
  and g_136087_(_046167_, _046339_, _046416_);
  or g_136088_(_046165_, _046338_, _046417_);
  and g_136089_(_046159_, _046338_, _046418_);
  or g_136090_(_046160_, _046339_, _046420_);
  and g_136091_(_046417_, _046420_, _046421_);
  or g_136092_(_046416_, _046418_, _046422_);
  and g_136093_(_046414_, _046421_, _046423_);
  or g_136094_(_046415_, _046422_, _046424_);
  and g_136095_(_046405_, _046410_, _046425_);
  or g_136096_(_046406_, _046411_, _046426_);
  and g_136097_(_046424_, _046426_, _046427_);
  or g_136098_(_046423_, _046425_, _046428_);
  and g_136099_(_046413_, _046427_, _046429_);
  or g_136100_(_046412_, _046428_, _046431_);
  xor g_136101_(out[707], _046348_, _046432_);
  xor g_136102_(_000318_, _046348_, _046433_);
  and g_136103_(_046149_, _046338_, _046434_);
  or g_136104_(_046148_, _046339_, _046435_);
  and g_136105_(_046156_, _046339_, _046436_);
  or g_136106_(_046154_, _046338_, _046437_);
  and g_136107_(_046435_, _046437_, _046438_);
  or g_136108_(_046434_, _046436_, _046439_);
  and g_136109_(_046432_, _046439_, _046440_);
  or g_136110_(_046433_, _046438_, _046442_);
  and g_136111_(_046415_, _046422_, _046443_);
  or g_136112_(_046414_, _046421_, _046444_);
  and g_136113_(_046442_, _046444_, _046445_);
  or g_136114_(_046440_, _046443_, _046446_);
  and g_136115_(_046431_, _046445_, _046447_);
  or g_136116_(_046429_, _046446_, _046448_);
  and g_136117_(_046433_, _046438_, _046449_);
  or g_136118_(_046432_, _046439_, _046450_);
  and g_136119_(_046382_, _046388_, _046451_);
  or g_136120_(_046381_, _046389_, _046453_);
  and g_136121_(_046450_, _046453_, _046454_);
  or g_136122_(_046449_, _046451_, _046455_);
  and g_136123_(_046448_, _046454_, _046456_);
  or g_136124_(_046447_, _046455_, _046457_);
  and g_136125_(_046391_, _046457_, _046458_);
  or g_136126_(_046390_, _046456_, _046459_);
  and g_136127_(_046380_, _046459_, _046460_);
  or g_136128_(_046379_, _046458_, _046461_);
  and g_136129_(_046360_, _046367_, _046462_);
  or g_136130_(_046359_, _046366_, _046464_);
  and g_136131_(_046370_, _046378_, _046465_);
  or g_136132_(_046371_, _046377_, _046466_);
  and g_136133_(_046464_, _046466_, _046467_);
  or g_136134_(_046462_, _046465_, _046468_);
  and g_136135_(_046461_, _046467_, _046469_);
  or g_136136_(_046460_, _046468_, _046470_);
  and g_136137_(_046369_, _046470_, _046471_);
  or g_136138_(_046368_, _046469_, _046472_);
  and g_136139_(_046358_, _046472_, _046473_);
  or g_136140_(_046357_, _046471_, _046475_);
  and g_136141_(out[712], _046354_, _046476_);
  or g_136142_(out[713], _046476_, _046477_);
  and g_136143_(out[714], _046477_, _046478_);
  xor g_136144_(out[714], _046477_, _046479_);
  xor g_136145_(_000351_, _046477_, _046480_);
  and g_136146_(_046264_, _046339_, _046481_);
  or g_136147_(_046263_, _046338_, _046482_);
  and g_136148_(_046258_, _046338_, _046483_);
  or g_136149_(_046257_, _046339_, _046484_);
  and g_136150_(_046482_, _046484_, _046486_);
  or g_136151_(_046481_, _046483_, _046487_);
  and g_136152_(_046479_, _046487_, _046488_);
  or g_136153_(_046480_, _046486_, _046489_);
  xor g_136154_(out[715], _046478_, _046490_);
  xor g_136155_(_000230_, _046478_, _046491_);
  and g_136156_(_046268_, _046270_, _046492_);
  or g_136157_(_046269_, _046271_, _046493_);
  and g_136158_(_046268_, _046272_, _046494_);
  or g_136159_(_046269_, _046273_, _046495_);
  and g_136160_(_046490_, _046495_, _046497_);
  or g_136161_(_046491_, _046494_, _046498_);
  and g_136162_(_046489_, _046498_, _046499_);
  or g_136163_(_046488_, _046497_, _046500_);
  and g_136164_(_046480_, _046486_, _046501_);
  or g_136165_(_046479_, _046487_, _046502_);
  and g_136166_(_046491_, _046492_, _046503_);
  or g_136167_(_046490_, _046493_, _046504_);
  and g_136168_(_046502_, _046504_, _046505_);
  or g_136169_(_046501_, _046503_, _046506_);
  and g_136170_(_046499_, _046505_, _046508_);
  or g_136171_(_046500_, _046506_, _046509_);
  xor g_136172_(out[713], _046476_, _046510_);
  xor g_136173_(_000340_, _046476_, _046511_);
  and g_136174_(_046306_, _046339_, _046512_);
  or g_136175_(_046305_, _046338_, _046513_);
  and g_136176_(_046299_, _046338_, _046514_);
  or g_136177_(_046300_, _046339_, _046515_);
  and g_136178_(_046513_, _046515_, _046516_);
  or g_136179_(_046512_, _046514_, _046517_);
  and g_136180_(_046511_, _046517_, _046519_);
  or g_136181_(_046510_, _046516_, _046520_);
  xor g_136182_(out[712], _046354_, _046521_);
  xor g_136183_(_000329_, _046354_, _046522_);
  and g_136184_(_046295_, _046339_, _046523_);
  or g_136185_(_046294_, _046338_, _046524_);
  and g_136186_(_046289_, _046338_, _046525_);
  or g_136187_(_046288_, _046339_, _046526_);
  and g_136188_(_046524_, _046526_, _046527_);
  or g_136189_(_046523_, _046525_, _046528_);
  and g_136190_(_046521_, _046528_, _046530_);
  or g_136191_(_046522_, _046527_, _046531_);
  and g_136192_(_046520_, _046531_, _046532_);
  or g_136193_(_046519_, _046530_, _046533_);
  and g_136194_(_046345_, _046356_, _046534_);
  or g_136195_(_046346_, _046355_, _046535_);
  and g_136196_(_046522_, _046527_, _046536_);
  or g_136197_(_046521_, _046528_, _046537_);
  and g_136198_(_046510_, _046516_, _046538_);
  or g_136199_(_046511_, _046517_, _046539_);
  and g_136200_(_046537_, _046539_, _046541_);
  or g_136201_(_046536_, _046538_, _046542_);
  and g_136202_(_046535_, _046541_, _046543_);
  or g_136203_(_046534_, _046542_, _046544_);
  and g_136204_(_046532_, _046543_, _046545_);
  or g_136205_(_046533_, _046544_, _046546_);
  and g_136206_(_046508_, _046545_, _046547_);
  or g_136207_(_046509_, _046546_, _046548_);
  and g_136208_(_046475_, _046547_, _046549_);
  or g_136209_(_046473_, _046548_, _046550_);
  and g_136210_(_046500_, _046504_, _046552_);
  or g_136211_(_046499_, _046503_, _046553_);
  and g_136212_(_046533_, _046539_, _046554_);
  or g_136213_(_046532_, _046538_, _046555_);
  and g_136214_(_046508_, _046554_, _046556_);
  or g_136215_(_046509_, _046555_, _046557_);
  and g_136216_(_046553_, _046557_, _046558_);
  or g_136217_(_046552_, _046556_, _046559_);
  and g_136218_(_046550_, _046558_, _046560_);
  or g_136219_(_046549_, _046559_, _046561_);
  and g_136220_(_046346_, _046561_, _046563_);
  or g_136221_(_046345_, _046560_, _046564_);
  and g_136222_(_046356_, _046560_, _046565_);
  or g_136223_(_046355_, _046561_, _046566_);
  and g_136224_(_046564_, _046566_, _046567_);
  or g_136225_(_046563_, _046565_, _046568_);
  or g_136226_(out[721], out[720], _046569_);
  or g_136227_(out[720], _000239_, _046570_);
  and g_136228_(out[723], _046570_, _046571_);
  xor g_136229_(out[723], _046570_, _046572_);
  xor g_136230_(_000450_, _046570_, _046574_);
  and g_136231_(_046433_, _046560_, _046575_);
  or g_136232_(_046432_, _046561_, _046576_);
  and g_136233_(_046439_, _046561_, _046577_);
  or g_136234_(_046438_, _046560_, _046578_);
  and g_136235_(_046576_, _046578_, _046579_);
  or g_136236_(_046575_, _046577_, _046580_);
  and g_136237_(_046572_, _046580_, _046581_);
  or g_136238_(_046574_, _046579_, _046582_);
  xor g_136239_(out[722], _046569_, _046583_);
  not g_136240_(_046583_, _046585_);
  and g_136241_(_046422_, _046561_, _046586_);
  or g_136242_(_046421_, _046560_, _046587_);
  and g_136243_(_046414_, _046560_, _046588_);
  or g_136244_(_046415_, _046561_, _046589_);
  and g_136245_(_046587_, _046589_, _046590_);
  or g_136246_(_046586_, _046588_, _046591_);
  and g_136247_(_046583_, _046590_, _046592_);
  or g_136248_(_046585_, _046591_, _046593_);
  and g_136249_(_046574_, _046579_, _046594_);
  or g_136250_(_046572_, _046580_, _046596_);
  and g_136251_(_046593_, _046596_, _046597_);
  or g_136252_(_046592_, _046594_, _046598_);
  and g_136253_(_046582_, _046598_, _046599_);
  or g_136254_(_046581_, _046597_, _046600_);
  xor g_136255_(out[721], out[720], _046601_);
  not g_136256_(_046601_, _046602_);
  and g_136257_(_046410_, _046560_, _046603_);
  or g_136258_(_046411_, _046561_, _046604_);
  and g_136259_(_046406_, _046561_, _046605_);
  or g_136260_(_046405_, _046560_, _046607_);
  and g_136261_(_046604_, _046607_, _046608_);
  or g_136262_(_046603_, _046605_, _046609_);
  and g_136263_(_046601_, _046608_, _046610_);
  or g_136264_(_046602_, _046609_, _046611_);
  and g_136265_(out[704], _046560_, _046612_);
  or g_136266_(_000296_, _046561_, _046613_);
  and g_136267_(_046398_, _046561_, _046614_);
  not g_136268_(_046614_, _046615_);
  and g_136269_(_046613_, _046615_, _046616_);
  or g_136270_(_046612_, _046614_, _046618_);
  and g_136271_(_000428_, _046618_, _046619_);
  or g_136272_(out[720], _046616_, _046620_);
  xor g_136273_(_046601_, _046608_, _046621_);
  xor g_136274_(_046602_, _046608_, _046622_);
  and g_136275_(_046620_, _046621_, _046623_);
  or g_136276_(_046619_, _046622_, _046624_);
  and g_136277_(_046611_, _046624_, _046625_);
  or g_136278_(_046610_, _046623_, _046626_);
  and g_136279_(_046582_, _046596_, _046627_);
  or g_136280_(_046581_, _046594_, _046629_);
  xor g_136281_(_046583_, _046590_, _046630_);
  xor g_136282_(_046585_, _046590_, _046631_);
  and g_136283_(_046627_, _046630_, _046632_);
  or g_136284_(_046629_, _046631_, _046633_);
  and g_136285_(_046626_, _046632_, _046634_);
  or g_136286_(_046625_, _046633_, _046635_);
  and g_136287_(_046600_, _046635_, _046636_);
  or g_136288_(_046599_, _046634_, _046637_);
  and g_136289_(_024554_, _046570_, _046638_);
  and g_136290_(out[725], _046638_, _046640_);
  or g_136291_(out[726], _046640_, _046641_);
  and g_136292_(out[727], _046641_, _046642_);
  and g_136293_(out[728], _046642_, _046643_);
  or g_136294_(out[729], _046643_, _046644_);
  xor g_136295_(out[729], _046643_, _046645_);
  xor g_136296_(_000472_, _046643_, _046646_);
  and g_136297_(_046517_, _046561_, _046647_);
  or g_136298_(_046516_, _046560_, _046648_);
  and g_136299_(_046510_, _046560_, _046649_);
  or g_136300_(_046511_, _046561_, _046651_);
  and g_136301_(_046648_, _046651_, _046652_);
  or g_136302_(_046647_, _046649_, _046653_);
  and g_136303_(_046646_, _046653_, _046654_);
  or g_136304_(_046645_, _046652_, _046655_);
  and g_136305_(out[730], _046644_, _046656_);
  xor g_136306_(out[731], _046656_, _046657_);
  xor g_136307_(_000362_, _046656_, _046658_);
  and g_136308_(_046490_, _046492_, _046659_);
  or g_136309_(_046491_, _046493_, _046660_);
  and g_136310_(_046490_, _046494_, _046662_);
  or g_136311_(_046491_, _046495_, _046663_);
  and g_136312_(_046657_, _046660_, _046664_);
  or g_136313_(_046658_, _046659_, _046665_);
  xor g_136314_(out[730], _046644_, _046666_);
  xor g_136315_(_000483_, _046644_, _046667_);
  and g_136316_(_046487_, _046561_, _046668_);
  or g_136317_(_046486_, _046560_, _046669_);
  and g_136318_(_046480_, _046560_, _046670_);
  or g_136319_(_046479_, _046561_, _046671_);
  and g_136320_(_046669_, _046671_, _046673_);
  or g_136321_(_046668_, _046670_, _046674_);
  and g_136322_(_046666_, _046674_, _046675_);
  or g_136323_(_046667_, _046673_, _046676_);
  xor g_136324_(out[728], _046642_, _046677_);
  xor g_136325_(_000461_, _046642_, _046678_);
  and g_136326_(_046528_, _046561_, _046679_);
  or g_136327_(_046527_, _046560_, _046680_);
  and g_136328_(_046522_, _046560_, _046681_);
  or g_136329_(_046521_, _046561_, _046682_);
  and g_136330_(_046680_, _046682_, _046684_);
  or g_136331_(_046679_, _046681_, _046685_);
  and g_136332_(_046677_, _046685_, _046686_);
  or g_136333_(_046678_, _046684_, _046687_);
  and g_136334_(_046678_, _046684_, _046688_);
  or g_136335_(_046677_, _046685_, _046689_);
  and g_136336_(_046645_, _046652_, _046690_);
  or g_136337_(_046646_, _046653_, _046691_);
  and g_136338_(_046689_, _046691_, _046692_);
  or g_136339_(_046688_, _046690_, _046693_);
  and g_136340_(_046667_, _046673_, _046695_);
  or g_136341_(_046666_, _046674_, _046696_);
  and g_136342_(_046658_, _046659_, _046697_);
  or g_136343_(_046657_, _046660_, _046698_);
  and g_136344_(_046696_, _046698_, _046699_);
  or g_136345_(_046695_, _046697_, _046700_);
  and g_136346_(_046665_, _046676_, _046701_);
  or g_136347_(_046664_, _046675_, _046702_);
  and g_136348_(_046699_, _046701_, _046703_);
  or g_136349_(_046700_, _046702_, _046704_);
  and g_136350_(_046655_, _046687_, _046706_);
  or g_136351_(_046654_, _046686_, _046707_);
  and g_136352_(_046692_, _046706_, _046708_);
  or g_136353_(_046693_, _046707_, _046709_);
  and g_136354_(_046703_, _046708_, _046710_);
  or g_136355_(_046704_, _046709_, _046711_);
  xor g_136356_(out[727], _046641_, _046712_);
  xor g_136357_(_000373_, _046641_, _046713_);
  and g_136358_(_046567_, _046713_, _046714_);
  or g_136359_(_046568_, _046712_, _046715_);
  xor g_136360_(out[726], _046640_, _046717_);
  xor g_136361_(_000384_, _046640_, _046718_);
  and g_136362_(_046367_, _046561_, _046719_);
  or g_136363_(_046366_, _046560_, _046720_);
  and g_136364_(_046359_, _046560_, _046721_);
  or g_136365_(_046360_, _046561_, _046722_);
  and g_136366_(_046720_, _046722_, _046723_);
  or g_136367_(_046719_, _046721_, _046724_);
  and g_136368_(_046717_, _046723_, _046725_);
  or g_136369_(_046718_, _046724_, _046726_);
  and g_136370_(_046715_, _046726_, _046728_);
  or g_136371_(_046714_, _046725_, _046729_);
  xor g_136372_(out[725], _046638_, _046730_);
  xor g_136373_(_000395_, _046638_, _046731_);
  and g_136374_(_046371_, _046560_, _046732_);
  or g_136375_(_046370_, _046561_, _046733_);
  and g_136376_(_046378_, _046561_, _046734_);
  or g_136377_(_046377_, _046560_, _046735_);
  and g_136378_(_046733_, _046735_, _046736_);
  or g_136379_(_046732_, _046734_, _046737_);
  and g_136380_(_046730_, _046737_, _046739_);
  or g_136381_(_046731_, _046736_, _046740_);
  xor g_136382_(out[724], _046571_, _046741_);
  xor g_136383_(_000406_, _046571_, _046742_);
  and g_136384_(_046382_, _046560_, _046743_);
  or g_136385_(_046381_, _046561_, _046744_);
  and g_136386_(_046389_, _046561_, _046745_);
  or g_136387_(_046388_, _046560_, _046746_);
  and g_136388_(_046744_, _046746_, _046747_);
  or g_136389_(_046743_, _046745_, _046748_);
  and g_136390_(_046741_, _046748_, _046750_);
  or g_136391_(_046742_, _046747_, _046751_);
  and g_136392_(_046740_, _046751_, _046752_);
  or g_136393_(_046739_, _046750_, _046753_);
  and g_136394_(_046731_, _046736_, _046754_);
  or g_136395_(_046730_, _046737_, _046755_);
  and g_136396_(_046742_, _046747_, _046756_);
  or g_136397_(_046741_, _046748_, _046757_);
  and g_136398_(_046755_, _046757_, _046758_);
  or g_136399_(_046754_, _046756_, _046759_);
  and g_136400_(_046718_, _046724_, _046761_);
  or g_136401_(_046717_, _046723_, _046762_);
  and g_136402_(_046568_, _046712_, _046763_);
  or g_136403_(_046567_, _046713_, _046764_);
  and g_136404_(_046762_, _046764_, _046765_);
  or g_136405_(_046761_, _046763_, _046766_);
  and g_136406_(_046728_, _046765_, _046767_);
  or g_136407_(_046729_, _046766_, _046768_);
  and g_136408_(_046752_, _046758_, _046769_);
  or g_136409_(_046753_, _046759_, _046770_);
  and g_136410_(_046767_, _046769_, _046772_);
  or g_136411_(_046768_, _046770_, _046773_);
  and g_136412_(_046710_, _046772_, _046774_);
  or g_136413_(_046711_, _046773_, _046775_);
  and g_136414_(_046637_, _046774_, _046776_);
  or g_136415_(_046636_, _046775_, _046777_);
  and g_136416_(_046655_, _046676_, _046778_);
  or g_136417_(_046654_, _046675_, _046779_);
  and g_136418_(_046693_, _046778_, _046780_);
  or g_136419_(_046692_, _046779_, _046781_);
  and g_136420_(_046699_, _046781_, _046783_);
  or g_136421_(_046700_, _046780_, _046784_);
  and g_136422_(_046665_, _046784_, _046785_);
  or g_136423_(_046664_, _046783_, _046786_);
  and g_136424_(_046729_, _046764_, _046787_);
  or g_136425_(_046728_, _046763_, _046788_);
  and g_136426_(_046740_, _046765_, _046789_);
  or g_136427_(_046739_, _046766_, _046790_);
  and g_136428_(_046759_, _046789_, _046791_);
  or g_136429_(_046758_, _046790_, _046792_);
  and g_136430_(_046788_, _046792_, _046794_);
  or g_136431_(_046787_, _046791_, _046795_);
  and g_136432_(_046710_, _046795_, _046796_);
  or g_136433_(_046711_, _046794_, _046797_);
  and g_136434_(_046786_, _046797_, _046798_);
  or g_136435_(_046785_, _046796_, _046799_);
  and g_136436_(_046777_, _046798_, _046800_);
  or g_136437_(_046776_, _046799_, _046801_);
  and g_136438_(out[720], _046616_, _046802_);
  or g_136439_(_000428_, _046618_, _046803_);
  and g_136440_(_046623_, _046632_, _046805_);
  or g_136441_(_046624_, _046633_, _046806_);
  and g_136442_(_046774_, _046805_, _046807_);
  or g_136443_(_046775_, _046806_, _046808_);
  and g_136444_(_046803_, _046807_, _046809_);
  or g_136445_(_046802_, _046808_, _046810_);
  and g_136446_(_046801_, _046810_, _046811_);
  or g_136447_(_046800_, _046809_, _046812_);
  and g_136448_(_046568_, _046812_, _046813_);
  or g_136449_(_046567_, _046811_, _046814_);
  and g_136450_(_046713_, _046811_, _046816_);
  or g_136451_(_046712_, _046812_, _046817_);
  and g_136452_(_046814_, _046817_, _046818_);
  or g_136453_(_046813_, _046816_, _046819_);
  and g_136454_(_043417_, _046819_, _046820_);
  or g_136455_(_043418_, _046818_, _046821_);
  xor g_136456_(out[742], _043408_, _046822_);
  xor g_136457_(_000516_, _043408_, _046823_);
  and g_136458_(_046724_, _046812_, _046824_);
  or g_136459_(_046723_, _046811_, _046825_);
  and g_136460_(_046717_, _046811_, _046827_);
  or g_136461_(_046718_, _046812_, _046828_);
  and g_136462_(_046825_, _046828_, _046829_);
  or g_136463_(_046824_, _046827_, _046830_);
  and g_136464_(_046822_, _046829_, _046831_);
  or g_136465_(_046823_, _046830_, _046832_);
  xor g_136466_(out[737], out[736], _046833_);
  xor g_136467_(_000549_, out[736], _046834_);
  and g_136468_(_046609_, _046812_, _046835_);
  or g_136469_(_046608_, _046811_, _046836_);
  and g_136470_(_046601_, _046811_, _046838_);
  or g_136471_(_046602_, _046812_, _046839_);
  and g_136472_(_046836_, _046839_, _046840_);
  or g_136473_(_046835_, _046838_, _046841_);
  and g_136474_(_046833_, _046840_, _046842_);
  or g_136475_(_046834_, _046841_, _046843_);
  and g_136476_(out[720], _046811_, _046844_);
  or g_136477_(_000428_, _046812_, _046845_);
  and g_136478_(_046618_, _046812_, _046846_);
  or g_136479_(_046616_, _046811_, _046847_);
  and g_136480_(_046845_, _046847_, _046849_);
  or g_136481_(_046844_, _046846_, _046850_);
  and g_136482_(out[736], _046849_, _046851_);
  or g_136483_(_000560_, _046850_, _046852_);
  and g_136484_(_046843_, _046852_, _046853_);
  or g_136485_(_046842_, _046851_, _046854_);
  xor g_136486_(out[738], _043403_, _046855_);
  xor g_136487_(_000571_, _043403_, _046856_);
  and g_136488_(_046583_, _046811_, _046857_);
  or g_136489_(_046585_, _046812_, _046858_);
  and g_136490_(_046591_, _046812_, _046860_);
  or g_136491_(_046590_, _046811_, _046861_);
  and g_136492_(_046858_, _046861_, _046862_);
  or g_136493_(_046857_, _046860_, _046863_);
  and g_136494_(_046856_, _046863_, _046864_);
  or g_136495_(_046855_, _046862_, _046865_);
  and g_136496_(out[737], _046841_, _046866_);
  or g_136497_(_000549_, _046840_, _046867_);
  and g_136498_(_046865_, _046867_, _046868_);
  or g_136499_(_046864_, _046866_, _046869_);
  and g_136500_(_046854_, _046868_, _046871_);
  or g_136501_(_046853_, _046869_, _046872_);
  xor g_136502_(out[739], _043404_, _046873_);
  xor g_136503_(_000582_, _043404_, _046874_);
  and g_136504_(_046574_, _046811_, _046875_);
  or g_136505_(_046572_, _046812_, _046876_);
  and g_136506_(_046580_, _046812_, _046877_);
  or g_136507_(_046579_, _046811_, _046878_);
  and g_136508_(_046876_, _046878_, _046879_);
  or g_136509_(_046875_, _046877_, _046880_);
  and g_136510_(_046874_, _046879_, _046882_);
  or g_136511_(_046873_, _046880_, _046883_);
  and g_136512_(_046855_, _046862_, _046884_);
  or g_136513_(_046856_, _046863_, _046885_);
  and g_136514_(_046883_, _046885_, _046886_);
  or g_136515_(_046882_, _046884_, _046887_);
  and g_136516_(_046872_, _046886_, _046888_);
  or g_136517_(_046871_, _046887_, _046889_);
  xor g_136518_(out[740], _043406_, _046890_);
  xor g_136519_(_000538_, _043406_, _046891_);
  and g_136520_(_046742_, _046811_, _046893_);
  or g_136521_(_046741_, _046812_, _046894_);
  and g_136522_(_046748_, _046812_, _046895_);
  or g_136523_(_046747_, _046811_, _046896_);
  and g_136524_(_046894_, _046896_, _046897_);
  or g_136525_(_046893_, _046895_, _046898_);
  and g_136526_(_046890_, _046898_, _046899_);
  or g_136527_(_046891_, _046897_, _046900_);
  and g_136528_(_046873_, _046880_, _046901_);
  or g_136529_(_046874_, _046879_, _046902_);
  and g_136530_(_046900_, _046902_, _046904_);
  or g_136531_(_046899_, _046901_, _046905_);
  and g_136532_(_046889_, _046904_, _046906_);
  or g_136533_(_046888_, _046905_, _046907_);
  xor g_136534_(out[741], _043407_, _046908_);
  xor g_136535_(_000527_, _043407_, _046909_);
  and g_136536_(_046737_, _046812_, _046910_);
  or g_136537_(_046736_, _046811_, _046911_);
  and g_136538_(_046731_, _046811_, _046912_);
  or g_136539_(_046730_, _046812_, _046913_);
  and g_136540_(_046911_, _046913_, _046915_);
  or g_136541_(_046910_, _046912_, _046916_);
  and g_136542_(_046909_, _046915_, _046917_);
  or g_136543_(_046908_, _046916_, _046918_);
  and g_136544_(_046891_, _046897_, _046919_);
  or g_136545_(_046890_, _046898_, _046920_);
  and g_136546_(_046918_, _046920_, _046921_);
  or g_136547_(_046917_, _046919_, _046922_);
  and g_136548_(_046907_, _046921_, _046923_);
  or g_136549_(_046906_, _046922_, _046924_);
  and g_136550_(_046823_, _046830_, _046926_);
  or g_136551_(_046822_, _046829_, _046927_);
  and g_136552_(_046908_, _046916_, _046928_);
  or g_136553_(_046909_, _046915_, _046929_);
  and g_136554_(_046927_, _046929_, _046930_);
  or g_136555_(_046926_, _046928_, _046931_);
  and g_136556_(_046924_, _046930_, _046932_);
  or g_136557_(_046923_, _046931_, _046933_);
  and g_136558_(_046832_, _046933_, _046934_);
  or g_136559_(_046831_, _046932_, _046935_);
  and g_136560_(_046821_, _046935_, _046937_);
  or g_136561_(_046820_, _046934_, _046938_);
  and g_136562_(_046674_, _046812_, _046939_);
  or g_136563_(_046673_, _046811_, _046940_);
  and g_136564_(_046667_, _046811_, _046941_);
  or g_136565_(_046666_, _046812_, _046942_);
  and g_136566_(_046940_, _046942_, _046943_);
  or g_136567_(_046939_, _046941_, _046944_);
  and g_136568_(_043414_, _046944_, _046945_);
  or g_136569_(_043415_, _046943_, _046946_);
  xor g_136570_(out[747], _043413_, _046948_);
  xor g_136571_(_000494_, _043413_, _046949_);
  and g_136572_(_046658_, _046811_, _046950_);
  or g_136573_(_046657_, _046812_, _046951_);
  and g_136574_(_046660_, _046812_, _046952_);
  or g_136575_(_046659_, _046811_, _046953_);
  and g_136576_(_046951_, _046953_, _046954_);
  or g_136577_(_046950_, _046952_, _046955_);
  and g_136578_(_046662_, _046812_, _046956_);
  or g_136579_(_046663_, _046811_, _046957_);
  and g_136580_(_046657_, _046811_, _046959_);
  or g_136581_(_046658_, _046812_, _046960_);
  and g_136582_(_046957_, _046960_, _046961_);
  or g_136583_(_046956_, _046959_, _046962_);
  and g_136584_(_046948_, _046961_, _046963_);
  or g_136585_(_046949_, _046962_, _046964_);
  and g_136586_(_046946_, _046964_, _046965_);
  or g_136587_(_046945_, _046963_, _046966_);
  and g_136588_(_043415_, _046943_, _046967_);
  or g_136589_(_043414_, _046944_, _046968_);
  and g_136590_(_046949_, _046954_, _046970_);
  or g_136591_(_046948_, _046955_, _046971_);
  and g_136592_(_046968_, _046971_, _046972_);
  or g_136593_(_046967_, _046970_, _046973_);
  and g_136594_(_046965_, _046972_, _046974_);
  or g_136595_(_046966_, _046973_, _046975_);
  xor g_136596_(out[744], _043410_, _046976_);
  xor g_136597_(_000593_, _043410_, _046977_);
  and g_136598_(_046685_, _046812_, _046978_);
  or g_136599_(_046684_, _046811_, _046979_);
  and g_136600_(_046678_, _046811_, _046981_);
  or g_136601_(_046677_, _046812_, _046982_);
  and g_136602_(_046979_, _046982_, _046983_);
  or g_136603_(_046978_, _046981_, _046984_);
  and g_136604_(_046976_, _046984_, _046985_);
  or g_136605_(_046977_, _046983_, _046986_);
  and g_136606_(_046653_, _046812_, _046987_);
  or g_136607_(_046652_, _046811_, _046988_);
  and g_136608_(_046645_, _046811_, _046989_);
  or g_136609_(_046646_, _046812_, _046990_);
  and g_136610_(_046988_, _046990_, _046992_);
  or g_136611_(_046987_, _046989_, _046993_);
  xor g_136612_(out[745], _043411_, _046994_);
  xor g_136613_(_000604_, _043411_, _046995_);
  and g_136614_(_046993_, _046995_, _046996_);
  or g_136615_(_046992_, _046994_, _046997_);
  and g_136616_(_046986_, _046997_, _046998_);
  or g_136617_(_046985_, _046996_, _046999_);
  and g_136618_(_046992_, _046994_, _047000_);
  or g_136619_(_046993_, _046995_, _047001_);
  and g_136620_(_046977_, _046983_, _047003_);
  or g_136621_(_046976_, _046984_, _047004_);
  and g_136622_(_047001_, _047004_, _047005_);
  or g_136623_(_047000_, _047003_, _047006_);
  and g_136624_(_043418_, _046818_, _047007_);
  or g_136625_(_043417_, _046819_, _047008_);
  and g_136626_(_047005_, _047008_, _047009_);
  or g_136627_(_047006_, _047007_, _047010_);
  and g_136628_(_046998_, _047009_, _047011_);
  or g_136629_(_046999_, _047010_, _047012_);
  and g_136630_(_046974_, _047011_, _047014_);
  or g_136631_(_046975_, _047012_, _047015_);
  and g_136632_(_046938_, _047014_, _047016_);
  or g_136633_(_046937_, _047015_, _047017_);
  and g_136634_(_046999_, _047001_, _047018_);
  or g_136635_(_046998_, _047000_, _047019_);
  and g_136636_(_046974_, _047018_, _047020_);
  or g_136637_(_046975_, _047019_, _047021_);
  and g_136638_(_046945_, _046971_, _047022_);
  or g_136639_(_046946_, _046970_, _047023_);
  and g_136640_(_046964_, _047023_, _047025_);
  or g_136641_(_046963_, _047022_, _047026_);
  and g_136642_(_047021_, _047025_, _047027_);
  or g_136643_(_047020_, _047026_, _047028_);
  and g_136644_(_047017_, _047027_, _047029_);
  or g_136645_(_047016_, _047028_, _047030_);
  or g_136646_(_043414_, _047030_, _047031_);
  not g_136647_(_047031_, _047032_);
  and g_136648_(_046944_, _047030_, _047033_);
  not g_136649_(_047033_, _047034_);
  and g_136650_(_047031_, _047034_, _047036_);
  or g_136651_(_047032_, _047033_, _047037_);
  or g_136652_(out[753], out[752], _047038_);
  or g_136653_(out[752], _000650_, _047039_);
  and g_136654_(out[755], _047039_, _047040_);
  and g_136655_(_025001_, _047039_, _047041_);
  and g_136656_(out[757], _047041_, _047042_);
  or g_136657_(out[758], _047042_, _047043_);
  and g_136658_(out[759], _047043_, _047044_);
  xor g_136659_(out[759], _047043_, _047045_);
  xor g_136660_(_000637_, _047043_, _047047_);
  or g_136661_(_043417_, _047030_, _047048_);
  not g_136662_(_047048_, _047049_);
  and g_136663_(_046819_, _047030_, _047050_);
  not g_136664_(_047050_, _047051_);
  and g_136665_(_047048_, _047051_, _047052_);
  or g_136666_(_047049_, _047050_, _047053_);
  and g_136667_(_047045_, _047053_, _047054_);
  or g_136668_(_047047_, _047052_, _047055_);
  xor g_136669_(out[757], _047041_, _047056_);
  xor g_136670_(_000659_, _047041_, _047058_);
  and g_136671_(_046916_, _047030_, _047059_);
  not g_136672_(_047059_, _047060_);
  or g_136673_(_046908_, _047030_, _047061_);
  not g_136674_(_047061_, _047062_);
  and g_136675_(_047060_, _047061_, _047063_);
  or g_136676_(_047059_, _047062_, _047064_);
  and g_136677_(_047058_, _047063_, _047065_);
  or g_136678_(_047056_, _047064_, _047066_);
  xor g_136679_(out[756], _047040_, _047067_);
  xor g_136680_(_000670_, _047040_, _047069_);
  or g_136681_(_046890_, _047030_, _047070_);
  not g_136682_(_047070_, _047071_);
  and g_136683_(_046898_, _047030_, _047072_);
  not g_136684_(_047072_, _047073_);
  and g_136685_(_047070_, _047073_, _047074_);
  or g_136686_(_047071_, _047072_, _047075_);
  and g_136687_(_047067_, _047075_, _047076_);
  or g_136688_(_047069_, _047074_, _047077_);
  xor g_136689_(out[754], _047038_, _047078_);
  xor g_136690_(_000703_, _047038_, _047080_);
  and g_136691_(_046863_, _047030_, _047081_);
  not g_136692_(_047081_, _047082_);
  or g_136693_(_046856_, _047030_, _047083_);
  not g_136694_(_047083_, _047084_);
  and g_136695_(_047082_, _047083_, _047085_);
  or g_136696_(_047081_, _047084_, _047086_);
  and g_136697_(_047078_, _047085_, _047087_);
  or g_136698_(_047080_, _047086_, _047088_);
  and g_136699_(_046833_, _047029_, _047089_);
  or g_136700_(_046834_, _047030_, _047091_);
  and g_136701_(_046841_, _047030_, _047092_);
  or g_136702_(_046840_, _047029_, _047093_);
  and g_136703_(_047091_, _047093_, _047094_);
  or g_136704_(_047089_, _047092_, _047095_);
  and g_136705_(out[753], _047095_, _047096_);
  not g_136706_(_047096_, _047097_);
  xor g_136707_(out[753], out[752], _047098_);
  xor g_136708_(_000681_, out[752], _047099_);
  and g_136709_(_047094_, _047098_, _047100_);
  or g_136710_(_047095_, _047099_, _047102_);
  and g_136711_(out[736], _047029_, _047103_);
  or g_136712_(_000560_, _047030_, _047104_);
  and g_136713_(_046850_, _047030_, _047105_);
  or g_136714_(_046849_, _047029_, _047106_);
  and g_136715_(_047104_, _047106_, _047107_);
  or g_136716_(_047103_, _047105_, _047108_);
  and g_136717_(out[752], _047107_, _047109_);
  or g_136718_(_000692_, _047108_, _047110_);
  and g_136719_(_047102_, _047110_, _047111_);
  or g_136720_(_047100_, _047109_, _047113_);
  and g_136721_(_047097_, _047113_, _047114_);
  or g_136722_(_047096_, _047111_, _047115_);
  and g_136723_(_047088_, _047115_, _047116_);
  or g_136724_(_047087_, _047114_, _047117_);
  and g_136725_(_047080_, _047086_, _047118_);
  or g_136726_(_047078_, _047085_, _047119_);
  xor g_136727_(out[755], _047039_, _047120_);
  xor g_136728_(_000714_, _047039_, _047121_);
  or g_136729_(_046873_, _047030_, _047122_);
  not g_136730_(_047122_, _047124_);
  and g_136731_(_046880_, _047030_, _047125_);
  not g_136732_(_047125_, _047126_);
  and g_136733_(_047122_, _047126_, _047127_);
  or g_136734_(_047124_, _047125_, _047128_);
  and g_136735_(_047120_, _047128_, _047129_);
  or g_136736_(_047121_, _047127_, _047130_);
  and g_136737_(_047119_, _047130_, _047131_);
  or g_136738_(_047118_, _047129_, _047132_);
  and g_136739_(_047117_, _047131_, _047133_);
  or g_136740_(_047116_, _047132_, _047135_);
  and g_136741_(_047069_, _047074_, _047136_);
  or g_136742_(_047067_, _047075_, _047137_);
  and g_136743_(_047121_, _047127_, _047138_);
  or g_136744_(_047120_, _047128_, _047139_);
  and g_136745_(_047137_, _047139_, _047140_);
  or g_136746_(_047136_, _047138_, _047141_);
  and g_136747_(_047135_, _047140_, _047142_);
  or g_136748_(_047133_, _047141_, _047143_);
  and g_136749_(_047077_, _047143_, _047144_);
  or g_136750_(_047076_, _047142_, _047146_);
  and g_136751_(_047066_, _047146_, _047147_);
  or g_136752_(_047065_, _047144_, _047148_);
  xor g_136753_(out[758], _047042_, _047149_);
  xor g_136754_(_000648_, _047042_, _047150_);
  or g_136755_(_046823_, _047030_, _047151_);
  not g_136756_(_047151_, _047152_);
  and g_136757_(_046830_, _047030_, _047153_);
  not g_136758_(_047153_, _047154_);
  and g_136759_(_047151_, _047154_, _047155_);
  or g_136760_(_047152_, _047153_, _047157_);
  and g_136761_(_047150_, _047157_, _047158_);
  or g_136762_(_047149_, _047155_, _047159_);
  and g_136763_(_047056_, _047064_, _047160_);
  or g_136764_(_047058_, _047063_, _047161_);
  and g_136765_(_047159_, _047161_, _047162_);
  or g_136766_(_047158_, _047160_, _047163_);
  and g_136767_(_047148_, _047162_, _047164_);
  or g_136768_(_047147_, _047163_, _047165_);
  and g_136769_(_047047_, _047052_, _047166_);
  or g_136770_(_047045_, _047053_, _047168_);
  and g_136771_(_047149_, _047155_, _047169_);
  or g_136772_(_047150_, _047157_, _047170_);
  and g_136773_(_047168_, _047170_, _047171_);
  or g_136774_(_047166_, _047169_, _047172_);
  and g_136775_(_047165_, _047171_, _047173_);
  or g_136776_(_047164_, _047172_, _047174_);
  and g_136777_(_047055_, _047174_, _047175_);
  or g_136778_(_047054_, _047173_, _047176_);
  and g_136779_(out[760], _047044_, _047177_);
  or g_136780_(out[761], _047177_, _047179_);
  and g_136781_(out[762], _047179_, _047180_);
  xor g_136782_(out[762], _047179_, _047181_);
  xor g_136783_(_000747_, _047179_, _047182_);
  and g_136784_(_047037_, _047181_, _047183_);
  or g_136785_(_047036_, _047182_, _047184_);
  xor g_136786_(out[763], _047180_, _047185_);
  xor g_136787_(_000626_, _047180_, _047186_);
  and g_136788_(_046948_, _046954_, _047187_);
  or g_136789_(_046949_, _046955_, _047188_);
  and g_136790_(_046948_, _046962_, _047190_);
  or g_136791_(_046949_, _046961_, _047191_);
  and g_136792_(_047185_, _047191_, _047192_);
  or g_136793_(_047186_, _047190_, _047193_);
  and g_136794_(_047184_, _047193_, _047194_);
  or g_136795_(_047183_, _047192_, _047195_);
  xor g_136796_(out[761], _047177_, _047196_);
  xor g_136797_(_000736_, _047177_, _047197_);
  or g_136798_(_046995_, _047030_, _047198_);
  not g_136799_(_047198_, _047199_);
  and g_136800_(_046993_, _047030_, _047201_);
  not g_136801_(_047201_, _047202_);
  and g_136802_(_047198_, _047202_, _047203_);
  or g_136803_(_047199_, _047201_, _047204_);
  and g_136804_(_047196_, _047203_, _047205_);
  or g_136805_(_047197_, _047204_, _047206_);
  and g_136806_(_047036_, _047182_, _047207_);
  or g_136807_(_047037_, _047181_, _047208_);
  and g_136808_(_047186_, _047187_, _047209_);
  or g_136809_(_047185_, _047188_, _047210_);
  and g_136810_(_047208_, _047210_, _047212_);
  or g_136811_(_047207_, _047209_, _047213_);
  and g_136812_(_047194_, _047212_, _047214_);
  or g_136813_(_047195_, _047213_, _047215_);
  and g_136814_(_047206_, _047214_, _047216_);
  or g_136815_(_047205_, _047215_, _047217_);
  xor g_136816_(out[760], _047044_, _047218_);
  xor g_136817_(_000725_, _047044_, _047219_);
  or g_136818_(_046976_, _047030_, _047220_);
  not g_136819_(_047220_, _047221_);
  and g_136820_(_046984_, _047030_, _047223_);
  not g_136821_(_047223_, _047224_);
  and g_136822_(_047220_, _047224_, _047225_);
  or g_136823_(_047221_, _047223_, _047226_);
  and g_136824_(_047218_, _047226_, _047227_);
  or g_136825_(_047219_, _047225_, _047228_);
  and g_136826_(_047197_, _047204_, _047229_);
  or g_136827_(_047196_, _047203_, _047230_);
  and g_136828_(_047228_, _047230_, _047231_);
  or g_136829_(_047227_, _047229_, _047232_);
  and g_136830_(_047219_, _047225_, _047234_);
  or g_136831_(_047218_, _047226_, _047235_);
  and g_136832_(_047231_, _047235_, _047236_);
  or g_136833_(_047232_, _047234_, _047237_);
  and g_136834_(_047216_, _047236_, _047238_);
  or g_136835_(_047217_, _047237_, _047239_);
  and g_136836_(_047176_, _047238_, _047240_);
  or g_136837_(_047175_, _047239_, _047241_);
  and g_136838_(_047216_, _047232_, _047242_);
  or g_136839_(_047217_, _047231_, _047243_);
  and g_136840_(_047195_, _047210_, _047245_);
  or g_136841_(_047194_, _047209_, _047246_);
  and g_136842_(_047243_, _047246_, _047247_);
  or g_136843_(_047242_, _047245_, _047248_);
  and g_136844_(_047241_, _047247_, _047249_);
  or g_136845_(_047240_, _047248_, _047250_);
  and g_136846_(_047037_, _047250_, _047251_);
  not g_136847_(_047251_, _047252_);
  or g_136848_(_047181_, _047250_, _047253_);
  not g_136849_(_047253_, _047254_);
  and g_136850_(_047252_, _047253_, _047256_);
  or g_136851_(_047251_, _047254_, _047257_);
  or g_136852_(out[769], out[768], _047258_);
  or g_136853_(out[768], _000827_, _047259_);
  and g_136854_(out[771], _047259_, _047260_);
  and g_136855_(_025187_, _047259_, _047261_);
  and g_136856_(out[773], _047261_, _047262_);
  or g_136857_(out[774], _047262_, _047263_);
  and g_136858_(out[775], _047263_, _047264_);
  xor g_136859_(out[775], _047263_, _047265_);
  xor g_136860_(_000769_, _047263_, _047267_);
  and g_136861_(_047053_, _047250_, _047268_);
  not g_136862_(_047268_, _047269_);
  or g_136863_(_047045_, _047250_, _047270_);
  not g_136864_(_047270_, _047271_);
  and g_136865_(_047269_, _047270_, _047272_);
  or g_136866_(_047268_, _047271_, _047273_);
  and g_136867_(_047265_, _047273_, _047274_);
  or g_136868_(_047267_, _047272_, _047275_);
  xor g_136869_(out[774], _047262_, _047276_);
  xor g_136870_(_000780_, _047262_, _047278_);
  and g_136871_(_047157_, _047250_, _047279_);
  not g_136872_(_047279_, _047280_);
  or g_136873_(_047150_, _047250_, _047281_);
  not g_136874_(_047281_, _047282_);
  and g_136875_(_047280_, _047281_, _047283_);
  or g_136876_(_047279_, _047282_, _047284_);
  and g_136877_(_047278_, _047284_, _047285_);
  or g_136878_(_047276_, _047283_, _047286_);
  xor g_136879_(out[773], _047261_, _047287_);
  xor g_136880_(_000791_, _047261_, _047289_);
  or g_136881_(_047056_, _047250_, _047290_);
  not g_136882_(_047290_, _047291_);
  and g_136883_(_047064_, _047250_, _047292_);
  not g_136884_(_047292_, _047293_);
  and g_136885_(_047290_, _047293_, _047294_);
  or g_136886_(_047291_, _047292_, _047295_);
  and g_136887_(_047289_, _047294_, _047296_);
  or g_136888_(_047287_, _047295_, _047297_);
  xor g_136889_(out[770], _047258_, _047298_);
  xor g_136890_(_000835_, _047258_, _047300_);
  and g_136891_(_047086_, _047250_, _047301_);
  not g_136892_(_047301_, _047302_);
  or g_136893_(_047080_, _047250_, _047303_);
  not g_136894_(_047303_, _047304_);
  and g_136895_(_047302_, _047303_, _047305_);
  or g_136896_(_047301_, _047304_, _047306_);
  and g_136897_(_047298_, _047305_, _047307_);
  or g_136898_(_047300_, _047306_, _047308_);
  and g_136899_(_047098_, _047249_, _047309_);
  or g_136900_(_047099_, _047250_, _047311_);
  and g_136901_(_047095_, _047250_, _047312_);
  or g_136902_(_047094_, _047249_, _047313_);
  and g_136903_(_047311_, _047313_, _047314_);
  or g_136904_(_047309_, _047312_, _047315_);
  and g_136905_(out[769], _047315_, _047316_);
  not g_136906_(_047316_, _047317_);
  xor g_136907_(_000813_, out[768], _047318_);
  not g_136908_(_047318_, _047319_);
  and g_136909_(_047314_, _047319_, _047320_);
  or g_136910_(_047315_, _047318_, _047322_);
  and g_136911_(out[752], _047249_, _047323_);
  or g_136912_(_000692_, _047250_, _047324_);
  and g_136913_(_047108_, _047250_, _047325_);
  or g_136914_(_047107_, _047249_, _047326_);
  and g_136915_(_047324_, _047326_, _047327_);
  or g_136916_(_047323_, _047325_, _047328_);
  and g_136917_(out[768], _047327_, _047329_);
  or g_136918_(_000824_, _047328_, _047330_);
  and g_136919_(_047322_, _047330_, _047331_);
  or g_136920_(_047320_, _047329_, _047333_);
  and g_136921_(_047317_, _047333_, _047334_);
  or g_136922_(_047316_, _047331_, _047335_);
  and g_136923_(_047308_, _047335_, _047336_);
  or g_136924_(_047307_, _047334_, _047337_);
  and g_136925_(_047300_, _047306_, _047338_);
  or g_136926_(_047298_, _047305_, _047339_);
  xor g_136927_(out[771], _047259_, _047340_);
  xor g_136928_(_000846_, _047259_, _047341_);
  or g_136929_(_047120_, _047250_, _047342_);
  not g_136930_(_047342_, _047344_);
  and g_136931_(_047128_, _047250_, _047345_);
  not g_136932_(_047345_, _047346_);
  and g_136933_(_047342_, _047346_, _047347_);
  or g_136934_(_047344_, _047345_, _047348_);
  and g_136935_(_047340_, _047348_, _047349_);
  or g_136936_(_047341_, _047347_, _047350_);
  and g_136937_(_047339_, _047350_, _047351_);
  or g_136938_(_047338_, _047349_, _047352_);
  and g_136939_(_047337_, _047351_, _047353_);
  or g_136940_(_047336_, _047352_, _047355_);
  xor g_136941_(out[772], _047260_, _047356_);
  xor g_136942_(_000802_, _047260_, _047357_);
  and g_136943_(_047075_, _047250_, _047358_);
  not g_136944_(_047358_, _047359_);
  or g_136945_(_047067_, _047250_, _047360_);
  not g_136946_(_047360_, _047361_);
  and g_136947_(_047359_, _047360_, _047362_);
  or g_136948_(_047358_, _047361_, _047363_);
  and g_136949_(_047357_, _047362_, _047364_);
  or g_136950_(_047356_, _047363_, _047366_);
  and g_136951_(_047341_, _047347_, _047367_);
  or g_136952_(_047340_, _047348_, _047368_);
  and g_136953_(_047366_, _047368_, _047369_);
  or g_136954_(_047364_, _047367_, _047370_);
  and g_136955_(_047355_, _047369_, _047371_);
  or g_136956_(_047353_, _047370_, _047372_);
  and g_136957_(_047287_, _047295_, _047373_);
  or g_136958_(_047289_, _047294_, _047374_);
  and g_136959_(_047356_, _047363_, _047375_);
  or g_136960_(_047357_, _047362_, _047377_);
  and g_136961_(_047374_, _047377_, _047378_);
  or g_136962_(_047373_, _047375_, _047379_);
  and g_136963_(_047372_, _047378_, _047380_);
  or g_136964_(_047371_, _047379_, _047381_);
  and g_136965_(_047297_, _047381_, _047382_);
  or g_136966_(_047296_, _047380_, _047383_);
  and g_136967_(_047286_, _047383_, _047384_);
  or g_136968_(_047285_, _047382_, _047385_);
  and g_136969_(_047267_, _047272_, _047386_);
  or g_136970_(_047265_, _047273_, _047388_);
  and g_136971_(_047276_, _047283_, _047389_);
  or g_136972_(_047278_, _047284_, _047390_);
  and g_136973_(_047388_, _047390_, _047391_);
  or g_136974_(_047386_, _047389_, _047392_);
  and g_136975_(_047385_, _047391_, _047393_);
  or g_136976_(_047384_, _047392_, _047394_);
  and g_136977_(_047275_, _047394_, _047395_);
  or g_136978_(_047274_, _047393_, _047396_);
  and g_136979_(out[776], _047264_, _047397_);
  or g_136980_(out[777], _047397_, _047399_);
  and g_136981_(out[778], _047399_, _047400_);
  xor g_136982_(out[778], _047399_, _047401_);
  xor g_136983_(_000879_, _047399_, _047402_);
  and g_136984_(_047257_, _047401_, _047403_);
  or g_136985_(_047256_, _047402_, _047404_);
  xor g_136986_(out[779], _047400_, _047405_);
  xor g_136987_(_000758_, _047400_, _047406_);
  and g_136988_(_047185_, _047187_, _047407_);
  or g_136989_(_047186_, _047188_, _047408_);
  and g_136990_(_047185_, _047190_, _047410_);
  or g_136991_(_047186_, _047191_, _047411_);
  and g_136992_(_047405_, _047411_, _047412_);
  or g_136993_(_047406_, _047410_, _047413_);
  and g_136994_(_047404_, _047413_, _047414_);
  or g_136995_(_047403_, _047412_, _047415_);
  and g_136996_(_047256_, _047402_, _047416_);
  or g_136997_(_047257_, _047401_, _047417_);
  and g_136998_(_047406_, _047407_, _047418_);
  or g_136999_(_047405_, _047408_, _047419_);
  and g_137000_(_047417_, _047419_, _047421_);
  or g_137001_(_047416_, _047418_, _047422_);
  and g_137002_(_047414_, _047421_, _047423_);
  or g_137003_(_047415_, _047422_, _047424_);
  xor g_137004_(out[776], _047264_, _047425_);
  xor g_137005_(_000857_, _047264_, _047426_);
  and g_137006_(_047226_, _047250_, _047427_);
  not g_137007_(_047427_, _047428_);
  or g_137008_(_047218_, _047250_, _047429_);
  not g_137009_(_047429_, _047430_);
  and g_137010_(_047428_, _047429_, _047432_);
  or g_137011_(_047427_, _047430_, _047433_);
  and g_137012_(_047426_, _047432_, _047434_);
  or g_137013_(_047425_, _047433_, _047435_);
  xor g_137014_(out[777], _047397_, _047436_);
  xor g_137015_(_000868_, _047397_, _047437_);
  and g_137016_(_047204_, _047250_, _047438_);
  not g_137017_(_047438_, _047439_);
  or g_137018_(_047197_, _047250_, _047440_);
  not g_137019_(_047440_, _047441_);
  and g_137020_(_047439_, _047440_, _047443_);
  or g_137021_(_047438_, _047441_, _047444_);
  and g_137022_(_047436_, _047443_, _047445_);
  or g_137023_(_047437_, _047444_, _047446_);
  and g_137024_(_047435_, _047446_, _047447_);
  or g_137025_(_047434_, _047445_, _047448_);
  and g_137026_(_047437_, _047444_, _047449_);
  or g_137027_(_047436_, _047443_, _047450_);
  and g_137028_(_047425_, _047433_, _047451_);
  or g_137029_(_047426_, _047432_, _047452_);
  and g_137030_(_047450_, _047452_, _047454_);
  or g_137031_(_047449_, _047451_, _047455_);
  and g_137032_(_047447_, _047454_, _047456_);
  or g_137033_(_047448_, _047455_, _047457_);
  and g_137034_(_047423_, _047456_, _047458_);
  or g_137035_(_047424_, _047457_, _047459_);
  and g_137036_(_047396_, _047458_, _047460_);
  or g_137037_(_047395_, _047459_, _047461_);
  and g_137038_(_047415_, _047419_, _047462_);
  or g_137039_(_047414_, _047418_, _047463_);
  and g_137040_(_047446_, _047455_, _047465_);
  or g_137041_(_047445_, _047454_, _047466_);
  and g_137042_(_047423_, _047465_, _047467_);
  or g_137043_(_047424_, _047466_, _047468_);
  and g_137044_(_047463_, _047468_, _047469_);
  or g_137045_(_047462_, _047467_, _047470_);
  and g_137046_(_047461_, _047469_, _047471_);
  or g_137047_(_047460_, _047470_, _047472_);
  and g_137048_(_047257_, _047472_, _047473_);
  not g_137049_(_047473_, _047474_);
  or g_137050_(_047401_, _047472_, _047476_);
  not g_137051_(_047476_, _047477_);
  and g_137052_(_047474_, _047476_, _047478_);
  or g_137053_(_047473_, _047477_, _047479_);
  or g_137054_(_043402_, _047479_, _047480_);
  xor g_137055_(out[795], _043401_, _047481_);
  xor g_137056_(_000890_, _043401_, _047482_);
  and g_137057_(_047405_, _047407_, _047483_);
  or g_137058_(_047406_, _047408_, _047484_);
  or g_137059_(_047481_, _047484_, _047485_);
  and g_137060_(_047480_, _047485_, _047487_);
  and g_137061_(_047405_, _047410_, _047488_);
  or g_137062_(_047406_, _047411_, _047489_);
  and g_137063_(_047481_, _047484_, _047490_);
  xor g_137064_(out[793], _043399_, _047491_);
  xor g_137065_(_001000_, _043399_, _047492_);
  and g_137066_(_047444_, _047472_, _047493_);
  not g_137067_(_047493_, _047494_);
  and g_137068_(_047436_, _047471_, _047495_);
  or g_137069_(_047437_, _047472_, _047496_);
  and g_137070_(_047494_, _047496_, _047498_);
  or g_137071_(_047493_, _047495_, _047499_);
  and g_137072_(_047492_, _047499_, _047500_);
  or g_137073_(_047491_, _047498_, _047501_);
  xor g_137074_(_047482_, _047488_, _047502_);
  xor g_137075_(_047481_, _047488_, _047503_);
  xor g_137076_(_043402_, _047479_, _047504_);
  xor g_137077_(_043402_, _047478_, _047505_);
  and g_137078_(_047502_, _047504_, _047506_);
  or g_137079_(_047503_, _047505_, _047507_);
  and g_137080_(_047501_, _047506_, _047509_);
  or g_137081_(_047500_, _047507_, _047510_);
  and g_137082_(_047491_, _047498_, _047511_);
  or g_137083_(_047492_, _047499_, _047512_);
  xor g_137084_(out[792], _043398_, _047513_);
  xor g_137085_(_000989_, _043398_, _047514_);
  and g_137086_(_047433_, _047472_, _047515_);
  not g_137087_(_047515_, _047516_);
  or g_137088_(_047425_, _047472_, _047517_);
  not g_137089_(_047517_, _047518_);
  and g_137090_(_047516_, _047517_, _047520_);
  or g_137091_(_047515_, _047518_, _047521_);
  and g_137092_(_047514_, _047520_, _047522_);
  or g_137093_(_047513_, _047521_, _047523_);
  and g_137094_(_047512_, _047523_, _047524_);
  or g_137095_(_047511_, _047522_, _047525_);
  and g_137096_(_047513_, _047521_, _047526_);
  or g_137097_(_047514_, _047520_, _047527_);
  and g_137098_(_047524_, _047527_, _047528_);
  or g_137099_(_047525_, _047526_, _047529_);
  and g_137100_(_047509_, _047528_, _047531_);
  or g_137101_(_047510_, _047529_, _047532_);
  xor g_137102_(out[790], _043396_, _047533_);
  xor g_137103_(_000912_, _043396_, _047534_);
  and g_137104_(_047284_, _047472_, _047535_);
  or g_137105_(_047283_, _047471_, _047536_);
  and g_137106_(_047276_, _047471_, _047537_);
  or g_137107_(_047278_, _047472_, _047538_);
  and g_137108_(_047536_, _047538_, _047539_);
  or g_137109_(_047535_, _047537_, _047540_);
  and g_137110_(_047533_, _047539_, _047542_);
  or g_137111_(_047534_, _047540_, _047543_);
  xor g_137112_(out[791], _043397_, _047544_);
  xor g_137113_(_000901_, _043397_, _047545_);
  and g_137114_(_047273_, _047472_, _047546_);
  or g_137115_(_047272_, _047471_, _047547_);
  and g_137116_(_047267_, _047471_, _047548_);
  or g_137117_(_047265_, _047472_, _047549_);
  and g_137118_(_047547_, _047549_, _047550_);
  or g_137119_(_047546_, _047548_, _047551_);
  and g_137120_(_047545_, _047550_, _047553_);
  or g_137121_(_047544_, _047551_, _047554_);
  and g_137122_(_047543_, _047554_, _047555_);
  or g_137123_(_047542_, _047553_, _047556_);
  and g_137124_(_047544_, _047551_, _047557_);
  or g_137125_(_047545_, _047550_, _047558_);
  and g_137126_(_047534_, _047540_, _047559_);
  or g_137127_(_047533_, _047539_, _047560_);
  and g_137128_(_047558_, _047560_, _047561_);
  or g_137129_(_047557_, _047559_, _047562_);
  xor g_137130_(out[789], _043392_, _047564_);
  xor g_137131_(_000923_, _043392_, _047565_);
  or g_137132_(_047287_, _047472_, _047566_);
  not g_137133_(_047566_, _047567_);
  and g_137134_(_047295_, _047472_, _047568_);
  not g_137135_(_047568_, _047569_);
  and g_137136_(_047566_, _047569_, _047570_);
  or g_137137_(_047567_, _047568_, _047571_);
  and g_137138_(_047564_, _047571_, _047572_);
  or g_137139_(_047565_, _047570_, _047573_);
  and g_137140_(_047555_, _047561_, _047575_);
  or g_137141_(_047556_, _047562_, _047576_);
  and g_137142_(_047573_, _047575_, _047577_);
  or g_137143_(_047572_, _047576_, _047578_);
  and g_137144_(_047565_, _047570_, _047579_);
  or g_137145_(_047564_, _047571_, _047580_);
  or g_137146_(_047356_, _047472_, _047581_);
  not g_137147_(_047581_, _047582_);
  and g_137148_(_047363_, _047472_, _047583_);
  not g_137149_(_047583_, _047584_);
  and g_137150_(_047581_, _047584_, _047586_);
  or g_137151_(_047582_, _047583_, _047587_);
  and g_137152_(_043395_, _047586_, _047588_);
  or g_137153_(_043393_, _047587_, _047589_);
  and g_137154_(_047580_, _047589_, _047590_);
  or g_137155_(_047579_, _047588_, _047591_);
  and g_137156_(_043393_, _047587_, _047592_);
  or g_137157_(_043395_, _047586_, _047593_);
  and g_137158_(_047590_, _047593_, _047594_);
  or g_137159_(_047591_, _047592_, _047595_);
  and g_137160_(_047577_, _047594_, _047597_);
  or g_137161_(_047578_, _047595_, _047598_);
  xor g_137162_(out[787], _043390_, _047599_);
  xor g_137163_(_000978_, _043390_, _047600_);
  or g_137164_(_047340_, _047472_, _047601_);
  not g_137165_(_047601_, _047602_);
  and g_137166_(_047348_, _047472_, _047603_);
  not g_137167_(_047603_, _047604_);
  and g_137168_(_047601_, _047604_, _047605_);
  or g_137169_(_047602_, _047603_, _047606_);
  and g_137170_(_047599_, _047606_, _047608_);
  or g_137171_(_047600_, _047605_, _047609_);
  and g_137172_(_047600_, _047605_, _047610_);
  or g_137173_(_047599_, _047606_, _047611_);
  xor g_137174_(out[786], _043389_, _047612_);
  xor g_137175_(_000967_, _043389_, _047613_);
  and g_137176_(_047298_, _047471_, _047614_);
  or g_137177_(_047300_, _047472_, _047615_);
  and g_137178_(_047306_, _047472_, _047616_);
  not g_137179_(_047616_, _047617_);
  and g_137180_(_047615_, _047617_, _047619_);
  or g_137181_(_047614_, _047616_, _047620_);
  and g_137182_(_047612_, _047619_, _047621_);
  or g_137183_(_047613_, _047620_, _047622_);
  and g_137184_(_047611_, _047622_, _047623_);
  or g_137185_(_047610_, _047621_, _047624_);
  and g_137186_(_047609_, _047624_, _047625_);
  or g_137187_(_047608_, _047623_, _047626_);
  xor g_137188_(out[785], out[784], _047627_);
  not g_137189_(_047627_, _047628_);
  or g_137190_(_047318_, _047472_, _047630_);
  or g_137191_(_047314_, _047471_, _047631_);
  and g_137192_(_047630_, _047631_, _047632_);
  not g_137193_(_047632_, _047633_);
  and g_137194_(_047627_, _047632_, _047634_);
  not g_137195_(_047634_, _047635_);
  and g_137196_(out[768], _047471_, _047636_);
  or g_137197_(_000824_, _047472_, _047637_);
  and g_137198_(_047328_, _047472_, _047638_);
  or g_137199_(_047327_, _047471_, _047639_);
  and g_137200_(_047637_, _047639_, _047641_);
  or g_137201_(_047636_, _047638_, _047642_);
  and g_137202_(_000956_, _047642_, _047643_);
  or g_137203_(out[784], _047641_, _047644_);
  xor g_137204_(_047627_, _047632_, _047645_);
  xor g_137205_(_047628_, _047632_, _047646_);
  and g_137206_(_047644_, _047645_, _047647_);
  or g_137207_(_047643_, _047646_, _047648_);
  and g_137208_(_047635_, _047648_, _047649_);
  or g_137209_(_047634_, _047647_, _047650_);
  and g_137210_(_047613_, _047620_, _047652_);
  or g_137211_(_047612_, _047619_, _047653_);
  and g_137212_(_047609_, _047653_, _047654_);
  or g_137213_(_047608_, _047652_, _047655_);
  and g_137214_(_047650_, _047654_, _047656_);
  or g_137215_(_047649_, _047655_, _047657_);
  and g_137216_(_047626_, _047657_, _047658_);
  or g_137217_(_047625_, _047656_, _047659_);
  and g_137218_(_047597_, _047659_, _047660_);
  or g_137219_(_047598_, _047658_, _047661_);
  and g_137220_(_047577_, _047591_, _047663_);
  or g_137221_(_047578_, _047590_, _047664_);
  and g_137222_(_047556_, _047558_, _047665_);
  or g_137223_(_047555_, _047557_, _047666_);
  and g_137224_(_047664_, _047666_, _047667_);
  or g_137225_(_047663_, _047665_, _047668_);
  and g_137226_(_047661_, _047667_, _047669_);
  or g_137227_(_047660_, _047668_, _047670_);
  and g_137228_(_047531_, _047670_, _047671_);
  or g_137229_(_047532_, _047669_, _047672_);
  and g_137230_(_047509_, _047525_, _047674_);
  or g_137231_(_047510_, _047524_, _047675_);
  or g_137232_(_047487_, _047490_, _047676_);
  not g_137233_(_047676_, _047677_);
  and g_137234_(_047675_, _047676_, _047678_);
  or g_137235_(_047674_, _047677_, _047679_);
  and g_137236_(_047672_, _047678_, _047680_);
  or g_137237_(_047671_, _047679_, _047681_);
  and g_137238_(out[784], _047641_, _047682_);
  or g_137239_(_000956_, _047642_, _047683_);
  and g_137240_(_047623_, _047654_, _047685_);
  or g_137241_(_047624_, _047655_, _047686_);
  and g_137242_(_047683_, _047685_, _047687_);
  or g_137243_(_047682_, _047686_, _047688_);
  and g_137244_(_047647_, _047687_, _047689_);
  or g_137245_(_047648_, _047688_, _047690_);
  and g_137246_(_047531_, _047689_, _047691_);
  or g_137247_(_047532_, _047690_, _047692_);
  and g_137248_(_047597_, _047691_, _047693_);
  or g_137249_(_047598_, _047692_, _047694_);
  and g_137250_(_047681_, _047694_, _047696_);
  or g_137251_(_047680_, _047693_, _047697_);
  and g_137252_(_043395_, _047696_, _047698_);
  or g_137253_(_043393_, _047697_, _047699_);
  and g_137254_(_047587_, _047697_, _047700_);
  or g_137255_(_047586_, _047696_, _047701_);
  and g_137256_(_047699_, _047701_, _047702_);
  or g_137257_(_047698_, _047700_, _047703_);
  or g_137258_(out[801], out[800], _047704_);
  or g_137259_(out[800], _001210_, _047705_);
  and g_137260_(out[803], _047705_, _047707_);
  and g_137261_(_025554_, _047705_, _047708_);
  and g_137262_(out[805], _047708_, _047709_);
  or g_137263_(out[806], _047709_, _047710_);
  and g_137264_(out[807], _047710_, _047711_);
  and g_137265_(out[808], _047711_, _047712_);
  or g_137266_(out[809], _047712_, _047713_);
  and g_137267_(out[810], _047713_, _047714_);
  xor g_137268_(out[810], _047713_, _047715_);
  or g_137269_(_043402_, _047697_, _047716_);
  not g_137270_(_047716_, _047718_);
  and g_137271_(_047479_, _047697_, _047719_);
  or g_137272_(_047478_, _047696_, _047720_);
  and g_137273_(_047716_, _047720_, _047721_);
  or g_137274_(_047718_, _047719_, _047722_);
  and g_137275_(_047715_, _047722_, _047723_);
  xor g_137276_(out[811], _047714_, _047724_);
  xor g_137277_(_001022_, _047714_, _047725_);
  and g_137278_(_047482_, _047696_, _047726_);
  or g_137279_(_047481_, _047697_, _047727_);
  and g_137280_(_047484_, _047697_, _047729_);
  or g_137281_(_047483_, _047696_, _047730_);
  and g_137282_(_047727_, _047730_, _047731_);
  or g_137283_(_047726_, _047729_, _047732_);
  and g_137284_(_047488_, _047697_, _047733_);
  or g_137285_(_047489_, _047696_, _047734_);
  and g_137286_(_047481_, _047696_, _047735_);
  or g_137287_(_047482_, _047697_, _047736_);
  and g_137288_(_047734_, _047736_, _047737_);
  or g_137289_(_047733_, _047735_, _047738_);
  and g_137290_(_047724_, _047732_, _047740_);
  or g_137291_(_047723_, _047740_, _047741_);
  or g_137292_(_047724_, _047732_, _047742_);
  and g_137293_(_047741_, _047742_, _047743_);
  not g_137294_(_047743_, _047744_);
  xor g_137295_(out[809], _047712_, _047745_);
  xor g_137296_(_001132_, _047712_, _047746_);
  and g_137297_(_047491_, _047696_, _047747_);
  or g_137298_(_047492_, _047697_, _047748_);
  and g_137299_(_047499_, _047697_, _047749_);
  or g_137300_(_047498_, _047696_, _047751_);
  and g_137301_(_047748_, _047751_, _047752_);
  or g_137302_(_047747_, _047749_, _047753_);
  and g_137303_(_047746_, _047753_, _047754_);
  or g_137304_(_047745_, _047752_, _047755_);
  xor g_137305_(out[808], _047711_, _047756_);
  xor g_137306_(_001121_, _047711_, _047757_);
  and g_137307_(_047514_, _047696_, _047758_);
  or g_137308_(_047513_, _047697_, _047759_);
  and g_137309_(_047521_, _047697_, _047760_);
  or g_137310_(_047520_, _047696_, _047762_);
  and g_137311_(_047759_, _047762_, _047763_);
  or g_137312_(_047758_, _047760_, _047764_);
  and g_137313_(_047756_, _047764_, _047765_);
  or g_137314_(_047757_, _047763_, _047766_);
  and g_137315_(_047755_, _047766_, _047767_);
  or g_137316_(_047754_, _047765_, _047768_);
  xor g_137317_(out[807], _047710_, _047769_);
  xor g_137318_(_001033_, _047710_, _047770_);
  and g_137319_(_047545_, _047696_, _047771_);
  or g_137320_(_047544_, _047697_, _047773_);
  and g_137321_(_047551_, _047697_, _047774_);
  or g_137322_(_047550_, _047696_, _047775_);
  and g_137323_(_047773_, _047775_, _047776_);
  or g_137324_(_047771_, _047774_, _047777_);
  and g_137325_(_047769_, _047777_, _047778_);
  or g_137326_(_047770_, _047776_, _047779_);
  xor g_137327_(out[801], out[800], _047780_);
  xor g_137328_(_001077_, out[800], _047781_);
  and g_137329_(_047633_, _047697_, _047782_);
  or g_137330_(_047632_, _047696_, _047784_);
  and g_137331_(_047627_, _047696_, _047785_);
  or g_137332_(_047628_, _047697_, _047786_);
  and g_137333_(_047784_, _047786_, _047787_);
  or g_137334_(_047782_, _047785_, _047788_);
  and g_137335_(_047780_, _047787_, _047789_);
  or g_137336_(_047781_, _047788_, _047790_);
  and g_137337_(out[784], _047696_, _047791_);
  or g_137338_(_000956_, _047697_, _047792_);
  and g_137339_(_047642_, _047697_, _047793_);
  or g_137340_(_047641_, _047696_, _047795_);
  and g_137341_(_047792_, _047795_, _047796_);
  or g_137342_(_047791_, _047793_, _047797_);
  and g_137343_(out[800], _047796_, _047798_);
  or g_137344_(_001088_, _047797_, _047799_);
  and g_137345_(_047790_, _047799_, _047800_);
  or g_137346_(_047789_, _047798_, _047801_);
  xor g_137347_(out[802], _047704_, _047802_);
  xor g_137348_(_001099_, _047704_, _047803_);
  and g_137349_(_047612_, _047696_, _047804_);
  or g_137350_(_047613_, _047697_, _047806_);
  and g_137351_(_047620_, _047697_, _047807_);
  or g_137352_(_047619_, _047696_, _047808_);
  and g_137353_(_047806_, _047808_, _047809_);
  or g_137354_(_047804_, _047807_, _047810_);
  and g_137355_(_047803_, _047810_, _047811_);
  or g_137356_(_047802_, _047809_, _047812_);
  and g_137357_(out[801], _047788_, _047813_);
  or g_137358_(_001077_, _047787_, _047814_);
  and g_137359_(_047812_, _047814_, _047815_);
  or g_137360_(_047811_, _047813_, _047817_);
  and g_137361_(_047801_, _047815_, _047818_);
  or g_137362_(_047800_, _047817_, _047819_);
  xor g_137363_(out[803], _047705_, _047820_);
  xor g_137364_(_001110_, _047705_, _047821_);
  and g_137365_(_047600_, _047696_, _047822_);
  or g_137366_(_047599_, _047697_, _047823_);
  and g_137367_(_047606_, _047697_, _047824_);
  or g_137368_(_047605_, _047696_, _047825_);
  and g_137369_(_047823_, _047825_, _047826_);
  or g_137370_(_047822_, _047824_, _047828_);
  and g_137371_(_047821_, _047826_, _047829_);
  or g_137372_(_047820_, _047828_, _047830_);
  and g_137373_(_047802_, _047809_, _047831_);
  or g_137374_(_047803_, _047810_, _047832_);
  and g_137375_(_047830_, _047832_, _047833_);
  or g_137376_(_047829_, _047831_, _047834_);
  and g_137377_(_047819_, _047833_, _047835_);
  or g_137378_(_047818_, _047834_, _047836_);
  and g_137379_(_047820_, _047828_, _047837_);
  or g_137380_(_047821_, _047826_, _047839_);
  xor g_137381_(out[804], _047707_, _047840_);
  xor g_137382_(_001066_, _047707_, _047841_);
  and g_137383_(_047703_, _047840_, _047842_);
  or g_137384_(_047702_, _047841_, _047843_);
  and g_137385_(_047839_, _047843_, _047844_);
  or g_137386_(_047837_, _047842_, _047845_);
  and g_137387_(_047836_, _047844_, _047846_);
  or g_137388_(_047835_, _047845_, _047847_);
  xor g_137389_(out[805], _047708_, _047848_);
  xor g_137390_(_001055_, _047708_, _047850_);
  and g_137391_(_047565_, _047696_, _047851_);
  or g_137392_(_047564_, _047697_, _047852_);
  and g_137393_(_047571_, _047697_, _047853_);
  or g_137394_(_047570_, _047696_, _047854_);
  and g_137395_(_047852_, _047854_, _047855_);
  or g_137396_(_047851_, _047853_, _047856_);
  and g_137397_(_047850_, _047855_, _047857_);
  or g_137398_(_047848_, _047856_, _047858_);
  and g_137399_(_047702_, _047841_, _047859_);
  or g_137400_(_047703_, _047840_, _047861_);
  and g_137401_(_047858_, _047861_, _047862_);
  or g_137402_(_047857_, _047859_, _047863_);
  and g_137403_(_047847_, _047862_, _047864_);
  or g_137404_(_047846_, _047863_, _047865_);
  xor g_137405_(out[806], _047709_, _047866_);
  xor g_137406_(_001044_, _047709_, _047867_);
  and g_137407_(_047533_, _047696_, _047868_);
  or g_137408_(_047534_, _047697_, _047869_);
  and g_137409_(_047540_, _047697_, _047870_);
  or g_137410_(_047539_, _047696_, _047872_);
  and g_137411_(_047869_, _047872_, _047873_);
  or g_137412_(_047868_, _047870_, _047874_);
  and g_137413_(_047867_, _047874_, _047875_);
  or g_137414_(_047866_, _047873_, _047876_);
  and g_137415_(_047848_, _047856_, _047877_);
  or g_137416_(_047850_, _047855_, _047878_);
  and g_137417_(_047876_, _047878_, _047879_);
  or g_137418_(_047875_, _047877_, _047880_);
  and g_137419_(_047865_, _047879_, _047881_);
  or g_137420_(_047864_, _047880_, _047883_);
  and g_137421_(_047770_, _047776_, _047884_);
  or g_137422_(_047769_, _047777_, _047885_);
  and g_137423_(_047866_, _047873_, _047886_);
  or g_137424_(_047867_, _047874_, _047887_);
  and g_137425_(_047885_, _047887_, _047888_);
  or g_137426_(_047884_, _047886_, _047889_);
  and g_137427_(_047883_, _047888_, _047890_);
  or g_137428_(_047881_, _047889_, _047891_);
  and g_137429_(_047779_, _047891_, _047892_);
  or g_137430_(_047778_, _047890_, _047894_);
  and g_137431_(_047757_, _047763_, _047895_);
  or g_137432_(_047756_, _047764_, _047896_);
  and g_137433_(_047745_, _047752_, _047897_);
  or g_137434_(_047746_, _047753_, _047898_);
  xor g_137435_(_047715_, _047722_, _047899_);
  xor g_137436_(_047715_, _047721_, _047900_);
  xor g_137437_(_047724_, _047737_, _047901_);
  xor g_137438_(_047725_, _047737_, _047902_);
  and g_137439_(_047899_, _047901_, _047903_);
  or g_137440_(_047900_, _047902_, _047905_);
  and g_137441_(_047768_, _047903_, _047906_);
  or g_137442_(_047767_, _047905_, _047907_);
  and g_137443_(_047898_, _047906_, _047908_);
  or g_137444_(_047897_, _047907_, _047909_);
  and g_137445_(_047766_, _047898_, _047910_);
  or g_137446_(_047765_, _047897_, _047911_);
  and g_137447_(_047755_, _047896_, _047912_);
  or g_137448_(_047754_, _047895_, _047913_);
  and g_137449_(_047903_, _047912_, _047914_);
  or g_137450_(_047905_, _047913_, _047916_);
  and g_137451_(_047910_, _047914_, _047917_);
  or g_137452_(_047911_, _047916_, _047918_);
  and g_137453_(_047894_, _047917_, _047919_);
  or g_137454_(_047892_, _047918_, _047920_);
  and g_137455_(_047744_, _047920_, _047921_);
  or g_137456_(_047743_, _047919_, _047922_);
  and g_137457_(_047909_, _047921_, _047923_);
  or g_137458_(_047908_, _047922_, _047924_);
  and g_137459_(_047703_, _047924_, _047925_);
  not g_137460_(_047925_, _047927_);
  or g_137461_(_047840_, _047924_, _047928_);
  not g_137462_(_047928_, _047929_);
  and g_137463_(_047927_, _047928_, _047930_);
  or g_137464_(_047925_, _047929_, _047931_);
  and g_137465_(_043388_, _047930_, _047932_);
  or g_137466_(_043387_, _047931_, _047933_);
  xor g_137467_(out[819], _043378_, _047934_);
  xor g_137468_(_001242_, _043378_, _047935_);
  and g_137469_(_047828_, _047924_, _047936_);
  or g_137470_(_047826_, _047923_, _047938_);
  and g_137471_(_047821_, _047923_, _047939_);
  or g_137472_(_047820_, _047924_, _047940_);
  and g_137473_(_047938_, _047940_, _047941_);
  or g_137474_(_047936_, _047939_, _047942_);
  and g_137475_(_047934_, _047942_, _047943_);
  or g_137476_(_047935_, _047941_, _047944_);
  xor g_137477_(out[817], out[816], _047945_);
  xor g_137478_(_001209_, out[816], _047946_);
  and g_137479_(_047780_, _047923_, _047947_);
  or g_137480_(_047781_, _047924_, _047949_);
  and g_137481_(_047788_, _047924_, _047950_);
  or g_137482_(_047787_, _047923_, _047951_);
  and g_137483_(_047949_, _047951_, _047952_);
  or g_137484_(_047947_, _047950_, _047953_);
  and g_137485_(_047945_, _047952_, _047954_);
  or g_137486_(_047946_, _047953_, _047955_);
  and g_137487_(_047797_, _047924_, _047956_);
  or g_137488_(_047796_, _047923_, _047957_);
  and g_137489_(out[800], _047923_, _047958_);
  or g_137490_(_001088_, _047924_, _047960_);
  and g_137491_(_047957_, _047960_, _047961_);
  or g_137492_(_047956_, _047958_, _047962_);
  and g_137493_(out[816], _047961_, _047963_);
  or g_137494_(_001220_, _047962_, _047964_);
  and g_137495_(_047955_, _047964_, _047965_);
  or g_137496_(_047954_, _047963_, _047966_);
  xor g_137497_(out[818], _043377_, _047967_);
  xor g_137498_(_001231_, _043377_, _047968_);
  and g_137499_(_047810_, _047924_, _047969_);
  or g_137500_(_047809_, _047923_, _047971_);
  and g_137501_(_047802_, _047923_, _047972_);
  or g_137502_(_047803_, _047924_, _047973_);
  and g_137503_(_047971_, _047973_, _047974_);
  or g_137504_(_047969_, _047972_, _047975_);
  and g_137505_(_047968_, _047975_, _047976_);
  or g_137506_(_047967_, _047974_, _047977_);
  and g_137507_(out[817], _047953_, _047978_);
  or g_137508_(_001209_, _047952_, _047979_);
  and g_137509_(_047977_, _047979_, _047980_);
  or g_137510_(_047976_, _047978_, _047982_);
  and g_137511_(_047966_, _047980_, _047983_);
  or g_137512_(_047965_, _047982_, _047984_);
  and g_137513_(_047935_, _047941_, _047985_);
  or g_137514_(_047934_, _047942_, _047986_);
  and g_137515_(_047967_, _047974_, _047987_);
  or g_137516_(_047968_, _047975_, _047988_);
  and g_137517_(_047986_, _047988_, _047989_);
  or g_137518_(_047985_, _047987_, _047990_);
  and g_137519_(_047984_, _047989_, _047991_);
  or g_137520_(_047983_, _047990_, _047993_);
  and g_137521_(_047944_, _047993_, _047994_);
  or g_137522_(_047943_, _047991_, _047995_);
  and g_137523_(_047933_, _047995_, _047996_);
  or g_137524_(_047932_, _047994_, _047997_);
  xor g_137525_(out[821], _043380_, _047998_);
  xor g_137526_(_001187_, _043380_, _047999_);
  or g_137527_(_047848_, _047924_, _048000_);
  not g_137528_(_048000_, _048001_);
  and g_137529_(_047856_, _047924_, _048002_);
  not g_137530_(_048002_, _048004_);
  and g_137531_(_048000_, _048004_, _048005_);
  or g_137532_(_048001_, _048002_, _048006_);
  and g_137533_(_047998_, _048006_, _048007_);
  or g_137534_(_047999_, _048005_, _048008_);
  and g_137535_(_043387_, _047931_, _048009_);
  or g_137536_(_043388_, _047930_, _048010_);
  and g_137537_(_048008_, _048010_, _048011_);
  or g_137538_(_048007_, _048009_, _048012_);
  and g_137539_(_047997_, _048011_, _048013_);
  or g_137540_(_047996_, _048012_, _048015_);
  xor g_137541_(out[822], _043381_, _048016_);
  xor g_137542_(_001176_, _043381_, _048017_);
  or g_137543_(_047867_, _047924_, _048018_);
  or g_137544_(_047873_, _047923_, _048019_);
  and g_137545_(_048018_, _048019_, _048020_);
  not g_137546_(_048020_, _048021_);
  and g_137547_(_048016_, _048020_, _048022_);
  or g_137548_(_048017_, _048021_, _048023_);
  and g_137549_(_047999_, _048005_, _048024_);
  or g_137550_(_047998_, _048006_, _048026_);
  and g_137551_(_048023_, _048026_, _048027_);
  or g_137552_(_048022_, _048024_, _048028_);
  and g_137553_(_048015_, _048027_, _048029_);
  or g_137554_(_048013_, _048028_, _048030_);
  or g_137555_(_047769_, _047924_, _048031_);
  or g_137556_(_047776_, _047923_, _048032_);
  and g_137557_(_048031_, _048032_, _048033_);
  not g_137558_(_048033_, _048034_);
  and g_137559_(_043385_, _048034_, _048035_);
  or g_137560_(_043386_, _048033_, _048037_);
  and g_137561_(_048017_, _048021_, _048038_);
  or g_137562_(_048016_, _048020_, _048039_);
  and g_137563_(_048037_, _048039_, _048040_);
  or g_137564_(_048035_, _048038_, _048041_);
  and g_137565_(_048030_, _048040_, _048042_);
  or g_137566_(_048029_, _048041_, _048043_);
  and g_137567_(out[824], _043384_, _048044_);
  xor g_137568_(out[824], _043384_, _048045_);
  xor g_137569_(_001253_, _043384_, _048046_);
  or g_137570_(_047756_, _047924_, _048048_);
  not g_137571_(_048048_, _048049_);
  and g_137572_(_047764_, _047924_, _048050_);
  not g_137573_(_048050_, _048051_);
  and g_137574_(_048048_, _048051_, _048052_);
  or g_137575_(_048049_, _048050_, _048053_);
  and g_137576_(_048046_, _048052_, _048054_);
  or g_137577_(_048045_, _048053_, _048055_);
  or g_137578_(out[825], _048044_, _048056_);
  and g_137579_(out[826], _048056_, _048057_);
  xor g_137580_(out[827], _048057_, _048059_);
  xor g_137581_(_001154_, _048057_, _048060_);
  and g_137582_(_047724_, _047731_, _048061_);
  or g_137583_(_047725_, _047732_, _048062_);
  and g_137584_(_048060_, _048061_, _048063_);
  or g_137585_(_048059_, _048062_, _048064_);
  and g_137586_(_043386_, _048033_, _048065_);
  or g_137587_(_043385_, _048034_, _048066_);
  and g_137588_(_048064_, _048066_, _048067_);
  or g_137589_(_048063_, _048065_, _048068_);
  and g_137590_(_048055_, _048067_, _048070_);
  or g_137591_(_048054_, _048068_, _048071_);
  xor g_137592_(out[825], _048044_, _048072_);
  xor g_137593_(_001264_, _048044_, _048073_);
  and g_137594_(_047753_, _047924_, _048074_);
  not g_137595_(_048074_, _048075_);
  or g_137596_(_047746_, _047924_, _048076_);
  not g_137597_(_048076_, _048077_);
  and g_137598_(_048075_, _048076_, _048078_);
  or g_137599_(_048074_, _048077_, _048079_);
  and g_137600_(_048073_, _048079_, _048081_);
  or g_137601_(_048072_, _048078_, _048082_);
  and g_137602_(_048045_, _048053_, _048083_);
  or g_137603_(_048046_, _048052_, _048084_);
  and g_137604_(_048082_, _048084_, _048085_);
  or g_137605_(_048081_, _048083_, _048086_);
  xor g_137606_(out[826], _048056_, _048087_);
  xor g_137607_(_001275_, _048056_, _048088_);
  or g_137608_(_047715_, _047924_, _048089_);
  not g_137609_(_048089_, _048090_);
  and g_137610_(_047722_, _047924_, _048092_);
  not g_137611_(_048092_, _048093_);
  and g_137612_(_048089_, _048093_, _048094_);
  or g_137613_(_048090_, _048092_, _048095_);
  and g_137614_(_048087_, _048095_, _048096_);
  or g_137615_(_048088_, _048094_, _048097_);
  and g_137616_(_047724_, _047738_, _048098_);
  or g_137617_(_047725_, _047737_, _048099_);
  and g_137618_(_048059_, _048062_, _048100_);
  or g_137619_(_048060_, _048061_, _048101_);
  and g_137620_(_048097_, _048101_, _048103_);
  or g_137621_(_048096_, _048100_, _048104_);
  and g_137622_(_048088_, _048094_, _048105_);
  or g_137623_(_048087_, _048095_, _048106_);
  and g_137624_(_048072_, _048078_, _048107_);
  or g_137625_(_048073_, _048079_, _048108_);
  and g_137626_(_048106_, _048108_, _048109_);
  or g_137627_(_048105_, _048107_, _048110_);
  and g_137628_(_048103_, _048109_, _048111_);
  or g_137629_(_048104_, _048110_, _048112_);
  and g_137630_(_048085_, _048111_, _048114_);
  or g_137631_(_048086_, _048112_, _048115_);
  and g_137632_(_048070_, _048114_, _048116_);
  or g_137633_(_048071_, _048115_, _048117_);
  and g_137634_(_048043_, _048116_, _048118_);
  or g_137635_(_048042_, _048117_, _048119_);
  and g_137636_(_048086_, _048109_, _048120_);
  or g_137637_(_048085_, _048110_, _048121_);
  and g_137638_(_048103_, _048121_, _048122_);
  or g_137639_(_048104_, _048120_, _048123_);
  and g_137640_(_048064_, _048123_, _048125_);
  or g_137641_(_048063_, _048122_, _048126_);
  and g_137642_(_048119_, _048126_, _048127_);
  or g_137643_(_048118_, _048125_, _048128_);
  or g_137644_(_043385_, _048128_, _048129_);
  or g_137645_(_048033_, _048127_, _048130_);
  and g_137646_(_048129_, _048130_, _048131_);
  not g_137647_(_048131_, _048132_);
  and g_137648_(_043375_, _048132_, _048133_);
  or g_137649_(_043376_, _048131_, _048134_);
  xor g_137650_(out[837], _043370_, _048136_);
  xor g_137651_(_001319_, _043370_, _048137_);
  and g_137652_(_048006_, _048128_, _048138_);
  or g_137653_(_048005_, _048127_, _048139_);
  and g_137654_(_047999_, _048127_, _048140_);
  or g_137655_(_047998_, _048128_, _048141_);
  and g_137656_(_048139_, _048141_, _048142_);
  or g_137657_(_048138_, _048140_, _048143_);
  and g_137658_(_048137_, _048142_, _048144_);
  or g_137659_(_048136_, _048143_, _048145_);
  xor g_137660_(out[836], _043367_, _048147_);
  xor g_137661_(_001330_, _043367_, _048148_);
  and g_137662_(_043388_, _048127_, _048149_);
  or g_137663_(_043387_, _048128_, _048150_);
  and g_137664_(_047931_, _048128_, _048151_);
  or g_137665_(_047930_, _048127_, _048152_);
  and g_137666_(_048150_, _048152_, _048153_);
  or g_137667_(_048149_, _048151_, _048154_);
  and g_137668_(_048147_, _048154_, _048155_);
  or g_137669_(_048148_, _048153_, _048156_);
  xor g_137670_(out[834], _043365_, _048158_);
  xor g_137671_(_001363_, _043365_, _048159_);
  and g_137672_(_047975_, _048128_, _048160_);
  or g_137673_(_047974_, _048127_, _048161_);
  and g_137674_(_047967_, _048127_, _048162_);
  or g_137675_(_047968_, _048128_, _048163_);
  and g_137676_(_048161_, _048163_, _048164_);
  or g_137677_(_048160_, _048162_, _048165_);
  and g_137678_(_048158_, _048164_, _048166_);
  or g_137679_(_048159_, _048165_, _048167_);
  and g_137680_(_047945_, _048127_, _048169_);
  or g_137681_(_047946_, _048128_, _048170_);
  and g_137682_(_047953_, _048128_, _048171_);
  or g_137683_(_047952_, _048127_, _048172_);
  and g_137684_(_048170_, _048172_, _048173_);
  or g_137685_(_048169_, _048171_, _048174_);
  and g_137686_(out[833], _048174_, _048175_);
  not g_137687_(_048175_, _048176_);
  xor g_137688_(out[833], out[832], _048177_);
  xor g_137689_(_001341_, out[832], _048178_);
  and g_137690_(_048173_, _048177_, _048180_);
  or g_137691_(_048174_, _048178_, _048181_);
  and g_137692_(out[816], _048127_, _048182_);
  or g_137693_(_001220_, _048128_, _048183_);
  and g_137694_(_047962_, _048128_, _048184_);
  or g_137695_(_047961_, _048127_, _048185_);
  and g_137696_(_048183_, _048185_, _048186_);
  or g_137697_(_048182_, _048184_, _048187_);
  and g_137698_(out[832], _048186_, _048188_);
  or g_137699_(_001352_, _048187_, _048189_);
  and g_137700_(_048181_, _048189_, _048191_);
  or g_137701_(_048180_, _048188_, _048192_);
  and g_137702_(_048176_, _048192_, _048193_);
  or g_137703_(_048175_, _048191_, _048194_);
  and g_137704_(_048167_, _048194_, _048195_);
  or g_137705_(_048166_, _048193_, _048196_);
  and g_137706_(_048159_, _048165_, _048197_);
  or g_137707_(_048158_, _048164_, _048198_);
  and g_137708_(_047942_, _048128_, _048199_);
  or g_137709_(_047941_, _048127_, _048200_);
  and g_137710_(_047935_, _048127_, _048202_);
  or g_137711_(_047934_, _048128_, _048203_);
  and g_137712_(_048200_, _048203_, _048204_);
  or g_137713_(_048199_, _048202_, _048205_);
  and g_137714_(_043368_, _048205_, _048206_);
  or g_137715_(_043369_, _048204_, _048207_);
  and g_137716_(_048198_, _048207_, _048208_);
  or g_137717_(_048197_, _048206_, _048209_);
  and g_137718_(_048196_, _048208_, _048210_);
  or g_137719_(_048195_, _048209_, _048211_);
  and g_137720_(_048148_, _048153_, _048213_);
  or g_137721_(_048147_, _048154_, _048214_);
  and g_137722_(_043369_, _048204_, _048215_);
  or g_137723_(_043368_, _048205_, _048216_);
  and g_137724_(_048214_, _048216_, _048217_);
  or g_137725_(_048213_, _048215_, _048218_);
  and g_137726_(_048211_, _048217_, _048219_);
  or g_137727_(_048210_, _048218_, _048220_);
  and g_137728_(_048156_, _048220_, _048221_);
  or g_137729_(_048155_, _048219_, _048222_);
  and g_137730_(_048145_, _048222_, _048224_);
  or g_137731_(_048144_, _048221_, _048225_);
  xor g_137732_(out[838], _043371_, _048226_);
  xor g_137733_(_001308_, _043371_, _048227_);
  or g_137734_(_048017_, _048128_, _048228_);
  or g_137735_(_048020_, _048127_, _048229_);
  and g_137736_(_048228_, _048229_, _048230_);
  not g_137737_(_048230_, _048231_);
  and g_137738_(_048227_, _048231_, _048232_);
  or g_137739_(_048226_, _048230_, _048233_);
  and g_137740_(_048136_, _048143_, _048235_);
  or g_137741_(_048137_, _048142_, _048236_);
  and g_137742_(_048233_, _048236_, _048237_);
  or g_137743_(_048232_, _048235_, _048238_);
  and g_137744_(_048225_, _048237_, _048239_);
  or g_137745_(_048224_, _048238_, _048240_);
  and g_137746_(_043376_, _048131_, _048241_);
  or g_137747_(_043375_, _048132_, _048242_);
  and g_137748_(_048226_, _048230_, _048243_);
  or g_137749_(_048227_, _048231_, _048244_);
  and g_137750_(_048242_, _048244_, _048246_);
  or g_137751_(_048241_, _048243_, _048247_);
  and g_137752_(_048240_, _048246_, _048248_);
  or g_137753_(_048239_, _048247_, _048249_);
  and g_137754_(_048134_, _048249_, _048250_);
  or g_137755_(_048133_, _048248_, _048251_);
  and g_137756_(out[840], _043374_, _048252_);
  or g_137757_(out[841], _048252_, _048253_);
  and g_137758_(out[842], _048253_, _048254_);
  xor g_137759_(out[842], _048253_, _048255_);
  xor g_137760_(_001407_, _048253_, _048257_);
  and g_137761_(_048088_, _048127_, _048258_);
  or g_137762_(_048087_, _048128_, _048259_);
  and g_137763_(_048095_, _048128_, _048260_);
  or g_137764_(_048094_, _048127_, _048261_);
  and g_137765_(_048259_, _048261_, _048262_);
  or g_137766_(_048258_, _048260_, _048263_);
  and g_137767_(_048255_, _048263_, _048264_);
  or g_137768_(_048257_, _048262_, _048265_);
  xor g_137769_(out[843], _048254_, _048266_);
  xor g_137770_(_001286_, _048254_, _048268_);
  and g_137771_(_048059_, _048061_, _048269_);
  and g_137772_(_048059_, _048098_, _048270_);
  or g_137773_(_048060_, _048099_, _048271_);
  and g_137774_(_048266_, _048271_, _048272_);
  or g_137775_(_048268_, _048269_, _048273_);
  and g_137776_(_048265_, _048273_, _048274_);
  or g_137777_(_048264_, _048272_, _048275_);
  and g_137778_(_048257_, _048262_, _048276_);
  or g_137779_(_048255_, _048263_, _048277_);
  and g_137780_(_048268_, _048270_, _048279_);
  or g_137781_(_048266_, _048271_, _048280_);
  and g_137782_(_048277_, _048280_, _048281_);
  or g_137783_(_048276_, _048279_, _048282_);
  xor g_137784_(out[841], _048252_, _048283_);
  xor g_137785_(_001396_, _048252_, _048284_);
  and g_137786_(_048072_, _048127_, _048285_);
  or g_137787_(_048073_, _048128_, _048286_);
  and g_137788_(_048079_, _048128_, _048287_);
  or g_137789_(_048078_, _048127_, _048288_);
  and g_137790_(_048286_, _048288_, _048290_);
  or g_137791_(_048285_, _048287_, _048291_);
  and g_137792_(_048283_, _048290_, _048292_);
  or g_137793_(_048284_, _048291_, _048293_);
  and g_137794_(_048281_, _048293_, _048294_);
  or g_137795_(_048282_, _048292_, _048295_);
  and g_137796_(_048274_, _048294_, _048296_);
  or g_137797_(_048275_, _048295_, _048297_);
  and g_137798_(_048284_, _048291_, _048298_);
  or g_137799_(_048283_, _048290_, _048299_);
  xor g_137800_(out[840], _043374_, _048301_);
  xor g_137801_(_001385_, _043374_, _048302_);
  and g_137802_(_048046_, _048127_, _048303_);
  or g_137803_(_048045_, _048128_, _048304_);
  and g_137804_(_048053_, _048128_, _048305_);
  or g_137805_(_048052_, _048127_, _048306_);
  and g_137806_(_048304_, _048306_, _048307_);
  or g_137807_(_048303_, _048305_, _048308_);
  and g_137808_(_048301_, _048308_, _048309_);
  or g_137809_(_048302_, _048307_, _048310_);
  and g_137810_(_048299_, _048310_, _048312_);
  or g_137811_(_048298_, _048309_, _048313_);
  and g_137812_(_048302_, _048307_, _048314_);
  or g_137813_(_048301_, _048308_, _048315_);
  and g_137814_(_048312_, _048315_, _048316_);
  or g_137815_(_048313_, _048314_, _048317_);
  and g_137816_(_048296_, _048316_, _048318_);
  or g_137817_(_048297_, _048317_, _048319_);
  and g_137818_(_048251_, _048318_, _048320_);
  or g_137819_(_048250_, _048319_, _048321_);
  and g_137820_(_048296_, _048313_, _048323_);
  or g_137821_(_048297_, _048312_, _048324_);
  and g_137822_(_048275_, _048280_, _048325_);
  or g_137823_(_048274_, _048279_, _048326_);
  and g_137824_(_048324_, _048326_, _048327_);
  or g_137825_(_048323_, _048325_, _048328_);
  and g_137826_(_048321_, _048327_, _048329_);
  or g_137827_(_048320_, _048328_, _048330_);
  or g_137828_(_043368_, _048330_, _048331_);
  not g_137829_(_048331_, _048332_);
  and g_137830_(_048205_, _048330_, _048334_);
  not g_137831_(_048334_, _048335_);
  and g_137832_(_048331_, _048335_, _048336_);
  or g_137833_(_048332_, _048334_, _048337_);
  and g_137834_(_043363_, _048337_, _048338_);
  or g_137835_(_043364_, _048336_, _048339_);
  and g_137836_(_043364_, _048336_, _048340_);
  or g_137837_(_043363_, _048337_, _048341_);
  xor g_137838_(out[850], _043353_, _048342_);
  not g_137839_(_048342_, _048343_);
  and g_137840_(_048165_, _048330_, _048345_);
  not g_137841_(_048345_, _048346_);
  or g_137842_(_048159_, _048330_, _048347_);
  not g_137843_(_048347_, _048348_);
  and g_137844_(_048346_, _048347_, _048349_);
  or g_137845_(_048345_, _048348_, _048350_);
  and g_137846_(_048342_, _048349_, _048351_);
  or g_137847_(_048343_, _048350_, _048352_);
  and g_137848_(_048341_, _048352_, _048353_);
  or g_137849_(_048340_, _048351_, _048354_);
  and g_137850_(_048339_, _048354_, _048356_);
  or g_137851_(_048338_, _048353_, _048357_);
  xor g_137852_(out[849], out[848], _048358_);
  xor g_137853_(_001473_, out[848], _048359_);
  and g_137854_(_048177_, _048329_, _048360_);
  and g_137855_(_048174_, _048330_, _048361_);
  or g_137856_(_048360_, _048361_, _048362_);
  not g_137857_(_048362_, _048363_);
  or g_137858_(_048359_, _048362_, _048364_);
  not g_137859_(_048364_, _048365_);
  and g_137860_(out[832], _048329_, _048367_);
  or g_137861_(_001352_, _048330_, _048368_);
  and g_137862_(_048187_, _048330_, _048369_);
  or g_137863_(_048186_, _048329_, _048370_);
  and g_137864_(_048368_, _048370_, _048371_);
  or g_137865_(_048367_, _048369_, _048372_);
  and g_137866_(_001484_, _048372_, _048373_);
  or g_137867_(out[848], _048371_, _048374_);
  xor g_137868_(_048359_, _048362_, _048375_);
  xor g_137869_(_048358_, _048362_, _048376_);
  and g_137870_(_048374_, _048375_, _048378_);
  or g_137871_(_048373_, _048376_, _048379_);
  and g_137872_(_048364_, _048379_, _048380_);
  or g_137873_(_048365_, _048378_, _048381_);
  and g_137874_(_048343_, _048350_, _048382_);
  or g_137875_(_048342_, _048349_, _048383_);
  and g_137876_(_048339_, _048383_, _048384_);
  or g_137877_(_048338_, _048382_, _048385_);
  and g_137878_(_048381_, _048384_, _048386_);
  or g_137879_(_048380_, _048385_, _048387_);
  and g_137880_(_048357_, _048387_, _048389_);
  or g_137881_(_048356_, _048386_, _048390_);
  and g_137882_(out[856], _043359_, _048391_);
  or g_137883_(out[857], _048391_, _048392_);
  xor g_137884_(out[857], _048391_, _048393_);
  not g_137885_(_048393_, _048394_);
  and g_137886_(_048291_, _048330_, _048395_);
  or g_137887_(_048290_, _048329_, _048396_);
  and g_137888_(_048283_, _048329_, _048397_);
  or g_137889_(_048284_, _048330_, _048398_);
  and g_137890_(_048396_, _048398_, _048400_);
  or g_137891_(_048395_, _048397_, _048401_);
  and g_137892_(_048393_, _048400_, _048402_);
  or g_137893_(_048394_, _048401_, _048403_);
  xor g_137894_(out[856], _043359_, _048404_);
  xor g_137895_(_001517_, _043359_, _048405_);
  and g_137896_(_048308_, _048330_, _048406_);
  or g_137897_(_048307_, _048329_, _048407_);
  and g_137898_(_048302_, _048329_, _048408_);
  or g_137899_(_048301_, _048330_, _048409_);
  and g_137900_(_048407_, _048409_, _048411_);
  or g_137901_(_048406_, _048408_, _048412_);
  and g_137902_(_048405_, _048411_, _048413_);
  or g_137903_(_048404_, _048412_, _048414_);
  and g_137904_(_048403_, _048414_, _048415_);
  or g_137905_(_048402_, _048413_, _048416_);
  and g_137906_(out[858], _048392_, _048417_);
  xor g_137907_(out[859], _048417_, _048418_);
  xor g_137908_(_001418_, _048417_, _048419_);
  and g_137909_(_048266_, _048269_, _048420_);
  or g_137910_(_048268_, _048271_, _048422_);
  and g_137911_(_048418_, _048422_, _048423_);
  or g_137912_(_048419_, _048420_, _048424_);
  and g_137913_(_048404_, _048412_, _048425_);
  or g_137914_(_048405_, _048411_, _048426_);
  and g_137915_(_048424_, _048426_, _048427_);
  or g_137916_(_048423_, _048425_, _048428_);
  and g_137917_(_048415_, _048427_, _048429_);
  or g_137918_(_048416_, _048428_, _048430_);
  xor g_137919_(out[858], _048392_, _048431_);
  xor g_137920_(_001539_, _048392_, _048433_);
  and g_137921_(_048263_, _048330_, _048434_);
  or g_137922_(_048262_, _048329_, _048435_);
  and g_137923_(_048257_, _048329_, _048436_);
  or g_137924_(_048255_, _048330_, _048437_);
  and g_137925_(_048435_, _048437_, _048438_);
  or g_137926_(_048434_, _048436_, _048439_);
  and g_137927_(_048433_, _048438_, _048440_);
  or g_137928_(_048431_, _048439_, _048441_);
  or g_137929_(_048418_, _048422_, _048442_);
  not g_137930_(_048442_, _048444_);
  and g_137931_(_048441_, _048442_, _048445_);
  or g_137932_(_048440_, _048444_, _048446_);
  and g_137933_(_048431_, _048439_, _048447_);
  or g_137934_(_048433_, _048438_, _048448_);
  and g_137935_(_048394_, _048401_, _048449_);
  or g_137936_(_048393_, _048400_, _048450_);
  and g_137937_(_048448_, _048450_, _048451_);
  or g_137938_(_048447_, _048449_, _048452_);
  and g_137939_(_048445_, _048451_, _048453_);
  or g_137940_(_048446_, _048452_, _048455_);
  and g_137941_(_048429_, _048453_, _048456_);
  or g_137942_(_048430_, _048455_, _048457_);
  or g_137943_(_048131_, _048329_, _048458_);
  or g_137944_(_043375_, _048330_, _048459_);
  and g_137945_(_048458_, _048459_, _048460_);
  and g_137946_(_043360_, _048460_, _048461_);
  or g_137947_(_043360_, _048460_, _048462_);
  xor g_137948_(_043360_, _048460_, _048463_);
  xor g_137949_(_043362_, _048460_, _048464_);
  xor g_137950_(out[854], _043357_, _048466_);
  not g_137951_(_048466_, _048467_);
  or g_137952_(_048230_, _048329_, _048468_);
  or g_137953_(_048227_, _048330_, _048469_);
  and g_137954_(_048468_, _048469_, _048470_);
  and g_137955_(_048466_, _048470_, _048471_);
  xor g_137956_(_048466_, _048470_, _048472_);
  xor g_137957_(_048467_, _048470_, _048473_);
  and g_137958_(_048463_, _048472_, _048474_);
  or g_137959_(_048464_, _048473_, _048475_);
  xor g_137960_(out[852], _043355_, _048477_);
  xor g_137961_(_001462_, _043355_, _048478_);
  and g_137962_(_048148_, _048329_, _048479_);
  or g_137963_(_048147_, _048330_, _048480_);
  and g_137964_(_048154_, _048330_, _048481_);
  or g_137965_(_048153_, _048329_, _048482_);
  and g_137966_(_048480_, _048482_, _048483_);
  or g_137967_(_048479_, _048481_, _048484_);
  and g_137968_(_048478_, _048483_, _048485_);
  or g_137969_(_048477_, _048484_, _048486_);
  xor g_137970_(out[853], _043356_, _048488_);
  xor g_137971_(_001451_, _043356_, _048489_);
  and g_137972_(_048137_, _048329_, _048490_);
  or g_137973_(_048136_, _048330_, _048491_);
  and g_137974_(_048143_, _048330_, _048492_);
  or g_137975_(_048142_, _048329_, _048493_);
  and g_137976_(_048491_, _048493_, _048494_);
  or g_137977_(_048490_, _048492_, _048495_);
  and g_137978_(_048489_, _048494_, _048496_);
  or g_137979_(_048488_, _048495_, _048497_);
  and g_137980_(_048486_, _048497_, _048499_);
  or g_137981_(_048485_, _048496_, _048500_);
  or g_137982_(_048489_, _048494_, _048501_);
  not g_137983_(_048501_, _048502_);
  or g_137984_(_048478_, _048483_, _048503_);
  and g_137985_(_048501_, _048503_, _048504_);
  not g_137986_(_048504_, _048505_);
  and g_137987_(_048499_, _048504_, _048506_);
  or g_137988_(_048500_, _048505_, _048507_);
  and g_137989_(_048474_, _048506_, _048508_);
  or g_137990_(_048457_, _048507_, _048510_);
  and g_137991_(_048456_, _048508_, _048511_);
  or g_137992_(_048475_, _048510_, _048512_);
  and g_137993_(_048390_, _048511_, _048513_);
  or g_137994_(_048389_, _048512_, _048514_);
  and g_137995_(_048474_, _048500_, _048515_);
  or g_137996_(_048475_, _048499_, _048516_);
  and g_137997_(_048501_, _048515_, _048517_);
  or g_137998_(_048502_, _048516_, _048518_);
  and g_137999_(_048462_, _048471_, _048519_);
  or g_138000_(_048461_, _048519_, _048521_);
  not g_138001_(_048521_, _048522_);
  and g_138002_(_048518_, _048522_, _048523_);
  or g_138003_(_048517_, _048521_, _048524_);
  and g_138004_(_048456_, _048524_, _048525_);
  or g_138005_(_048457_, _048523_, _048526_);
  and g_138006_(_048416_, _048451_, _048527_);
  or g_138007_(_048415_, _048452_, _048528_);
  and g_138008_(_048445_, _048528_, _048529_);
  or g_138009_(_048446_, _048527_, _048530_);
  and g_138010_(_048424_, _048530_, _048532_);
  or g_138011_(_048423_, _048529_, _048533_);
  and g_138012_(_048526_, _048533_, _048534_);
  or g_138013_(_048525_, _048532_, _048535_);
  and g_138014_(_048514_, _048534_, _048536_);
  or g_138015_(_048513_, _048535_, _048537_);
  and g_138016_(out[848], _048371_, _048538_);
  or g_138017_(_001484_, _048372_, _048539_);
  and g_138018_(_048353_, _048384_, _048540_);
  or g_138019_(_048354_, _048385_, _048541_);
  and g_138020_(_048539_, _048540_, _048543_);
  or g_138021_(_048538_, _048541_, _048544_);
  or g_138022_(_048379_, _048544_, _048545_);
  and g_138023_(_048511_, _048543_, _048546_);
  and g_138024_(_048378_, _048546_, _048547_);
  or g_138025_(_048512_, _048545_, _048548_);
  and g_138026_(_048537_, _048548_, _048549_);
  or g_138027_(_048536_, _048547_, _048550_);
  and g_138028_(_043360_, _048549_, _048551_);
  not g_138029_(_048551_, _048552_);
  or g_138030_(_048460_, _048549_, _048554_);
  not g_138031_(_048554_, _048555_);
  and g_138032_(_048552_, _048554_, _048556_);
  or g_138033_(_048551_, _048555_, _048557_);
  and g_138034_(_043351_, _048557_, _048558_);
  or g_138035_(_043352_, _048556_, _048559_);
  and g_138036_(_048466_, _048549_, _048560_);
  not g_138037_(_048560_, _048561_);
  or g_138038_(_048470_, _048549_, _048562_);
  not g_138039_(_048562_, _048563_);
  and g_138040_(_048561_, _048562_, _048565_);
  or g_138041_(_048560_, _048563_, _048566_);
  and g_138042_(_043348_, _048566_, _048567_);
  or g_138043_(_043347_, _048565_, _048568_);
  xor g_138044_(out[869], _043344_, _048569_);
  xor g_138045_(_001583_, _043344_, _048570_);
  or g_138046_(_048494_, _048549_, _048571_);
  not g_138047_(_048571_, _048572_);
  and g_138048_(_048489_, _048549_, _048573_);
  not g_138049_(_048573_, _048574_);
  and g_138050_(_048571_, _048574_, _048576_);
  or g_138051_(_048572_, _048573_, _048577_);
  and g_138052_(_048570_, _048576_, _048578_);
  or g_138053_(_048569_, _048577_, _048579_);
  xor g_138054_(out[866], _043341_, _048580_);
  xor g_138055_(_001627_, _043341_, _048581_);
  or g_138056_(_048349_, _048549_, _048582_);
  not g_138057_(_048582_, _048583_);
  and g_138058_(_048342_, _048549_, _048584_);
  not g_138059_(_048584_, _048585_);
  and g_138060_(_048582_, _048585_, _048587_);
  or g_138061_(_048583_, _048584_, _048588_);
  and g_138062_(_048580_, _048587_, _048589_);
  or g_138063_(_048581_, _048588_, _048590_);
  and g_138064_(_048362_, _048550_, _048591_);
  or g_138065_(_048363_, _048549_, _048592_);
  and g_138066_(_048358_, _048549_, _048593_);
  or g_138067_(_048359_, _048550_, _048594_);
  and g_138068_(_048592_, _048594_, _048595_);
  or g_138069_(_048591_, _048593_, _048596_);
  and g_138070_(out[865], _048596_, _048598_);
  not g_138071_(_048598_, _048599_);
  xor g_138072_(out[865], out[864], _048600_);
  xor g_138073_(_001605_, out[864], _048601_);
  and g_138074_(_048595_, _048600_, _048602_);
  or g_138075_(_048596_, _048601_, _048603_);
  and g_138076_(out[848], _048549_, _048604_);
  or g_138077_(_001484_, _048550_, _048605_);
  and g_138078_(_048372_, _048550_, _048606_);
  or g_138079_(_048371_, _048549_, _048607_);
  and g_138080_(_048605_, _048607_, _048609_);
  or g_138081_(_048604_, _048606_, _048610_);
  and g_138082_(out[864], _048609_, _048611_);
  or g_138083_(_001616_, _048610_, _048612_);
  and g_138084_(_048603_, _048612_, _048613_);
  or g_138085_(_048602_, _048611_, _048614_);
  and g_138086_(_048599_, _048614_, _048615_);
  or g_138087_(_048598_, _048613_, _048616_);
  and g_138088_(_048590_, _048616_, _048617_);
  or g_138089_(_048589_, _048615_, _048618_);
  and g_138090_(_048581_, _048588_, _048620_);
  or g_138091_(_048580_, _048587_, _048621_);
  xor g_138092_(out[867], _043342_, _048622_);
  xor g_138093_(_001638_, _043342_, _048623_);
  or g_138094_(_048336_, _048549_, _048624_);
  not g_138095_(_048624_, _048625_);
  and g_138096_(_043364_, _048549_, _048626_);
  not g_138097_(_048626_, _048627_);
  and g_138098_(_048624_, _048627_, _048628_);
  or g_138099_(_048625_, _048626_, _048629_);
  and g_138100_(_048622_, _048629_, _048631_);
  or g_138101_(_048623_, _048628_, _048632_);
  and g_138102_(_048621_, _048632_, _048633_);
  or g_138103_(_048620_, _048631_, _048634_);
  and g_138104_(_048618_, _048633_, _048635_);
  or g_138105_(_048617_, _048634_, _048636_);
  and g_138106_(_048623_, _048628_, _048637_);
  or g_138107_(_048622_, _048629_, _048638_);
  xor g_138108_(out[868], _043343_, _048639_);
  xor g_138109_(_001594_, _043343_, _048640_);
  and g_138110_(_048478_, _048549_, _048642_);
  not g_138111_(_048642_, _048643_);
  or g_138112_(_048483_, _048549_, _048644_);
  not g_138113_(_048644_, _048645_);
  and g_138114_(_048643_, _048644_, _048646_);
  or g_138115_(_048642_, _048645_, _048647_);
  and g_138116_(_048640_, _048646_, _048648_);
  or g_138117_(_048639_, _048647_, _048649_);
  and g_138118_(_048638_, _048649_, _048650_);
  or g_138119_(_048637_, _048648_, _048651_);
  and g_138120_(_048636_, _048650_, _048653_);
  or g_138121_(_048635_, _048651_, _048654_);
  and g_138122_(_048569_, _048577_, _048655_);
  or g_138123_(_048570_, _048576_, _048656_);
  and g_138124_(_048639_, _048647_, _048657_);
  or g_138125_(_048640_, _048646_, _048658_);
  and g_138126_(_048656_, _048658_, _048659_);
  or g_138127_(_048655_, _048657_, _048660_);
  and g_138128_(_048654_, _048659_, _048661_);
  or g_138129_(_048653_, _048660_, _048662_);
  and g_138130_(_048579_, _048662_, _048664_);
  or g_138131_(_048578_, _048661_, _048665_);
  and g_138132_(_048568_, _048665_, _048666_);
  or g_138133_(_048567_, _048664_, _048667_);
  and g_138134_(_043352_, _048556_, _048668_);
  or g_138135_(_043351_, _048557_, _048669_);
  and g_138136_(_043347_, _048565_, _048670_);
  or g_138137_(_043348_, _048566_, _048671_);
  and g_138138_(_048669_, _048671_, _048672_);
  or g_138139_(_048668_, _048670_, _048673_);
  and g_138140_(_048667_, _048672_, _048675_);
  or g_138141_(_048666_, _048673_, _048676_);
  and g_138142_(_048559_, _048676_, _048677_);
  or g_138143_(_048558_, _048675_, _048678_);
  and g_138144_(_048433_, _048549_, _048679_);
  not g_138145_(_048679_, _048680_);
  or g_138146_(_048438_, _048549_, _048681_);
  not g_138147_(_048681_, _048682_);
  and g_138148_(_048680_, _048681_, _048683_);
  or g_138149_(_048679_, _048682_, _048684_);
  and g_138150_(out[872], _043349_, _048686_);
  or g_138151_(out[873], _048686_, _048687_);
  and g_138152_(out[874], _048687_, _048688_);
  xor g_138153_(out[874], _048687_, _048689_);
  and g_138154_(_048684_, _048689_, _048690_);
  xor g_138155_(out[875], _048688_, _048691_);
  xor g_138156_(_001550_, _048688_, _048692_);
  and g_138157_(_048419_, _048549_, _048693_);
  not g_138158_(_048693_, _048694_);
  or g_138159_(_048420_, _048549_, _048695_);
  not g_138160_(_048695_, _048697_);
  and g_138161_(_048694_, _048695_, _048698_);
  or g_138162_(_048693_, _048697_, _048699_);
  or g_138163_(_048422_, _048549_, _048700_);
  not g_138164_(_048700_, _048701_);
  and g_138165_(_048418_, _048549_, _048702_);
  not g_138166_(_048702_, _048703_);
  and g_138167_(_048700_, _048703_, _048704_);
  or g_138168_(_048701_, _048702_, _048705_);
  and g_138169_(_048691_, _048704_, _048706_);
  or g_138170_(_048691_, _048699_, _048708_);
  xor g_138171_(_048684_, _048689_, _048709_);
  xor g_138172_(_048683_, _048689_, _048710_);
  xor g_138173_(_048691_, _048704_, _048711_);
  xor g_138174_(_048692_, _048704_, _048712_);
  and g_138175_(_048709_, _048711_, _048713_);
  or g_138176_(_048710_, _048712_, _048714_);
  xor g_138177_(out[873], _048686_, _048715_);
  xor g_138178_(_001660_, _048686_, _048716_);
  and g_138179_(_048393_, _048549_, _048717_);
  not g_138180_(_048717_, _048719_);
  or g_138181_(_048400_, _048549_, _048720_);
  not g_138182_(_048720_, _048721_);
  and g_138183_(_048719_, _048720_, _048722_);
  or g_138184_(_048717_, _048721_, _048723_);
  and g_138185_(_048716_, _048723_, _048724_);
  or g_138186_(_048715_, _048722_, _048725_);
  xor g_138187_(out[872], _043349_, _048726_);
  xor g_138188_(_001649_, _043349_, _048727_);
  and g_138189_(_048405_, _048549_, _048728_);
  not g_138190_(_048728_, _048730_);
  or g_138191_(_048411_, _048549_, _048731_);
  not g_138192_(_048731_, _048732_);
  and g_138193_(_048730_, _048731_, _048733_);
  or g_138194_(_048728_, _048732_, _048734_);
  and g_138195_(_048726_, _048734_, _048735_);
  or g_138196_(_048727_, _048733_, _048736_);
  and g_138197_(_048725_, _048736_, _048737_);
  or g_138198_(_048724_, _048735_, _048738_);
  and g_138199_(_048715_, _048722_, _048739_);
  or g_138200_(_048716_, _048723_, _048741_);
  and g_138201_(_048727_, _048733_, _048742_);
  or g_138202_(_048726_, _048734_, _048743_);
  and g_138203_(_048741_, _048743_, _048744_);
  or g_138204_(_048739_, _048742_, _048745_);
  and g_138205_(_048737_, _048744_, _048746_);
  or g_138206_(_048738_, _048745_, _048747_);
  and g_138207_(_048713_, _048746_, _048748_);
  or g_138208_(_048714_, _048747_, _048749_);
  and g_138209_(_048678_, _048748_, _048750_);
  or g_138210_(_048677_, _048749_, _048752_);
  and g_138211_(_048713_, _048738_, _048753_);
  or g_138212_(_048714_, _048737_, _048754_);
  and g_138213_(_048741_, _048753_, _048755_);
  or g_138214_(_048739_, _048754_, _048756_);
  and g_138215_(_048690_, _048708_, _048757_);
  or g_138216_(_048706_, _048757_, _048758_);
  not g_138217_(_048758_, _048759_);
  and g_138218_(_048756_, _048759_, _048760_);
  or g_138219_(_048755_, _048758_, _048761_);
  and g_138220_(_048752_, _048760_, _048763_);
  or g_138221_(_048750_, _048761_, _048764_);
  or g_138222_(_043348_, _048764_, _048765_);
  not g_138223_(_048765_, _048766_);
  and g_138224_(_048566_, _048764_, _048767_);
  not g_138225_(_048767_, _048768_);
  and g_138226_(_048765_, _048768_, _048769_);
  or g_138227_(_048766_, _048767_, _048770_);
  or g_138228_(out[881], out[880], _048771_);
  or g_138229_(out[880], _002075_, _048772_);
  and g_138230_(out[883], _048772_, _048774_);
  and g_138231_(_026535_, _048772_, _048775_);
  and g_138232_(out[885], _048775_, _048776_);
  or g_138233_(out[886], _048776_, _048777_);
  and g_138234_(out[887], _048777_, _048778_);
  xor g_138235_(out[887], _048777_, _048779_);
  xor g_138236_(_001693_, _048777_, _048780_);
  or g_138237_(_043351_, _048764_, _048781_);
  not g_138238_(_048781_, _048782_);
  and g_138239_(_048557_, _048764_, _048783_);
  not g_138240_(_048783_, _048785_);
  and g_138241_(_048781_, _048785_, _048786_);
  or g_138242_(_048782_, _048783_, _048787_);
  and g_138243_(_048779_, _048787_, _048788_);
  or g_138244_(_048780_, _048786_, _048789_);
  xor g_138245_(out[886], _048776_, _048790_);
  xor g_138246_(_001704_, _048776_, _048791_);
  and g_138247_(_048770_, _048791_, _048792_);
  or g_138248_(_048769_, _048790_, _048793_);
  xor g_138249_(out[885], _048775_, _048794_);
  xor g_138250_(_001715_, _048775_, _048796_);
  and g_138251_(_048577_, _048764_, _048797_);
  not g_138252_(_048797_, _048798_);
  or g_138253_(_048569_, _048764_, _048799_);
  not g_138254_(_048799_, _048800_);
  and g_138255_(_048798_, _048799_, _048801_);
  or g_138256_(_048797_, _048800_, _048802_);
  and g_138257_(_048796_, _048801_, _048803_);
  or g_138258_(_048794_, _048802_, _048804_);
  and g_138259_(out[864], _048763_, _048805_);
  or g_138260_(_001616_, _048764_, _048807_);
  and g_138261_(_048610_, _048764_, _048808_);
  or g_138262_(_048609_, _048763_, _048809_);
  and g_138263_(_048807_, _048809_, _048810_);
  or g_138264_(_048805_, _048808_, _048811_);
  and g_138265_(out[880], _048810_, _048812_);
  or g_138266_(_001748_, _048811_, _048813_);
  and g_138267_(_048600_, _048763_, _048814_);
  or g_138268_(_048601_, _048764_, _048815_);
  and g_138269_(_048596_, _048764_, _048816_);
  or g_138270_(_048595_, _048763_, _048818_);
  and g_138271_(_048815_, _048818_, _048819_);
  or g_138272_(_048814_, _048816_, _048820_);
  and g_138273_(out[881], _048820_, _048821_);
  or g_138274_(_001737_, _048819_, _048822_);
  xor g_138275_(out[881], out[880], _048823_);
  xor g_138276_(_001737_, out[880], _048824_);
  and g_138277_(_048812_, _048822_, _048825_);
  or g_138278_(_048813_, _048821_, _048826_);
  xor g_138279_(out[882], _048771_, _048827_);
  xor g_138280_(_001759_, _048771_, _048829_);
  and g_138281_(_048588_, _048764_, _048830_);
  or g_138282_(_048587_, _048763_, _048831_);
  and g_138283_(_048580_, _048763_, _048832_);
  or g_138284_(_048581_, _048764_, _048833_);
  and g_138285_(_048831_, _048833_, _048834_);
  or g_138286_(_048830_, _048832_, _048835_);
  and g_138287_(_048827_, _048834_, _048836_);
  or g_138288_(_048829_, _048835_, _048837_);
  and g_138289_(_048819_, _048823_, _048838_);
  or g_138290_(_048820_, _048824_, _048840_);
  and g_138291_(_048837_, _048840_, _048841_);
  or g_138292_(_048836_, _048838_, _048842_);
  and g_138293_(_048826_, _048841_, _048843_);
  or g_138294_(_048825_, _048842_, _048844_);
  xor g_138295_(out[883], _048772_, _048845_);
  xor g_138296_(_001770_, _048772_, _048846_);
  or g_138297_(_048622_, _048764_, _048847_);
  not g_138298_(_048847_, _048848_);
  and g_138299_(_048629_, _048764_, _048849_);
  not g_138300_(_048849_, _048851_);
  and g_138301_(_048847_, _048851_, _048852_);
  or g_138302_(_048848_, _048849_, _048853_);
  and g_138303_(_048845_, _048853_, _048854_);
  or g_138304_(_048846_, _048852_, _048855_);
  and g_138305_(_048829_, _048835_, _048856_);
  or g_138306_(_048827_, _048834_, _048857_);
  and g_138307_(_048855_, _048857_, _048858_);
  or g_138308_(_048854_, _048856_, _048859_);
  and g_138309_(_048844_, _048858_, _048860_);
  or g_138310_(_048843_, _048859_, _048862_);
  xor g_138311_(out[884], _048774_, _048863_);
  xor g_138312_(_001726_, _048774_, _048864_);
  and g_138313_(_048647_, _048764_, _048865_);
  not g_138314_(_048865_, _048866_);
  or g_138315_(_048639_, _048764_, _048867_);
  not g_138316_(_048867_, _048868_);
  and g_138317_(_048866_, _048867_, _048869_);
  or g_138318_(_048865_, _048868_, _048870_);
  and g_138319_(_048864_, _048869_, _048871_);
  or g_138320_(_048863_, _048870_, _048873_);
  and g_138321_(_048846_, _048852_, _048874_);
  or g_138322_(_048845_, _048853_, _048875_);
  and g_138323_(_048873_, _048875_, _048876_);
  or g_138324_(_048871_, _048874_, _048877_);
  and g_138325_(_048862_, _048876_, _048878_);
  or g_138326_(_048860_, _048877_, _048879_);
  and g_138327_(_048794_, _048802_, _048880_);
  or g_138328_(_048796_, _048801_, _048881_);
  and g_138329_(_048863_, _048870_, _048882_);
  or g_138330_(_048864_, _048869_, _048884_);
  and g_138331_(_048881_, _048884_, _048885_);
  or g_138332_(_048880_, _048882_, _048886_);
  and g_138333_(_048879_, _048885_, _048887_);
  or g_138334_(_048878_, _048886_, _048888_);
  and g_138335_(_048804_, _048888_, _048889_);
  or g_138336_(_048803_, _048887_, _048890_);
  and g_138337_(_048793_, _048890_, _048891_);
  or g_138338_(_048792_, _048889_, _048892_);
  and g_138339_(_048780_, _048786_, _048893_);
  or g_138340_(_048779_, _048787_, _048895_);
  and g_138341_(_048769_, _048790_, _048896_);
  or g_138342_(_048770_, _048791_, _048897_);
  and g_138343_(_048895_, _048897_, _048898_);
  or g_138344_(_048893_, _048896_, _048899_);
  and g_138345_(_048892_, _048898_, _048900_);
  or g_138346_(_048891_, _048899_, _048901_);
  and g_138347_(_048789_, _048901_, _048902_);
  or g_138348_(_048788_, _048900_, _048903_);
  and g_138349_(out[888], _048778_, _048904_);
  or g_138350_(out[889], _048904_, _048906_);
  and g_138351_(out[890], _048906_, _048907_);
  xor g_138352_(out[890], _048906_, _048908_);
  xor g_138353_(_001803_, _048906_, _048909_);
  or g_138354_(_048689_, _048764_, _048910_);
  not g_138355_(_048910_, _048911_);
  and g_138356_(_048684_, _048764_, _048912_);
  not g_138357_(_048912_, _048913_);
  and g_138358_(_048910_, _048913_, _048914_);
  or g_138359_(_048911_, _048912_, _048915_);
  and g_138360_(_048908_, _048915_, _048917_);
  or g_138361_(_048909_, _048914_, _048918_);
  xor g_138362_(out[891], _048907_, _048919_);
  xor g_138363_(_001682_, _048907_, _048920_);
  and g_138364_(_048691_, _048698_, _048921_);
  or g_138365_(_048692_, _048699_, _048922_);
  and g_138366_(_048691_, _048705_, _048923_);
  and g_138367_(_048919_, _048922_, _048924_);
  or g_138368_(_048920_, _048923_, _048925_);
  and g_138369_(_048918_, _048925_, _048926_);
  or g_138370_(_048917_, _048924_, _048928_);
  and g_138371_(_048909_, _048914_, _048929_);
  or g_138372_(_048908_, _048915_, _048930_);
  and g_138373_(_048920_, _048921_, _048931_);
  or g_138374_(_048919_, _048922_, _048932_);
  and g_138375_(_048930_, _048932_, _048933_);
  or g_138376_(_048929_, _048931_, _048934_);
  and g_138377_(_048926_, _048933_, _048935_);
  or g_138378_(_048928_, _048934_, _048936_);
  xor g_138379_(out[889], _048904_, _048937_);
  not g_138380_(_048937_, _048939_);
  or g_138381_(_048716_, _048764_, _048940_);
  not g_138382_(_048940_, _048941_);
  and g_138383_(_048723_, _048764_, _048942_);
  not g_138384_(_048942_, _048943_);
  and g_138385_(_048940_, _048943_, _048944_);
  or g_138386_(_048941_, _048942_, _048945_);
  and g_138387_(_048937_, _048944_, _048946_);
  or g_138388_(_048939_, _048945_, _048947_);
  xor g_138389_(out[888], _048778_, _048948_);
  not g_138390_(_048948_, _048950_);
  or g_138391_(_048726_, _048764_, _048951_);
  not g_138392_(_048951_, _048952_);
  and g_138393_(_048734_, _048764_, _048953_);
  not g_138394_(_048953_, _048954_);
  and g_138395_(_048951_, _048954_, _048955_);
  or g_138396_(_048952_, _048953_, _048956_);
  and g_138397_(_048950_, _048955_, _048957_);
  or g_138398_(_048948_, _048956_, _048958_);
  and g_138399_(_048947_, _048958_, _048959_);
  or g_138400_(_048946_, _048957_, _048961_);
  and g_138401_(_048939_, _048945_, _048962_);
  or g_138402_(_048937_, _048944_, _048963_);
  and g_138403_(_048948_, _048956_, _048964_);
  or g_138404_(_048950_, _048955_, _048965_);
  and g_138405_(_048963_, _048965_, _048966_);
  or g_138406_(_048962_, _048964_, _048967_);
  and g_138407_(_048959_, _048966_, _048968_);
  or g_138408_(_048961_, _048967_, _048969_);
  and g_138409_(_048935_, _048968_, _048970_);
  or g_138410_(_048936_, _048969_, _048972_);
  and g_138411_(_048903_, _048970_, _048973_);
  or g_138412_(_048902_, _048972_, _048974_);
  and g_138413_(_048947_, _048967_, _048975_);
  or g_138414_(_048946_, _048966_, _048976_);
  and g_138415_(_048935_, _048975_, _048977_);
  or g_138416_(_048936_, _048976_, _048978_);
  and g_138417_(_048928_, _048932_, _048979_);
  or g_138418_(_048926_, _048931_, _048980_);
  and g_138419_(_048978_, _048980_, _048981_);
  or g_138420_(_048977_, _048979_, _048983_);
  and g_138421_(_048974_, _048981_, _048984_);
  or g_138422_(_048973_, _048983_, _048985_);
  and g_138423_(_048770_, _048985_, _048986_);
  not g_138424_(_048986_, _048987_);
  or g_138425_(_048791_, _048985_, _048988_);
  not g_138426_(_048988_, _048989_);
  and g_138427_(_048987_, _048988_, _048990_);
  or g_138428_(_048986_, _048989_, _048991_);
  and g_138429_(out[880], _048984_, _048992_);
  or g_138430_(_001748_, _048985_, _048994_);
  and g_138431_(_048811_, _048985_, _048995_);
  or g_138432_(_048810_, _048984_, _048996_);
  and g_138433_(_048994_, _048996_, _048997_);
  or g_138434_(_048992_, _048995_, _048998_);
  and g_138435_(out[896], _048997_, _048999_);
  or g_138436_(_001880_, _048998_, _049000_);
  and g_138437_(_048823_, _048984_, _049001_);
  or g_138438_(_048824_, _048985_, _049002_);
  and g_138439_(_048820_, _048985_, _049003_);
  or g_138440_(_048819_, _048984_, _049005_);
  and g_138441_(_049002_, _049005_, _049006_);
  or g_138442_(_049001_, _049003_, _049007_);
  and g_138443_(out[897], _049007_, _049008_);
  or g_138444_(_001869_, _049006_, _049009_);
  or g_138445_(out[897], out[896], _049010_);
  xor g_138446_(_001869_, out[896], _049011_);
  not g_138447_(_049011_, _049012_);
  and g_138448_(_048999_, _049009_, _049013_);
  or g_138449_(_049000_, _049008_, _049014_);
  or g_138450_(out[896], _002332_, _049016_);
  xor g_138451_(out[898], _049010_, _049017_);
  xor g_138452_(_001891_, _049010_, _049018_);
  and g_138453_(_048827_, _048984_, _049019_);
  or g_138454_(_048829_, _048985_, _049020_);
  and g_138455_(_048835_, _048985_, _049021_);
  or g_138456_(_048834_, _048984_, _049022_);
  and g_138457_(_049020_, _049022_, _049023_);
  or g_138458_(_049019_, _049021_, _049024_);
  and g_138459_(_049017_, _049023_, _049025_);
  or g_138460_(_049018_, _049024_, _049027_);
  and g_138461_(_049006_, _049012_, _049028_);
  or g_138462_(_049007_, _049011_, _049029_);
  and g_138463_(_049027_, _049029_, _049030_);
  or g_138464_(_049025_, _049028_, _049031_);
  and g_138465_(_049014_, _049030_, _049032_);
  or g_138466_(_049013_, _049031_, _049033_);
  and g_138467_(out[899], _049016_, _049034_);
  xor g_138468_(out[899], _049016_, _049035_);
  xor g_138469_(_001902_, _049016_, _049036_);
  or g_138470_(_048845_, _048985_, _049038_);
  not g_138471_(_049038_, _049039_);
  and g_138472_(_048853_, _048985_, _049040_);
  not g_138473_(_049040_, _049041_);
  and g_138474_(_049038_, _049041_, _049042_);
  or g_138475_(_049039_, _049040_, _049043_);
  and g_138476_(_049035_, _049043_, _049044_);
  or g_138477_(_049036_, _049042_, _049045_);
  and g_138478_(_049018_, _049024_, _049046_);
  or g_138479_(_049017_, _049023_, _049047_);
  and g_138480_(_049045_, _049047_, _049049_);
  or g_138481_(_049044_, _049046_, _049050_);
  and g_138482_(_049033_, _049049_, _049051_);
  or g_138483_(_049032_, _049050_, _049052_);
  and g_138484_(_026777_, _049016_, _049053_);
  xor g_138485_(out[900], _049034_, _049054_);
  xor g_138486_(_001858_, _049034_, _049055_);
  or g_138487_(_048863_, _048985_, _049056_);
  not g_138488_(_049056_, _049057_);
  and g_138489_(_048870_, _048985_, _049058_);
  not g_138490_(_049058_, _049060_);
  and g_138491_(_049056_, _049060_, _049061_);
  or g_138492_(_049057_, _049058_, _049062_);
  and g_138493_(_049055_, _049061_, _049063_);
  or g_138494_(_049054_, _049062_, _049064_);
  and g_138495_(_049036_, _049042_, _049065_);
  or g_138496_(_049035_, _049043_, _049066_);
  and g_138497_(_049064_, _049066_, _049067_);
  or g_138498_(_049063_, _049065_, _049068_);
  and g_138499_(_049052_, _049067_, _049069_);
  or g_138500_(_049051_, _049068_, _049071_);
  and g_138501_(out[901], _049053_, _049072_);
  xor g_138502_(out[901], _049053_, _049073_);
  xor g_138503_(_001847_, _049053_, _049074_);
  or g_138504_(_048794_, _048985_, _049075_);
  not g_138505_(_049075_, _049076_);
  and g_138506_(_048802_, _048985_, _049077_);
  not g_138507_(_049077_, _049078_);
  and g_138508_(_049075_, _049078_, _049079_);
  or g_138509_(_049076_, _049077_, _049080_);
  and g_138510_(_049073_, _049080_, _049082_);
  or g_138511_(_049074_, _049079_, _049083_);
  and g_138512_(_049054_, _049062_, _049084_);
  or g_138513_(_049055_, _049061_, _049085_);
  and g_138514_(_049083_, _049085_, _049086_);
  or g_138515_(_049082_, _049084_, _049087_);
  and g_138516_(_049071_, _049086_, _049088_);
  or g_138517_(_049069_, _049087_, _049089_);
  or g_138518_(out[902], _049072_, _049090_);
  xor g_138519_(out[902], _049072_, _049091_);
  xor g_138520_(_001836_, _049072_, _049093_);
  and g_138521_(_048990_, _049091_, _049094_);
  or g_138522_(_048991_, _049093_, _049095_);
  and g_138523_(_049074_, _049079_, _049096_);
  or g_138524_(_049073_, _049080_, _049097_);
  and g_138525_(_049095_, _049097_, _049098_);
  or g_138526_(_049094_, _049096_, _049099_);
  and g_138527_(_049089_, _049098_, _049100_);
  or g_138528_(_049088_, _049099_, _049101_);
  and g_138529_(out[903], _049090_, _049102_);
  xor g_138530_(out[903], _049090_, _049104_);
  xor g_138531_(_001825_, _049090_, _049105_);
  and g_138532_(_048787_, _048985_, _049106_);
  not g_138533_(_049106_, _049107_);
  or g_138534_(_048779_, _048985_, _049108_);
  not g_138535_(_049108_, _049109_);
  and g_138536_(_049107_, _049108_, _049110_);
  or g_138537_(_049106_, _049109_, _049111_);
  and g_138538_(_049104_, _049111_, _049112_);
  or g_138539_(_049105_, _049110_, _049113_);
  and g_138540_(_048991_, _049093_, _049115_);
  or g_138541_(_048990_, _049091_, _049116_);
  and g_138542_(_049113_, _049116_, _049117_);
  or g_138543_(_049112_, _049115_, _049118_);
  and g_138544_(_049101_, _049117_, _049119_);
  or g_138545_(_049100_, _049118_, _049120_);
  and g_138546_(out[904], _049102_, _049121_);
  or g_138547_(out[905], _049121_, _049122_);
  and g_138548_(out[906], _049122_, _049123_);
  xor g_138549_(out[906], _049122_, _049124_);
  xor g_138550_(_001935_, _049122_, _049126_);
  and g_138551_(_048915_, _048985_, _049127_);
  not g_138552_(_049127_, _049128_);
  or g_138553_(_048908_, _048985_, _049129_);
  not g_138554_(_049129_, _049130_);
  and g_138555_(_049128_, _049129_, _049131_);
  or g_138556_(_049127_, _049130_, _049132_);
  and g_138557_(_049126_, _049131_, _049133_);
  or g_138558_(_049124_, _049132_, _049134_);
  xor g_138559_(out[905], _049121_, _049135_);
  xor g_138560_(_001924_, _049121_, _049137_);
  and g_138561_(_048945_, _048985_, _049138_);
  not g_138562_(_049138_, _049139_);
  or g_138563_(_048939_, _048985_, _049140_);
  not g_138564_(_049140_, _049141_);
  and g_138565_(_049139_, _049140_, _049142_);
  or g_138566_(_049138_, _049141_, _049143_);
  and g_138567_(_049137_, _049143_, _049144_);
  or g_138568_(_049135_, _049142_, _049145_);
  xor g_138569_(out[904], _049102_, _049146_);
  xor g_138570_(_001913_, _049102_, _049148_);
  and g_138571_(_048956_, _048985_, _049149_);
  not g_138572_(_049149_, _049150_);
  or g_138573_(_048948_, _048985_, _049151_);
  not g_138574_(_049151_, _049152_);
  and g_138575_(_049150_, _049151_, _049153_);
  or g_138576_(_049149_, _049152_, _049154_);
  and g_138577_(_049148_, _049153_, _049155_);
  or g_138578_(_049146_, _049154_, _049156_);
  and g_138579_(_049145_, _049156_, _049157_);
  or g_138580_(_049144_, _049155_, _049159_);
  and g_138581_(_049134_, _049157_, _049160_);
  or g_138582_(_049133_, _049159_, _049161_);
  and g_138583_(_049124_, _049132_, _049162_);
  or g_138584_(_049126_, _049131_, _049163_);
  xor g_138585_(out[907], _049123_, _049164_);
  xor g_138586_(_001814_, _049123_, _049165_);
  and g_138587_(_048919_, _048921_, _049166_);
  or g_138588_(_048920_, _048922_, _049167_);
  and g_138589_(_048919_, _048923_, _049168_);
  and g_138590_(_049164_, _049167_, _049170_);
  or g_138591_(_049165_, _049168_, _049171_);
  and g_138592_(_049163_, _049171_, _049172_);
  or g_138593_(_049162_, _049170_, _049173_);
  and g_138594_(_049135_, _049142_, _049174_);
  or g_138595_(_049137_, _049143_, _049175_);
  and g_138596_(_049146_, _049154_, _049176_);
  or g_138597_(_049148_, _049153_, _049177_);
  and g_138598_(_049175_, _049177_, _049178_);
  or g_138599_(_049174_, _049176_, _049179_);
  and g_138600_(_049165_, _049166_, _049181_);
  or g_138601_(_049164_, _049167_, _049182_);
  and g_138602_(_049105_, _049110_, _049183_);
  or g_138603_(_049104_, _049111_, _049184_);
  and g_138604_(_049182_, _049184_, _049185_);
  or g_138605_(_049181_, _049183_, _049186_);
  and g_138606_(_049178_, _049185_, _049187_);
  or g_138607_(_049179_, _049186_, _049188_);
  and g_138608_(_049172_, _049187_, _049189_);
  or g_138609_(_049173_, _049188_, _049190_);
  and g_138610_(_049160_, _049189_, _049192_);
  or g_138611_(_049161_, _049190_, _049193_);
  and g_138612_(_049120_, _049192_, _049194_);
  or g_138613_(_049119_, _049193_, _049195_);
  and g_138614_(_049175_, _049176_, _049196_);
  or g_138615_(_049174_, _049177_, _049197_);
  and g_138616_(_049145_, _049197_, _049198_);
  or g_138617_(_049144_, _049196_, _049199_);
  and g_138618_(_049134_, _049199_, _049200_);
  or g_138619_(_049133_, _049198_, _049201_);
  and g_138620_(_049172_, _049201_, _049203_);
  or g_138621_(_049173_, _049200_, _049204_);
  and g_138622_(_049182_, _049204_, _049205_);
  or g_138623_(_049181_, _049203_, _049206_);
  and g_138624_(_049195_, _049206_, _049207_);
  or g_138625_(_049194_, _049205_, _049208_);
  and g_138626_(_048991_, _049208_, _049209_);
  or g_138627_(_048990_, _049207_, _049210_);
  and g_138628_(_049091_, _049207_, _049211_);
  or g_138629_(_049093_, _049208_, _049212_);
  and g_138630_(_049210_, _049212_, _049214_);
  or g_138631_(_049209_, _049211_, _049215_);
  or g_138632_(out[913], out[912], _049216_);
  or g_138633_(out[912], _002528_, _049217_);
  and g_138634_(out[915], _049217_, _049218_);
  and g_138635_(_026932_, _049217_, _049219_);
  and g_138636_(out[917], _049219_, _049220_);
  or g_138637_(out[918], _049220_, _049221_);
  and g_138638_(out[919], _049221_, _049222_);
  and g_138639_(out[920], _049222_, _049223_);
  or g_138640_(out[921], _049223_, _049225_);
  and g_138641_(out[922], _049225_, _049226_);
  xor g_138642_(out[923], _049226_, _049227_);
  not g_138643_(_049227_, _049228_);
  and g_138644_(_049164_, _049166_, _049229_);
  not g_138645_(_049229_, _049230_);
  and g_138646_(_049164_, _049168_, _049231_);
  and g_138647_(_049227_, _049230_, _049232_);
  or g_138648_(_049228_, _049229_, _049233_);
  and g_138649_(_049228_, _049229_, _049234_);
  or g_138650_(_049227_, _049230_, _049236_);
  xor g_138651_(out[922], _049225_, _049237_);
  xor g_138652_(_002067_, _049225_, _049238_);
  or g_138653_(_049131_, _049207_, _049239_);
  not g_138654_(_049239_, _049240_);
  and g_138655_(_049126_, _049207_, _049241_);
  not g_138656_(_049241_, _049242_);
  and g_138657_(_049239_, _049242_, _049243_);
  or g_138658_(_049240_, _049241_, _049244_);
  and g_138659_(_049238_, _049243_, _049245_);
  or g_138660_(_049237_, _049244_, _049247_);
  and g_138661_(_049236_, _049247_, _049248_);
  or g_138662_(_049234_, _049245_, _049249_);
  and g_138663_(_049233_, _049249_, _049250_);
  or g_138664_(_049232_, _049248_, _049251_);
  xor g_138665_(out[921], _049223_, _049252_);
  not g_138666_(_049252_, _049253_);
  and g_138667_(_049143_, _049208_, _049254_);
  and g_138668_(_049135_, _049207_, _049255_);
  or g_138669_(_049254_, _049255_, _049256_);
  not g_138670_(_049256_, _049258_);
  and g_138671_(_049252_, _049258_, _049259_);
  or g_138672_(_049253_, _049256_, _049260_);
  xor g_138673_(out[920], _049222_, _049261_);
  not g_138674_(_049261_, _049262_);
  or g_138675_(_049153_, _049207_, _049263_);
  or g_138676_(_049146_, _049208_, _049264_);
  and g_138677_(_049263_, _049264_, _049265_);
  not g_138678_(_049265_, _049266_);
  and g_138679_(_049262_, _049265_, _049267_);
  or g_138680_(_049261_, _049266_, _049269_);
  and g_138681_(_049260_, _049269_, _049270_);
  or g_138682_(_049259_, _049267_, _049271_);
  and g_138683_(_049253_, _049256_, _049272_);
  or g_138684_(_049252_, _049258_, _049273_);
  and g_138685_(_049261_, _049266_, _049274_);
  or g_138686_(_049262_, _049265_, _049275_);
  and g_138687_(_049273_, _049275_, _049276_);
  or g_138688_(_049272_, _049274_, _049277_);
  and g_138689_(_049270_, _049276_, _049278_);
  or g_138690_(_049271_, _049277_, _049280_);
  xor g_138691_(out[918], _049220_, _049281_);
  not g_138692_(_049281_, _049282_);
  and g_138693_(_049214_, _049281_, _049283_);
  or g_138694_(_049215_, _049282_, _049284_);
  xor g_138695_(out[919], _049221_, _049285_);
  xor g_138696_(_001957_, _049221_, _049286_);
  and g_138697_(_049111_, _049208_, _049287_);
  or g_138698_(_049110_, _049207_, _049288_);
  and g_138699_(_049105_, _049207_, _049289_);
  or g_138700_(_049104_, _049208_, _049291_);
  and g_138701_(_049288_, _049291_, _049292_);
  or g_138702_(_049287_, _049289_, _049293_);
  and g_138703_(_049286_, _049292_, _049294_);
  or g_138704_(_049285_, _049293_, _049295_);
  and g_138705_(_049284_, _049295_, _049296_);
  or g_138706_(_049283_, _049294_, _049297_);
  and g_138707_(_049285_, _049293_, _049298_);
  or g_138708_(_049286_, _049292_, _049299_);
  and g_138709_(_049215_, _049282_, _049300_);
  or g_138710_(_049214_, _049281_, _049302_);
  and g_138711_(_049299_, _049302_, _049303_);
  or g_138712_(_049298_, _049300_, _049304_);
  xor g_138713_(out[917], _049219_, _049305_);
  xor g_138714_(_001979_, _049219_, _049306_);
  and g_138715_(_049074_, _049207_, _049307_);
  not g_138716_(_049307_, _049308_);
  or g_138717_(_049079_, _049207_, _049309_);
  not g_138718_(_049309_, _049310_);
  and g_138719_(_049308_, _049309_, _049311_);
  or g_138720_(_049307_, _049310_, _049313_);
  and g_138721_(_049305_, _049313_, _049314_);
  or g_138722_(_049306_, _049311_, _049315_);
  and g_138723_(_049296_, _049303_, _049316_);
  or g_138724_(_049297_, _049304_, _049317_);
  and g_138725_(_049315_, _049316_, _049318_);
  or g_138726_(_049314_, _049317_, _049319_);
  and g_138727_(_049306_, _049311_, _049320_);
  or g_138728_(_049305_, _049313_, _049321_);
  xor g_138729_(out[916], _049218_, _049322_);
  xor g_138730_(_001990_, _049218_, _049324_);
  or g_138731_(_049061_, _049207_, _049325_);
  not g_138732_(_049325_, _049326_);
  and g_138733_(_049055_, _049207_, _049327_);
  not g_138734_(_049327_, _049328_);
  and g_138735_(_049325_, _049328_, _049329_);
  or g_138736_(_049326_, _049327_, _049330_);
  and g_138737_(_049324_, _049329_, _049331_);
  or g_138738_(_049322_, _049330_, _049332_);
  and g_138739_(_049321_, _049332_, _049333_);
  or g_138740_(_049320_, _049331_, _049335_);
  and g_138741_(_049322_, _049330_, _049336_);
  or g_138742_(_049324_, _049329_, _049337_);
  and g_138743_(_049333_, _049337_, _049338_);
  or g_138744_(_049335_, _049336_, _049339_);
  and g_138745_(_049318_, _049338_, _049340_);
  or g_138746_(_049319_, _049339_, _049341_);
  xor g_138747_(out[914], _049216_, _049342_);
  not g_138748_(_049342_, _049343_);
  or g_138749_(_049023_, _049207_, _049344_);
  not g_138750_(_049344_, _049346_);
  and g_138751_(_049017_, _049207_, _049347_);
  not g_138752_(_049347_, _049348_);
  and g_138753_(_049344_, _049348_, _049349_);
  or g_138754_(_049346_, _049347_, _049350_);
  and g_138755_(_049342_, _049349_, _049351_);
  or g_138756_(_049343_, _049350_, _049352_);
  xor g_138757_(out[915], _049217_, _049353_);
  xor g_138758_(_002034_, _049217_, _049354_);
  and g_138759_(_049036_, _049207_, _049355_);
  not g_138760_(_049355_, _049357_);
  or g_138761_(_049042_, _049207_, _049358_);
  not g_138762_(_049358_, _049359_);
  and g_138763_(_049357_, _049358_, _049360_);
  or g_138764_(_049355_, _049359_, _049361_);
  and g_138765_(_049354_, _049360_, _049362_);
  or g_138766_(_049353_, _049361_, _049363_);
  and g_138767_(_049352_, _049363_, _049364_);
  or g_138768_(_049351_, _049362_, _049365_);
  and g_138769_(_049353_, _049361_, _049366_);
  or g_138770_(_049354_, _049360_, _049368_);
  xor g_138771_(_049342_, _049349_, _049369_);
  xor g_138772_(_049343_, _049349_, _049370_);
  xor g_138773_(_049354_, _049360_, _049371_);
  xor g_138774_(_049353_, _049360_, _049372_);
  and g_138775_(_049369_, _049371_, _049373_);
  or g_138776_(_049370_, _049372_, _049374_);
  xor g_138777_(out[913], out[912], _049375_);
  not g_138778_(_049375_, _049376_);
  or g_138779_(_049011_, _049208_, _049377_);
  or g_138780_(_049006_, _049207_, _049379_);
  and g_138781_(_049377_, _049379_, _049380_);
  not g_138782_(_049380_, _049381_);
  and g_138783_(_049375_, _049380_, _049382_);
  not g_138784_(_049382_, _049383_);
  and g_138785_(out[896], _049207_, _049384_);
  or g_138786_(_001880_, _049208_, _049385_);
  and g_138787_(_048998_, _049208_, _049386_);
  or g_138788_(_048997_, _049207_, _049387_);
  and g_138789_(_049385_, _049387_, _049388_);
  or g_138790_(_049384_, _049386_, _049390_);
  and g_138791_(_002012_, _049390_, _049391_);
  or g_138792_(out[912], _049388_, _049392_);
  xor g_138793_(_049375_, _049380_, _049393_);
  xor g_138794_(_049376_, _049380_, _049394_);
  and g_138795_(_049392_, _049393_, _049395_);
  or g_138796_(_049391_, _049394_, _049396_);
  and g_138797_(_049383_, _049396_, _049397_);
  or g_138798_(_049382_, _049395_, _049398_);
  and g_138799_(_049373_, _049398_, _049399_);
  or g_138800_(_049374_, _049397_, _049401_);
  and g_138801_(_049365_, _049368_, _049402_);
  or g_138802_(_049364_, _049366_, _049403_);
  and g_138803_(_049401_, _049403_, _049404_);
  or g_138804_(_049399_, _049402_, _049405_);
  and g_138805_(_049340_, _049405_, _049406_);
  or g_138806_(_049341_, _049404_, _049407_);
  and g_138807_(_049318_, _049335_, _049408_);
  or g_138808_(_049319_, _049333_, _049409_);
  or g_138809_(_049296_, _049298_, _049410_);
  not g_138810_(_049410_, _049412_);
  and g_138811_(_049409_, _049410_, _049413_);
  or g_138812_(_049408_, _049412_, _049414_);
  and g_138813_(_049407_, _049413_, _049415_);
  or g_138814_(_049406_, _049414_, _049416_);
  and g_138815_(_049278_, _049416_, _049417_);
  or g_138816_(_049280_, _049415_, _049418_);
  and g_138817_(_049271_, _049273_, _049419_);
  or g_138818_(_049270_, _049272_, _049420_);
  and g_138819_(_049418_, _049420_, _049421_);
  or g_138820_(_049417_, _049419_, _049423_);
  and g_138821_(_049237_, _049244_, _049424_);
  or g_138822_(_049238_, _049243_, _049425_);
  and g_138823_(_049233_, _049425_, _049426_);
  or g_138824_(_049232_, _049424_, _049427_);
  and g_138825_(_049423_, _049426_, _049428_);
  or g_138826_(_049421_, _049427_, _049429_);
  or g_138827_(_049249_, _049427_, _049430_);
  and g_138828_(_049251_, _049429_, _049431_);
  or g_138829_(_049250_, _049428_, _049432_);
  and g_138830_(out[912], _049388_, _049434_);
  or g_138831_(_049430_, _049434_, _049435_);
  or g_138832_(_049396_, _049435_, _049436_);
  or g_138833_(_049341_, _049436_, _049437_);
  not g_138834_(_049437_, _049438_);
  and g_138835_(_049278_, _049438_, _049439_);
  or g_138836_(_049280_, _049437_, _049440_);
  and g_138837_(_049373_, _049439_, _049441_);
  or g_138838_(_049374_, _049440_, _049442_);
  and g_138839_(_049432_, _049442_, _049443_);
  or g_138840_(_049431_, _049441_, _049445_);
  and g_138841_(_049215_, _049445_, _049446_);
  and g_138842_(_049281_, _049443_, _049447_);
  or g_138843_(_049446_, _049447_, _049448_);
  not g_138844_(_049448_, _049449_);
  or g_138845_(out[929], out[928], _049450_);
  or g_138846_(out[928], _002719_, _049451_);
  and g_138847_(out[931], _049451_, _049452_);
  and g_138848_(_027088_, _049451_, _049453_);
  and g_138849_(out[933], _049453_, _049454_);
  or g_138850_(out[934], _049454_, _049456_);
  and g_138851_(out[935], _049456_, _049457_);
  xor g_138852_(out[935], _049456_, _049458_);
  xor g_138853_(_002078_, _049456_, _049459_);
  and g_138854_(_049293_, _049445_, _049460_);
  and g_138855_(_049286_, _049443_, _049461_);
  or g_138856_(_049460_, _049461_, _049462_);
  not g_138857_(_049462_, _049463_);
  and g_138858_(_049458_, _049462_, _049464_);
  or g_138859_(_049459_, _049463_, _049465_);
  xor g_138860_(out[934], _049454_, _049467_);
  not g_138861_(_049467_, _049468_);
  and g_138862_(_049449_, _049467_, _049469_);
  or g_138863_(_049448_, _049468_, _049470_);
  and g_138864_(_049381_, _049445_, _049471_);
  or g_138865_(_049380_, _049443_, _049472_);
  and g_138866_(_049375_, _049443_, _049473_);
  or g_138867_(_049376_, _049445_, _049474_);
  and g_138868_(_049472_, _049474_, _049475_);
  or g_138869_(_049471_, _049473_, _049476_);
  xor g_138870_(out[929], out[928], _049478_);
  xor g_138871_(_002111_, out[928], _049479_);
  and g_138872_(_049475_, _049478_, _049480_);
  or g_138873_(_049476_, _049479_, _049481_);
  and g_138874_(out[912], _049443_, _049482_);
  or g_138875_(_002012_, _049445_, _049483_);
  and g_138876_(_049390_, _049445_, _049484_);
  or g_138877_(_049388_, _049443_, _049485_);
  and g_138878_(_049483_, _049485_, _049486_);
  or g_138879_(_049482_, _049484_, _049487_);
  and g_138880_(out[928], _049486_, _049489_);
  or g_138881_(_002122_, _049487_, _049490_);
  and g_138882_(_049481_, _049490_, _049491_);
  or g_138883_(_049480_, _049489_, _049492_);
  xor g_138884_(out[930], _049450_, _049493_);
  xor g_138885_(_002133_, _049450_, _049494_);
  and g_138886_(_049350_, _049445_, _049495_);
  or g_138887_(_049349_, _049443_, _049496_);
  and g_138888_(_049342_, _049443_, _049497_);
  or g_138889_(_049343_, _049445_, _049498_);
  and g_138890_(_049496_, _049498_, _049500_);
  or g_138891_(_049495_, _049497_, _049501_);
  and g_138892_(_049494_, _049501_, _049502_);
  or g_138893_(_049493_, _049500_, _049503_);
  and g_138894_(out[929], _049476_, _049504_);
  or g_138895_(_002111_, _049475_, _049505_);
  and g_138896_(_049503_, _049505_, _049506_);
  or g_138897_(_049502_, _049504_, _049507_);
  and g_138898_(_049492_, _049506_, _049508_);
  or g_138899_(_049491_, _049507_, _049509_);
  xor g_138900_(out[931], _049451_, _049511_);
  xor g_138901_(_002144_, _049451_, _049512_);
  or g_138902_(_049353_, _049445_, _049513_);
  not g_138903_(_049513_, _049514_);
  and g_138904_(_049361_, _049445_, _049515_);
  or g_138905_(_049360_, _049443_, _049516_);
  and g_138906_(_049513_, _049516_, _049517_);
  or g_138907_(_049514_, _049515_, _049518_);
  and g_138908_(_049512_, _049517_, _049519_);
  or g_138909_(_049511_, _049518_, _049520_);
  and g_138910_(_049493_, _049500_, _049522_);
  or g_138911_(_049494_, _049501_, _049523_);
  and g_138912_(_049520_, _049523_, _049524_);
  or g_138913_(_049519_, _049522_, _049525_);
  and g_138914_(_049509_, _049524_, _049526_);
  or g_138915_(_049508_, _049525_, _049527_);
  xor g_138916_(out[932], _049452_, _049528_);
  and g_138917_(_049324_, _049443_, _049529_);
  and g_138918_(_049330_, _049445_, _049530_);
  or g_138919_(_049529_, _049530_, _049531_);
  and g_138920_(_049528_, _049531_, _049533_);
  and g_138921_(_049511_, _049518_, _049534_);
  or g_138922_(_049533_, _049534_, _049535_);
  not g_138923_(_049535_, _049536_);
  and g_138924_(_049527_, _049536_, _049537_);
  or g_138925_(_049526_, _049535_, _049538_);
  xor g_138926_(out[933], _049453_, _049539_);
  xor g_138927_(_002089_, _049453_, _049540_);
  and g_138928_(_049313_, _049445_, _049541_);
  and g_138929_(_049306_, _049443_, _049542_);
  or g_138930_(_049541_, _049542_, _049544_);
  not g_138931_(_049544_, _049545_);
  or g_138932_(_049539_, _049544_, _049546_);
  or g_138933_(_049528_, _049531_, _049547_);
  and g_138934_(_049546_, _049547_, _049548_);
  not g_138935_(_049548_, _049549_);
  and g_138936_(_049538_, _049548_, _049550_);
  or g_138937_(_049537_, _049549_, _049551_);
  and g_138938_(_049448_, _049468_, _049552_);
  or g_138939_(_049449_, _049467_, _049553_);
  and g_138940_(_049539_, _049544_, _049555_);
  or g_138941_(_049540_, _049545_, _049556_);
  and g_138942_(_049553_, _049556_, _049557_);
  or g_138943_(_049552_, _049555_, _049558_);
  and g_138944_(_049551_, _049557_, _049559_);
  or g_138945_(_049550_, _049558_, _049560_);
  and g_138946_(_049470_, _049560_, _049561_);
  or g_138947_(_049469_, _049559_, _049562_);
  and g_138948_(_049465_, _049562_, _049563_);
  or g_138949_(_049464_, _049561_, _049564_);
  and g_138950_(out[936], _049457_, _049566_);
  or g_138951_(out[937], _049566_, _049567_);
  and g_138952_(out[938], _049567_, _049568_);
  xor g_138953_(out[938], _049567_, _049569_);
  not g_138954_(_049569_, _049570_);
  and g_138955_(_049244_, _049445_, _049571_);
  or g_138956_(_049243_, _049443_, _049572_);
  or g_138957_(_049237_, _049445_, _049573_);
  not g_138958_(_049573_, _049574_);
  and g_138959_(_049572_, _049573_, _049575_);
  or g_138960_(_049571_, _049574_, _049577_);
  and g_138961_(_049569_, _049577_, _049578_);
  or g_138962_(_049570_, _049575_, _049579_);
  xor g_138963_(out[939], _049568_, _049580_);
  not g_138964_(_049580_, _049581_);
  or g_138965_(_049227_, _049445_, _049582_);
  or g_138966_(_049229_, _049443_, _049583_);
  and g_138967_(_049582_, _049583_, _049584_);
  not g_138968_(_049584_, _049585_);
  and g_138969_(_049231_, _049445_, _049586_);
  and g_138970_(_049227_, _049443_, _049588_);
  or g_138971_(_049586_, _049588_, _049589_);
  and g_138972_(_049580_, _049585_, _049590_);
  or g_138973_(_049581_, _049589_, _049591_);
  or g_138974_(_049578_, _049590_, _049592_);
  and g_138975_(_049570_, _049575_, _049593_);
  and g_138976_(_049581_, _049584_, _049594_);
  or g_138977_(_049580_, _049585_, _049595_);
  or g_138978_(_049593_, _049594_, _049596_);
  xor g_138979_(_049570_, _049575_, _049597_);
  and g_138980_(_049591_, _049595_, _049599_);
  and g_138981_(_049597_, _049599_, _049600_);
  or g_138982_(_049592_, _049596_, _049601_);
  xor g_138983_(out[936], _049457_, _049602_);
  not g_138984_(_049602_, _049603_);
  or g_138985_(_049265_, _049443_, _049604_);
  or g_138986_(_049261_, _049445_, _049605_);
  and g_138987_(_049604_, _049605_, _049606_);
  not g_138988_(_049606_, _049607_);
  and g_138989_(_049602_, _049607_, _049608_);
  or g_138990_(_049603_, _049606_, _049610_);
  xor g_138991_(out[937], _049566_, _049611_);
  not g_138992_(_049611_, _049612_);
  and g_138993_(_049256_, _049445_, _049613_);
  and g_138994_(_049252_, _049443_, _049614_);
  or g_138995_(_049613_, _049614_, _049615_);
  not g_138996_(_049615_, _049616_);
  and g_138997_(_049612_, _049615_, _049617_);
  or g_138998_(_049611_, _049616_, _049618_);
  and g_138999_(_049610_, _049618_, _049619_);
  or g_139000_(_049608_, _049617_, _049621_);
  and g_139001_(_049611_, _049616_, _049622_);
  or g_139002_(_049612_, _049615_, _049623_);
  and g_139003_(_049603_, _049606_, _049624_);
  or g_139004_(_049602_, _049607_, _049625_);
  and g_139005_(_049623_, _049625_, _049626_);
  or g_139006_(_049622_, _049624_, _049627_);
  and g_139007_(_049459_, _049463_, _049628_);
  or g_139008_(_049458_, _049462_, _049629_);
  and g_139009_(_049626_, _049629_, _049630_);
  or g_139010_(_049627_, _049628_, _049632_);
  and g_139011_(_049619_, _049630_, _049633_);
  or g_139012_(_049621_, _049632_, _049634_);
  and g_139013_(_049600_, _049633_, _049635_);
  or g_139014_(_049601_, _049634_, _049636_);
  and g_139015_(_049564_, _049635_, _049637_);
  or g_139016_(_049563_, _049636_, _049638_);
  and g_139017_(_049621_, _049623_, _049639_);
  or g_139018_(_049619_, _049622_, _049640_);
  and g_139019_(_049600_, _049639_, _049641_);
  or g_139020_(_049601_, _049640_, _049643_);
  and g_139021_(_049578_, _049595_, _049644_);
  or g_139022_(_049579_, _049594_, _049645_);
  and g_139023_(_049591_, _049645_, _049646_);
  or g_139024_(_049590_, _049644_, _049647_);
  and g_139025_(_049643_, _049646_, _049648_);
  or g_139026_(_049641_, _049647_, _049649_);
  and g_139027_(_049638_, _049648_, _049650_);
  or g_139028_(_049637_, _049649_, _049651_);
  and g_139029_(_049448_, _049651_, _049652_);
  and g_139030_(_049467_, _049650_, _049654_);
  or g_139031_(_049652_, _049654_, _049655_);
  not g_139032_(_049655_, _049656_);
  and g_139033_(_043338_, _049656_, _049657_);
  or g_139034_(_043340_, _049655_, _049658_);
  xor g_139035_(out[949], _043329_, _049659_);
  xor g_139036_(_002210_, _043329_, _049660_);
  and g_139037_(_049544_, _049651_, _049661_);
  and g_139038_(_049540_, _049650_, _049662_);
  or g_139039_(_049661_, _049662_, _049663_);
  and g_139040_(_049659_, _049663_, _049665_);
  not g_139041_(_049665_, _049666_);
  and g_139042_(_049478_, _049650_, _049667_);
  or g_139043_(_049479_, _049651_, _049668_);
  and g_139044_(_049476_, _049651_, _049669_);
  or g_139045_(_049475_, _049650_, _049670_);
  and g_139046_(_049668_, _049670_, _049671_);
  or g_139047_(_049667_, _049669_, _049672_);
  xor g_139048_(_054336_, out[944], _049673_);
  not g_139049_(_049673_, _049674_);
  and g_139050_(_049671_, _049674_, _049676_);
  or g_139051_(_049672_, _049673_, _049677_);
  and g_139052_(out[928], _049650_, _049678_);
  or g_139053_(_002122_, _049651_, _049679_);
  and g_139054_(_049487_, _049651_, _049680_);
  or g_139055_(_049486_, _049650_, _049681_);
  and g_139056_(_049679_, _049681_, _049682_);
  or g_139057_(_049678_, _049680_, _049683_);
  and g_139058_(out[944], _049682_, _049684_);
  or g_139059_(_002232_, _049683_, _049685_);
  and g_139060_(_049677_, _049685_, _049687_);
  or g_139061_(_049676_, _049684_, _049688_);
  xor g_139062_(out[946], _043325_, _049689_);
  xor g_139063_(_002243_, _043325_, _049690_);
  and g_139064_(_049493_, _049650_, _049691_);
  or g_139065_(_049494_, _049651_, _049692_);
  and g_139066_(_049501_, _049651_, _049693_);
  or g_139067_(_049500_, _049650_, _049694_);
  and g_139068_(_049692_, _049694_, _049695_);
  or g_139069_(_049691_, _049693_, _049696_);
  and g_139070_(_049690_, _049696_, _049698_);
  or g_139071_(_049689_, _049695_, _049699_);
  and g_139072_(out[945], _049672_, _049700_);
  or g_139073_(_054336_, _049671_, _049701_);
  and g_139074_(_049699_, _049701_, _049702_);
  or g_139075_(_049698_, _049700_, _049703_);
  and g_139076_(_049688_, _049702_, _049704_);
  or g_139077_(_049687_, _049703_, _049705_);
  xor g_139078_(out[947], _043326_, _049706_);
  and g_139079_(_049512_, _049650_, _049707_);
  and g_139080_(_049518_, _049651_, _049709_);
  or g_139081_(_049707_, _049709_, _049710_);
  or g_139082_(_049706_, _049710_, _049711_);
  not g_139083_(_049711_, _049712_);
  and g_139084_(_049689_, _049695_, _049713_);
  not g_139085_(_049713_, _049714_);
  and g_139086_(_049711_, _049714_, _049715_);
  or g_139087_(_049712_, _049713_, _049716_);
  and g_139088_(_049705_, _049715_, _049717_);
  or g_139089_(_049704_, _049716_, _049718_);
  and g_139090_(_049706_, _049710_, _049720_);
  xor g_139091_(out[948], _043327_, _049721_);
  not g_139092_(_049721_, _049722_);
  or g_139093_(_049528_, _049651_, _049723_);
  not g_139094_(_049723_, _049724_);
  and g_139095_(_049531_, _049651_, _049725_);
  or g_139096_(_049724_, _049725_, _049726_);
  and g_139097_(_049721_, _049726_, _049727_);
  or g_139098_(_049720_, _049727_, _049728_);
  not g_139099_(_049728_, _049729_);
  and g_139100_(_049718_, _049729_, _049731_);
  or g_139101_(_049717_, _049728_, _049732_);
  or g_139102_(_049659_, _049663_, _049733_);
  or g_139103_(_049721_, _049726_, _049734_);
  and g_139104_(_049733_, _049734_, _049735_);
  not g_139105_(_049735_, _049736_);
  and g_139106_(_049732_, _049735_, _049737_);
  or g_139107_(_049731_, _049736_, _049738_);
  and g_139108_(_049666_, _049738_, _049739_);
  or g_139109_(_049665_, _049737_, _049740_);
  and g_139110_(_049658_, _049740_, _049742_);
  or g_139111_(_049657_, _049739_, _049743_);
  xor g_139112_(out[951], _043331_, _049744_);
  xor g_139113_(_002188_, _043331_, _049745_);
  and g_139114_(_049462_, _049651_, _049746_);
  and g_139115_(_049459_, _049650_, _049747_);
  or g_139116_(_049746_, _049747_, _049748_);
  not g_139117_(_049748_, _049749_);
  and g_139118_(_049744_, _049748_, _049750_);
  or g_139119_(_049745_, _049749_, _049751_);
  and g_139120_(_043340_, _049655_, _049753_);
  or g_139121_(_043338_, _049656_, _049754_);
  and g_139122_(_049751_, _049754_, _049755_);
  or g_139123_(_049750_, _049753_, _049756_);
  and g_139124_(_049743_, _049755_, _049757_);
  or g_139125_(_049742_, _049756_, _049758_);
  xor g_139126_(out[952], _043332_, _049759_);
  not g_139127_(_049759_, _049760_);
  or g_139128_(_049606_, _049650_, _049761_);
  or g_139129_(_049602_, _049651_, _049762_);
  and g_139130_(_049761_, _049762_, _049764_);
  not g_139131_(_049764_, _049765_);
  and g_139132_(_049760_, _049764_, _049766_);
  or g_139133_(_049759_, _049765_, _049767_);
  and g_139134_(_049759_, _049765_, _049768_);
  or g_139135_(_049760_, _049764_, _049769_);
  xor g_139136_(out[953], _043333_, _049770_);
  not g_139137_(_049770_, _049771_);
  and g_139138_(_049615_, _049651_, _049772_);
  and g_139139_(_049611_, _049650_, _049773_);
  or g_139140_(_049772_, _049773_, _049775_);
  not g_139141_(_049775_, _049776_);
  and g_139142_(_049771_, _049775_, _049777_);
  or g_139143_(_049770_, _049776_, _049778_);
  and g_139144_(_049769_, _049778_, _049779_);
  or g_139145_(_049768_, _049777_, _049780_);
  and g_139146_(_049767_, _049779_, _049781_);
  or g_139147_(_049766_, _049780_, _049782_);
  and g_139148_(_049580_, _049584_, _049783_);
  not g_139149_(_049783_, _049784_);
  and g_139150_(_043337_, _049783_, _049786_);
  or g_139151_(_043336_, _049784_, _049787_);
  xor g_139152_(out[954], _043334_, _049788_);
  xor g_139153_(_002287_, _043334_, _049789_);
  and g_139154_(_049577_, _049651_, _049790_);
  or g_139155_(_049569_, _049651_, _049791_);
  not g_139156_(_049791_, _049792_);
  or g_139157_(_049790_, _049792_, _049793_);
  not g_139158_(_049793_, _049794_);
  and g_139159_(_049789_, _049794_, _049795_);
  or g_139160_(_049788_, _049793_, _049797_);
  and g_139161_(_049787_, _049797_, _049798_);
  or g_139162_(_049786_, _049795_, _049799_);
  and g_139163_(_049788_, _049793_, _049800_);
  or g_139164_(_049789_, _049794_, _049801_);
  and g_139165_(_049580_, _049589_, _049802_);
  and g_139166_(_043336_, _049784_, _049803_);
  or g_139167_(_043337_, _049802_, _049804_);
  and g_139168_(_049801_, _049804_, _049805_);
  or g_139169_(_049800_, _049803_, _049806_);
  and g_139170_(_049745_, _049749_, _049808_);
  or g_139171_(_049744_, _049748_, _049809_);
  and g_139172_(_049770_, _049776_, _049810_);
  or g_139173_(_049771_, _049775_, _049811_);
  and g_139174_(_049809_, _049811_, _049812_);
  or g_139175_(_049808_, _049810_, _049813_);
  and g_139176_(_049805_, _049812_, _049814_);
  or g_139177_(_049806_, _049813_, _049815_);
  and g_139178_(_049798_, _049814_, _049816_);
  or g_139179_(_049799_, _049815_, _049817_);
  and g_139180_(_049781_, _049816_, _049819_);
  or g_139181_(_049782_, _049817_, _049820_);
  and g_139182_(_049758_, _049819_, _049821_);
  or g_139183_(_049757_, _049820_, _049822_);
  and g_139184_(_049787_, _049806_, _049823_);
  or g_139185_(_049786_, _049805_, _049824_);
  and g_139186_(_049798_, _049811_, _049825_);
  or g_139187_(_049799_, _049810_, _049826_);
  and g_139188_(_049780_, _049825_, _049827_);
  or g_139189_(_049779_, _049826_, _049828_);
  and g_139190_(_049824_, _049828_, _049830_);
  or g_139191_(_049823_, _049827_, _049831_);
  and g_139192_(_049822_, _049830_, _049832_);
  or g_139193_(_049821_, _049831_, _049833_);
  xor g_139194_(out[469], _038245_, _049834_);
  not g_139195_(_049834_, _049835_);
  and g_139196_(_043087_, _043304_, _049836_);
  or g_139197_(_043088_, _043303_, _049837_);
  and g_139198_(_038346_, _043303_, _049838_);
  or g_139199_(_038347_, _043304_, _049839_);
  and g_139200_(_049837_, _049839_, _049841_);
  or g_139201_(_049836_, _049838_, _049842_);
  and g_139202_(_038332_, _049842_, _049843_);
  or g_139203_(_038333_, _049841_, _049844_);
  and g_139204_(_038319_, _049843_, _049845_);
  or g_139205_(_038320_, _049844_, _049846_);
  and g_139206_(_038306_, _049845_, _049847_);
  or g_139207_(_038307_, _049846_, _049848_);
  or g_139208_(_038294_, _049848_, _049849_);
  or g_139209_(_038281_, _049849_, _049850_);
  or g_139210_(_038267_, _049850_, _049852_);
  and g_139211_(_038253_, _049852_, _049853_);
  or g_139212_(_038254_, _043323_, _049854_);
  xor g_139213_(out[458], _038264_, _049855_);
  not g_139214_(_049855_, _049856_);
  and g_139215_(_038267_, _043321_, _049857_);
  or g_139216_(_038266_, _043322_, _049858_);
  xor g_139217_(out[442], _038277_, _049859_);
  xor g_139218_(_004784_, _038277_, _049860_);
  xor g_139219_(_054105_, _038269_, _049861_);
  xor g_139220_(out[418], _038282_, _049863_);
  not g_139221_(_049863_, _049864_);
  xor g_139222_(out[426], _038291_, _049865_);
  not g_139223_(_049865_, _049866_);
  xor g_139224_(out[394], _038317_, _049867_);
  xor g_139225_(_004685_, _038317_, _049868_);
  or g_139226_(_038348_, _043304_, _049869_);
  or g_139227_(_043080_, _043303_, _049870_);
  and g_139228_(_049869_, _049870_, _049871_);
  not g_139229_(_049871_, _049872_);
  and g_139230_(_043098_, _043303_, _049874_);
  or g_139231_(_043099_, _043304_, _049875_);
  and g_139232_(_043105_, _043304_, _049876_);
  or g_139233_(_043104_, _043303_, _049877_);
  and g_139234_(_049875_, _049877_, _049878_);
  or g_139235_(_049874_, _049876_, _049879_);
  xor g_139236_(out[377], _038329_, _049880_);
  xor g_139237_(_053731_, _038329_, _049881_);
  and g_139238_(_049879_, _049881_, _049882_);
  or g_139239_(_049878_, _049880_, _049883_);
  xor g_139240_(out[376], _038328_, _049885_);
  xor g_139241_(_053654_, _038328_, _049886_);
  and g_139242_(_043116_, _043303_, _049887_);
  or g_139243_(_043115_, _043304_, _049888_);
  and g_139244_(_043123_, _043304_, _049889_);
  or g_139245_(_043122_, _043303_, _049890_);
  and g_139246_(_049888_, _049890_, _049891_);
  or g_139247_(_049887_, _049889_, _049892_);
  and g_139248_(_049885_, _049892_, _049893_);
  or g_139249_(_049886_, _049891_, _049894_);
  and g_139250_(_049883_, _049894_, _049896_);
  or g_139251_(_049882_, _049893_, _049897_);
  and g_139252_(out[352], _043303_, _049898_);
  or g_139253_(_004608_, _043304_, _049899_);
  and g_139254_(_043180_, _043304_, _049900_);
  or g_139255_(_043179_, _043303_, _049901_);
  and g_139256_(_049899_, _049901_, _049902_);
  or g_139257_(_049898_, _049900_, _049903_);
  and g_139258_(out[368], _049902_, _049904_);
  or g_139259_(_004641_, _049903_, _049905_);
  and g_139260_(_043171_, _043304_, _049907_);
  or g_139261_(_043170_, _043303_, _049908_);
  and g_139262_(_043164_, _043303_, _049909_);
  or g_139263_(_043165_, _043304_, _049910_);
  and g_139264_(_049908_, _049910_, _049911_);
  or g_139265_(_049907_, _049909_, _049912_);
  and g_139266_(out[369], _049912_, _049913_);
  or g_139267_(_053720_, _049911_, _049914_);
  xor g_139268_(out[369], out[368], _049915_);
  xor g_139269_(_053720_, out[368], _049916_);
  and g_139270_(_049904_, _049914_, _049918_);
  or g_139271_(_049905_, _049913_, _049919_);
  and g_139272_(_043145_, _043304_, _049920_);
  or g_139273_(_043144_, _043303_, _049921_);
  and g_139274_(_043137_, _043303_, _049922_);
  or g_139275_(_043138_, _043304_, _049923_);
  and g_139276_(_049921_, _049923_, _049924_);
  or g_139277_(_049920_, _049922_, _049925_);
  xor g_139278_(out[370], _038321_, _049926_);
  xor g_139279_(_053709_, _038321_, _049927_);
  and g_139280_(_049924_, _049926_, _049929_);
  or g_139281_(_049925_, _049927_, _049930_);
  and g_139282_(_049911_, _049915_, _049931_);
  or g_139283_(_049912_, _049916_, _049932_);
  and g_139284_(_049930_, _049932_, _049933_);
  or g_139285_(_049929_, _049931_, _049934_);
  and g_139286_(_049919_, _049933_, _049935_);
  or g_139287_(_049918_, _049934_, _049936_);
  xor g_139288_(out[371], _038322_, _049937_);
  xor g_139289_(_053687_, _038322_, _049938_);
  and g_139290_(_043149_, _043303_, _049940_);
  or g_139291_(_043148_, _043304_, _049941_);
  and g_139292_(_043156_, _043304_, _049942_);
  or g_139293_(_043155_, _043303_, _049943_);
  and g_139294_(_049941_, _049943_, _049944_);
  or g_139295_(_049940_, _049942_, _049945_);
  and g_139296_(_049937_, _049945_, _049946_);
  or g_139297_(_049938_, _049944_, _049947_);
  and g_139298_(_049925_, _049927_, _049948_);
  or g_139299_(_049924_, _049926_, _049949_);
  and g_139300_(_049947_, _049949_, _049951_);
  or g_139301_(_049946_, _049948_, _049952_);
  and g_139302_(_049936_, _049951_, _049953_);
  or g_139303_(_049935_, _049952_, _049954_);
  xor g_139304_(out[372], _038324_, _049955_);
  xor g_139305_(_053698_, _038324_, _049956_);
  and g_139306_(_043242_, _043303_, _049957_);
  or g_139307_(_043241_, _043304_, _049958_);
  and g_139308_(_043248_, _043304_, _049959_);
  or g_139309_(_043247_, _043303_, _049960_);
  and g_139310_(_049958_, _049960_, _049962_);
  or g_139311_(_049957_, _049959_, _049963_);
  and g_139312_(_049956_, _049962_, _049964_);
  or g_139313_(_049955_, _049963_, _049965_);
  and g_139314_(_049938_, _049944_, _049966_);
  or g_139315_(_049937_, _049945_, _049967_);
  and g_139316_(_049965_, _049967_, _049968_);
  or g_139317_(_049964_, _049966_, _049969_);
  and g_139318_(_049954_, _049968_, _049970_);
  or g_139319_(_049953_, _049969_, _049971_);
  xor g_139320_(out[373], _038325_, _049973_);
  xor g_139321_(_053665_, _038325_, _049974_);
  and g_139322_(_043226_, _043304_, _049975_);
  or g_139323_(_043225_, _043303_, _049976_);
  and g_139324_(_043220_, _043303_, _049977_);
  or g_139325_(_043219_, _043304_, _049978_);
  and g_139326_(_049976_, _049978_, _049979_);
  or g_139327_(_049975_, _049977_, _049980_);
  and g_139328_(_049973_, _049980_, _049981_);
  or g_139329_(_049974_, _049979_, _049982_);
  and g_139330_(_049955_, _049963_, _049984_);
  or g_139331_(_049956_, _049962_, _049985_);
  and g_139332_(_049982_, _049985_, _049986_);
  or g_139333_(_049981_, _049984_, _049987_);
  and g_139334_(_049971_, _049986_, _049988_);
  or g_139335_(_049970_, _049987_, _049989_);
  xor g_139336_(out[374], _038326_, _049990_);
  xor g_139337_(_053676_, _038326_, _049991_);
  and g_139338_(_043194_, _043303_, _049992_);
  or g_139339_(_043195_, _043304_, _049993_);
  and g_139340_(_043202_, _043304_, _049995_);
  or g_139341_(_043201_, _043303_, _049996_);
  and g_139342_(_049993_, _049996_, _049997_);
  or g_139343_(_049992_, _049995_, _049998_);
  and g_139344_(_049990_, _049997_, _049999_);
  or g_139345_(_049991_, _049998_, _050000_);
  and g_139346_(_049974_, _049979_, _050001_);
  or g_139347_(_049973_, _049980_, _050002_);
  and g_139348_(_050000_, _050002_, _050003_);
  or g_139349_(_049999_, _050001_, _050004_);
  and g_139350_(_049989_, _050003_, _050006_);
  or g_139351_(_049988_, _050004_, _050007_);
  xor g_139352_(out[375], _038327_, _050008_);
  xor g_139353_(_053643_, _038327_, _050009_);
  and g_139354_(_043206_, _043303_, _050010_);
  or g_139355_(_043205_, _043304_, _050011_);
  and g_139356_(_043213_, _043304_, _050012_);
  or g_139357_(_043212_, _043303_, _050013_);
  and g_139358_(_050011_, _050013_, _050014_);
  or g_139359_(_050010_, _050012_, _050015_);
  and g_139360_(_050008_, _050015_, _050017_);
  or g_139361_(_050009_, _050014_, _050018_);
  and g_139362_(_049991_, _049998_, _050019_);
  or g_139363_(_049990_, _049997_, _050020_);
  and g_139364_(_050018_, _050020_, _050021_);
  or g_139365_(_050017_, _050019_, _050022_);
  and g_139366_(_050007_, _050021_, _050023_);
  or g_139367_(_050006_, _050022_, _050024_);
  and g_139368_(_049886_, _049891_, _050025_);
  or g_139369_(_049885_, _049892_, _050026_);
  and g_139370_(_050009_, _050014_, _050028_);
  or g_139371_(_050008_, _050015_, _050029_);
  and g_139372_(_050026_, _050029_, _050030_);
  or g_139373_(_050025_, _050028_, _050031_);
  xor g_139374_(out[378], _038330_, _050032_);
  not g_139375_(_050032_, _050033_);
  and g_139376_(_038332_, _049841_, _050034_);
  or g_139377_(_038333_, _049842_, _050035_);
  and g_139378_(_049872_, _050032_, _050036_);
  or g_139379_(_049871_, _050033_, _050037_);
  and g_139380_(_049878_, _049880_, _050039_);
  or g_139381_(_049879_, _049881_, _050040_);
  and g_139382_(_038333_, _043310_, _050041_);
  or g_139383_(_038332_, _043311_, _050042_);
  xor g_139384_(_049871_, _050033_, _050043_);
  xor g_139385_(_049871_, _050032_, _050044_);
  and g_139386_(_050035_, _050042_, _050045_);
  or g_139387_(_050034_, _050041_, _050046_);
  and g_139388_(_050043_, _050045_, _050047_);
  or g_139389_(_050044_, _050046_, _050048_);
  and g_139390_(_049896_, _050040_, _050050_);
  or g_139391_(_049897_, _050039_, _050051_);
  and g_139392_(_050030_, _050050_, _050052_);
  or g_139393_(_050031_, _050051_, _050053_);
  and g_139394_(_050036_, _050042_, _050054_);
  or g_139395_(_050037_, _050041_, _050055_);
  and g_139396_(_050047_, _050052_, _050056_);
  or g_139397_(_050048_, _050053_, _050057_);
  and g_139398_(_050024_, _050056_, _050058_);
  or g_139399_(_050023_, _050057_, _050059_);
  and g_139400_(_049897_, _050047_, _050061_);
  or g_139401_(_049896_, _050048_, _050062_);
  and g_139402_(_050040_, _050061_, _050063_);
  or g_139403_(_050039_, _050062_, _050064_);
  and g_139404_(_050035_, _050064_, _050065_);
  or g_139405_(_050034_, _050063_, _050066_);
  and g_139406_(_050055_, _050065_, _050067_);
  or g_139407_(_050054_, _050066_, _050068_);
  and g_139408_(_050059_, _050067_, _050069_);
  or g_139409_(_050058_, _050068_, _050070_);
  and g_139410_(_049872_, _050070_, _050072_);
  or g_139411_(_049871_, _050069_, _050073_);
  and g_139412_(_050033_, _050069_, _050074_);
  or g_139413_(_050032_, _050070_, _050075_);
  and g_139414_(_050073_, _050075_, _050076_);
  or g_139415_(_050072_, _050074_, _050077_);
  and g_139416_(_049868_, _050076_, _050078_);
  or g_139417_(_049867_, _050077_, _050079_);
  and g_139418_(_038320_, _043312_, _050080_);
  or g_139419_(_038319_, _043313_, _050081_);
  and g_139420_(_050079_, _050081_, _050083_);
  or g_139421_(_050078_, _050080_, _050084_);
  or g_139422_(_050033_, _050070_, _050085_);
  or g_139423_(_049872_, _050069_, _050086_);
  and g_139424_(_050085_, _050086_, _050087_);
  and g_139425_(_049867_, _050077_, _050088_);
  or g_139426_(_049868_, _050076_, _050089_);
  and g_139427_(_038319_, _049844_, _050090_);
  or g_139428_(_038320_, _049843_, _050091_);
  xor g_139429_(out[393], _038316_, _050092_);
  xor g_139430_(_053830_, _038316_, _050094_);
  and g_139431_(_049879_, _050070_, _050095_);
  or g_139432_(_049878_, _050069_, _050096_);
  and g_139433_(_049880_, _050069_, _050097_);
  or g_139434_(_049881_, _050070_, _050098_);
  and g_139435_(_050096_, _050098_, _050099_);
  or g_139436_(_050095_, _050097_, _050100_);
  and g_139437_(_050094_, _050100_, _050101_);
  or g_139438_(_050092_, _050099_, _050102_);
  xor g_139439_(out[392], _038315_, _050103_);
  xor g_139440_(_053753_, _038315_, _050105_);
  and g_139441_(_049892_, _050070_, _050106_);
  or g_139442_(_049891_, _050069_, _050107_);
  and g_139443_(_049886_, _050069_, _050108_);
  or g_139444_(_049885_, _050070_, _050109_);
  and g_139445_(_050107_, _050109_, _050110_);
  or g_139446_(_050106_, _050108_, _050111_);
  and g_139447_(_050103_, _050111_, _050112_);
  or g_139448_(_050105_, _050110_, _050113_);
  and g_139449_(_050092_, _050099_, _050114_);
  or g_139450_(_050094_, _050100_, _050116_);
  and g_139451_(_050105_, _050110_, _050117_);
  or g_139452_(_050103_, _050111_, _050118_);
  and g_139453_(_050116_, _050118_, _050119_);
  or g_139454_(_050114_, _050117_, _050120_);
  and g_139455_(_050102_, _050119_, _050121_);
  or g_139456_(_050101_, _050120_, _050122_);
  and g_139457_(_050083_, _050089_, _050123_);
  or g_139458_(_050084_, _050088_, _050124_);
  and g_139459_(_050091_, _050123_, _050125_);
  or g_139460_(_050090_, _050124_, _050127_);
  and g_139461_(_050113_, _050125_, _050128_);
  or g_139462_(_050112_, _050127_, _050129_);
  and g_139463_(_050121_, _050128_, _050130_);
  or g_139464_(_050122_, _050129_, _050131_);
  xor g_139465_(out[390], _038313_, _050132_);
  xor g_139466_(_053775_, _038313_, _050133_);
  and g_139467_(_049998_, _050070_, _050134_);
  or g_139468_(_049997_, _050069_, _050135_);
  and g_139469_(_049990_, _050069_, _050136_);
  or g_139470_(_049991_, _050070_, _050138_);
  and g_139471_(_050135_, _050138_, _050139_);
  or g_139472_(_050134_, _050136_, _050140_);
  and g_139473_(_050132_, _050139_, _050141_);
  or g_139474_(_050133_, _050140_, _050142_);
  xor g_139475_(out[391], _038314_, _050143_);
  xor g_139476_(_053742_, _038314_, _050144_);
  and g_139477_(_050015_, _050070_, _050145_);
  or g_139478_(_050014_, _050069_, _050146_);
  and g_139479_(_050009_, _050069_, _050147_);
  or g_139480_(_050008_, _050070_, _050149_);
  and g_139481_(_050146_, _050149_, _050150_);
  or g_139482_(_050145_, _050147_, _050151_);
  and g_139483_(_050144_, _050150_, _050152_);
  or g_139484_(_050143_, _050151_, _050153_);
  and g_139485_(_050142_, _050153_, _050154_);
  or g_139486_(_050141_, _050152_, _050155_);
  and g_139487_(_050133_, _050140_, _050156_);
  or g_139488_(_050132_, _050139_, _050157_);
  and g_139489_(_050143_, _050151_, _050158_);
  or g_139490_(_050144_, _050150_, _050160_);
  xor g_139491_(out[389], _038311_, _050161_);
  xor g_139492_(_053764_, _038311_, _050162_);
  and g_139493_(_049974_, _050069_, _050163_);
  or g_139494_(_049973_, _050070_, _050164_);
  and g_139495_(_049980_, _050070_, _050165_);
  or g_139496_(_049979_, _050069_, _050166_);
  and g_139497_(_050164_, _050166_, _050167_);
  or g_139498_(_050163_, _050165_, _050168_);
  and g_139499_(_050161_, _050168_, _050169_);
  or g_139500_(_050162_, _050167_, _050171_);
  and g_139501_(_050160_, _050171_, _050172_);
  or g_139502_(_050158_, _050169_, _050173_);
  and g_139503_(_050157_, _050172_, _050174_);
  or g_139504_(_050156_, _050173_, _050175_);
  and g_139505_(_050154_, _050174_, _050176_);
  or g_139506_(_050155_, _050175_, _050177_);
  xor g_139507_(out[388], _038310_, _050178_);
  xor g_139508_(_053797_, _038310_, _050179_);
  and g_139509_(_049956_, _050069_, _050180_);
  or g_139510_(_049955_, _050070_, _050182_);
  and g_139511_(_049963_, _050070_, _050183_);
  or g_139512_(_049962_, _050069_, _050184_);
  and g_139513_(_050182_, _050184_, _050185_);
  or g_139514_(_050180_, _050183_, _050186_);
  and g_139515_(_050178_, _050186_, _050187_);
  or g_139516_(_050179_, _050185_, _050188_);
  and g_139517_(_050179_, _050185_, _050189_);
  or g_139518_(_050178_, _050186_, _050190_);
  and g_139519_(_050162_, _050167_, _050191_);
  or g_139520_(_050161_, _050168_, _050193_);
  and g_139521_(_050190_, _050193_, _050194_);
  or g_139522_(_050189_, _050191_, _050195_);
  and g_139523_(_050188_, _050194_, _050196_);
  or g_139524_(_050187_, _050195_, _050197_);
  and g_139525_(_050176_, _050196_, _050198_);
  or g_139526_(_050177_, _050197_, _050199_);
  xor g_139527_(out[387], _038309_, _050200_);
  xor g_139528_(_053786_, _038309_, _050201_);
  and g_139529_(_049945_, _050070_, _050202_);
  or g_139530_(_049944_, _050069_, _050204_);
  and g_139531_(_049938_, _050069_, _050205_);
  or g_139532_(_049937_, _050070_, _050206_);
  and g_139533_(_050204_, _050206_, _050207_);
  or g_139534_(_050202_, _050205_, _050208_);
  and g_139535_(_050201_, _050207_, _050209_);
  or g_139536_(_050200_, _050208_, _050210_);
  and g_139537_(_049925_, _050070_, _050211_);
  or g_139538_(_049924_, _050069_, _050212_);
  and g_139539_(_049926_, _050069_, _050213_);
  or g_139540_(_049927_, _050070_, _050215_);
  and g_139541_(_050212_, _050215_, _050216_);
  or g_139542_(_050211_, _050213_, _050217_);
  xor g_139543_(out[386], _038308_, _050218_);
  not g_139544_(_050218_, _050219_);
  and g_139545_(_050216_, _050218_, _050220_);
  or g_139546_(_050217_, _050219_, _050221_);
  and g_139547_(_050210_, _050221_, _050222_);
  or g_139548_(_050209_, _050220_, _050223_);
  and g_139549_(_050200_, _050208_, _050224_);
  or g_139550_(_050201_, _050207_, _050226_);
  and g_139551_(_050217_, _050219_, _050227_);
  or g_139552_(_050216_, _050218_, _050228_);
  and g_139553_(_050226_, _050228_, _050229_);
  or g_139554_(_050224_, _050227_, _050230_);
  and g_139555_(_050222_, _050229_, _050231_);
  or g_139556_(_050223_, _050230_, _050232_);
  xor g_139557_(out[385], out[384], _050233_);
  not g_139558_(_050233_, _050234_);
  and g_139559_(_049915_, _050069_, _050235_);
  or g_139560_(_049916_, _050070_, _050237_);
  and g_139561_(_049912_, _050070_, _050238_);
  or g_139562_(_049911_, _050069_, _050239_);
  and g_139563_(_050237_, _050239_, _050240_);
  or g_139564_(_050235_, _050238_, _050241_);
  and g_139565_(_050233_, _050240_, _050242_);
  or g_139566_(_050234_, _050241_, _050243_);
  and g_139567_(out[368], _050069_, _050244_);
  or g_139568_(_004641_, _050070_, _050245_);
  and g_139569_(_049903_, _050070_, _050246_);
  or g_139570_(_049902_, _050069_, _050248_);
  and g_139571_(_050245_, _050248_, _050249_);
  or g_139572_(_050244_, _050246_, _050250_);
  and g_139573_(_004674_, _050250_, _050251_);
  or g_139574_(out[384], _050249_, _050252_);
  xor g_139575_(_050233_, _050240_, _050253_);
  xor g_139576_(_050234_, _050240_, _050254_);
  and g_139577_(_050252_, _050253_, _050255_);
  or g_139578_(_050251_, _050254_, _050256_);
  and g_139579_(_050243_, _050256_, _050257_);
  or g_139580_(_050242_, _050255_, _050259_);
  and g_139581_(_050231_, _050259_, _050260_);
  or g_139582_(_050232_, _050257_, _050261_);
  and g_139583_(_050223_, _050226_, _050262_);
  or g_139584_(_050222_, _050224_, _050263_);
  and g_139585_(_050261_, _050263_, _050264_);
  or g_139586_(_050260_, _050262_, _050265_);
  and g_139587_(_050198_, _050265_, _050266_);
  or g_139588_(_050199_, _050264_, _050267_);
  and g_139589_(_050155_, _050160_, _050268_);
  or g_139590_(_050154_, _050158_, _050270_);
  and g_139591_(_050176_, _050195_, _050271_);
  or g_139592_(_050177_, _050194_, _050272_);
  and g_139593_(_050270_, _050272_, _050273_);
  or g_139594_(_050268_, _050271_, _050274_);
  and g_139595_(_050267_, _050273_, _050275_);
  or g_139596_(_050266_, _050274_, _050276_);
  and g_139597_(_050130_, _050276_, _050277_);
  or g_139598_(_050131_, _050275_, _050278_);
  and g_139599_(_050102_, _050120_, _050279_);
  or g_139600_(_050101_, _050119_, _050281_);
  and g_139601_(_050125_, _050279_, _050282_);
  or g_139602_(_050127_, _050281_, _050283_);
  and g_139603_(_050084_, _050091_, _050284_);
  or g_139604_(_050083_, _050090_, _050285_);
  and g_139605_(_050283_, _050285_, _050286_);
  or g_139606_(_050282_, _050284_, _050287_);
  and g_139607_(_050278_, _050286_, _050288_);
  or g_139608_(_050277_, _050287_, _050289_);
  and g_139609_(out[384], _050249_, _050290_);
  or g_139610_(_004674_, _050250_, _050292_);
  and g_139611_(_050231_, _050255_, _050293_);
  or g_139612_(_050232_, _050256_, _050294_);
  and g_139613_(_050292_, _050293_, _050295_);
  or g_139614_(_050290_, _050294_, _050296_);
  and g_139615_(_050198_, _050295_, _050297_);
  or g_139616_(_050199_, _050296_, _050298_);
  and g_139617_(_050130_, _050297_, _050299_);
  or g_139618_(_050131_, _050298_, _050300_);
  and g_139619_(_050289_, _050300_, _050301_);
  or g_139620_(_050288_, _050299_, _050303_);
  and g_139621_(_049868_, _050301_, _050304_);
  or g_139622_(_049867_, _050303_, _050305_);
  and g_139623_(_050077_, _050303_, _050306_);
  or g_139624_(_050076_, _050301_, _050307_);
  and g_139625_(_050305_, _050307_, _050308_);
  or g_139626_(_050304_, _050306_, _050309_);
  xor g_139627_(out[407], _038300_, _050310_);
  xor g_139628_(_053841_, _038300_, _050311_);
  and g_139629_(_050144_, _050301_, _050312_);
  or g_139630_(_050143_, _050303_, _050314_);
  and g_139631_(_050151_, _050303_, _050315_);
  or g_139632_(_050150_, _050301_, _050316_);
  and g_139633_(_050314_, _050316_, _050317_);
  or g_139634_(_050312_, _050315_, _050318_);
  and g_139635_(_050310_, _050318_, _050319_);
  or g_139636_(_050311_, _050317_, _050320_);
  xor g_139637_(out[406], _038299_, _050321_);
  xor g_139638_(_053874_, _038299_, _050322_);
  and g_139639_(_050132_, _050301_, _050323_);
  or g_139640_(_050133_, _050303_, _050325_);
  and g_139641_(_050140_, _050303_, _050326_);
  or g_139642_(_050139_, _050301_, _050327_);
  and g_139643_(_050325_, _050327_, _050328_);
  or g_139644_(_050323_, _050326_, _050329_);
  and g_139645_(_050321_, _050328_, _050330_);
  or g_139646_(_050322_, _050329_, _050331_);
  xor g_139647_(out[405], _038298_, _050332_);
  xor g_139648_(_053863_, _038298_, _050333_);
  and g_139649_(_050162_, _050301_, _050334_);
  or g_139650_(_050161_, _050303_, _050336_);
  and g_139651_(_050168_, _050303_, _050337_);
  or g_139652_(_050167_, _050301_, _050338_);
  and g_139653_(_050336_, _050338_, _050339_);
  or g_139654_(_050334_, _050337_, _050340_);
  and g_139655_(_050333_, _050339_, _050341_);
  or g_139656_(_050332_, _050340_, _050342_);
  xor g_139657_(out[404], _038297_, _050343_);
  xor g_139658_(_053896_, _038297_, _050344_);
  and g_139659_(_050186_, _050303_, _050345_);
  or g_139660_(_050185_, _050301_, _050347_);
  and g_139661_(_050179_, _050301_, _050348_);
  or g_139662_(_050178_, _050303_, _050349_);
  and g_139663_(_050347_, _050349_, _050350_);
  or g_139664_(_050345_, _050348_, _050351_);
  and g_139665_(_050343_, _050351_, _050352_);
  or g_139666_(_050344_, _050350_, _050353_);
  and g_139667_(_050217_, _050303_, _050354_);
  or g_139668_(_050216_, _050301_, _050355_);
  and g_139669_(_050218_, _050301_, _050356_);
  not g_139670_(_050356_, _050358_);
  and g_139671_(_050355_, _050358_, _050359_);
  or g_139672_(_050354_, _050356_, _050360_);
  xor g_139673_(out[402], _038295_, _050361_);
  xor g_139674_(_053907_, _038295_, _050362_);
  and g_139675_(_050359_, _050361_, _050363_);
  or g_139676_(_050360_, _050362_, _050364_);
  and g_139677_(_050241_, _050303_, _050365_);
  or g_139678_(_050240_, _050301_, _050366_);
  and g_139679_(_050233_, _050301_, _050367_);
  or g_139680_(_050234_, _050303_, _050369_);
  and g_139681_(_050366_, _050369_, _050370_);
  or g_139682_(_050365_, _050367_, _050371_);
  and g_139683_(out[401], _050371_, _050372_);
  not g_139684_(_050372_, _050373_);
  xor g_139685_(out[401], out[400], _050374_);
  xor g_139686_(_053918_, out[400], _050375_);
  and g_139687_(_050370_, _050374_, _050376_);
  or g_139688_(_050371_, _050375_, _050377_);
  and g_139689_(_050250_, _050303_, _050378_);
  or g_139690_(_050249_, _050301_, _050380_);
  and g_139691_(out[384], _050301_, _050381_);
  or g_139692_(_004674_, _050303_, _050382_);
  and g_139693_(_050380_, _050382_, _050383_);
  or g_139694_(_050378_, _050381_, _050384_);
  and g_139695_(out[400], _050383_, _050385_);
  or g_139696_(_004707_, _050384_, _050386_);
  and g_139697_(_050377_, _050386_, _050387_);
  or g_139698_(_050376_, _050385_, _050388_);
  and g_139699_(_050373_, _050388_, _050389_);
  or g_139700_(_050372_, _050387_, _050391_);
  and g_139701_(_050364_, _050391_, _050392_);
  or g_139702_(_050363_, _050389_, _050393_);
  and g_139703_(_050360_, _050362_, _050394_);
  or g_139704_(_050359_, _050361_, _050395_);
  xor g_139705_(out[403], _038296_, _050396_);
  xor g_139706_(_053885_, _038296_, _050397_);
  and g_139707_(_050208_, _050303_, _050398_);
  or g_139708_(_050207_, _050301_, _050399_);
  and g_139709_(_050201_, _050301_, _050400_);
  or g_139710_(_050200_, _050303_, _050402_);
  and g_139711_(_050399_, _050402_, _050403_);
  or g_139712_(_050398_, _050400_, _050404_);
  and g_139713_(_050396_, _050404_, _050405_);
  or g_139714_(_050397_, _050403_, _050406_);
  and g_139715_(_050395_, _050406_, _050407_);
  or g_139716_(_050394_, _050405_, _050408_);
  and g_139717_(_050393_, _050407_, _050409_);
  or g_139718_(_050392_, _050408_, _050410_);
  and g_139719_(_050344_, _050350_, _050411_);
  or g_139720_(_050343_, _050351_, _050413_);
  and g_139721_(_050397_, _050403_, _050414_);
  or g_139722_(_050396_, _050404_, _050415_);
  and g_139723_(_050413_, _050415_, _050416_);
  or g_139724_(_050411_, _050414_, _050417_);
  and g_139725_(_050410_, _050416_, _050418_);
  or g_139726_(_050409_, _050417_, _050419_);
  and g_139727_(_050353_, _050419_, _050420_);
  or g_139728_(_050352_, _050418_, _050421_);
  and g_139729_(_050342_, _050421_, _050422_);
  or g_139730_(_050341_, _050420_, _050424_);
  and g_139731_(_050322_, _050329_, _050425_);
  or g_139732_(_050321_, _050328_, _050426_);
  and g_139733_(_050332_, _050340_, _050427_);
  or g_139734_(_050333_, _050339_, _050428_);
  and g_139735_(_050426_, _050428_, _050429_);
  or g_139736_(_050425_, _050427_, _050430_);
  and g_139737_(_050424_, _050429_, _050431_);
  or g_139738_(_050422_, _050430_, _050432_);
  and g_139739_(_050331_, _050432_, _050433_);
  or g_139740_(_050330_, _050431_, _050435_);
  and g_139741_(_050320_, _050435_, _050436_);
  or g_139742_(_050319_, _050433_, _050437_);
  and g_139743_(_038306_, _049846_, _050438_);
  or g_139744_(_038307_, _049845_, _050439_);
  xor g_139745_(out[410], _038304_, _050440_);
  xor g_139746_(_004718_, _038304_, _050441_);
  or g_139747_(_049868_, _050303_, _050442_);
  or g_139748_(_050087_, _050301_, _050443_);
  and g_139749_(_050442_, _050443_, _050444_);
  and g_139750_(_050309_, _050440_, _050446_);
  or g_139751_(_050308_, _050441_, _050447_);
  and g_139752_(_050439_, _050447_, _050448_);
  or g_139753_(_050438_, _050446_, _050449_);
  and g_139754_(_050308_, _050441_, _050450_);
  or g_139755_(_050309_, _050440_, _050451_);
  and g_139756_(_038307_, _043314_, _050452_);
  or g_139757_(_038306_, _043315_, _050453_);
  xor g_139758_(out[409], _038303_, _050454_);
  xor g_139759_(_053929_, _038303_, _050455_);
  and g_139760_(_050092_, _050301_, _050457_);
  or g_139761_(_050094_, _050303_, _050458_);
  and g_139762_(_050100_, _050303_, _050459_);
  or g_139763_(_050099_, _050301_, _050460_);
  and g_139764_(_050458_, _050460_, _050461_);
  or g_139765_(_050457_, _050459_, _050462_);
  and g_139766_(_050454_, _050461_, _050463_);
  or g_139767_(_050455_, _050462_, _050464_);
  and g_139768_(_050453_, _050464_, _050465_);
  or g_139769_(_050452_, _050463_, _050466_);
  and g_139770_(_050451_, _050465_, _050468_);
  or g_139771_(_050450_, _050466_, _050469_);
  and g_139772_(_050448_, _050468_, _050470_);
  or g_139773_(_050449_, _050469_, _050471_);
  xor g_139774_(out[408], _038302_, _050472_);
  xor g_139775_(_053852_, _038302_, _050473_);
  and g_139776_(_050105_, _050301_, _050474_);
  or g_139777_(_050103_, _050303_, _050475_);
  and g_139778_(_050111_, _050303_, _050476_);
  or g_139779_(_050110_, _050301_, _050477_);
  and g_139780_(_050475_, _050477_, _050479_);
  or g_139781_(_050474_, _050476_, _050480_);
  and g_139782_(_050473_, _050479_, _050481_);
  or g_139783_(_050472_, _050480_, _050482_);
  and g_139784_(_050311_, _050317_, _050483_);
  or g_139785_(_050310_, _050318_, _050484_);
  and g_139786_(_050482_, _050484_, _050485_);
  or g_139787_(_050481_, _050483_, _050486_);
  and g_139788_(_050472_, _050480_, _050487_);
  or g_139789_(_050473_, _050479_, _050488_);
  and g_139790_(_050455_, _050462_, _050490_);
  or g_139791_(_050454_, _050461_, _050491_);
  and g_139792_(_050488_, _050491_, _050492_);
  or g_139793_(_050487_, _050490_, _050493_);
  and g_139794_(_050485_, _050492_, _050494_);
  or g_139795_(_050486_, _050493_, _050495_);
  and g_139796_(_050470_, _050494_, _050496_);
  or g_139797_(_050471_, _050495_, _050497_);
  and g_139798_(_050437_, _050496_, _050498_);
  or g_139799_(_050436_, _050497_, _050499_);
  and g_139800_(_050470_, _050493_, _050501_);
  or g_139801_(_050471_, _050492_, _050502_);
  and g_139802_(_050449_, _050453_, _050503_);
  or g_139803_(_050448_, _050452_, _050504_);
  and g_139804_(_050502_, _050504_, _050505_);
  or g_139805_(_050501_, _050503_, _050506_);
  and g_139806_(_050499_, _050505_, _050507_);
  or g_139807_(_050498_, _050506_, _050508_);
  and g_139808_(_050309_, _050508_, _050509_);
  not g_139809_(_050509_, _050510_);
  or g_139810_(_050440_, _050508_, _050512_);
  not g_139811_(_050512_, _050513_);
  and g_139812_(_050510_, _050512_, _050514_);
  or g_139813_(_050509_, _050513_, _050515_);
  or g_139814_(_050441_, _050508_, _050516_);
  or g_139815_(_050444_, _050507_, _050517_);
  and g_139816_(_050516_, _050517_, _050518_);
  and g_139817_(_049865_, _050518_, _050519_);
  or g_139818_(_049866_, _050514_, _050520_);
  and g_139819_(_038293_, _049848_, _050521_);
  or g_139820_(_038294_, _049847_, _050523_);
  and g_139821_(_038294_, _049847_, _050524_);
  or g_139822_(_038293_, _049848_, _050525_);
  and g_139823_(_050523_, _050525_, _050526_);
  or g_139824_(_050521_, _050524_, _050527_);
  xor g_139825_(_049866_, _050514_, _050528_);
  xor g_139826_(_049865_, _050514_, _050529_);
  and g_139827_(_050526_, _050528_, _050530_);
  or g_139828_(_050527_, _050529_, _050531_);
  and g_139829_(_050360_, _050508_, _050532_);
  and g_139830_(_050361_, _050507_, _050534_);
  or g_139831_(_050532_, _050534_, _050535_);
  not g_139832_(_050535_, _050536_);
  and g_139833_(_049863_, _050536_, _050537_);
  or g_139834_(_049864_, _050535_, _050538_);
  and g_139835_(_050374_, _050507_, _050539_);
  or g_139836_(_050375_, _050508_, _050540_);
  and g_139837_(_050371_, _050508_, _050541_);
  or g_139838_(_050370_, _050507_, _050542_);
  and g_139839_(_050540_, _050542_, _050543_);
  or g_139840_(_050539_, _050541_, _050545_);
  and g_139841_(out[417], _050545_, _050546_);
  not g_139842_(_050546_, _050547_);
  xor g_139843_(out[417], out[416], _050548_);
  not g_139844_(_050548_, _050549_);
  and g_139845_(_050543_, _050548_, _050550_);
  or g_139846_(_050545_, _050549_, _050551_);
  and g_139847_(out[400], _050507_, _050552_);
  or g_139848_(_004707_, _050508_, _050553_);
  and g_139849_(_050384_, _050508_, _050554_);
  or g_139850_(_050383_, _050507_, _050556_);
  and g_139851_(_050553_, _050556_, _050557_);
  or g_139852_(_050552_, _050554_, _050558_);
  and g_139853_(out[416], _050557_, _050559_);
  or g_139854_(_004740_, _050558_, _050560_);
  and g_139855_(_050551_, _050560_, _050561_);
  or g_139856_(_050550_, _050559_, _050562_);
  and g_139857_(_050547_, _050562_, _050563_);
  or g_139858_(_050546_, _050561_, _050564_);
  and g_139859_(_050538_, _050564_, _050565_);
  or g_139860_(_050537_, _050563_, _050567_);
  and g_139861_(_049864_, _050535_, _050568_);
  or g_139862_(_049863_, _050536_, _050569_);
  xor g_139863_(out[419], _038283_, _050570_);
  xor g_139864_(_053984_, _038283_, _050571_);
  or g_139865_(_050396_, _050508_, _050572_);
  not g_139866_(_050572_, _050573_);
  and g_139867_(_050404_, _050508_, _050574_);
  not g_139868_(_050574_, _050575_);
  and g_139869_(_050572_, _050575_, _050576_);
  or g_139870_(_050573_, _050574_, _050578_);
  and g_139871_(_050570_, _050578_, _050579_);
  or g_139872_(_050571_, _050576_, _050580_);
  and g_139873_(_050569_, _050580_, _050581_);
  or g_139874_(_050568_, _050579_, _050582_);
  and g_139875_(_050567_, _050581_, _050583_);
  or g_139876_(_050565_, _050582_, _050584_);
  xor g_139877_(out[420], _038284_, _050585_);
  and g_139878_(_050344_, _050507_, _050586_);
  and g_139879_(_050351_, _050508_, _050587_);
  or g_139880_(_050586_, _050587_, _050589_);
  or g_139881_(_050585_, _050589_, _050590_);
  or g_139882_(_050570_, _050578_, _050591_);
  and g_139883_(_050590_, _050591_, _050592_);
  not g_139884_(_050592_, _050593_);
  and g_139885_(_050584_, _050592_, _050594_);
  or g_139886_(_050583_, _050593_, _050595_);
  xor g_139887_(out[421], _038285_, _050596_);
  xor g_139888_(_053962_, _038285_, _050597_);
  or g_139889_(_050332_, _050508_, _050598_);
  not g_139890_(_050598_, _050600_);
  and g_139891_(_050340_, _050508_, _050601_);
  not g_139892_(_050601_, _050602_);
  and g_139893_(_050598_, _050602_, _050603_);
  or g_139894_(_050600_, _050601_, _050604_);
  and g_139895_(_050596_, _050604_, _050605_);
  and g_139896_(_050585_, _050589_, _050606_);
  or g_139897_(_050605_, _050606_, _050607_);
  not g_139898_(_050607_, _050608_);
  and g_139899_(_050595_, _050608_, _050609_);
  or g_139900_(_050594_, _050607_, _050611_);
  xor g_139901_(out[422], _038286_, _050612_);
  xor g_139902_(_053973_, _038286_, _050613_);
  and g_139903_(_050329_, _050508_, _050614_);
  not g_139904_(_050614_, _050615_);
  or g_139905_(_050322_, _050508_, _050616_);
  not g_139906_(_050616_, _050617_);
  and g_139907_(_050615_, _050616_, _050618_);
  or g_139908_(_050614_, _050617_, _050619_);
  and g_139909_(_050612_, _050618_, _050620_);
  or g_139910_(_050613_, _050619_, _050622_);
  and g_139911_(_050597_, _050603_, _050623_);
  or g_139912_(_050596_, _050604_, _050624_);
  and g_139913_(_050622_, _050624_, _050625_);
  or g_139914_(_050620_, _050623_, _050626_);
  and g_139915_(_050611_, _050625_, _050627_);
  or g_139916_(_050609_, _050626_, _050628_);
  xor g_139917_(out[423], _038287_, _050629_);
  not g_139918_(_050629_, _050630_);
  and g_139919_(_050318_, _050508_, _050631_);
  not g_139920_(_050631_, _050633_);
  or g_139921_(_050310_, _050508_, _050634_);
  not g_139922_(_050634_, _050635_);
  and g_139923_(_050633_, _050634_, _050636_);
  or g_139924_(_050631_, _050635_, _050637_);
  and g_139925_(_050629_, _050637_, _050638_);
  or g_139926_(_050630_, _050636_, _050639_);
  and g_139927_(_050613_, _050619_, _050640_);
  or g_139928_(_050612_, _050618_, _050641_);
  and g_139929_(_050639_, _050641_, _050642_);
  or g_139930_(_050638_, _050640_, _050644_);
  and g_139931_(_050628_, _050642_, _050645_);
  or g_139932_(_050627_, _050644_, _050646_);
  xor g_139933_(out[424], _038288_, _050647_);
  not g_139934_(_050647_, _050648_);
  and g_139935_(_050480_, _050508_, _050649_);
  not g_139936_(_050649_, _050650_);
  or g_139937_(_050472_, _050508_, _050651_);
  not g_139938_(_050651_, _050652_);
  and g_139939_(_050650_, _050651_, _050653_);
  or g_139940_(_050649_, _050652_, _050655_);
  and g_139941_(_050647_, _050655_, _050656_);
  or g_139942_(_050648_, _050653_, _050657_);
  xor g_139943_(out[425], _038289_, _050658_);
  xor g_139944_(_054028_, _038289_, _050659_);
  and g_139945_(_050462_, _050508_, _050660_);
  not g_139946_(_050660_, _050661_);
  or g_139947_(_050455_, _050508_, _050662_);
  not g_139948_(_050662_, _050663_);
  and g_139949_(_050661_, _050662_, _050664_);
  or g_139950_(_050660_, _050663_, _050666_);
  and g_139951_(_050658_, _050664_, _050667_);
  or g_139952_(_050659_, _050666_, _050668_);
  and g_139953_(_050630_, _050636_, _050669_);
  or g_139954_(_050629_, _050637_, _050670_);
  xor g_139955_(_050648_, _050653_, _050671_);
  xor g_139956_(_050647_, _050653_, _050672_);
  and g_139957_(_050670_, _050671_, _050673_);
  or g_139958_(_050669_, _050672_, _050674_);
  and g_139959_(_050668_, _050673_, _050675_);
  or g_139960_(_050667_, _050674_, _050677_);
  and g_139961_(_050646_, _050675_, _050678_);
  or g_139962_(_050645_, _050677_, _050679_);
  and g_139963_(_050659_, _050666_, _050680_);
  or g_139964_(_050658_, _050664_, _050681_);
  and g_139965_(_050656_, _050668_, _050682_);
  or g_139966_(_050657_, _050667_, _050683_);
  and g_139967_(_050681_, _050683_, _050684_);
  or g_139968_(_050680_, _050682_, _050685_);
  and g_139969_(_050679_, _050684_, _050686_);
  or g_139970_(_050678_, _050685_, _050688_);
  and g_139971_(_050530_, _050688_, _050689_);
  or g_139972_(_050531_, _050686_, _050690_);
  and g_139973_(_050519_, _050525_, _050691_);
  or g_139974_(_050520_, _050524_, _050692_);
  and g_139975_(_050523_, _050692_, _050693_);
  or g_139976_(_050521_, _050691_, _050694_);
  and g_139977_(_050690_, _050693_, _050695_);
  or g_139978_(_050689_, _050694_, _050696_);
  and g_139979_(_049863_, _050695_, _050697_);
  and g_139980_(_050535_, _050696_, _050699_);
  or g_139981_(_050697_, _050699_, _050700_);
  or g_139982_(_049861_, _050700_, _050701_);
  and g_139983_(_050548_, _050695_, _050702_);
  and g_139984_(_050545_, _050696_, _050703_);
  or g_139985_(_050702_, _050703_, _050704_);
  and g_139986_(out[433], _050704_, _050705_);
  xor g_139987_(_054116_, out[432], _050706_);
  not g_139988_(_050706_, _050707_);
  or g_139989_(_050704_, _050706_, _050708_);
  and g_139990_(out[416], _050695_, _050710_);
  and g_139991_(_050558_, _050696_, _050711_);
  or g_139992_(_050710_, _050711_, _050712_);
  not g_139993_(_050712_, _050713_);
  or g_139994_(_004773_, _050712_, _050714_);
  and g_139995_(_050708_, _050714_, _050715_);
  or g_139996_(_050705_, _050715_, _050716_);
  and g_139997_(_050701_, _050716_, _050717_);
  and g_139998_(_049861_, _050700_, _050718_);
  xor g_139999_(out[435], _038270_, _050719_);
  and g_140000_(_050578_, _050696_, _050721_);
  and g_140001_(_050571_, _050695_, _050722_);
  or g_140002_(_050721_, _050722_, _050723_);
  and g_140003_(_050719_, _050723_, _050724_);
  or g_140004_(_050718_, _050724_, _050725_);
  or g_140005_(_050717_, _050725_, _050726_);
  xor g_140006_(out[436], _038271_, _050727_);
  or g_140007_(_050585_, _050696_, _050728_);
  not g_140008_(_050728_, _050729_);
  and g_140009_(_050589_, _050696_, _050730_);
  or g_140010_(_050729_, _050730_, _050732_);
  not g_140011_(_050732_, _050733_);
  or g_140012_(_050727_, _050732_, _050734_);
  or g_140013_(_050719_, _050723_, _050735_);
  and g_140014_(_050734_, _050735_, _050736_);
  and g_140015_(_050726_, _050736_, _050737_);
  xor g_140016_(out[437], _038272_, _050738_);
  not g_140017_(_050738_, _050739_);
  or g_140018_(_050596_, _050696_, _050740_);
  not g_140019_(_050740_, _050741_);
  and g_140020_(_050604_, _050696_, _050743_);
  not g_140021_(_050743_, _050744_);
  and g_140022_(_050740_, _050744_, _050745_);
  or g_140023_(_050741_, _050743_, _050746_);
  and g_140024_(_050738_, _050746_, _050747_);
  and g_140025_(_050727_, _050732_, _050748_);
  or g_140026_(_050747_, _050748_, _050749_);
  or g_140027_(_050737_, _050749_, _050750_);
  not g_140028_(_050750_, _050751_);
  xor g_140029_(out[438], _038273_, _050752_);
  xor g_140030_(_054072_, _038273_, _050754_);
  and g_140031_(_050619_, _050696_, _050755_);
  not g_140032_(_050755_, _050756_);
  or g_140033_(_050613_, _050696_, _050757_);
  not g_140034_(_050757_, _050758_);
  and g_140035_(_050756_, _050757_, _050759_);
  or g_140036_(_050755_, _050758_, _050760_);
  and g_140037_(_050752_, _050759_, _050761_);
  or g_140038_(_050754_, _050760_, _050762_);
  and g_140039_(_050739_, _050745_, _050763_);
  or g_140040_(_050738_, _050746_, _050765_);
  and g_140041_(_050762_, _050765_, _050766_);
  or g_140042_(_050761_, _050763_, _050767_);
  and g_140043_(_050750_, _050766_, _050768_);
  or g_140044_(_050751_, _050767_, _050769_);
  xor g_140045_(out[439], _038274_, _050770_);
  xor g_140046_(_054039_, _038274_, _050771_);
  and g_140047_(_050637_, _050696_, _050772_);
  not g_140048_(_050772_, _050773_);
  or g_140049_(_050629_, _050696_, _050774_);
  not g_140050_(_050774_, _050776_);
  and g_140051_(_050773_, _050774_, _050777_);
  or g_140052_(_050772_, _050776_, _050778_);
  and g_140053_(_050770_, _050778_, _050779_);
  or g_140054_(_050771_, _050777_, _050780_);
  and g_140055_(_050754_, _050760_, _050781_);
  or g_140056_(_050752_, _050759_, _050782_);
  and g_140057_(_050780_, _050782_, _050783_);
  or g_140058_(_050779_, _050781_, _050784_);
  and g_140059_(_050769_, _050783_, _050785_);
  or g_140060_(_050768_, _050784_, _050787_);
  and g_140061_(_050771_, _050777_, _050788_);
  or g_140062_(_050770_, _050778_, _050789_);
  and g_140063_(_050515_, _050696_, _050790_);
  not g_140064_(_050790_, _050791_);
  or g_140065_(_049865_, _050696_, _050792_);
  not g_140066_(_050792_, _050793_);
  and g_140067_(_050791_, _050792_, _050794_);
  or g_140068_(_050790_, _050793_, _050795_);
  and g_140069_(_049860_, _050794_, _050796_);
  or g_140070_(_049859_, _050795_, _050798_);
  xor g_140071_(out[440], _038275_, _050799_);
  not g_140072_(_050799_, _050800_);
  and g_140073_(_050655_, _050696_, _050801_);
  not g_140074_(_050801_, _050802_);
  or g_140075_(_050647_, _050696_, _050803_);
  not g_140076_(_050803_, _050804_);
  and g_140077_(_050802_, _050803_, _050805_);
  or g_140078_(_050801_, _050804_, _050806_);
  or g_140079_(_050799_, _050806_, _050807_);
  or g_140080_(_049866_, _050696_, _050809_);
  or g_140081_(_050518_, _050695_, _050810_);
  and g_140082_(_050809_, _050810_, _050811_);
  and g_140083_(_049859_, _050811_, _050812_);
  or g_140084_(_049860_, _050794_, _050813_);
  and g_140085_(_038280_, _049849_, _050814_);
  or g_140086_(_038281_, _043319_, _050815_);
  and g_140087_(_050813_, _050815_, _050816_);
  or g_140088_(_050812_, _050814_, _050817_);
  xor g_140089_(out[441], _038276_, _050818_);
  and g_140090_(_050666_, _050696_, _050820_);
  not g_140091_(_050820_, _050821_);
  or g_140092_(_050659_, _050696_, _050822_);
  not g_140093_(_050822_, _050823_);
  and g_140094_(_050821_, _050822_, _050824_);
  or g_140095_(_050820_, _050823_, _050825_);
  or g_140096_(_050818_, _050824_, _050826_);
  and g_140097_(_038281_, _043319_, _050827_);
  or g_140098_(_038280_, _043320_, _050828_);
  and g_140099_(_050818_, _050824_, _050829_);
  or g_140100_(_050800_, _050805_, _050831_);
  or g_140101_(_050817_, _050827_, _050832_);
  not g_140102_(_050832_, _050833_);
  and g_140103_(_050798_, _050833_, _050834_);
  or g_140104_(_050796_, _050832_, _050835_);
  xor g_140105_(_050818_, _050824_, _050836_);
  xor g_140106_(_050818_, _050825_, _050837_);
  and g_140107_(_050789_, _050807_, _050838_);
  and g_140108_(_050836_, _050838_, _050839_);
  and g_140109_(_050834_, _050839_, _050840_);
  and g_140110_(_050831_, _050840_, _050842_);
  xor g_140111_(_050799_, _050805_, _050843_);
  or g_140112_(_050788_, _050837_, _050844_);
  or g_140113_(_050835_, _050844_, _050845_);
  or g_140114_(_050785_, _050845_, _050846_);
  and g_140115_(_050787_, _050842_, _050847_);
  or g_140116_(_050843_, _050846_, _050848_);
  and g_140117_(_050826_, _050831_, _050849_);
  or g_140118_(_050829_, _050849_, _050850_);
  not g_140119_(_050850_, _050851_);
  and g_140120_(_050798_, _050851_, _050853_);
  or g_140121_(_050796_, _050850_, _050854_);
  and g_140122_(_050816_, _050854_, _050855_);
  or g_140123_(_050817_, _050853_, _050856_);
  and g_140124_(_050828_, _050856_, _050857_);
  or g_140125_(_050827_, _050855_, _050858_);
  and g_140126_(_050848_, _050858_, _050859_);
  or g_140127_(_050847_, _050857_, _050860_);
  or g_140128_(_049859_, _050860_, _050861_);
  or g_140129_(_050794_, _050859_, _050862_);
  and g_140130_(_050861_, _050862_, _050864_);
  and g_140131_(_049856_, _050864_, _050865_);
  not g_140132_(_050865_, _050866_);
  and g_140133_(_049858_, _050866_, _050867_);
  or g_140134_(_049857_, _050865_, _050868_);
  and g_140135_(_038266_, _049850_, _050869_);
  or g_140136_(_038267_, _043321_, _050870_);
  or g_140137_(_049860_, _050860_, _050871_);
  or g_140138_(_050811_, _050859_, _050872_);
  and g_140139_(_050871_, _050872_, _050873_);
  and g_140140_(_049855_, _050873_, _050875_);
  or g_140141_(_049856_, _050864_, _050876_);
  and g_140142_(_050870_, _050876_, _050877_);
  or g_140143_(_050869_, _050875_, _050878_);
  xor g_140144_(out[457], _038263_, _050879_);
  xor g_140145_(_054226_, _038263_, _050880_);
  and g_140146_(_050818_, _050859_, _050881_);
  not g_140147_(_050881_, _050882_);
  or g_140148_(_050824_, _050859_, _050883_);
  not g_140149_(_050883_, _050884_);
  and g_140150_(_050882_, _050883_, _050886_);
  or g_140151_(_050881_, _050884_, _050887_);
  and g_140152_(_050880_, _050887_, _050888_);
  or g_140153_(_050879_, _050886_, _050889_);
  and g_140154_(_050877_, _050889_, _050890_);
  or g_140155_(_050878_, _050888_, _050891_);
  and g_140156_(_050867_, _050890_, _050892_);
  or g_140157_(_050868_, _050891_, _050893_);
  xor g_140158_(out[456], _038262_, _050894_);
  xor g_140159_(_054149_, _038262_, _050895_);
  and g_140160_(_050806_, _050860_, _050897_);
  and g_140161_(_050800_, _050859_, _050898_);
  or g_140162_(_050897_, _050898_, _050899_);
  not g_140163_(_050899_, _050900_);
  and g_140164_(_050895_, _050900_, _050901_);
  or g_140165_(_050894_, _050899_, _050902_);
  and g_140166_(_050879_, _050886_, _050903_);
  not g_140167_(_050903_, _050904_);
  and g_140168_(_050902_, _050904_, _050905_);
  or g_140169_(_050901_, _050903_, _050906_);
  and g_140170_(_050894_, _050899_, _050908_);
  or g_140171_(_050895_, _050900_, _050909_);
  or g_140172_(_050906_, _050908_, _050910_);
  and g_140173_(_050892_, _050909_, _050911_);
  and g_140174_(_050905_, _050911_, _050912_);
  or g_140175_(_050893_, _050910_, _050913_);
  xor g_140176_(out[454], _038260_, _050914_);
  xor g_140177_(_054171_, _038260_, _050915_);
  and g_140178_(_050752_, _050859_, _050916_);
  or g_140179_(_050754_, _050860_, _050917_);
  and g_140180_(_050760_, _050860_, _050919_);
  or g_140181_(_050759_, _050859_, _050920_);
  and g_140182_(_050917_, _050920_, _050921_);
  or g_140183_(_050916_, _050919_, _050922_);
  and g_140184_(_050914_, _050921_, _050923_);
  or g_140185_(_050915_, _050922_, _050924_);
  xor g_140186_(out[455], _038261_, _050925_);
  not g_140187_(_050925_, _050926_);
  and g_140188_(_050771_, _050859_, _050927_);
  or g_140189_(_050770_, _050860_, _050928_);
  and g_140190_(_050778_, _050860_, _050930_);
  or g_140191_(_050777_, _050859_, _050931_);
  and g_140192_(_050928_, _050931_, _050932_);
  or g_140193_(_050927_, _050930_, _050933_);
  and g_140194_(_050926_, _050932_, _050934_);
  or g_140195_(_050925_, _050933_, _050935_);
  and g_140196_(_050924_, _050935_, _050936_);
  or g_140197_(_050923_, _050934_, _050937_);
  or g_140198_(_050926_, _050932_, _050938_);
  or g_140199_(_050914_, _050921_, _050939_);
  and g_140200_(_050938_, _050939_, _050941_);
  not g_140201_(_050941_, _050942_);
  and g_140202_(_050936_, _050941_, _050943_);
  or g_140203_(_050937_, _050942_, _050944_);
  xor g_140204_(out[452], _038258_, _050945_);
  not g_140205_(_050945_, _050946_);
  or g_140206_(_050727_, _050860_, _050947_);
  or g_140207_(_050733_, _050859_, _050948_);
  and g_140208_(_050947_, _050948_, _050949_);
  not g_140209_(_050949_, _050950_);
  and g_140210_(_050946_, _050949_, _050952_);
  or g_140211_(_050945_, _050950_, _050953_);
  xor g_140212_(out[453], _038259_, _050954_);
  not g_140213_(_050954_, _050955_);
  or g_140214_(_050745_, _050859_, _050956_);
  or g_140215_(_050738_, _050860_, _050957_);
  and g_140216_(_050956_, _050957_, _050958_);
  not g_140217_(_050958_, _050959_);
  and g_140218_(_050955_, _050958_, _050960_);
  or g_140219_(_050954_, _050959_, _050961_);
  and g_140220_(_050953_, _050961_, _050963_);
  or g_140221_(_050952_, _050960_, _050964_);
  and g_140222_(_050954_, _050959_, _050965_);
  or g_140223_(_050955_, _050958_, _050966_);
  and g_140224_(_050945_, _050950_, _050967_);
  or g_140225_(_050946_, _050949_, _050968_);
  and g_140226_(_050966_, _050968_, _050969_);
  or g_140227_(_050965_, _050967_, _050970_);
  and g_140228_(_050963_, _050969_, _050971_);
  or g_140229_(_050964_, _050970_, _050972_);
  and g_140230_(_050943_, _050971_, _050974_);
  or g_140231_(_050944_, _050972_, _050975_);
  and g_140232_(_050912_, _050974_, _050976_);
  or g_140233_(_050913_, _050975_, _050977_);
  xor g_140234_(out[451], _038256_, _050978_);
  xor g_140235_(_054182_, _038256_, _050979_);
  and g_140236_(_050719_, _050859_, _050980_);
  or g_140237_(_050723_, _050859_, _050981_);
  not g_140238_(_050981_, _050982_);
  or g_140239_(_050980_, _050982_, _050983_);
  not g_140240_(_050983_, _050985_);
  and g_140241_(_050979_, _050983_, _050986_);
  or g_140242_(_050978_, _050985_, _050987_);
  xor g_140243_(out[450], _038255_, _050988_);
  not g_140244_(_050988_, _050989_);
  or g_140245_(_050700_, _050859_, _050990_);
  and g_140246_(_049861_, _050859_, _050991_);
  not g_140247_(_050991_, _050992_);
  and g_140248_(_050990_, _050992_, _050993_);
  not g_140249_(_050993_, _050994_);
  and g_140250_(_050988_, _050994_, _050996_);
  or g_140251_(_050989_, _050993_, _050997_);
  and g_140252_(_050987_, _050997_, _050998_);
  or g_140253_(_050986_, _050996_, _050999_);
  and g_140254_(_050978_, _050985_, _051000_);
  or g_140255_(_050979_, _050983_, _051001_);
  xor g_140256_(_050978_, _050983_, _051002_);
  xor g_140257_(_050988_, _050993_, _051003_);
  or g_140258_(_051002_, _051003_, _051004_);
  not g_140259_(_051004_, _051005_);
  xor g_140260_(out[449], out[448], _051007_);
  not g_140261_(_051007_, _051008_);
  and g_140262_(_050707_, _050859_, _051009_);
  not g_140263_(_051009_, _051010_);
  and g_140264_(_050704_, _050860_, _051011_);
  not g_140265_(_051011_, _051012_);
  and g_140266_(_051010_, _051012_, _051013_);
  or g_140267_(_051009_, _051011_, _051014_);
  and g_140268_(_051007_, _051013_, _051015_);
  or g_140269_(_051008_, _051014_, _051016_);
  or g_140270_(_004773_, _050860_, _051018_);
  or g_140271_(_050713_, _050859_, _051019_);
  and g_140272_(_051018_, _051019_, _051020_);
  not g_140273_(_051020_, _051021_);
  or g_140274_(out[448], _051020_, _051022_);
  not g_140275_(_051022_, _051023_);
  xor g_140276_(_051008_, _051014_, _051024_);
  xor g_140277_(_051007_, _051014_, _051025_);
  and g_140278_(_051022_, _051024_, _051026_);
  or g_140279_(_051023_, _051025_, _051027_);
  and g_140280_(_051016_, _051027_, _051029_);
  or g_140281_(_051015_, _051026_, _051030_);
  and g_140282_(_051005_, _051030_, _051031_);
  or g_140283_(_051004_, _051029_, _051032_);
  and g_140284_(_050999_, _051001_, _051033_);
  or g_140285_(_050998_, _051000_, _051034_);
  and g_140286_(_051032_, _051034_, _051035_);
  or g_140287_(_051031_, _051033_, _051036_);
  and g_140288_(_050976_, _051036_, _051037_);
  or g_140289_(_050977_, _051035_, _051038_);
  and g_140290_(_050964_, _050966_, _051040_);
  or g_140291_(_050963_, _050965_, _051041_);
  and g_140292_(_050943_, _051040_, _051042_);
  or g_140293_(_050944_, _051041_, _051043_);
  and g_140294_(_050937_, _050938_, _051044_);
  not g_140295_(_051044_, _051045_);
  and g_140296_(_051043_, _051045_, _051046_);
  or g_140297_(_051042_, _051044_, _051047_);
  and g_140298_(_050912_, _051047_, _051048_);
  or g_140299_(_050913_, _051046_, _051049_);
  and g_140300_(_050892_, _050906_, _051051_);
  and g_140301_(_050868_, _050870_, _051052_);
  or g_140302_(_051051_, _051052_, _051053_);
  not g_140303_(_051053_, _051054_);
  and g_140304_(_051049_, _051054_, _051055_);
  or g_140305_(_051048_, _051053_, _051056_);
  and g_140306_(_051038_, _051055_, _051057_);
  or g_140307_(_051037_, _051056_, _051058_);
  and g_140308_(out[448], _051020_, _051059_);
  or g_140309_(_051004_, _051059_, _051060_);
  or g_140310_(_051027_, _051060_, _051062_);
  or g_140311_(_050977_, _051062_, _051063_);
  not g_140312_(_051063_, _051064_);
  and g_140313_(_051058_, _051063_, _051065_);
  or g_140314_(_051057_, _051064_, _051066_);
  or g_140315_(_049855_, _051066_, _051067_);
  or g_140316_(_050864_, _051065_, _051068_);
  and g_140317_(_051067_, _051068_, _051069_);
  not g_140318_(_051069_, _051070_);
  xor g_140319_(out[474], _038251_, _051071_);
  not g_140320_(_051071_, _051073_);
  and g_140321_(_038254_, _043323_, _051074_);
  or g_140322_(_038253_, _043324_, _051075_);
  or g_140323_(_051073_, _051074_, _051076_);
  or g_140324_(_051069_, _051076_, _051077_);
  or g_140325_(_050873_, _051065_, _051078_);
  or g_140326_(_049856_, _051066_, _051079_);
  and g_140327_(_051078_, _051079_, _051080_);
  and g_140328_(_051071_, _051080_, _051081_);
  or g_140329_(_049853_, _051081_, _051082_);
  and g_140330_(_049854_, _051077_, _051084_);
  and g_140331_(_051075_, _051082_, _051085_);
  and g_140332_(out[448], _051065_, _051086_);
  or g_140333_(_004806_, _051066_, _051087_);
  and g_140334_(_051021_, _051066_, _051088_);
  or g_140335_(_051020_, _051065_, _051089_);
  and g_140336_(_051087_, _051089_, _051090_);
  or g_140337_(_051086_, _051088_, _051091_);
  and g_140338_(out[464], _051090_, _051092_);
  or g_140339_(_004839_, _051091_, _051093_);
  and g_140340_(_051007_, _051065_, _051095_);
  or g_140341_(_051008_, _051066_, _051096_);
  and g_140342_(_051014_, _051066_, _051097_);
  or g_140343_(_051013_, _051065_, _051098_);
  and g_140344_(_051096_, _051098_, _051099_);
  or g_140345_(_051095_, _051097_, _051100_);
  and g_140346_(out[465], _051100_, _051101_);
  or g_140347_(_054314_, _051099_, _051102_);
  xor g_140348_(out[465], out[464], _051103_);
  not g_140349_(_051103_, _051104_);
  and g_140350_(_051092_, _051102_, _051106_);
  or g_140351_(_051093_, _051101_, _051107_);
  xor g_140352_(out[466], _038242_, _051108_);
  not g_140353_(_051108_, _051109_);
  and g_140354_(_050988_, _051065_, _051110_);
  and g_140355_(_050993_, _051066_, _051111_);
  or g_140356_(_051110_, _051111_, _051112_);
  not g_140357_(_051112_, _051113_);
  and g_140358_(_051108_, _051113_, _051114_);
  or g_140359_(_051109_, _051112_, _051115_);
  or g_140360_(_051100_, _051104_, _051117_);
  not g_140361_(_051117_, _051118_);
  and g_140362_(_051115_, _051117_, _051119_);
  or g_140363_(_051106_, _051118_, _051120_);
  and g_140364_(_051107_, _051119_, _051121_);
  or g_140365_(_051114_, _051120_, _051122_);
  xor g_140366_(_054281_, _038243_, _051123_);
  or g_140367_(_050978_, _051066_, _051124_);
  or g_140368_(_050983_, _051065_, _051125_);
  and g_140369_(_051124_, _051125_, _051126_);
  or g_140370_(_051123_, _051126_, _051128_);
  not g_140371_(_051128_, _051129_);
  and g_140372_(_051109_, _051112_, _051130_);
  or g_140373_(_051108_, _051113_, _051131_);
  and g_140374_(_051128_, _051131_, _051132_);
  or g_140375_(_051129_, _051130_, _051133_);
  and g_140376_(_051122_, _051132_, _051134_);
  or g_140377_(_051121_, _051133_, _051135_);
  xor g_140378_(out[468], _038244_, _051136_);
  xor g_140379_(_054292_, _038244_, _051137_);
  or g_140380_(_050945_, _051066_, _051139_);
  or g_140381_(_050949_, _051065_, _051140_);
  and g_140382_(_051139_, _051140_, _051141_);
  not g_140383_(_051141_, _051142_);
  and g_140384_(_051137_, _051141_, _051143_);
  and g_140385_(_051123_, _051126_, _051144_);
  or g_140386_(_051143_, _051144_, _051145_);
  not g_140387_(_051145_, _051146_);
  and g_140388_(_051135_, _051146_, _051147_);
  or g_140389_(_051134_, _051145_, _051148_);
  or g_140390_(_050954_, _051066_, _051150_);
  or g_140391_(_050958_, _051065_, _051151_);
  and g_140392_(_051150_, _051151_, _051152_);
  not g_140393_(_051152_, _051153_);
  and g_140394_(_049834_, _051153_, _051154_);
  or g_140395_(_049835_, _051152_, _051155_);
  and g_140396_(_051136_, _051142_, _051156_);
  or g_140397_(_051137_, _051141_, _051157_);
  and g_140398_(_051155_, _051157_, _051158_);
  or g_140399_(_051154_, _051156_, _051159_);
  and g_140400_(_051148_, _051158_, _051161_);
  or g_140401_(_051147_, _051159_, _051162_);
  xor g_140402_(out[470], _038247_, _051163_);
  xor g_140403_(_054270_, _038247_, _051164_);
  or g_140404_(_050915_, _051066_, _051165_);
  or g_140405_(_050921_, _051065_, _051166_);
  and g_140406_(_051165_, _051166_, _051167_);
  not g_140407_(_051167_, _051168_);
  and g_140408_(_051163_, _051167_, _051169_);
  or g_140409_(_051164_, _051168_, _051170_);
  and g_140410_(_049835_, _051152_, _051172_);
  or g_140411_(_049834_, _051153_, _051173_);
  and g_140412_(_051170_, _051173_, _051174_);
  or g_140413_(_051169_, _051172_, _051175_);
  and g_140414_(_051162_, _051174_, _051176_);
  or g_140415_(_051161_, _051175_, _051177_);
  xor g_140416_(out[471], _038248_, _051178_);
  not g_140417_(_051178_, _051179_);
  or g_140418_(_050925_, _051066_, _051180_);
  or g_140419_(_050932_, _051065_, _051181_);
  and g_140420_(_051180_, _051181_, _051183_);
  not g_140421_(_051183_, _051184_);
  and g_140422_(_051178_, _051184_, _051185_);
  or g_140423_(_051179_, _051183_, _051186_);
  and g_140424_(_051164_, _051168_, _051187_);
  or g_140425_(_051163_, _051167_, _051188_);
  and g_140426_(_051186_, _051188_, _051189_);
  or g_140427_(_051185_, _051187_, _051190_);
  and g_140428_(_051177_, _051189_, _051191_);
  or g_140429_(_051176_, _051190_, _051192_);
  and g_140430_(_051179_, _051183_, _051194_);
  or g_140431_(_051178_, _051184_, _051195_);
  xor g_140432_(out[472], _038249_, _051196_);
  xor g_140433_(_054248_, _038249_, _051197_);
  and g_140434_(_050895_, _051065_, _051198_);
  and g_140435_(_050899_, _051066_, _051199_);
  or g_140436_(_051198_, _051199_, _051200_);
  not g_140437_(_051200_, _051201_);
  and g_140438_(_051197_, _051201_, _051202_);
  or g_140439_(_051196_, _051200_, _051203_);
  and g_140440_(_051195_, _051203_, _051205_);
  or g_140441_(_051194_, _051202_, _051206_);
  and g_140442_(_051196_, _051200_, _051207_);
  or g_140443_(_051197_, _051201_, _051208_);
  xor g_140444_(out[473], _038250_, _051209_);
  xor g_140445_(_054325_, _038250_, _051210_);
  or g_140446_(_050880_, _051066_, _051211_);
  or g_140447_(_050886_, _051065_, _051212_);
  and g_140448_(_051211_, _051212_, _051213_);
  not g_140449_(_051213_, _051214_);
  and g_140450_(_051209_, _051213_, _051216_);
  or g_140451_(_051210_, _051214_, _051217_);
  and g_140452_(_051208_, _051217_, _051218_);
  or g_140453_(_051207_, _051216_, _051219_);
  and g_140454_(_051205_, _051218_, _051220_);
  or g_140455_(_051206_, _051219_, _051221_);
  and g_140456_(_051192_, _051220_, _051222_);
  or g_140457_(_051191_, _051221_, _051223_);
  and g_140458_(_051210_, _051214_, _051224_);
  or g_140459_(_051209_, _051213_, _051225_);
  and g_140460_(_051207_, _051217_, _051227_);
  or g_140461_(_051208_, _051216_, _051228_);
  and g_140462_(_051225_, _051228_, _051229_);
  or g_140463_(_051224_, _051227_, _051230_);
  and g_140464_(_051223_, _051229_, _051231_);
  or g_140465_(_051222_, _051230_, _051232_);
  and g_140466_(_051069_, _051073_, _051233_);
  or g_140467_(_051070_, _051071_, _051234_);
  and g_140468_(_051075_, _051234_, _051235_);
  or g_140469_(_051074_, _051233_, _051236_);
  and g_140470_(_051232_, _051235_, _051238_);
  or g_140471_(_051231_, _051236_, _051239_);
  and g_140472_(_051084_, _051239_, _051240_);
  or g_140473_(_051085_, _051238_, _051241_);
  or g_140474_(_049834_, _051241_, _051242_);
  or g_140475_(_051152_, _051240_, _051243_);
  and g_140476_(_051242_, _051243_, _051244_);
  or g_140477_(_049660_, _049833_, _051245_);
  or g_140478_(_049663_, _049832_, _051246_);
  and g_140479_(_051245_, _051246_, _051247_);
  or g_140480_(_049794_, _049832_, _051249_);
  or g_140481_(_049788_, _049833_, _051250_);
  and g_140482_(_051249_, _051250_, _051251_);
  or g_140483_(_051141_, _051240_, _051252_);
  or g_140484_(_051136_, _051241_, _051253_);
  and g_140485_(_051252_, _051253_, _051254_);
  or g_140486_(_049722_, _049833_, _051255_);
  or g_140487_(_049726_, _049832_, _051256_);
  and g_140488_(_051255_, _051256_, _051257_);
  xor g_140489_(_051254_, _051257_, _051258_);
  and g_140490_(out[464], _051240_, _051260_);
  and g_140491_(_051091_, _051241_, _051261_);
  or g_140492_(_051260_, _051261_, _051262_);
  or g_140493_(_002232_, _049833_, _051263_);
  or g_140494_(_049682_, _049832_, _051264_);
  and g_140495_(_051263_, _051264_, _051265_);
  xor g_140496_(_051262_, _051265_, _051266_);
  or g_140497_(_051126_, _051240_, _051267_);
  and g_140498_(_051123_, _051240_, _051268_);
  not g_140499_(_051268_, _051269_);
  and g_140500_(_051267_, _051269_, _051271_);
  and g_140501_(_049706_, _049832_, _051272_);
  not g_140502_(_051272_, _051273_);
  or g_140503_(_049710_, _049832_, _051274_);
  and g_140504_(_051273_, _051274_, _051275_);
  xor g_140505_(_051271_, _051275_, _051276_);
  or g_140506_(_051210_, _051241_, _051277_);
  or g_140507_(_051213_, _051240_, _051278_);
  and g_140508_(_051277_, _051278_, _051279_);
  or g_140509_(_049775_, _049832_, _051280_);
  or g_140510_(_049770_, _049833_, _051282_);
  and g_140511_(_051280_, _051282_, _051283_);
  or g_140512_(_051178_, _051241_, _051284_);
  or g_140513_(_051183_, _051240_, _051285_);
  and g_140514_(_051284_, _051285_, _051286_);
  or g_140515_(_049745_, _049833_, _051287_);
  or g_140516_(_049748_, _049832_, _051288_);
  and g_140517_(_051287_, _051288_, _051289_);
  and g_140518_(_051197_, _051240_, _051290_);
  and g_140519_(_051200_, _051241_, _051291_);
  or g_140520_(_051290_, _051291_, _051293_);
  or g_140521_(_049764_, _049832_, _051294_);
  or g_140522_(_049759_, _049833_, _051295_);
  and g_140523_(_051294_, _051295_, _051296_);
  and g_140524_(_051108_, _051240_, _051297_);
  and g_140525_(_051112_, _051241_, _051298_);
  or g_140526_(_051297_, _051298_, _051299_);
  or g_140527_(_049695_, _049832_, _051300_);
  or g_140528_(_049690_, _049833_, _051301_);
  and g_140529_(_051300_, _051301_, _051302_);
  and g_140530_(_051103_, _051240_, _051304_);
  and g_140531_(_051100_, _051241_, _051305_);
  or g_140532_(_051304_, _051305_, _051306_);
  or g_140533_(_049673_, _049833_, _051307_);
  or g_140534_(_049671_, _049832_, _051308_);
  and g_140535_(_051307_, _051308_, _051309_);
  or g_140536_(_051164_, _051241_, _051310_);
  or g_140537_(_051167_, _051240_, _051311_);
  and g_140538_(_051310_, _051311_, _051312_);
  or g_140539_(_049655_, _049832_, _051313_);
  or g_140540_(_043338_, _049833_, _051315_);
  and g_140541_(_051313_, _051315_, _051316_);
  xor g_140542_(_051312_, _051316_, _051317_);
  xor g_140543_(_051244_, _051247_, _051318_);
  xor g_140544_(_051293_, _051296_, _051319_);
  xor g_140545_(_051279_, _051283_, _051320_);
  xor g_140546_(_051299_, _051302_, _051321_);
  xor g_140547_(_051306_, _051309_, _051322_);
  and g_140548_(_051317_, _051318_, _051323_);
  and g_140549_(_051322_, _051323_, _051324_);
  and g_140550_(_051258_, _051320_, _051326_);
  and g_140551_(_051276_, _051326_, _051327_);
  and g_140552_(_051324_, _051327_, _051328_);
  xor g_140553_(_051286_, _051289_, _051329_);
  and g_140554_(_051319_, _051329_, _051330_);
  or g_140555_(_051073_, _051241_, _051331_);
  or g_140556_(_051080_, _051240_, _051332_);
  and g_140557_(_051331_, _051332_, _051333_);
  xor g_140558_(_051251_, _051333_, _051334_);
  and g_140559_(_051330_, _051334_, _051335_);
  and g_140560_(_051266_, _051321_, _051337_);
  or g_140561_(_038254_, _049852_, _051338_);
  and g_140562_(_049802_, _049833_, _051339_);
  and g_140563_(_043336_, _049832_, _051340_);
  or g_140564_(_051339_, _051340_, _051341_);
  xor g_140565_(_051338_, _051341_, _051342_);
  and g_140566_(_051337_, _051342_, _051343_);
  and g_140567_(_051335_, _051343_, _051344_);
  and g_140568_(_051328_, _051344_, _051345_);
  and g_140569_(_038241_, _051345_, _051346_);
  or g_140570_(_038241_, _051345_, _051348_);
  xor g_140571_(_038241_, _051345_, _051349_);
  xor g_140572_(_027659_, _051349_, _051350_);
  xor g_140573_(_027658_, _051349_, _051351_);
  and g_140574_(_015554_, _051350_, _051352_);
  and g_140575_(_015555_, _051351_, _051353_);
  not g_140576_(_051353_, _051354_);
  xor g_140577_(_015554_, _051350_, _051355_);
  xor g_140578_(_003120_, _051355_, out[960]);
  or g_140579_(_027659_, _051346_, _051356_);
  and g_140580_(_051348_, _051356_, _051358_);
  or g_140581_(_003120_, _051352_, _051359_);
  and g_140582_(_051354_, _051359_, _051360_);
  and g_140583_(_051358_, _051360_, out[962]);
  xor g_140584_(_051358_, _051360_, out[961]);
  czero b_0_(out[974]);
  czero b_1_(out[973]);
  czero b_2_(out[972]);
  czero b_3_(out[971]);
  czero b_4_(out[970]);
  czero b_5_(out[969]);
  czero b_6_(out[968]);
  czero b_7_(out[967]);
  czero b_8_(out[966]);
  czero b_9_(out[965]);
  czero b_10_(out[970]);
  buf b_11_(set1[432], out[912]);
  buf b_12_(set1[341], out[821]);
  buf b_13_(set2[31], out[31]);
  buf b_14_(set2[94], out[94]);
  buf b_15_(set1[92], out[572]);
  buf b_16_(set1[164], out[644]);
  buf b_17_(set1[317], out[797]);
  buf b_18_(set1[340], out[820]);
  buf b_19_(set2[309], out[309]);
  buf b_20_(set1[458], out[938]);
  buf b_21_(set2[26], out[26]);
  buf b_22_(set2[285], out[285]);
  buf b_23_(set2[470], out[470]);
  buf b_24_(set1[61], out[541]);
  buf b_25_(set2[452], out[452]);
  buf b_26_(set1[277], out[757]);
  buf b_27_(set2[204], out[204]);
  buf b_28_(set2[446], out[446]);
  buf b_29_(set2[290], out[290]);
  buf b_30_(set2[40], out[40]);
  buf b_31_(set1[447], out[927]);
  buf b_32_(set1[188], out[668]);
  buf b_33_(set2[326], out[326]);
  buf b_34_(set2[352], out[352]);
  buf b_35_(set1[59], out[539]);
  buf b_36_(set2[272], out[272]);
  buf b_37_(set1[283], out[763]);
  buf b_38_(set2[107], out[107]);
  buf b_39_(set1[184], out[664]);
  buf b_40_(set2[353], out[353]);
  buf b_41_(set1[154], out[634]);
  buf b_42_(set1[58], out[538]);
  buf b_43_(set2[410], out[410]);
  buf b_44_(set1[450], out[930]);
  buf b_45_(set2[424], out[424]);
  buf b_46_(set2[280], out[280]);
  buf b_47_(set2[173], out[173]);
  buf b_48_(set2[228], out[228]);
  buf b_49_(set1[134], out[614]);
  buf b_50_(set2[115], out[115]);
  czero b_51_(out[963]);
  buf b_52_(set1[147], out[627]);
  buf b_53_(set1[388], out[868]);
  buf b_54_(set2[82], out[82]);
  buf b_55_(set1[457], out[937]);
  buf b_56_(set2[46], out[46]);
  buf b_57_(set2[44], out[44]);
  buf b_58_(set2[229], out[229]);
  buf b_59_(set2[209], out[209]);
  buf b_60_(set1[409], out[889]);
  buf b_61_(set1[270], out[750]);
  buf b_62_(set1[53], out[533]);
  buf b_63_(set1[473], out[953]);
  buf b_64_(set2[235], out[235]);
  buf b_65_(set2[35], out[35]);
  buf b_66_(set2[51], out[51]);
  buf b_67_(set1[195], out[675]);
  buf b_68_(set2[93], out[93]);
  buf b_69_(set1[404], out[884]);
  buf b_70_(set2[105], out[105]);
  buf b_71_(set1[374], out[854]);
  buf b_72_(set2[129], out[129]);
  buf b_73_(set2[170], out[170]);
  buf b_74_(set2[186], out[186]);
  buf b_75_(set1[379], out[859]);
  buf b_76_(set2[421], out[421]);
  buf b_77_(set2[251], out[251]);
  buf b_78_(set2[96], out[96]);
  buf b_79_(set1[181], out[661]);
  buf b_80_(set2[274], out[274]);
  buf b_81_(set1[167], out[647]);
  buf b_82_(set1[135], out[615]);
  buf b_83_(set1[299], out[779]);
  buf b_84_(set1[149], out[629]);
  buf b_85_(set1[470], out[950]);
  buf b_86_(set2[298], out[298]);
  buf b_87_(set2[238], out[238]);
  buf b_88_(set2[224], out[224]);
  buf b_89_(set2[183], out[183]);
  buf b_90_(set1[32], out[512]);
  buf b_91_(set1[67], out[547]);
  buf b_92_(set1[122], out[602]);
  czero b_93_(out[974]);
  buf b_94_(set1[419], out[899]);
  buf b_95_(set2[474], out[474]);
  buf b_96_(set1[336], out[816]);
  buf b_97_(set1[253], out[733]);
  buf b_98_(set2[350], out[350]);
  buf b_99_(set1[148], out[628]);
  buf b_100_(set1[227], out[707]);
  buf b_101_(set2[283], out[283]);
  buf b_102_(set2[125], out[125]);
  czero b_103_(out[964]);
  buf b_104_(set1[175], out[655]);
  buf b_105_(set1[23], out[503]);
  buf b_106_(set2[351], out[351]);
  buf b_107_(set1[151], out[631]);
  buf b_108_(set2[367], out[367]);
  buf b_109_(set2[136], out[136]);
  buf b_110_(set2[165], out[165]);
  buf b_111_(set1[49], out[529]);
  buf b_112_(set2[390], out[390]);
  buf b_113_(set2[258], out[258]);
  buf b_114_(set1[75], out[555]);
  buf b_115_(set1[267], out[747]);
  buf b_116_(set2[154], out[154]);
  buf b_117_(set2[210], out[210]);
  buf b_118_(set2[287], out[287]);
  buf b_119_(set1[256], out[736]);
  buf b_120_(set2[479], out[479]);
  buf b_121_(set2[69], out[69]);
  buf b_122_(set1[98], out[578]);
  buf b_123_(set2[341], out[341]);
  buf b_124_(set1[133], out[613]);
  buf b_125_(set2[260], out[260]);
  buf b_126_(set1[290], out[770]);
  buf b_127_(set2[412], out[412]);
  buf b_128_(set1[165], out[645]);
  buf b_129_(set2[132], out[132]);
  buf b_130_(set2[180], out[180]);
  buf b_131_(set1[315], out[795]);
  buf b_132_(set2[118], out[118]);
  buf b_133_(set2[244], out[244]);
  buf b_134_(set1[334], out[814]);
  buf b_135_(set1[6], out[486]);
  buf b_136_(set1[116], out[596]);
  buf b_137_(set1[251], out[731]);
  buf b_138_(set1[348], out[828]);
  buf b_139_(set1[7], out[487]);
  buf b_140_(set2[414], out[414]);
  buf b_141_(set1[180], out[660]);
  buf b_142_(set1[124], out[604]);
  buf b_143_(set1[51], out[531]);
  buf b_144_(set1[179], out[659]);
  buf b_145_(set2[162], out[162]);
  buf b_146_(set1[130], out[610]);
  buf b_147_(set1[249], out[729]);
  buf b_148_(set2[380], out[380]);
  buf b_149_(set2[9], out[9]);
  buf b_150_(set1[220], out[700]);
  buf b_151_(set2[357], out[357]);
  buf b_152_(set2[192], out[192]);
  buf b_153_(set2[432], out[432]);
  buf b_154_(set2[208], out[208]);
  buf b_155_(set1[178], out[658]);
  buf b_156_(set1[361], out[841]);
  buf b_157_(set1[319], out[799]);
  buf b_158_(set1[434], out[914]);
  buf b_159_(set2[319], out[319]);
  buf b_160_(set1[132], out[612]);
  buf b_161_(set1[60], out[540]);
  buf b_162_(set1[398], out[878]);
  buf b_163_(set2[85], out[85]);
  buf b_164_(set1[97], out[577]);
  buf b_165_(set2[249], out[249]);
  buf b_166_(set2[84], out[84]);
  buf b_167_(set1[390], out[870]);
  buf b_168_(set2[72], out[72]);
  buf b_169_(set2[471], out[471]);
  buf b_170_(set1[187], out[667]);
  buf b_171_(set2[294], out[294]);
  buf b_172_(set1[369], out[849]);
  buf b_173_(set2[18], out[18]);
  buf b_174_(set1[197], out[677]);
  buf b_175_(set1[265], out[745]);
  buf b_176_(set1[320], out[800]);
  buf b_177_(set2[425], out[425]);
  buf b_178_(set1[5], out[485]);
  buf b_179_(set2[216], out[216]);
  buf b_180_(set2[130], out[130]);
  buf b_181_(set2[218], out[218]);
  buf b_182_(set2[20], out[20]);
  buf b_183_(set1[465], out[945]);
  buf b_184_(set2[41], out[41]);
  buf b_185_(set1[99], out[579]);
  buf b_186_(set2[413], out[413]);
  buf b_187_(set1[308], out[788]);
  buf b_188_(set2[318], out[318]);
  buf b_189_(set2[196], out[196]);
  buf b_190_(set1[426], out[906]);
  buf b_191_(set2[174], out[174]);
  buf b_192_(set2[215], out[215]);
  buf b_193_(set1[69], out[549]);
  buf b_194_(set2[159], out[159]);
  buf b_195_(set1[33], out[513]);
  buf b_196_(set1[259], out[739]);
  buf b_197_(set1[406], out[886]);
  buf b_198_(set2[101], out[101]);
  buf b_199_(set2[112], out[112]);
  buf b_200_(set2[276], out[276]);
  buf b_201_(set1[362], out[842]);
  buf b_202_(set1[264], out[744]);
  buf b_203_(set1[155], out[635]);
  buf b_204_(set1[427], out[907]);
  buf b_205_(set2[212], out[212]);
  buf b_206_(set1[186], out[666]);
  buf b_207_(set2[369], out[369]);
  buf b_208_(set1[242], out[722]);
  buf b_209_(set1[295], out[775]);
  buf b_210_(set1[262], out[742]);
  buf b_211_(set1[209], out[689]);
  buf b_212_(set1[248], out[728]);
  buf b_213_(set2[37], out[37]);
  buf b_214_(set2[372], out[372]);
  buf b_215_(set1[428], out[908]);
  buf b_216_(set2[289], out[289]);
  buf b_217_(set1[223], out[703]);
  buf b_218_(set2[360], out[360]);
  buf b_219_(set1[64], out[544]);
  buf b_220_(set2[429], out[429]);
  buf b_221_(set1[136], out[616]);
  buf b_222_(set1[373], out[853]);
  buf b_223_(set2[250], out[250]);
  buf b_224_(set2[296], out[296]);
  buf b_225_(set2[422], out[422]);
  buf b_226_(set2[275], out[275]);
  buf b_227_(set1[176], out[656]);
  buf b_228_(set2[393], out[393]);
  buf b_229_(set2[58], out[58]);
  buf b_230_(set2[430], out[430]);
  buf b_231_(set2[359], out[359]);
  buf b_232_(set2[0], out[0]);
  buf b_233_(set1[39], out[519]);
  buf b_234_(set1[289], out[769]);
  buf b_235_(set2[86], out[86]);
  buf b_236_(set1[453], out[933]);
  buf b_237_(set2[439], out[439]);
  buf b_238_(set1[237], out[717]);
  buf b_239_(set2[255], out[255]);
  buf b_240_(set2[418], out[418]);
  buf b_241_(set2[340], out[340]);
  buf b_242_(set1[217], out[697]);
  buf b_243_(set1[153], out[633]);
  buf b_244_(set2[362], out[362]);
  buf b_245_(set2[230], out[230]);
  buf b_246_(set2[199], out[199]);
  buf b_247_(set1[162], out[642]);
  buf b_248_(set1[441], out[921]);
  buf b_249_(set1[111], out[591]);
  buf b_250_(set2[111], out[111]);
  buf b_251_(set1[71], out[551]);
  buf b_252_(set2[329], out[329]);
  buf b_253_(set1[70], out[550]);
  buf b_254_(set2[449], out[449]);
  buf b_255_(set2[104], out[104]);
  buf b_256_(set1[94], out[574]);
  buf b_257_(set1[405], out[885]);
  buf b_258_(set2[335], out[335]);
  buf b_259_(set2[15], out[15]);
  buf b_260_(set1[273], out[753]);
  buf b_261_(set2[197], out[197]);
  buf b_262_(set1[236], out[716]);
  buf b_263_(set1[93], out[573]);
  czero b_264_(_055969_);
  buf b_265_(set2[66], out[66]);
  buf b_266_(set1[211], out[691]);
  buf b_267_(set1[194], out[674]);
  buf b_268_(set1[439], out[919]);
  buf b_269_(set2[193], out[193]);
  buf b_270_(set2[273], out[273]);
  buf b_271_(set2[160], out[160]);
  buf b_272_(set1[174], out[654]);
  buf b_273_(set1[119], out[599]);
  buf b_274_(set2[465], out[465]);
  buf b_275_(set2[399], out[399]);
  buf b_276_(set2[311], out[311]);
  buf b_277_(set1[198], out[678]);
  buf b_278_(set2[417], out[417]);
  buf b_279_(set2[293], out[293]);
  buf b_280_(set1[466], out[946]);
  buf b_281_(set2[371], out[371]);
  buf b_282_(set1[293], out[773]);
  buf b_283_(set2[223], out[223]);
  buf b_284_(set1[42], out[522]);
  buf b_285_(set2[12], out[12]);
  buf b_286_(set2[117], out[117]);
  buf b_287_(set1[471], out[951]);
  buf b_288_(set1[113], out[593]);
  buf b_289_(set2[376], out[376]);
  buf b_290_(set2[299], out[299]);
  buf b_291_(set2[288], out[288]);
  buf b_292_(set1[425], out[905]);
  buf b_293_(set2[38], out[38]);
  buf b_294_(set1[316], out[796]);
  buf b_295_(set2[139], out[139]);
  buf b_296_(set2[59], out[59]);
  buf b_297_(set1[456], out[936]);
  buf b_298_(set1[228], out[708]);
  buf b_299_(set2[247], out[247]);
  buf b_300_(set2[62], out[62]);
  buf b_301_(set1[86], out[566]);
  buf b_302_(set2[386], out[386]);
  buf b_303_(set2[151], out[151]);
  buf b_304_(set1[268], out[748]);
  buf b_305_(set1[323], out[803]);
  buf b_306_(set2[328], out[328]);
  buf b_307_(set2[450], out[450]);
  buf b_308_(set2[354], out[354]);
  buf b_309_(set1[79], out[559]);
  buf b_310_(set1[255], out[735]);
  buf b_311_(set2[77], out[77]);
  buf b_312_(set2[34], out[34]);
  buf b_313_(set2[71], out[71]);
  buf b_314_(set1[78], out[558]);
  buf b_315_(set2[442], out[442]);
  buf b_316_(set1[418], out[898]);
  buf b_317_(set2[195], out[195]);
  buf b_318_(set2[13], out[13]);
  buf b_319_(set1[18], out[498]);
  buf b_320_(set2[451], out[451]);
  buf b_321_(set1[260], out[740]);
  buf b_322_(set1[143], out[623]);
  buf b_323_(set2[327], out[327]);
  buf b_324_(set1[15], out[495]);
  buf b_325_(set2[458], out[458]);
  buf b_326_(set2[234], out[234]);
  buf b_327_(set2[25], out[25]);
  buf b_328_(set1[442], out[922]);
  buf b_329_(set1[313], out[793]);
  buf b_330_(set2[80], out[80]);
  buf b_331_(set1[382], out[862]);
  buf b_332_(set2[344], out[344]);
  buf b_333_(set2[8], out[8]);
  buf b_334_(set1[312], out[792]);
  buf b_335_(set2[468], out[468]);
  buf b_336_(set1[394], out[874]);
  buf b_337_(set2[403], out[403]);
  buf b_338_(set1[120], out[600]);
  buf b_339_(set1[46], out[526]);
  buf b_340_(set2[98], out[98]);
  buf b_341_(set2[100], out[100]);
  buf b_342_(set1[479], out[959]);
  buf b_343_(set2[145], out[145]);
  buf b_344_(set1[363], out[843]);
  buf b_345_(set1[392], out[872]);
  buf b_346_(set1[65], out[545]);
  buf b_347_(set2[253], out[253]);
  buf b_348_(set2[382], out[382]);
  czero b_349_(out[967]);
  czero b_350_(out[975]);
  buf b_351_(set1[372], out[852]);
  buf b_352_(set1[375], out[855]);
  buf b_353_(set2[211], out[211]);
  buf b_354_(set1[52], out[532]);
  buf b_355_(set2[473], out[473]);
  buf b_356_(set2[437], out[437]);
  buf b_357_(set1[169], out[649]);
  buf b_358_(set1[66], out[546]);
  buf b_359_(set1[127], out[607]);
  buf b_360_(set1[170], out[650]);
  buf b_361_(set1[415], out[895]);
  buf b_362_(set2[102], out[102]);
  buf b_363_(set2[264], out[264]);
  buf b_364_(set1[182], out[662]);
  buf b_365_(set2[441], out[441]);
  buf b_366_(set2[314], out[314]);
  buf b_367_(set1[475], out[955]);
  buf b_368_(set1[266], out[746]);
  buf b_369_(set2[198], out[198]);
  buf b_370_(set2[133], out[133]);
  buf b_371_(set1[444], out[924]);
  buf b_372_(set1[19], out[499]);
  buf b_373_(set2[175], out[175]);
  buf b_374_(set1[365], out[845]);
  buf b_375_(set2[236], out[236]);
  buf b_376_(set1[359], out[839]);
  buf b_377_(set1[422], out[902]);
  buf b_378_(set2[303], out[303]);
  buf b_379_(set1[13], out[493]);
  buf b_380_(set2[5], out[5]);
  buf b_381_(set1[81], out[561]);
  buf b_382_(set1[205], out[685]);
  buf b_383_(set1[63], out[543]);
  buf b_384_(set1[297], out[777]);
  buf b_385_(set1[292], out[772]);
  buf b_386_(set1[331], out[811]);
  buf b_387_(set2[268], out[268]);
  buf b_388_(set2[6], out[6]);
  buf b_389_(set2[391], out[391]);
  buf b_390_(set1[100], out[580]);
  buf b_391_(set1[367], out[847]);
  buf b_392_(set1[417], out[897]);
  buf b_393_(set1[214], out[694]);
  buf b_394_(set1[114], out[594]);
  buf b_395_(set2[281], out[281]);
  buf b_396_(set2[1], out[1]);
  buf b_397_(set2[237], out[237]);
  buf b_398_(set1[396], out[876]);
  buf b_399_(set1[254], out[734]);
  buf b_400_(set2[144], out[144]);
  buf b_401_(set1[430], out[910]);
  buf b_402_(set2[466], out[466]);
  buf b_403_(set2[53], out[53]);
  buf b_404_(set2[438], out[438]);
  buf b_405_(set1[280], out[760]);
  buf b_406_(set2[14], out[14]);
  buf b_407_(set1[103], out[583]);
  buf b_408_(set2[78], out[78]);
  buf b_409_(set2[334], out[334]);
  buf b_410_(set1[12], out[492]);
  buf b_411_(set2[396], out[396]);
  buf b_412_(set2[349], out[349]);
  buf b_413_(set1[269], out[749]);
  buf b_414_(set2[476], out[476]);
  buf b_415_(set1[50], out[530]);
  buf b_416_(set2[419], out[419]);
  buf b_417_(set2[149], out[149]);
  buf b_418_(set2[141], out[141]);
  buf b_419_(set2[333], out[333]);
  buf b_420_(set1[34], out[514]);
  buf b_421_(set2[323], out[323]);
  buf b_422_(set1[327], out[807]);
  buf b_423_(set2[225], out[225]);
  buf b_424_(set2[191], out[191]);
  buf b_425_(set2[459], out[459]);
  buf b_426_(set1[244], out[724]);
  buf b_427_(set1[243], out[723]);
  buf b_428_(set1[343], out[823]);
  buf b_429_(set1[384], out[864]);
  buf b_430_(set1[429], out[909]);
  buf b_431_(set2[55], out[55]);
  buf b_432_(set2[291], out[291]);
  buf b_433_(set1[467], out[947]);
  buf b_434_(set2[407], out[407]);
  buf b_435_(set2[127], out[127]);
  buf b_436_(set1[204], out[684]);
  buf b_437_(set2[398], out[398]);
  buf b_438_(set2[79], out[79]);
  buf b_439_(set2[375], out[375]);
  buf b_440_(set1[96], out[576]);
  buf b_441_(set1[326], out[806]);
  buf b_442_(set1[278], out[758]);
  buf b_443_(set2[361], out[361]);
  buf b_444_(set1[462], out[942]);
  buf b_445_(set2[364], out[364]);
  buf b_446_(set2[74], out[74]);
  buf b_447_(set1[435], out[915]);
  buf b_448_(set2[214], out[214]);
  buf b_449_(set2[397], out[397]);
  buf b_450_(set1[352], out[832]);
  buf b_451_(set2[370], out[370]);
  buf b_452_(set1[189], out[669]);
  buf b_453_(set1[212], out[692]);
  buf b_454_(set1[448], out[928]);
  buf b_455_(set2[161], out[161]);
  buf b_456_(set2[406], out[406]);
  buf b_457_(set2[325], out[325]);
  buf b_458_(set1[74], out[554]);
  buf b_459_(set1[110], out[590]);
  buf b_460_(set2[348], out[348]);
  buf b_461_(set2[109], out[109]);
  buf b_462_(set2[124], out[124]);
  buf b_463_(set2[271], out[271]);
  buf b_464_(set1[377], out[857]);
  buf b_465_(set1[412], out[892]);
  buf b_466_(set2[39], out[39]);
  buf b_467_(set2[469], out[469]);
  buf b_468_(set2[90], out[90]);
  buf b_469_(set1[84], out[564]);
  buf b_470_(set2[363], out[363]);
  buf b_471_(set2[248], out[248]);
  buf b_472_(set2[445], out[445]);
  buf b_473_(set2[178], out[178]);
  buf b_474_(set2[241], out[241]);
  buf b_475_(set1[332], out[812]);
  buf b_476_(set2[36], out[36]);
  buf b_477_(set1[168], out[648]);
  buf b_478_(set2[240], out[240]);
  buf b_479_(set1[286], out[766]);
  buf b_480_(set2[453], out[453]);
  buf b_481_(set2[221], out[221]);
  buf b_482_(set2[239], out[239]);
  buf b_483_(set1[88], out[568]);
  buf b_484_(set2[436], out[436]);
  buf b_485_(set2[284], out[284]);
  buf b_486_(set2[324], out[324]);
  buf b_487_(set2[166], out[166]);
  buf b_488_(set1[213], out[693]);
  buf b_489_(set2[411], out[411]);
  buf b_490_(set2[188], out[188]);
  buf b_491_(set1[461], out[941]);
  buf b_492_(set2[143], out[143]);
  buf b_493_(set1[219], out[699]);
  buf b_494_(set2[300], out[300]);
  buf b_495_(set1[291], out[771]);
  buf b_496_(set2[404], out[404]);
  buf b_497_(set1[437], out[917]);
  buf b_498_(set1[224], out[704]);
  buf b_499_(set1[215], out[695]);
  buf b_500_(set1[309], out[789]);
  buf b_501_(set2[365], out[365]);
  buf b_502_(set2[279], out[279]);
  buf b_503_(set2[431], out[431]);
  buf b_504_(set1[172], out[652]);
  buf b_505_(set1[129], out[609]);
  buf b_506_(set1[173], out[653]);
  buf b_507_(set2[443], out[443]);
  buf b_508_(set1[395], out[875]);
  buf b_509_(set2[389], out[389]);
  buf b_510_(set1[196], out[676]);
  buf b_511_(set2[10], out[10]);
  buf b_512_(set2[17], out[17]);
  buf b_513_(set2[270], out[270]);
  buf b_514_(set1[218], out[698]);
  buf b_515_(set2[343], out[343]);
  buf b_516_(set2[83], out[83]);
  buf b_517_(set2[29], out[29]);
  buf b_518_(set1[210], out[690]);
  buf b_519_(set1[386], out[866]);
  buf b_520_(set1[337], out[817]);
  buf b_521_(set1[2], out[482]);
  buf b_522_(set2[60], out[60]);
  buf b_523_(set2[168], out[168]);
  buf b_524_(set2[152], out[152]);
  buf b_525_(set1[62], out[542]);
  czero b_526_(out[969]);
  buf b_527_(set2[310], out[310]);
  buf b_528_(set2[89], out[89]);
  buf b_529_(set2[475], out[475]);
  buf b_530_(set1[391], out[871]);
  buf b_531_(set2[50], out[50]);
  buf b_532_(set2[312], out[312]);
  buf b_533_(set1[183], out[663]);
  buf b_534_(set1[328], out[808]);
  buf b_535_(set2[27], out[27]);
  buf b_536_(set1[383], out[863]);
  buf b_537_(set2[400], out[400]);
  buf b_538_(set1[306], out[786]);
  buf b_539_(set2[73], out[73]);
  buf b_540_(set1[285], out[765]);
  buf b_541_(set2[30], out[30]);
  buf b_542_(set1[30], out[510]);
  buf b_543_(set1[271], out[751]);
  buf b_544_(set2[219], out[219]);
  buf b_545_(set2[203], out[203]);
  buf b_546_(set1[344], out[824]);
  buf b_547_(set2[242], out[242]);
  buf b_548_(set2[320], out[320]);
  buf b_549_(set2[409], out[409]);
  buf b_550_(set2[415], out[415]);
  buf b_551_(set2[434], out[434]);
  buf b_552_(set1[303], out[783]);
  buf b_553_(set1[3], out[483]);
  buf b_554_(set1[131], out[611]);
  buf b_555_(set1[357], out[837]);
  buf b_556_(set1[272], out[752]);
  buf b_557_(set2[356], out[356]);
  buf b_558_(set1[1], out[481]);
  buf b_559_(set2[301], out[301]);
  buf b_560_(set1[125], out[605]);
  buf b_561_(set2[330], out[330]);
  buf b_562_(set2[63], out[63]);
  buf b_563_(set1[226], out[706]);
  buf b_564_(set1[460], out[940]);
  buf b_565_(set1[177], out[657]);
  buf b_566_(set2[97], out[97]);
  buf b_567_(set2[266], out[266]);
  buf b_568_(set2[163], out[163]);
  buf b_569_(set1[443], out[923]);
  buf b_570_(set1[360], out[840]);
  buf b_571_(set1[241], out[721]);
  buf b_572_(set1[424], out[904]);
  buf b_573_(set2[402], out[402]);
  buf b_574_(set1[302], out[782]);
  buf b_575_(set1[347], out[827]);
  buf b_576_(set1[376], out[856]);
  buf b_577_(set2[91], out[91]);
  buf b_578_(set2[394], out[394]);
  buf b_579_(set2[28], out[28]);
  buf b_580_(set2[164], out[164]);
  buf b_581_(set1[330], out[810]);
  buf b_582_(set2[269], out[269]);
  buf b_583_(set1[106], out[586]);
  buf b_584_(set1[288], out[768]);
  buf b_585_(set2[295], out[295]);
  buf b_586_(set2[57], out[57]);
  buf b_587_(set1[221], out[701]);
  buf b_588_(set1[25], out[505]);
  buf b_589_(set1[9], out[489]);
  buf b_590_(set1[68], out[548]);
  buf b_591_(set2[454], out[454]);
  buf b_592_(set1[22], out[502]);
  czero b_593_(out[964]);
  buf b_594_(set2[246], out[246]);
  buf b_595_(set1[311], out[791]);
  buf b_596_(set1[150], out[630]);
  buf b_597_(set1[137], out[617]);
  buf b_598_(set1[231], out[711]);
  buf b_599_(set2[277], out[277]);
  buf b_600_(set2[190], out[190]);
  buf b_601_(set2[232], out[232]);
  buf b_602_(set1[190], out[670]);
  buf b_603_(set2[332], out[332]);
  buf b_604_(set2[463], out[463]);
  buf b_605_(set1[451], out[931]);
  buf b_606_(set1[411], out[891]);
  czero b_607_(out[968]);
  buf b_608_(set2[43], out[43]);
  buf b_609_(set1[163], out[643]);
  buf b_610_(set2[416], out[416]);
  buf b_611_(set1[477], out[957]);
  buf b_612_(set2[435], out[435]);
  buf b_613_(set1[449], out[929]);
  buf b_614_(set1[200], out[680]);
  buf b_615_(set1[385], out[865]);
  buf b_616_(set1[207], out[687]);
  buf b_617_(set1[239], out[719]);
  buf b_618_(set1[322], out[802]);
  buf b_619_(set1[123], out[603]);
  buf b_620_(set1[354], out[834]);
  buf b_621_(set1[105], out[585]);
  buf b_622_(set1[104], out[584]);
  buf b_623_(set2[448], out[448]);
  buf b_624_(set2[21], out[21]);
  czero b_625_(out[965]);
  buf b_626_(set2[337], out[337]);
  buf b_627_(set1[325], out[805]);
  buf b_628_(set1[356], out[836]);
  buf b_629_(set2[346], out[346]);
  buf b_630_(set2[304], out[304]);
  buf b_631_(set1[350], out[830]);
  buf b_632_(set2[202], out[202]);
  buf b_633_(set1[342], out[822]);
  buf b_634_(set1[307], out[787]);
  buf b_635_(set2[114], out[114]);
  buf b_636_(set2[207], out[207]);
  buf b_637_(set1[324], out[804]);
  buf b_638_(set2[373], out[373]);
  buf b_639_(set2[128], out[128]);
  buf b_640_(set1[192], out[672]);
  buf b_641_(set1[222], out[702]);
  buf b_642_(set2[261], out[261]);
  buf b_643_(set2[70], out[70]);
  buf b_644_(set1[145], out[625]);
  czero b_645_(out[973]);
  buf b_646_(set1[233], out[713]);
  buf b_647_(set2[205], out[205]);
  buf b_648_(set2[213], out[213]);
  buf b_649_(set2[131], out[131]);
  buf b_650_(set2[33], out[33]);
  buf b_651_(set2[278], out[278]);
  buf b_652_(set1[21], out[501]);
  buf b_653_(set2[220], out[220]);
  buf b_654_(set1[159], out[639]);
  buf b_655_(set1[0], out[480]);
  buf b_656_(set1[247], out[727]);
  buf b_657_(set2[126], out[126]);
  buf b_658_(set1[401], out[881]);
  buf b_659_(set1[77], out[557]);
  buf b_660_(set1[413], out[893]);
  buf b_661_(set2[377], out[377]);
  buf b_662_(set1[349], out[829]);
  buf b_663_(set2[405], out[405]);
  buf b_664_(set2[472], out[472]);
  buf b_665_(set1[420], out[900]);
  buf b_666_(set1[85], out[565]);
  buf b_667_(set1[216], out[696]);
  buf b_668_(set2[460], out[460]);
  buf b_669_(set1[321], out[801]);
  czero b_670_(_055968_);
  buf b_671_(set1[351], out[831]);
  buf b_672_(set2[456], out[456]);
  buf b_673_(set1[29], out[509]);
  buf b_674_(set1[76], out[556]);
  buf b_675_(set2[243], out[243]);
  buf b_676_(set1[57], out[537]);
  buf b_677_(set1[139], out[619]);
  buf b_678_(set1[229], out[709]);
  buf b_679_(set1[474], out[954]);
  buf b_680_(set2[245], out[245]);
  buf b_681_(set1[478], out[958]);
  buf b_682_(set2[321], out[321]);
  buf b_683_(set1[225], out[705]);
  buf b_684_(set1[345], out[825]);
  buf b_685_(set1[140], out[620]);
  buf b_686_(set2[99], out[99]);
  buf b_687_(set2[428], out[428]);
  buf b_688_(set1[423], out[903]);
  buf b_689_(set1[48], out[528]);
  buf b_690_(set1[44], out[524]);
  buf b_691_(set2[47], out[47]);
  buf b_692_(set2[169], out[169]);
  buf b_693_(set2[358], out[358]);
  buf b_694_(set1[407], out[887]);
  buf b_695_(set1[314], out[794]);
  buf b_696_(set2[148], out[148]);
  buf b_697_(set1[37], out[517]);
  buf b_698_(set1[41], out[521]);
  buf b_699_(set1[166], out[646]);
  buf b_700_(set1[431], out[911]);
  buf b_701_(set1[472], out[952]);
  buf b_702_(set1[240], out[720]);
  buf b_703_(set2[384], out[384]);
  buf b_704_(set2[345], out[345]);
  buf b_705_(set2[267], out[267]);
  buf b_706_(set2[22], out[22]);
  czero b_707_(out[975]);
  buf b_708_(set2[7], out[7]);
  buf b_709_(set2[305], out[305]);
  buf b_710_(set2[426], out[426]);
  buf b_711_(set2[123], out[123]);
  buf b_712_(set2[282], out[282]);
  buf b_713_(set2[11], out[11]);
  buf b_714_(set1[402], out[882]);
  buf b_715_(set2[257], out[257]);
  buf b_716_(set1[366], out[846]);
  buf b_717_(set2[336], out[336]);
  buf b_718_(set1[440], out[920]);
  buf b_719_(set2[331], out[331]);
  buf b_720_(set2[347], out[347]);
  buf b_721_(set1[115], out[595]);
  buf b_722_(set2[392], out[392]);
  buf b_723_(set1[80], out[560]);
  buf b_724_(set2[233], out[233]);
  buf b_725_(set1[191], out[671]);
  buf b_726_(set2[378], out[378]);
  buf b_727_(set1[160], out[640]);
  buf b_728_(set2[147], out[147]);
  buf b_729_(set2[462], out[462]);
  buf b_730_(set1[258], out[738]);
  buf b_731_(set2[315], out[315]);
  buf b_732_(set2[49], out[49]);
  buf b_733_(set1[378], out[858]);
  buf b_734_(set1[305], out[785]);
  buf b_735_(set2[222], out[222]);
  buf b_736_(set2[227], out[227]);
  buf b_737_(set1[371], out[851]);
  buf b_738_(set2[322], out[322]);
  buf b_739_(set2[184], out[184]);
  buf b_740_(set1[380], out[860]);
  buf b_741_(set2[134], out[134]);
  buf b_742_(set2[217], out[217]);
  buf b_743_(set2[226], out[226]);
  buf b_744_(set1[421], out[901]);
  buf b_745_(set2[64], out[64]);
  buf b_746_(set2[381], out[381]);
  buf b_747_(set1[28], out[508]);
  buf b_748_(set2[286], out[286]);
  buf b_749_(set1[261], out[741]);
  buf b_750_(set2[103], out[103]);
  buf b_751_(set1[83], out[563]);
  buf b_752_(set1[20], out[500]);
  buf b_753_(set1[468], out[948]);
  buf b_754_(set2[387], out[387]);
  buf b_755_(set2[206], out[206]);
  buf b_756_(set2[187], out[187]);
  buf b_757_(set1[235], out[715]);
  buf b_758_(set2[464], out[464]);
  buf b_759_(set1[201], out[681]);
  czero b_760_(out[972]);
  buf b_761_(set1[142], out[622]);
  buf b_762_(set2[172], out[172]);
  buf b_763_(set1[185], out[665]);
  buf b_764_(set1[55], out[535]);
  buf b_765_(set2[200], out[200]);
  buf b_766_(set1[296], out[776]);
  buf b_767_(set2[87], out[87]);
  buf b_768_(set2[427], out[427]);
  buf b_769_(set2[455], out[455]);
  buf b_770_(set2[16], out[16]);
  buf b_771_(set2[262], out[262]);
  buf b_772_(set1[128], out[608]);
  buf b_773_(set1[157], out[637]);
  buf b_774_(set1[43], out[523]);
  buf b_775_(set1[16], out[496]);
  buf b_776_(set2[167], out[167]);
  buf b_777_(set2[447], out[447]);
  buf b_778_(set2[457], out[457]);
  buf b_779_(set2[231], out[231]);
  buf b_780_(set1[338], out[818]);
  buf b_781_(set2[2], out[2]);
  buf b_782_(set1[358], out[838]);
  buf b_783_(set1[171], out[651]);
  buf b_784_(set2[355], out[355]);
  buf b_785_(set2[265], out[265]);
  buf b_786_(set2[368], out[368]);
  buf b_787_(set1[263], out[743]);
  buf b_788_(set2[444], out[444]);
  buf b_789_(set1[36], out[516]);
  buf b_790_(set2[420], out[420]);
  buf b_791_(set2[252], out[252]);
  buf b_792_(set1[414], out[894]);
  buf b_793_(set2[158], out[158]);
  buf b_794_(set2[48], out[48]);
  buf b_795_(set1[353], out[833]);
  buf b_796_(set1[138], out[618]);
  buf b_797_(set1[199], out[679]);
  buf b_798_(set2[189], out[189]);
  buf b_799_(set2[106], out[106]);
  buf b_800_(set2[150], out[150]);
  buf b_801_(set1[284], out[764]);
  buf b_802_(set1[408], out[888]);
  buf b_803_(set2[56], out[56]);
  buf b_804_(set1[87], out[567]);
  buf b_805_(set1[230], out[710]);
  buf b_806_(set1[282], out[762]);
  buf b_807_(set1[436], out[916]);
  buf b_808_(set1[368], out[848]);
  buf b_809_(set1[387], out[867]);
  buf b_810_(set2[306], out[306]);
  buf b_811_(set1[238], out[718]);
  buf b_812_(set1[304], out[784]);
  buf b_813_(set2[19], out[19]);
  buf b_814_(set1[126], out[606]);
  buf b_815_(set2[137], out[137]);
  buf b_816_(set1[452], out[932]);
  buf b_817_(set1[27], out[507]);
  buf b_818_(set2[54], out[54]);
  buf b_819_(set2[302], out[302]);
  buf b_820_(set1[257], out[737]);
  buf b_821_(set1[11], out[491]);
  buf b_822_(set2[76], out[76]);
  buf b_823_(set2[88], out[88]);
  buf b_824_(set2[388], out[388]);
  buf b_825_(set2[395], out[395]);
  buf b_826_(set1[279], out[759]);
  buf b_827_(set1[38], out[518]);
  buf b_828_(set1[72], out[552]);
  buf b_829_(set2[467], out[467]);
  buf b_830_(set1[275], out[755]);
  buf b_831_(set2[138], out[138]);
  buf b_832_(set2[4], out[4]);
  buf b_833_(set1[438], out[918]);
  buf b_834_(set2[338], out[338]);
  buf b_835_(set2[385], out[385]);
  buf b_836_(set2[119], out[119]);
  buf b_837_(set2[113], out[113]);
  buf b_838_(set2[68], out[68]);
  buf b_839_(set2[339], out[339]);
  buf b_840_(set1[141], out[621]);
  buf b_841_(set1[202], out[682]);
  buf b_842_(set2[342], out[342]);
  buf b_843_(set2[176], out[176]);
  buf b_844_(set1[234], out[714]);
  buf b_845_(set2[3], out[3]);
  buf b_846_(set1[82], out[562]);
  buf b_847_(set2[313], out[313]);
  buf b_848_(set2[45], out[45]);
  buf b_849_(set1[274], out[754]);
  buf b_850_(set1[54], out[534]);
  buf b_851_(set1[397], out[877]);
  buf b_852_(set1[459], out[939]);
  buf b_853_(set2[461], out[461]);
  buf b_854_(set2[142], out[142]);
  buf b_855_(set1[355], out[835]);
  buf b_856_(set1[464], out[944]);
  buf b_857_(set2[440], out[440]);
  buf b_858_(set2[67], out[67]);
  buf b_859_(set2[374], out[374]);
  buf b_860_(set1[364], out[844]);
  buf b_861_(set2[307], out[307]);
  buf b_862_(set2[401], out[401]);
  buf b_863_(set2[81], out[81]);
  buf b_864_(set1[118], out[598]);
  buf b_865_(set1[298], out[778]);
  buf b_866_(set2[308], out[308]);
  buf b_867_(set1[31], out[511]);
  buf b_868_(set1[193], out[673]);
  buf b_869_(set1[208], out[688]);
  buf b_870_(set1[463], out[943]);
  buf b_871_(set1[476], out[956]);
  buf b_872_(set1[158], out[638]);
  buf b_873_(set1[91], out[571]);
  buf b_874_(set1[101], out[581]);
  buf b_875_(set1[112], out[592]);
  buf b_876_(set1[310], out[790]);
  buf b_877_(set1[318], out[798]);
  buf b_878_(set1[433], out[913]);
  buf b_879_(set2[297], out[297]);
  buf b_880_(set2[201], out[201]);
  buf b_881_(set2[408], out[408]);
  buf b_882_(set2[153], out[153]);
  buf b_883_(set1[335], out[815]);
  buf b_884_(set2[478], out[478]);
  buf b_885_(set2[32], out[32]);
  buf b_886_(set2[383], out[383]);
  buf b_887_(set1[245], out[725]);
  buf b_888_(set1[117], out[597]);
  buf b_889_(set1[95], out[575]);
  buf b_890_(set1[203], out[683]);
  buf b_891_(set2[24], out[24]);
  buf b_892_(set1[206], out[686]);
  buf b_893_(set1[109], out[589]);
  buf b_894_(set2[171], out[171]);
  buf b_895_(set2[317], out[317]);
  buf b_896_(set1[152], out[632]);
  buf b_897_(set1[276], out[756]);
  buf b_898_(set2[122], out[122]);
  buf b_899_(set1[370], out[850]);
  buf b_900_(set1[108], out[588]);
  buf b_901_(set2[157], out[157]);
  buf b_902_(set2[52], out[52]);
  buf b_903_(set1[329], out[809]);
  buf b_904_(set1[24], out[504]);
  buf b_905_(set2[92], out[92]);
  buf b_906_(set2[116], out[116]);
  buf b_907_(set2[316], out[316]);
  buf b_908_(set1[107], out[587]);
  buf b_909_(set1[26], out[506]);
  buf b_910_(set1[445], out[925]);
  buf b_911_(set1[389], out[869]);
  buf b_912_(set1[156], out[636]);
  buf b_913_(set1[161], out[641]);
  buf b_914_(set1[333], out[813]);
  buf b_915_(set1[8], out[488]);
  buf b_916_(set1[252], out[732]);
  buf b_917_(set1[399], out[879]);
  buf b_918_(set1[250], out[730]);
  buf b_919_(set1[287], out[767]);
  buf b_920_(set2[95], out[95]);
  buf b_921_(set2[179], out[179]);
  buf b_922_(set1[381], out[861]);
  buf b_923_(set2[110], out[110]);
  buf b_924_(set1[4], out[484]);
  buf b_925_(set2[23], out[23]);
  buf b_926_(set2[135], out[135]);
  buf b_927_(set1[40], out[520]);
  buf b_928_(set2[65], out[65]);
  buf b_929_(set1[14], out[494]);
  buf b_930_(set2[259], out[259]);
  buf b_931_(set1[90], out[570]);
  buf b_932_(set1[89], out[569]);
  buf b_933_(set1[102], out[582]);
  buf b_934_(set1[47], out[527]);
  buf b_935_(set2[263], out[263]);
  buf b_936_(set1[400], out[880]);
  buf b_937_(set1[300], out[780]);
  buf b_938_(set1[10], out[490]);
  buf b_939_(set2[155], out[155]);
  buf b_940_(set2[477], out[477]);
  buf b_941_(set2[146], out[146]);
  buf b_942_(set2[423], out[423]);
  buf b_943_(set2[75], out[75]);
  buf b_944_(set1[301], out[781]);
  buf b_945_(set1[246], out[726]);
  buf b_946_(set2[42], out[42]);
  buf b_947_(set1[403], out[883]);
  czero b_948_(out[971]);
  buf b_949_(set1[294], out[774]);
  buf b_950_(set2[121], out[121]);
  buf b_951_(set1[45], out[525]);
  buf b_952_(set1[232], out[712]);
  buf b_953_(set2[61], out[61]);
  buf b_954_(set2[366], out[366]);
  buf b_955_(set1[56], out[536]);
  buf b_956_(set1[35], out[515]);
  buf b_957_(set2[292], out[292]);
  buf b_958_(set2[254], out[254]);
  buf b_959_(set1[339], out[819]);
  buf b_960_(set2[156], out[156]);
  buf b_961_(set2[181], out[181]);
  buf b_962_(set2[177], out[177]);
  buf b_963_(set1[455], out[935]);
  buf b_964_(set1[454], out[934]);
  buf b_965_(set1[393], out[873]);
  buf b_966_(set2[194], out[194]);
  buf b_967_(set2[120], out[120]);
  buf b_968_(set2[433], out[433]);
  buf b_969_(set1[416], out[896]);
  buf b_970_(set2[140], out[140]);
  buf b_971_(set1[469], out[949]);
  buf b_972_(set1[17], out[497]);
  buf b_973_(set1[410], out[890]);
  buf b_974_(set1[121], out[601]);
  buf b_975_(set1[346], out[826]);
  buf b_976_(set2[108], out[108]);
  buf b_977_(set2[379], out[379]);
  buf b_978_(set2[256], out[256]);
  buf b_979_(set1[146], out[626]);
  czero b_980_(out[966]);
  buf b_981_(set1[144], out[624]);
  buf b_982_(set2[185], out[185]);
  buf b_983_(set2[182], out[182]);
  buf b_984_(set1[446], out[926]);
  buf b_985_(set1[73], out[553]);
  buf b_986_(set1[281], out[761]);

endmodule
