module min_hash(
  input wire [479:0] set1,
  input wire [479:0] set2,
  output wire [975:0] out
);
  // lint_off MULTIPLY
  function automatic [21:0] umul22b_16b_x_6b (input reg [15:0] lhs, input reg [5:0] rhs);
    begin
      umul22b_16b_x_6b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [22:0] umul23b_16b_x_7b (input reg [15:0] lhs, input reg [6:0] rhs);
    begin
      umul23b_16b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [15:0] set1_unflattened[30];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  wire [15:0] set2_unflattened[30];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  wire [15:0] array_index_52333;
  wire [15:0] array_index_52335;
  wire [21:0] umul_52337;
  wire [21:0] umul_52338;
  wire [21:0] umul_52347;
  wire [21:0] umul_52348;
  wire [15:0] array_index_52349;
  wire [15:0] array_index_52353;
  wire [21:0] umul_52361;
  wire [15:0] add_52363;
  wire [21:0] umul_52365;
  wire [15:0] add_52367;
  wire [21:0] umul_52387;
  wire [21:0] umul_52388;
  wire [21:0] umul_52389;
  wire [21:0] add_52391;
  wire [21:0] umul_52393;
  wire [21:0] add_52395;
  wire [15:0] array_index_52397;
  wire [31:0] smod_52401;
  wire [15:0] array_index_52402;
  wire [31:0] smod_52406;
  wire [21:0] umul_52419;
  wire [15:0] add_52421;
  wire [21:0] umul_52425;
  wire [15:0] add_52427;
  wire [31:0] smod_52442;
  wire [31:0] smod_52446;
  wire [22:0] umul_52461;
  wire [22:0] umul_52462;
  wire [21:0] umul_52463;
  wire [20:0] add_52465;
  wire [21:0] umul_52467;
  wire [20:0] add_52469;
  wire [21:0] umul_52471;
  wire [21:0] add_52473;
  wire [21:0] umul_52477;
  wire [21:0] add_52479;
  wire [15:0] array_index_52483;
  wire [31:0] smod_52487;
  wire [15:0] array_index_52490;
  wire [31:0] smod_52494;
  wire [21:0] umul_52521;
  wire [15:0] add_52523;
  wire [15:0] sel_52528;
  wire [21:0] umul_52529;
  wire [15:0] add_52531;
  wire [15:0] sel_52536;
  wire [31:0] smod_52548;
  wire [31:0] smod_52552;
  wire [31:0] smod_52556;
  wire [31:0] smod_52562;
  wire [22:0] umul_52579;
  wire [22:0] umul_52580;
  wire [22:0] umul_52581;
  wire [22:0] add_52583;
  wire [22:0] umul_52585;
  wire [22:0] add_52587;
  wire [21:0] umul_52589;
  wire [20:0] add_52591;
  wire [21:0] umul_52595;
  wire [20:0] add_52597;
  wire [21:0] umul_52601;
  wire [21:0] add_52603;
  wire [15:0] sel_52608;
  wire [21:0] umul_52609;
  wire [21:0] add_52611;
  wire [15:0] sel_52616;
  wire [15:0] array_index_52617;
  wire [31:0] smod_52621;
  wire [15:0] array_index_52623;
  wire [31:0] smod_52627;
  wire [21:0] umul_52665;
  wire [15:0] add_52667;
  wire [15:0] sel_52672;
  wire [21:0] umul_52673;
  wire [15:0] add_52675;
  wire [15:0] sel_52680;
  wire [31:0] smod_52690;
  wire [31:0] smod_52694;
  wire [31:0] smod_52698;
  wire [31:0] smod_52704;
  wire [31:0] smod_52710;
  wire [31:0] smod_52715;
  wire [22:0] umul_52731;
  wire [20:0] add_52733;
  wire [22:0] umul_52735;
  wire [20:0] add_52737;
  wire [22:0] umul_52739;
  wire [22:0] add_52741;
  wire [22:0] umul_52745;
  wire [22:0] add_52747;
  wire [21:0] umul_52751;
  wire [20:0] add_52753;
  wire [15:0] sel_52758;
  wire [21:0] umul_52759;
  wire [20:0] add_52761;
  wire [15:0] sel_52766;
  wire [21:0] umul_52767;
  wire [21:0] add_52769;
  wire [15:0] sel_52774;
  wire [21:0] umul_52775;
  wire [21:0] add_52777;
  wire [15:0] sel_52782;
  wire [15:0] array_index_52783;
  wire [31:0] smod_52787;
  wire [15:0] array_index_52789;
  wire [31:0] smod_52793;
  wire [21:0] umul_52839;
  wire [15:0] add_52841;
  wire [15:0] sel_52846;
  wire [21:0] umul_52847;
  wire [15:0] add_52849;
  wire [15:0] sel_52854;
  wire [31:0] smod_52858;
  wire [31:0] smod_52862;
  wire [31:0] smod_52866;
  wire [31:0] smod_52872;
  wire [31:0] smod_52878;
  wire [31:0] smod_52883;
  wire [31:0] smod_52888;
  wire [31:0] smod_52893;
  wire [22:0] umul_52909;
  wire [20:0] add_52911;
  wire [22:0] umul_52915;
  wire [20:0] add_52917;
  wire [22:0] umul_52921;
  wire [22:0] add_52923;
  wire [15:0] sel_52928;
  wire [22:0] umul_52929;
  wire [22:0] add_52931;
  wire [15:0] sel_52936;
  wire [21:0] umul_52937;
  wire [20:0] add_52939;
  wire [15:0] sel_52944;
  wire [21:0] umul_52945;
  wire [20:0] add_52947;
  wire [15:0] sel_52952;
  wire [21:0] umul_52953;
  wire [21:0] add_52955;
  wire [15:0] sel_52960;
  wire [21:0] umul_52961;
  wire [21:0] add_52963;
  wire [15:0] sel_52968;
  wire [15:0] array_index_52969;
  wire [31:0] smod_52973;
  wire [15:0] array_index_52975;
  wire [31:0] smod_52979;
  wire [21:0] umul_53029;
  wire [15:0] add_53031;
  wire [15:0] sel_53036;
  wire [21:0] umul_53037;
  wire [15:0] add_53039;
  wire [15:0] sel_53044;
  wire [31:0] smod_53048;
  wire [31:0] smod_53054;
  wire [31:0] smod_53060;
  wire [31:0] smod_53065;
  wire [31:0] smod_53070;
  wire [31:0] smod_53075;
  wire [31:0] smod_53080;
  wire [31:0] smod_53085;
  wire [22:0] umul_53101;
  wire [20:0] add_53103;
  wire [15:0] sel_53108;
  wire [22:0] umul_53109;
  wire [20:0] add_53111;
  wire [15:0] sel_53116;
  wire [22:0] umul_53117;
  wire [22:0] add_53119;
  wire [15:0] sel_53124;
  wire [22:0] umul_53125;
  wire [22:0] add_53127;
  wire [15:0] sel_53132;
  wire [21:0] umul_53133;
  wire [20:0] add_53135;
  wire [15:0] sel_53140;
  wire [21:0] umul_53141;
  wire [20:0] add_53143;
  wire [15:0] sel_53148;
  wire [21:0] umul_53149;
  wire [21:0] add_53151;
  wire [15:0] sel_53156;
  wire [21:0] umul_53157;
  wire [21:0] add_53159;
  wire [15:0] sel_53164;
  wire [15:0] array_index_53165;
  wire [31:0] smod_53169;
  wire [15:0] array_index_53171;
  wire [31:0] smod_53175;
  wire [21:0] umul_53225;
  wire [15:0] add_53227;
  wire [15:0] sel_53232;
  wire [21:0] umul_53233;
  wire [15:0] add_53235;
  wire [15:0] sel_53240;
  wire [31:0] smod_53244;
  wire [31:0] smod_53249;
  wire [31:0] smod_53254;
  wire [31:0] smod_53259;
  wire [31:0] smod_53264;
  wire [31:0] smod_53269;
  wire [31:0] smod_53274;
  wire [31:0] smod_53279;
  wire [22:0] umul_53295;
  wire [20:0] add_53297;
  wire [15:0] sel_53302;
  wire [22:0] umul_53303;
  wire [20:0] add_53305;
  wire [15:0] sel_53310;
  wire [22:0] umul_53311;
  wire [22:0] add_53313;
  wire [15:0] sel_53318;
  wire [22:0] umul_53319;
  wire [22:0] add_53321;
  wire [15:0] sel_53326;
  wire [21:0] umul_53327;
  wire [20:0] add_53329;
  wire [15:0] sel_53334;
  wire [21:0] umul_53335;
  wire [20:0] add_53337;
  wire [15:0] sel_53342;
  wire [21:0] umul_53343;
  wire [21:0] add_53345;
  wire [15:0] sel_53350;
  wire [21:0] umul_53351;
  wire [21:0] add_53353;
  wire [15:0] sel_53358;
  wire [15:0] array_index_53359;
  wire [31:0] smod_53363;
  wire [15:0] array_index_53365;
  wire [31:0] smod_53369;
  wire [21:0] umul_53419;
  wire [15:0] add_53421;
  wire [15:0] sel_53426;
  wire [21:0] umul_53427;
  wire [15:0] add_53429;
  wire [15:0] sel_53434;
  wire [31:0] smod_53438;
  wire [31:0] smod_53443;
  wire [31:0] smod_53448;
  wire [31:0] smod_53453;
  wire [31:0] smod_53458;
  wire [31:0] smod_53463;
  wire [31:0] smod_53468;
  wire [31:0] smod_53473;
  wire [22:0] umul_53489;
  wire [20:0] add_53491;
  wire [15:0] sel_53496;
  wire [22:0] umul_53497;
  wire [20:0] add_53499;
  wire [15:0] sel_53504;
  wire [22:0] umul_53505;
  wire [22:0] add_53507;
  wire [15:0] sel_53512;
  wire [22:0] umul_53513;
  wire [22:0] add_53515;
  wire [15:0] sel_53520;
  wire [21:0] umul_53521;
  wire [20:0] add_53523;
  wire [15:0] sel_53528;
  wire [21:0] umul_53529;
  wire [20:0] add_53531;
  wire [15:0] sel_53536;
  wire [21:0] umul_53537;
  wire [21:0] add_53539;
  wire [15:0] sel_53544;
  wire [21:0] umul_53545;
  wire [21:0] add_53547;
  wire [15:0] sel_53552;
  wire [15:0] array_index_53553;
  wire [31:0] smod_53557;
  wire [15:0] array_index_53559;
  wire [31:0] smod_53563;
  wire [21:0] umul_53613;
  wire [15:0] add_53615;
  wire [15:0] sel_53620;
  wire [21:0] umul_53621;
  wire [15:0] add_53623;
  wire [15:0] sel_53628;
  wire [31:0] smod_53632;
  wire [31:0] smod_53637;
  wire [31:0] smod_53642;
  wire [31:0] smod_53647;
  wire [31:0] smod_53652;
  wire [31:0] smod_53657;
  wire [31:0] smod_53662;
  wire [31:0] smod_53667;
  wire [22:0] umul_53683;
  wire [20:0] add_53685;
  wire [15:0] sel_53690;
  wire [22:0] umul_53691;
  wire [20:0] add_53693;
  wire [15:0] sel_53698;
  wire [22:0] umul_53699;
  wire [22:0] add_53701;
  wire [15:0] sel_53706;
  wire [22:0] umul_53707;
  wire [22:0] add_53709;
  wire [15:0] sel_53714;
  wire [21:0] umul_53715;
  wire [20:0] add_53717;
  wire [15:0] sel_53722;
  wire [21:0] umul_53723;
  wire [20:0] add_53725;
  wire [15:0] sel_53730;
  wire [21:0] umul_53731;
  wire [21:0] add_53733;
  wire [15:0] sel_53738;
  wire [21:0] umul_53739;
  wire [21:0] add_53741;
  wire [15:0] sel_53746;
  wire [15:0] array_index_53747;
  wire [31:0] smod_53751;
  wire [15:0] array_index_53753;
  wire [31:0] smod_53757;
  wire [21:0] umul_53807;
  wire [15:0] add_53809;
  wire [15:0] sel_53814;
  wire [21:0] umul_53815;
  wire [15:0] add_53817;
  wire [15:0] sel_53822;
  wire [31:0] smod_53826;
  wire [31:0] smod_53831;
  wire [31:0] smod_53836;
  wire [31:0] smod_53841;
  wire [31:0] smod_53846;
  wire [31:0] smod_53851;
  wire [31:0] smod_53856;
  wire [31:0] smod_53861;
  wire [22:0] umul_53877;
  wire [20:0] add_53879;
  wire [15:0] sel_53884;
  wire [22:0] umul_53885;
  wire [20:0] add_53887;
  wire [15:0] sel_53892;
  wire [22:0] umul_53893;
  wire [22:0] add_53895;
  wire [15:0] sel_53900;
  wire [22:0] umul_53901;
  wire [22:0] add_53903;
  wire [15:0] sel_53908;
  wire [21:0] umul_53909;
  wire [20:0] add_53911;
  wire [15:0] sel_53916;
  wire [21:0] umul_53917;
  wire [20:0] add_53919;
  wire [15:0] sel_53924;
  wire [21:0] umul_53925;
  wire [21:0] add_53927;
  wire [15:0] sel_53932;
  wire [21:0] umul_53933;
  wire [21:0] add_53935;
  wire [15:0] sel_53940;
  wire [15:0] array_index_53941;
  wire [31:0] smod_53945;
  wire [15:0] array_index_53947;
  wire [31:0] smod_53951;
  wire [21:0] umul_54001;
  wire [15:0] add_54003;
  wire [15:0] sel_54008;
  wire [21:0] umul_54009;
  wire [15:0] add_54011;
  wire [15:0] sel_54016;
  wire [31:0] smod_54020;
  wire [31:0] smod_54025;
  wire [31:0] smod_54030;
  wire [31:0] smod_54035;
  wire [31:0] smod_54040;
  wire [31:0] smod_54045;
  wire [31:0] smod_54050;
  wire [31:0] smod_54055;
  wire [22:0] umul_54071;
  wire [20:0] add_54073;
  wire [15:0] sel_54078;
  wire [22:0] umul_54079;
  wire [20:0] add_54081;
  wire [15:0] sel_54086;
  wire [22:0] umul_54087;
  wire [22:0] add_54089;
  wire [15:0] sel_54094;
  wire [22:0] umul_54095;
  wire [22:0] add_54097;
  wire [15:0] sel_54102;
  wire [21:0] umul_54103;
  wire [20:0] add_54105;
  wire [15:0] sel_54110;
  wire [21:0] umul_54111;
  wire [20:0] add_54113;
  wire [15:0] sel_54118;
  wire [21:0] umul_54119;
  wire [21:0] add_54121;
  wire [15:0] sel_54126;
  wire [21:0] umul_54127;
  wire [21:0] add_54129;
  wire [15:0] sel_54134;
  wire [15:0] array_index_54135;
  wire [31:0] smod_54139;
  wire [15:0] array_index_54141;
  wire [31:0] smod_54145;
  wire [21:0] umul_54195;
  wire [15:0] add_54197;
  wire [15:0] sel_54202;
  wire [21:0] umul_54203;
  wire [15:0] add_54205;
  wire [15:0] sel_54210;
  wire [31:0] smod_54214;
  wire [31:0] smod_54219;
  wire [31:0] smod_54224;
  wire [31:0] smod_54229;
  wire [31:0] smod_54234;
  wire [31:0] smod_54239;
  wire [31:0] smod_54244;
  wire [31:0] smod_54249;
  wire [22:0] umul_54265;
  wire [20:0] add_54267;
  wire [15:0] sel_54272;
  wire [22:0] umul_54273;
  wire [20:0] add_54275;
  wire [15:0] sel_54280;
  wire [22:0] umul_54281;
  wire [22:0] add_54283;
  wire [15:0] sel_54288;
  wire [22:0] umul_54289;
  wire [22:0] add_54291;
  wire [15:0] sel_54296;
  wire [21:0] umul_54297;
  wire [20:0] add_54299;
  wire [15:0] sel_54304;
  wire [21:0] umul_54305;
  wire [20:0] add_54307;
  wire [15:0] sel_54312;
  wire [21:0] umul_54313;
  wire [21:0] add_54315;
  wire [15:0] sel_54320;
  wire [21:0] umul_54321;
  wire [21:0] add_54323;
  wire [15:0] sel_54328;
  wire [15:0] array_index_54329;
  wire [31:0] smod_54333;
  wire [15:0] array_index_54335;
  wire [31:0] smod_54339;
  wire [21:0] umul_54389;
  wire [15:0] add_54391;
  wire [15:0] sel_54396;
  wire [21:0] umul_54397;
  wire [15:0] add_54399;
  wire [15:0] sel_54404;
  wire [31:0] smod_54408;
  wire [31:0] smod_54413;
  wire [31:0] smod_54418;
  wire [31:0] smod_54423;
  wire [31:0] smod_54428;
  wire [31:0] smod_54433;
  wire [31:0] smod_54438;
  wire [31:0] smod_54443;
  wire [22:0] umul_54459;
  wire [20:0] add_54461;
  wire [15:0] sel_54466;
  wire [22:0] umul_54467;
  wire [20:0] add_54469;
  wire [15:0] sel_54474;
  wire [22:0] umul_54475;
  wire [22:0] add_54477;
  wire [15:0] sel_54482;
  wire [22:0] umul_54483;
  wire [22:0] add_54485;
  wire [15:0] sel_54490;
  wire [21:0] umul_54491;
  wire [20:0] add_54493;
  wire [15:0] sel_54498;
  wire [21:0] umul_54499;
  wire [20:0] add_54501;
  wire [15:0] sel_54506;
  wire [21:0] umul_54507;
  wire [21:0] add_54509;
  wire [15:0] sel_54514;
  wire [21:0] umul_54515;
  wire [21:0] add_54517;
  wire [15:0] sel_54522;
  wire [15:0] array_index_54523;
  wire [31:0] smod_54527;
  wire [15:0] array_index_54529;
  wire [31:0] smod_54533;
  wire [21:0] umul_54583;
  wire [15:0] add_54585;
  wire [15:0] sel_54590;
  wire [21:0] umul_54591;
  wire [15:0] add_54593;
  wire [15:0] sel_54598;
  wire [31:0] smod_54602;
  wire [31:0] smod_54607;
  wire [31:0] smod_54612;
  wire [31:0] smod_54617;
  wire [31:0] smod_54622;
  wire [31:0] smod_54627;
  wire [31:0] smod_54632;
  wire [31:0] smod_54637;
  wire [22:0] umul_54653;
  wire [20:0] add_54655;
  wire [15:0] sel_54660;
  wire [22:0] umul_54661;
  wire [20:0] add_54663;
  wire [15:0] sel_54668;
  wire [22:0] umul_54669;
  wire [22:0] add_54671;
  wire [15:0] sel_54676;
  wire [22:0] umul_54677;
  wire [22:0] add_54679;
  wire [15:0] sel_54684;
  wire [21:0] umul_54685;
  wire [20:0] add_54687;
  wire [15:0] sel_54692;
  wire [21:0] umul_54693;
  wire [20:0] add_54695;
  wire [15:0] sel_54700;
  wire [21:0] umul_54701;
  wire [21:0] add_54703;
  wire [15:0] sel_54708;
  wire [21:0] umul_54709;
  wire [21:0] add_54711;
  wire [15:0] sel_54716;
  wire [15:0] array_index_54717;
  wire [31:0] smod_54721;
  wire [15:0] array_index_54723;
  wire [31:0] smod_54727;
  wire [21:0] umul_54777;
  wire [15:0] add_54779;
  wire [15:0] sel_54784;
  wire [21:0] umul_54785;
  wire [15:0] add_54787;
  wire [15:0] sel_54792;
  wire [31:0] smod_54796;
  wire [31:0] smod_54801;
  wire [31:0] smod_54806;
  wire [31:0] smod_54811;
  wire [31:0] smod_54816;
  wire [31:0] smod_54821;
  wire [31:0] smod_54826;
  wire [31:0] smod_54831;
  wire [22:0] umul_54847;
  wire [20:0] add_54849;
  wire [15:0] sel_54854;
  wire [22:0] umul_54855;
  wire [20:0] add_54857;
  wire [15:0] sel_54862;
  wire [22:0] umul_54863;
  wire [22:0] add_54865;
  wire [15:0] sel_54870;
  wire [22:0] umul_54871;
  wire [22:0] add_54873;
  wire [15:0] sel_54878;
  wire [21:0] umul_54879;
  wire [20:0] add_54881;
  wire [15:0] sel_54886;
  wire [21:0] umul_54887;
  wire [20:0] add_54889;
  wire [15:0] sel_54894;
  wire [21:0] umul_54895;
  wire [21:0] add_54897;
  wire [15:0] sel_54902;
  wire [21:0] umul_54903;
  wire [21:0] add_54905;
  wire [15:0] sel_54910;
  wire [15:0] array_index_54911;
  wire [31:0] smod_54915;
  wire [15:0] array_index_54917;
  wire [31:0] smod_54921;
  wire [21:0] umul_54971;
  wire [15:0] add_54973;
  wire [15:0] sel_54978;
  wire [21:0] umul_54979;
  wire [15:0] add_54981;
  wire [15:0] sel_54986;
  wire [31:0] smod_54990;
  wire [31:0] smod_54995;
  wire [31:0] smod_55000;
  wire [31:0] smod_55005;
  wire [31:0] smod_55010;
  wire [31:0] smod_55015;
  wire [31:0] smod_55020;
  wire [31:0] smod_55025;
  wire [22:0] umul_55041;
  wire [20:0] add_55043;
  wire [15:0] sel_55048;
  wire [22:0] umul_55049;
  wire [20:0] add_55051;
  wire [15:0] sel_55056;
  wire [22:0] umul_55057;
  wire [22:0] add_55059;
  wire [15:0] sel_55064;
  wire [22:0] umul_55065;
  wire [22:0] add_55067;
  wire [15:0] sel_55072;
  wire [21:0] umul_55073;
  wire [20:0] add_55075;
  wire [15:0] sel_55080;
  wire [21:0] umul_55081;
  wire [20:0] add_55083;
  wire [15:0] sel_55088;
  wire [21:0] umul_55089;
  wire [21:0] add_55091;
  wire [15:0] sel_55096;
  wire [21:0] umul_55097;
  wire [21:0] add_55099;
  wire [15:0] sel_55104;
  wire [15:0] array_index_55105;
  wire [31:0] smod_55109;
  wire [15:0] array_index_55111;
  wire [31:0] smod_55115;
  wire [21:0] umul_55165;
  wire [15:0] add_55167;
  wire [15:0] sel_55172;
  wire [21:0] umul_55173;
  wire [15:0] add_55175;
  wire [15:0] sel_55180;
  wire [31:0] smod_55184;
  wire [31:0] smod_55189;
  wire [31:0] smod_55194;
  wire [31:0] smod_55199;
  wire [31:0] smod_55204;
  wire [31:0] smod_55209;
  wire [31:0] smod_55214;
  wire [31:0] smod_55219;
  wire [22:0] umul_55235;
  wire [20:0] add_55237;
  wire [15:0] sel_55242;
  wire [22:0] umul_55243;
  wire [20:0] add_55245;
  wire [15:0] sel_55250;
  wire [22:0] umul_55251;
  wire [22:0] add_55253;
  wire [15:0] sel_55258;
  wire [22:0] umul_55259;
  wire [22:0] add_55261;
  wire [15:0] sel_55266;
  wire [21:0] umul_55267;
  wire [20:0] add_55269;
  wire [15:0] sel_55274;
  wire [21:0] umul_55275;
  wire [20:0] add_55277;
  wire [15:0] sel_55282;
  wire [21:0] umul_55283;
  wire [21:0] add_55285;
  wire [15:0] sel_55290;
  wire [21:0] umul_55291;
  wire [21:0] add_55293;
  wire [15:0] sel_55298;
  wire [15:0] array_index_55299;
  wire [31:0] smod_55303;
  wire [15:0] array_index_55305;
  wire [31:0] smod_55309;
  wire [21:0] umul_55359;
  wire [15:0] add_55361;
  wire [15:0] sel_55366;
  wire [21:0] umul_55367;
  wire [15:0] add_55369;
  wire [15:0] sel_55374;
  wire [31:0] smod_55378;
  wire [31:0] smod_55383;
  wire [31:0] smod_55388;
  wire [31:0] smod_55393;
  wire [31:0] smod_55398;
  wire [31:0] smod_55403;
  wire [31:0] smod_55408;
  wire [31:0] smod_55413;
  wire [22:0] umul_55429;
  wire [20:0] add_55431;
  wire [15:0] sel_55436;
  wire [22:0] umul_55437;
  wire [20:0] add_55439;
  wire [15:0] sel_55444;
  wire [22:0] umul_55445;
  wire [22:0] add_55447;
  wire [15:0] sel_55452;
  wire [22:0] umul_55453;
  wire [22:0] add_55455;
  wire [15:0] sel_55460;
  wire [21:0] umul_55461;
  wire [20:0] add_55463;
  wire [15:0] sel_55468;
  wire [21:0] umul_55469;
  wire [20:0] add_55471;
  wire [15:0] sel_55476;
  wire [21:0] umul_55477;
  wire [21:0] add_55479;
  wire [15:0] sel_55484;
  wire [21:0] umul_55485;
  wire [21:0] add_55487;
  wire [15:0] sel_55492;
  wire [15:0] array_index_55493;
  wire [31:0] smod_55497;
  wire [15:0] array_index_55499;
  wire [31:0] smod_55503;
  wire [21:0] umul_55553;
  wire [15:0] add_55555;
  wire [15:0] sel_55560;
  wire [21:0] umul_55561;
  wire [15:0] add_55563;
  wire [15:0] sel_55568;
  wire [31:0] smod_55572;
  wire [31:0] smod_55577;
  wire [31:0] smod_55582;
  wire [31:0] smod_55587;
  wire [31:0] smod_55592;
  wire [31:0] smod_55597;
  wire [31:0] smod_55602;
  wire [31:0] smod_55607;
  wire [22:0] umul_55623;
  wire [20:0] add_55625;
  wire [15:0] sel_55630;
  wire [22:0] umul_55631;
  wire [20:0] add_55633;
  wire [15:0] sel_55638;
  wire [22:0] umul_55639;
  wire [22:0] add_55641;
  wire [15:0] sel_55646;
  wire [22:0] umul_55647;
  wire [22:0] add_55649;
  wire [15:0] sel_55654;
  wire [21:0] umul_55655;
  wire [20:0] add_55657;
  wire [15:0] sel_55662;
  wire [21:0] umul_55663;
  wire [20:0] add_55665;
  wire [15:0] sel_55670;
  wire [21:0] umul_55671;
  wire [21:0] add_55673;
  wire [15:0] sel_55678;
  wire [21:0] umul_55679;
  wire [21:0] add_55681;
  wire [15:0] sel_55686;
  wire [15:0] array_index_55687;
  wire [31:0] smod_55691;
  wire [15:0] array_index_55693;
  wire [31:0] smod_55697;
  wire [21:0] umul_55747;
  wire [15:0] add_55749;
  wire [15:0] sel_55754;
  wire [21:0] umul_55755;
  wire [15:0] add_55757;
  wire [15:0] sel_55762;
  wire [31:0] smod_55766;
  wire [31:0] smod_55771;
  wire [31:0] smod_55776;
  wire [31:0] smod_55781;
  wire [31:0] smod_55786;
  wire [31:0] smod_55791;
  wire [31:0] smod_55796;
  wire [31:0] smod_55801;
  wire [22:0] umul_55817;
  wire [20:0] add_55819;
  wire [15:0] sel_55824;
  wire [22:0] umul_55825;
  wire [20:0] add_55827;
  wire [15:0] sel_55832;
  wire [22:0] umul_55833;
  wire [22:0] add_55835;
  wire [15:0] sel_55840;
  wire [22:0] umul_55841;
  wire [22:0] add_55843;
  wire [15:0] sel_55848;
  wire [21:0] umul_55849;
  wire [20:0] add_55851;
  wire [15:0] sel_55856;
  wire [21:0] umul_55857;
  wire [20:0] add_55859;
  wire [15:0] sel_55864;
  wire [21:0] umul_55865;
  wire [21:0] add_55867;
  wire [15:0] sel_55872;
  wire [21:0] umul_55873;
  wire [21:0] add_55875;
  wire [15:0] sel_55880;
  wire [15:0] array_index_55881;
  wire [31:0] smod_55885;
  wire [15:0] array_index_55887;
  wire [31:0] smod_55891;
  wire [21:0] umul_55941;
  wire [15:0] add_55943;
  wire [15:0] sel_55948;
  wire [21:0] umul_55949;
  wire [15:0] add_55951;
  wire [15:0] sel_55956;
  wire [31:0] smod_55960;
  wire [31:0] smod_55965;
  wire [31:0] smod_55970;
  wire [31:0] smod_55975;
  wire [31:0] smod_55980;
  wire [31:0] smod_55985;
  wire [31:0] smod_55990;
  wire [31:0] smod_55995;
  wire [22:0] umul_56011;
  wire [20:0] add_56013;
  wire [15:0] sel_56018;
  wire [22:0] umul_56019;
  wire [20:0] add_56021;
  wire [15:0] sel_56026;
  wire [22:0] umul_56027;
  wire [22:0] add_56029;
  wire [15:0] sel_56034;
  wire [22:0] umul_56035;
  wire [22:0] add_56037;
  wire [15:0] sel_56042;
  wire [21:0] umul_56043;
  wire [20:0] add_56045;
  wire [15:0] sel_56050;
  wire [21:0] umul_56051;
  wire [20:0] add_56053;
  wire [15:0] sel_56058;
  wire [21:0] umul_56059;
  wire [21:0] add_56061;
  wire [15:0] sel_56066;
  wire [21:0] umul_56067;
  wire [21:0] add_56069;
  wire [15:0] sel_56074;
  wire [15:0] array_index_56075;
  wire [31:0] smod_56079;
  wire [15:0] array_index_56081;
  wire [31:0] smod_56085;
  wire [21:0] umul_56135;
  wire [15:0] add_56137;
  wire [15:0] sel_56142;
  wire [21:0] umul_56143;
  wire [15:0] add_56145;
  wire [15:0] sel_56150;
  wire [31:0] smod_56154;
  wire [31:0] smod_56159;
  wire [31:0] smod_56164;
  wire [31:0] smod_56169;
  wire [31:0] smod_56174;
  wire [31:0] smod_56179;
  wire [31:0] smod_56184;
  wire [31:0] smod_56189;
  wire [22:0] umul_56205;
  wire [20:0] add_56207;
  wire [15:0] sel_56212;
  wire [22:0] umul_56213;
  wire [20:0] add_56215;
  wire [15:0] sel_56220;
  wire [22:0] umul_56221;
  wire [22:0] add_56223;
  wire [15:0] sel_56228;
  wire [22:0] umul_56229;
  wire [22:0] add_56231;
  wire [15:0] sel_56236;
  wire [21:0] umul_56237;
  wire [20:0] add_56239;
  wire [15:0] sel_56244;
  wire [21:0] umul_56245;
  wire [20:0] add_56247;
  wire [15:0] sel_56252;
  wire [21:0] umul_56253;
  wire [21:0] add_56255;
  wire [15:0] sel_56260;
  wire [21:0] umul_56261;
  wire [21:0] add_56263;
  wire [15:0] sel_56268;
  wire [15:0] array_index_56269;
  wire [31:0] smod_56273;
  wire [15:0] array_index_56275;
  wire [31:0] smod_56279;
  wire [21:0] umul_56329;
  wire [15:0] add_56331;
  wire [15:0] sel_56336;
  wire [21:0] umul_56337;
  wire [15:0] add_56339;
  wire [15:0] sel_56344;
  wire [31:0] smod_56348;
  wire [31:0] smod_56353;
  wire [31:0] smod_56358;
  wire [31:0] smod_56363;
  wire [31:0] smod_56368;
  wire [31:0] smod_56373;
  wire [31:0] smod_56378;
  wire [31:0] smod_56383;
  wire [22:0] umul_56399;
  wire [20:0] add_56401;
  wire [15:0] sel_56406;
  wire [22:0] umul_56407;
  wire [20:0] add_56409;
  wire [15:0] sel_56414;
  wire [22:0] umul_56415;
  wire [22:0] add_56417;
  wire [15:0] sel_56422;
  wire [22:0] umul_56423;
  wire [22:0] add_56425;
  wire [15:0] sel_56430;
  wire [21:0] umul_56431;
  wire [20:0] add_56433;
  wire [15:0] sel_56438;
  wire [21:0] umul_56439;
  wire [20:0] add_56441;
  wire [15:0] sel_56446;
  wire [21:0] umul_56447;
  wire [21:0] add_56449;
  wire [15:0] sel_56454;
  wire [21:0] umul_56455;
  wire [21:0] add_56457;
  wire [15:0] sel_56462;
  wire [15:0] array_index_56463;
  wire [31:0] smod_56467;
  wire [15:0] array_index_56469;
  wire [31:0] smod_56473;
  wire [21:0] umul_56523;
  wire [15:0] add_56525;
  wire [15:0] sel_56530;
  wire [21:0] umul_56531;
  wire [15:0] add_56533;
  wire [15:0] sel_56538;
  wire [31:0] smod_56542;
  wire [31:0] smod_56547;
  wire [31:0] smod_56552;
  wire [31:0] smod_56557;
  wire [31:0] smod_56562;
  wire [31:0] smod_56567;
  wire [31:0] smod_56572;
  wire [31:0] smod_56577;
  wire [22:0] umul_56593;
  wire [20:0] add_56595;
  wire [15:0] sel_56600;
  wire [22:0] umul_56601;
  wire [20:0] add_56603;
  wire [15:0] sel_56608;
  wire [22:0] umul_56609;
  wire [22:0] add_56611;
  wire [15:0] sel_56616;
  wire [22:0] umul_56617;
  wire [22:0] add_56619;
  wire [15:0] sel_56624;
  wire [21:0] umul_56625;
  wire [20:0] add_56627;
  wire [15:0] sel_56632;
  wire [21:0] umul_56633;
  wire [20:0] add_56635;
  wire [15:0] sel_56640;
  wire [21:0] umul_56641;
  wire [21:0] add_56643;
  wire [15:0] sel_56648;
  wire [21:0] umul_56649;
  wire [21:0] add_56651;
  wire [15:0] sel_56656;
  wire [15:0] array_index_56657;
  wire [31:0] smod_56661;
  wire [15:0] array_index_56663;
  wire [31:0] smod_56667;
  wire [21:0] umul_56717;
  wire [15:0] add_56719;
  wire [15:0] sel_56724;
  wire [21:0] umul_56725;
  wire [15:0] add_56727;
  wire [15:0] sel_56732;
  wire [31:0] smod_56736;
  wire [31:0] smod_56741;
  wire [31:0] smod_56746;
  wire [31:0] smod_56751;
  wire [31:0] smod_56756;
  wire [31:0] smod_56761;
  wire [31:0] smod_56766;
  wire [31:0] smod_56771;
  wire [22:0] umul_56787;
  wire [20:0] add_56789;
  wire [15:0] sel_56794;
  wire [22:0] umul_56795;
  wire [20:0] add_56797;
  wire [15:0] sel_56802;
  wire [22:0] umul_56803;
  wire [22:0] add_56805;
  wire [15:0] sel_56810;
  wire [22:0] umul_56811;
  wire [22:0] add_56813;
  wire [15:0] sel_56818;
  wire [21:0] umul_56819;
  wire [20:0] add_56821;
  wire [15:0] sel_56826;
  wire [21:0] umul_56827;
  wire [20:0] add_56829;
  wire [15:0] sel_56834;
  wire [21:0] umul_56835;
  wire [21:0] add_56837;
  wire [15:0] sel_56842;
  wire [21:0] umul_56843;
  wire [21:0] add_56845;
  wire [15:0] sel_56850;
  wire [15:0] array_index_56851;
  wire [31:0] smod_56855;
  wire [15:0] array_index_56857;
  wire [31:0] smod_56861;
  wire [21:0] umul_56911;
  wire [15:0] add_56913;
  wire [15:0] sel_56918;
  wire [21:0] umul_56919;
  wire [15:0] add_56921;
  wire [15:0] sel_56926;
  wire [31:0] smod_56930;
  wire [31:0] smod_56935;
  wire [31:0] smod_56940;
  wire [31:0] smod_56945;
  wire [31:0] smod_56950;
  wire [31:0] smod_56955;
  wire [31:0] smod_56960;
  wire [31:0] smod_56965;
  wire [22:0] umul_56981;
  wire [20:0] add_56983;
  wire [15:0] sel_56988;
  wire [22:0] umul_56989;
  wire [20:0] add_56991;
  wire [15:0] sel_56996;
  wire [22:0] umul_56997;
  wire [22:0] add_56999;
  wire [15:0] sel_57004;
  wire [22:0] umul_57005;
  wire [22:0] add_57007;
  wire [15:0] sel_57012;
  wire [21:0] umul_57013;
  wire [20:0] add_57015;
  wire [15:0] sel_57020;
  wire [21:0] umul_57021;
  wire [20:0] add_57023;
  wire [15:0] sel_57028;
  wire [21:0] umul_57029;
  wire [21:0] add_57031;
  wire [15:0] sel_57036;
  wire [21:0] umul_57037;
  wire [21:0] add_57039;
  wire [15:0] sel_57044;
  wire [15:0] array_index_57045;
  wire [31:0] smod_57049;
  wire [15:0] array_index_57051;
  wire [31:0] smod_57055;
  wire [21:0] umul_57105;
  wire [15:0] add_57107;
  wire [15:0] sel_57112;
  wire [21:0] umul_57113;
  wire [15:0] add_57115;
  wire [15:0] sel_57120;
  wire [31:0] smod_57124;
  wire [31:0] smod_57129;
  wire [31:0] smod_57134;
  wire [31:0] smod_57139;
  wire [31:0] smod_57144;
  wire [31:0] smod_57149;
  wire [31:0] smod_57154;
  wire [31:0] smod_57159;
  wire [22:0] umul_57175;
  wire [20:0] add_57177;
  wire [15:0] sel_57182;
  wire [22:0] umul_57183;
  wire [20:0] add_57185;
  wire [15:0] sel_57190;
  wire [22:0] umul_57191;
  wire [22:0] add_57193;
  wire [15:0] sel_57198;
  wire [22:0] umul_57199;
  wire [22:0] add_57201;
  wire [15:0] sel_57206;
  wire [21:0] umul_57207;
  wire [20:0] add_57209;
  wire [15:0] sel_57214;
  wire [21:0] umul_57215;
  wire [20:0] add_57217;
  wire [15:0] sel_57222;
  wire [21:0] umul_57223;
  wire [21:0] add_57225;
  wire [15:0] sel_57230;
  wire [21:0] umul_57231;
  wire [21:0] add_57233;
  wire [15:0] sel_57238;
  wire [15:0] array_index_57239;
  wire [31:0] smod_57243;
  wire [15:0] array_index_57245;
  wire [31:0] smod_57249;
  wire [21:0] umul_57299;
  wire [15:0] add_57301;
  wire [15:0] sel_57306;
  wire [21:0] umul_57307;
  wire [15:0] add_57309;
  wire [15:0] sel_57314;
  wire [31:0] smod_57318;
  wire [31:0] smod_57323;
  wire [31:0] smod_57328;
  wire [31:0] smod_57333;
  wire [31:0] smod_57338;
  wire [31:0] smod_57343;
  wire [31:0] smod_57348;
  wire [31:0] smod_57353;
  wire [22:0] umul_57369;
  wire [20:0] add_57371;
  wire [15:0] sel_57376;
  wire [22:0] umul_57377;
  wire [20:0] add_57379;
  wire [15:0] sel_57384;
  wire [22:0] umul_57385;
  wire [22:0] add_57387;
  wire [15:0] sel_57392;
  wire [22:0] umul_57393;
  wire [22:0] add_57395;
  wire [15:0] sel_57400;
  wire [21:0] umul_57401;
  wire [20:0] add_57403;
  wire [15:0] sel_57408;
  wire [21:0] umul_57409;
  wire [20:0] add_57411;
  wire [15:0] sel_57416;
  wire [21:0] umul_57417;
  wire [21:0] add_57419;
  wire [15:0] sel_57424;
  wire [21:0] umul_57425;
  wire [21:0] add_57427;
  wire [15:0] sel_57432;
  wire [15:0] array_index_57433;
  wire [31:0] smod_57437;
  wire [15:0] array_index_57439;
  wire [31:0] smod_57443;
  wire [21:0] umul_57493;
  wire [15:0] add_57495;
  wire [15:0] sel_57500;
  wire [21:0] umul_57501;
  wire [15:0] add_57503;
  wire [15:0] sel_57508;
  wire [31:0] smod_57512;
  wire [31:0] smod_57517;
  wire [31:0] smod_57522;
  wire [31:0] smod_57527;
  wire [31:0] smod_57532;
  wire [31:0] smod_57537;
  wire [31:0] smod_57542;
  wire [31:0] smod_57547;
  wire [22:0] umul_57561;
  wire [20:0] add_57563;
  wire [15:0] sel_57568;
  wire [22:0] umul_57569;
  wire [20:0] add_57571;
  wire [15:0] sel_57576;
  wire [22:0] umul_57577;
  wire [22:0] add_57579;
  wire [15:0] sel_57584;
  wire [22:0] umul_57585;
  wire [22:0] add_57587;
  wire [15:0] sel_57592;
  wire [21:0] umul_57593;
  wire [20:0] add_57595;
  wire [15:0] sel_57600;
  wire [21:0] umul_57601;
  wire [20:0] add_57603;
  wire [15:0] sel_57608;
  wire [21:0] umul_57609;
  wire [21:0] add_57611;
  wire [15:0] sel_57616;
  wire [21:0] umul_57617;
  wire [21:0] add_57619;
  wire [15:0] sel_57624;
  wire [31:0] smod_57627;
  wire [31:0] smod_57631;
  wire [15:0] add_57682;
  wire [15:0] sel_57687;
  wire [15:0] add_57689;
  wire [15:0] sel_57694;
  wire [31:0] smod_57698;
  wire [31:0] smod_57703;
  wire [31:0] smod_57708;
  wire [31:0] smod_57713;
  wire [31:0] smod_57718;
  wire [31:0] smod_57723;
  wire [31:0] smod_57727;
  wire [31:0] smod_57731;
  wire [22:0] umul_57741;
  wire [20:0] add_57743;
  wire [15:0] sel_57748;
  wire [22:0] umul_57749;
  wire [20:0] add_57751;
  wire [15:0] sel_57756;
  wire [22:0] umul_57757;
  wire [22:0] add_57759;
  wire [15:0] sel_57764;
  wire [22:0] umul_57765;
  wire [22:0] add_57767;
  wire [15:0] sel_57772;
  wire [21:0] umul_57773;
  wire [20:0] add_57775;
  wire [15:0] sel_57780;
  wire [21:0] umul_57781;
  wire [20:0] add_57783;
  wire [15:0] sel_57788;
  wire [21:0] add_57790;
  wire [15:0] sel_57795;
  wire [21:0] add_57797;
  wire [15:0] sel_57802;
  wire [31:0] smod_57803;
  wire [31:0] smod_57805;
  wire [15:0] sel_57854;
  wire [15:0] sel_57858;
  wire [31:0] smod_57862;
  wire [31:0] smod_57867;
  wire [31:0] smod_57872;
  wire [31:0] smod_57877;
  wire [31:0] smod_57881;
  wire [31:0] smod_57885;
  wire [31:0] smod_57887;
  wire [31:0] smod_57889;
  wire [22:0] umul_57895;
  wire [20:0] add_57897;
  wire [15:0] sel_57902;
  wire [22:0] umul_57903;
  wire [20:0] add_57905;
  wire [15:0] sel_57910;
  wire [22:0] umul_57911;
  wire [22:0] add_57913;
  wire [15:0] sel_57918;
  wire [22:0] umul_57919;
  wire [22:0] add_57921;
  wire [15:0] sel_57926;
  wire [20:0] add_57928;
  wire [15:0] sel_57933;
  wire [20:0] add_57935;
  wire [15:0] sel_57940;
  wire [15:0] sel_57944;
  wire [15:0] sel_57948;
  wire [31:0] smod_57992;
  wire [31:0] smod_57997;
  wire [31:0] smod_58001;
  wire [31:0] smod_58005;
  wire [31:0] smod_58007;
  wire [31:0] smod_58009;
  wire [22:0] umul_58015;
  wire [20:0] add_58017;
  wire [15:0] sel_58022;
  wire [22:0] umul_58023;
  wire [20:0] add_58025;
  wire [15:0] sel_58030;
  wire [22:0] add_58032;
  wire [15:0] sel_58037;
  wire [22:0] add_58039;
  wire [15:0] sel_58044;
  wire [15:0] sel_58048;
  wire [15:0] sel_58052;
  wire [1:0] concat_58055;
  wire [1:0] add_58082;
  wire [31:0] smod_58085;
  wire [31:0] smod_58089;
  wire [31:0] smod_58091;
  wire [31:0] smod_58093;
  wire [20:0] add_58100;
  wire [15:0] sel_58105;
  wire [20:0] add_58107;
  wire [15:0] sel_58112;
  wire [15:0] sel_58116;
  wire [15:0] sel_58120;
  wire [2:0] concat_58123;
  wire [2:0] add_58138;
  wire [31:0] smod_58139;
  wire [31:0] smod_58141;
  wire [15:0] sel_58150;
  wire [15:0] sel_58154;
  wire [3:0] concat_58157;
  wire [3:0] add_58164;
  wire [4:0] concat_58171;
  wire [4:0] add_58174;
  assign array_index_52333 = set1_unflattened[5'h00];
  assign array_index_52335 = set2_unflattened[5'h00];
  assign umul_52337 = umul22b_16b_x_6b(array_index_52333, 6'h35);
  assign umul_52338 = umul22b_16b_x_6b(array_index_52335, 6'h35);
  assign umul_52347 = umul22b_16b_x_6b(array_index_52333, 6'h3b);
  assign umul_52348 = umul22b_16b_x_6b(array_index_52335, 6'h3b);
  assign array_index_52349 = set1_unflattened[5'h01];
  assign array_index_52353 = set2_unflattened[5'h01];
  assign umul_52361 = umul22b_16b_x_6b(array_index_52349, 6'h35);
  assign add_52363 = {1'h0, umul_52337[21:7]} + 16'h007d;
  assign umul_52365 = umul22b_16b_x_6b(array_index_52353, 6'h35);
  assign add_52367 = {1'h0, umul_52338[21:7]} + 16'h007d;
  assign umul_52387 = umul22b_16b_x_6b(array_index_52333, 6'h3d);
  assign umul_52388 = umul22b_16b_x_6b(array_index_52335, 6'h3d);
  assign umul_52389 = umul22b_16b_x_6b(array_index_52349, 6'h3b);
  assign add_52391 = {1'h0, umul_52347[21:1]} + 22'h00_1f59;
  assign umul_52393 = umul22b_16b_x_6b(array_index_52353, 6'h3b);
  assign add_52395 = {1'h0, umul_52348[21:1]} + 22'h00_1f59;
  assign array_index_52397 = set1_unflattened[5'h02];
  assign smod_52401 = $unsigned($signed({9'h000, add_52363, umul_52337[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_52402 = set2_unflattened[5'h02];
  assign smod_52406 = $unsigned($signed({9'h000, add_52367, umul_52338[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_52419 = umul22b_16b_x_6b(array_index_52397, 6'h35);
  assign add_52421 = {1'h0, umul_52361[21:7]} + 16'h007d;
  assign umul_52425 = umul22b_16b_x_6b(array_index_52402, 6'h35);
  assign add_52427 = {1'h0, umul_52365[21:7]} + 16'h007d;
  assign smod_52442 = $unsigned($signed({9'h000, add_52391, umul_52347[0]}) % $signed(32'h0000_3ffd));
  assign smod_52446 = $unsigned($signed({9'h000, add_52395, umul_52348[0]}) % $signed(32'h0000_3ffd));
  assign umul_52461 = umul23b_16b_x_7b(array_index_52333, 7'h47);
  assign umul_52462 = umul23b_16b_x_7b(array_index_52335, 7'h47);
  assign umul_52463 = umul22b_16b_x_6b(array_index_52349, 6'h3d);
  assign add_52465 = {1'h0, umul_52387[21:2]} + 21'h00_0fb9;
  assign umul_52467 = umul22b_16b_x_6b(array_index_52353, 6'h3d);
  assign add_52469 = {1'h0, umul_52388[21:2]} + 21'h00_0fb9;
  assign umul_52471 = umul22b_16b_x_6b(array_index_52397, 6'h3b);
  assign add_52473 = {1'h0, umul_52389[21:1]} + 22'h00_1f59;
  assign umul_52477 = umul22b_16b_x_6b(array_index_52402, 6'h3b);
  assign add_52479 = {1'h0, umul_52393[21:1]} + 22'h00_1f59;
  assign array_index_52483 = set1_unflattened[5'h03];
  assign smod_52487 = $unsigned($signed({9'h000, add_52421, umul_52361[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_52490 = set2_unflattened[5'h03];
  assign smod_52494 = $unsigned($signed({9'h000, add_52427, umul_52365[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_52521 = umul22b_16b_x_6b(array_index_52483, 6'h35);
  assign add_52523 = {1'h0, umul_52419[21:7]} + 16'h007d;
  assign sel_52528 = $signed({1'h0, smod_52401[15:0]}) < $signed(17'h0_3ffd) ? smod_52401[15:0] : 16'h3ffd;
  assign umul_52529 = umul22b_16b_x_6b(array_index_52490, 6'h35);
  assign add_52531 = {1'h0, umul_52425[21:7]} + 16'h007d;
  assign sel_52536 = $signed({1'h0, smod_52406[15:0]}) < $signed(17'h0_3ffd) ? smod_52406[15:0] : 16'h3ffd;
  assign smod_52548 = $unsigned($signed({9'h000, add_52465, umul_52387[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_52552 = $unsigned($signed({9'h000, add_52469, umul_52388[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_52556 = $unsigned($signed({9'h000, add_52473, umul_52389[0]}) % $signed(32'h0000_3ffd));
  assign smod_52562 = $unsigned($signed({9'h000, add_52479, umul_52393[0]}) % $signed(32'h0000_3ffd));
  assign umul_52579 = umul23b_16b_x_7b(array_index_52333, 7'h49);
  assign umul_52580 = umul23b_16b_x_7b(array_index_52335, 7'h49);
  assign umul_52581 = umul23b_16b_x_7b(array_index_52349, 7'h47);
  assign add_52583 = {1'h0, umul_52461[22:1]} + 23'h00_1f8b;
  assign umul_52585 = umul23b_16b_x_7b(array_index_52353, 7'h47);
  assign add_52587 = {1'h0, umul_52462[22:1]} + 23'h00_1f8b;
  assign umul_52589 = umul22b_16b_x_6b(array_index_52397, 6'h3d);
  assign add_52591 = {1'h0, umul_52463[21:2]} + 21'h00_0fb9;
  assign umul_52595 = umul22b_16b_x_6b(array_index_52402, 6'h3d);
  assign add_52597 = {1'h0, umul_52467[21:2]} + 21'h00_0fb9;
  assign umul_52601 = umul22b_16b_x_6b(array_index_52483, 6'h3b);
  assign add_52603 = {1'h0, umul_52471[21:1]} + 22'h00_1f59;
  assign sel_52608 = $signed({1'h0, smod_52442[15:0]}) < $signed(17'h0_3ffd) ? smod_52442[15:0] : 16'h3ffd;
  assign umul_52609 = umul22b_16b_x_6b(array_index_52490, 6'h3b);
  assign add_52611 = {1'h0, umul_52477[21:1]} + 22'h00_1f59;
  assign sel_52616 = $signed({1'h0, smod_52446[15:0]}) < $signed(17'h0_3ffd) ? smod_52446[15:0] : 16'h3ffd;
  assign array_index_52617 = set1_unflattened[5'h04];
  assign smod_52621 = $unsigned($signed({9'h000, add_52523, umul_52419[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_52623 = set2_unflattened[5'h04];
  assign smod_52627 = $unsigned($signed({9'h000, add_52531, umul_52425[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_52665 = umul22b_16b_x_6b(array_index_52617, 6'h35);
  assign add_52667 = {1'h0, umul_52521[21:7]} + 16'h007d;
  assign sel_52672 = $signed({1'h0, smod_52487[15:0]}) < $signed({1'h0, sel_52528}) ? smod_52487[15:0] : sel_52528;
  assign umul_52673 = umul22b_16b_x_6b(array_index_52623, 6'h35);
  assign add_52675 = {1'h0, umul_52529[21:7]} + 16'h007d;
  assign sel_52680 = $signed({1'h0, smod_52494[15:0]}) < $signed({1'h0, sel_52536}) ? smod_52494[15:0] : sel_52536;
  assign smod_52690 = $unsigned($signed({8'h00, add_52583, umul_52461[0]}) % $signed(32'h0000_3ffd));
  assign smod_52694 = $unsigned($signed({8'h00, add_52587, umul_52462[0]}) % $signed(32'h0000_3ffd));
  assign smod_52698 = $unsigned($signed({9'h000, add_52591, umul_52463[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_52704 = $unsigned($signed({9'h000, add_52597, umul_52467[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_52710 = $unsigned($signed({9'h000, add_52603, umul_52471[0]}) % $signed(32'h0000_3ffd));
  assign smod_52715 = $unsigned($signed({9'h000, add_52611, umul_52477[0]}) % $signed(32'h0000_3ffd));
  assign umul_52731 = umul23b_16b_x_7b(array_index_52349, 7'h49);
  assign add_52733 = {1'h0, umul_52579[22:3]} + 21'h00_07e9;
  assign umul_52735 = umul23b_16b_x_7b(array_index_52353, 7'h49);
  assign add_52737 = {1'h0, umul_52580[22:3]} + 21'h00_07e9;
  assign umul_52739 = umul23b_16b_x_7b(array_index_52397, 7'h47);
  assign add_52741 = {1'h0, umul_52581[22:1]} + 23'h00_1f8b;
  assign umul_52745 = umul23b_16b_x_7b(array_index_52402, 7'h47);
  assign add_52747 = {1'h0, umul_52585[22:1]} + 23'h00_1f8b;
  assign umul_52751 = umul22b_16b_x_6b(array_index_52483, 6'h3d);
  assign add_52753 = {1'h0, umul_52589[21:2]} + 21'h00_0fb9;
  assign sel_52758 = $signed({1'h0, smod_52548[15:0]}) < $signed(17'h0_3ffd) ? smod_52548[15:0] : 16'h3ffd;
  assign umul_52759 = umul22b_16b_x_6b(array_index_52490, 6'h3d);
  assign add_52761 = {1'h0, umul_52595[21:2]} + 21'h00_0fb9;
  assign sel_52766 = $signed({1'h0, smod_52552[15:0]}) < $signed(17'h0_3ffd) ? smod_52552[15:0] : 16'h3ffd;
  assign umul_52767 = umul22b_16b_x_6b(array_index_52617, 6'h3b);
  assign add_52769 = {1'h0, umul_52601[21:1]} + 22'h00_1f59;
  assign sel_52774 = $signed({1'h0, smod_52556[15:0]}) < $signed({1'h0, sel_52608}) ? smod_52556[15:0] : sel_52608;
  assign umul_52775 = umul22b_16b_x_6b(array_index_52623, 6'h3b);
  assign add_52777 = {1'h0, umul_52609[21:1]} + 22'h00_1f59;
  assign sel_52782 = $signed({1'h0, smod_52562[15:0]}) < $signed({1'h0, sel_52616}) ? smod_52562[15:0] : sel_52616;
  assign array_index_52783 = set1_unflattened[5'h05];
  assign smod_52787 = $unsigned($signed({9'h000, add_52667, umul_52521[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_52789 = set2_unflattened[5'h05];
  assign smod_52793 = $unsigned($signed({9'h000, add_52675, umul_52529[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_52839 = umul22b_16b_x_6b(array_index_52783, 6'h35);
  assign add_52841 = {1'h0, umul_52665[21:7]} + 16'h007d;
  assign sel_52846 = $signed({1'h0, smod_52621[15:0]}) < $signed({1'h0, sel_52672}) ? smod_52621[15:0] : sel_52672;
  assign umul_52847 = umul22b_16b_x_6b(array_index_52789, 6'h35);
  assign add_52849 = {1'h0, umul_52673[21:7]} + 16'h007d;
  assign sel_52854 = $signed({1'h0, smod_52627[15:0]}) < $signed({1'h0, sel_52680}) ? smod_52627[15:0] : sel_52680;
  assign smod_52858 = $unsigned($signed({8'h00, add_52733, umul_52579[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_52862 = $unsigned($signed({8'h00, add_52737, umul_52580[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_52866 = $unsigned($signed({8'h00, add_52741, umul_52581[0]}) % $signed(32'h0000_3ffd));
  assign smod_52872 = $unsigned($signed({8'h00, add_52747, umul_52585[0]}) % $signed(32'h0000_3ffd));
  assign smod_52878 = $unsigned($signed({9'h000, add_52753, umul_52589[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_52883 = $unsigned($signed({9'h000, add_52761, umul_52595[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_52888 = $unsigned($signed({9'h000, add_52769, umul_52601[0]}) % $signed(32'h0000_3ffd));
  assign smod_52893 = $unsigned($signed({9'h000, add_52777, umul_52609[0]}) % $signed(32'h0000_3ffd));
  assign umul_52909 = umul23b_16b_x_7b(array_index_52397, 7'h49);
  assign add_52911 = {1'h0, umul_52731[22:3]} + 21'h00_07e9;
  assign umul_52915 = umul23b_16b_x_7b(array_index_52402, 7'h49);
  assign add_52917 = {1'h0, umul_52735[22:3]} + 21'h00_07e9;
  assign umul_52921 = umul23b_16b_x_7b(array_index_52483, 7'h47);
  assign add_52923 = {1'h0, umul_52739[22:1]} + 23'h00_1f8b;
  assign sel_52928 = $signed({1'h0, smod_52690[15:0]}) < $signed(17'h0_3ffd) ? smod_52690[15:0] : 16'h3ffd;
  assign umul_52929 = umul23b_16b_x_7b(array_index_52490, 7'h47);
  assign add_52931 = {1'h0, umul_52745[22:1]} + 23'h00_1f8b;
  assign sel_52936 = $signed({1'h0, smod_52694[15:0]}) < $signed(17'h0_3ffd) ? smod_52694[15:0] : 16'h3ffd;
  assign umul_52937 = umul22b_16b_x_6b(array_index_52617, 6'h3d);
  assign add_52939 = {1'h0, umul_52751[21:2]} + 21'h00_0fb9;
  assign sel_52944 = $signed({1'h0, smod_52698[15:0]}) < $signed({1'h0, sel_52758}) ? smod_52698[15:0] : sel_52758;
  assign umul_52945 = umul22b_16b_x_6b(array_index_52623, 6'h3d);
  assign add_52947 = {1'h0, umul_52759[21:2]} + 21'h00_0fb9;
  assign sel_52952 = $signed({1'h0, smod_52704[15:0]}) < $signed({1'h0, sel_52766}) ? smod_52704[15:0] : sel_52766;
  assign umul_52953 = umul22b_16b_x_6b(array_index_52783, 6'h3b);
  assign add_52955 = {1'h0, umul_52767[21:1]} + 22'h00_1f59;
  assign sel_52960 = $signed({1'h0, smod_52710[15:0]}) < $signed({1'h0, sel_52774}) ? smod_52710[15:0] : sel_52774;
  assign umul_52961 = umul22b_16b_x_6b(array_index_52789, 6'h3b);
  assign add_52963 = {1'h0, umul_52775[21:1]} + 22'h00_1f59;
  assign sel_52968 = $signed({1'h0, smod_52715[15:0]}) < $signed({1'h0, sel_52782}) ? smod_52715[15:0] : sel_52782;
  assign array_index_52969 = set1_unflattened[5'h06];
  assign smod_52973 = $unsigned($signed({9'h000, add_52841, umul_52665[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_52975 = set2_unflattened[5'h06];
  assign smod_52979 = $unsigned($signed({9'h000, add_52849, umul_52673[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_53029 = umul22b_16b_x_6b(array_index_52969, 6'h35);
  assign add_53031 = {1'h0, umul_52839[21:7]} + 16'h007d;
  assign sel_53036 = $signed({1'h0, smod_52787[15:0]}) < $signed({1'h0, sel_52846}) ? smod_52787[15:0] : sel_52846;
  assign umul_53037 = umul22b_16b_x_6b(array_index_52975, 6'h35);
  assign add_53039 = {1'h0, umul_52847[21:7]} + 16'h007d;
  assign sel_53044 = $signed({1'h0, smod_52793[15:0]}) < $signed({1'h0, sel_52854}) ? smod_52793[15:0] : sel_52854;
  assign smod_53048 = $unsigned($signed({8'h00, add_52911, umul_52731[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53054 = $unsigned($signed({8'h00, add_52917, umul_52735[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53060 = $unsigned($signed({8'h00, add_52923, umul_52739[0]}) % $signed(32'h0000_3ffd));
  assign smod_53065 = $unsigned($signed({8'h00, add_52931, umul_52745[0]}) % $signed(32'h0000_3ffd));
  assign smod_53070 = $unsigned($signed({9'h000, add_52939, umul_52751[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53075 = $unsigned($signed({9'h000, add_52947, umul_52759[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53080 = $unsigned($signed({9'h000, add_52955, umul_52767[0]}) % $signed(32'h0000_3ffd));
  assign smod_53085 = $unsigned($signed({9'h000, add_52963, umul_52775[0]}) % $signed(32'h0000_3ffd));
  assign umul_53101 = umul23b_16b_x_7b(array_index_52483, 7'h49);
  assign add_53103 = {1'h0, umul_52909[22:3]} + 21'h00_07e9;
  assign sel_53108 = $signed({1'h0, smod_52858[15:0]}) < $signed(17'h0_3ffd) ? smod_52858[15:0] : 16'h3ffd;
  assign umul_53109 = umul23b_16b_x_7b(array_index_52490, 7'h49);
  assign add_53111 = {1'h0, umul_52915[22:3]} + 21'h00_07e9;
  assign sel_53116 = $signed({1'h0, smod_52862[15:0]}) < $signed(17'h0_3ffd) ? smod_52862[15:0] : 16'h3ffd;
  assign umul_53117 = umul23b_16b_x_7b(array_index_52617, 7'h47);
  assign add_53119 = {1'h0, umul_52921[22:1]} + 23'h00_1f8b;
  assign sel_53124 = $signed({1'h0, smod_52866[15:0]}) < $signed({1'h0, sel_52928}) ? smod_52866[15:0] : sel_52928;
  assign umul_53125 = umul23b_16b_x_7b(array_index_52623, 7'h47);
  assign add_53127 = {1'h0, umul_52929[22:1]} + 23'h00_1f8b;
  assign sel_53132 = $signed({1'h0, smod_52872[15:0]}) < $signed({1'h0, sel_52936}) ? smod_52872[15:0] : sel_52936;
  assign umul_53133 = umul22b_16b_x_6b(array_index_52783, 6'h3d);
  assign add_53135 = {1'h0, umul_52937[21:2]} + 21'h00_0fb9;
  assign sel_53140 = $signed({1'h0, smod_52878[15:0]}) < $signed({1'h0, sel_52944}) ? smod_52878[15:0] : sel_52944;
  assign umul_53141 = umul22b_16b_x_6b(array_index_52789, 6'h3d);
  assign add_53143 = {1'h0, umul_52945[21:2]} + 21'h00_0fb9;
  assign sel_53148 = $signed({1'h0, smod_52883[15:0]}) < $signed({1'h0, sel_52952}) ? smod_52883[15:0] : sel_52952;
  assign umul_53149 = umul22b_16b_x_6b(array_index_52969, 6'h3b);
  assign add_53151 = {1'h0, umul_52953[21:1]} + 22'h00_1f59;
  assign sel_53156 = $signed({1'h0, smod_52888[15:0]}) < $signed({1'h0, sel_52960}) ? smod_52888[15:0] : sel_52960;
  assign umul_53157 = umul22b_16b_x_6b(array_index_52975, 6'h3b);
  assign add_53159 = {1'h0, umul_52961[21:1]} + 22'h00_1f59;
  assign sel_53164 = $signed({1'h0, smod_52893[15:0]}) < $signed({1'h0, sel_52968}) ? smod_52893[15:0] : sel_52968;
  assign array_index_53165 = set1_unflattened[5'h07];
  assign smod_53169 = $unsigned($signed({9'h000, add_53031, umul_52839[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_53171 = set2_unflattened[5'h07];
  assign smod_53175 = $unsigned($signed({9'h000, add_53039, umul_52847[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_53225 = umul22b_16b_x_6b(array_index_53165, 6'h35);
  assign add_53227 = {1'h0, umul_53029[21:7]} + 16'h007d;
  assign sel_53232 = $signed({1'h0, smod_52973[15:0]}) < $signed({1'h0, sel_53036}) ? smod_52973[15:0] : sel_53036;
  assign umul_53233 = umul22b_16b_x_6b(array_index_53171, 6'h35);
  assign add_53235 = {1'h0, umul_53037[21:7]} + 16'h007d;
  assign sel_53240 = $signed({1'h0, smod_52979[15:0]}) < $signed({1'h0, sel_53044}) ? smod_52979[15:0] : sel_53044;
  assign smod_53244 = $unsigned($signed({8'h00, add_53103, umul_52909[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53249 = $unsigned($signed({8'h00, add_53111, umul_52915[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53254 = $unsigned($signed({8'h00, add_53119, umul_52921[0]}) % $signed(32'h0000_3ffd));
  assign smod_53259 = $unsigned($signed({8'h00, add_53127, umul_52929[0]}) % $signed(32'h0000_3ffd));
  assign smod_53264 = $unsigned($signed({9'h000, add_53135, umul_52937[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53269 = $unsigned($signed({9'h000, add_53143, umul_52945[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53274 = $unsigned($signed({9'h000, add_53151, umul_52953[0]}) % $signed(32'h0000_3ffd));
  assign smod_53279 = $unsigned($signed({9'h000, add_53159, umul_52961[0]}) % $signed(32'h0000_3ffd));
  assign umul_53295 = umul23b_16b_x_7b(array_index_52617, 7'h49);
  assign add_53297 = {1'h0, umul_53101[22:3]} + 21'h00_07e9;
  assign sel_53302 = $signed({1'h0, smod_53048[15:0]}) < $signed({1'h0, sel_53108}) ? smod_53048[15:0] : sel_53108;
  assign umul_53303 = umul23b_16b_x_7b(array_index_52623, 7'h49);
  assign add_53305 = {1'h0, umul_53109[22:3]} + 21'h00_07e9;
  assign sel_53310 = $signed({1'h0, smod_53054[15:0]}) < $signed({1'h0, sel_53116}) ? smod_53054[15:0] : sel_53116;
  assign umul_53311 = umul23b_16b_x_7b(array_index_52783, 7'h47);
  assign add_53313 = {1'h0, umul_53117[22:1]} + 23'h00_1f8b;
  assign sel_53318 = $signed({1'h0, smod_53060[15:0]}) < $signed({1'h0, sel_53124}) ? smod_53060[15:0] : sel_53124;
  assign umul_53319 = umul23b_16b_x_7b(array_index_52789, 7'h47);
  assign add_53321 = {1'h0, umul_53125[22:1]} + 23'h00_1f8b;
  assign sel_53326 = $signed({1'h0, smod_53065[15:0]}) < $signed({1'h0, sel_53132}) ? smod_53065[15:0] : sel_53132;
  assign umul_53327 = umul22b_16b_x_6b(array_index_52969, 6'h3d);
  assign add_53329 = {1'h0, umul_53133[21:2]} + 21'h00_0fb9;
  assign sel_53334 = $signed({1'h0, smod_53070[15:0]}) < $signed({1'h0, sel_53140}) ? smod_53070[15:0] : sel_53140;
  assign umul_53335 = umul22b_16b_x_6b(array_index_52975, 6'h3d);
  assign add_53337 = {1'h0, umul_53141[21:2]} + 21'h00_0fb9;
  assign sel_53342 = $signed({1'h0, smod_53075[15:0]}) < $signed({1'h0, sel_53148}) ? smod_53075[15:0] : sel_53148;
  assign umul_53343 = umul22b_16b_x_6b(array_index_53165, 6'h3b);
  assign add_53345 = {1'h0, umul_53149[21:1]} + 22'h00_1f59;
  assign sel_53350 = $signed({1'h0, smod_53080[15:0]}) < $signed({1'h0, sel_53156}) ? smod_53080[15:0] : sel_53156;
  assign umul_53351 = umul22b_16b_x_6b(array_index_53171, 6'h3b);
  assign add_53353 = {1'h0, umul_53157[21:1]} + 22'h00_1f59;
  assign sel_53358 = $signed({1'h0, smod_53085[15:0]}) < $signed({1'h0, sel_53164}) ? smod_53085[15:0] : sel_53164;
  assign array_index_53359 = set1_unflattened[5'h08];
  assign smod_53363 = $unsigned($signed({9'h000, add_53227, umul_53029[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_53365 = set2_unflattened[5'h08];
  assign smod_53369 = $unsigned($signed({9'h000, add_53235, umul_53037[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_53419 = umul22b_16b_x_6b(array_index_53359, 6'h35);
  assign add_53421 = {1'h0, umul_53225[21:7]} + 16'h007d;
  assign sel_53426 = $signed({1'h0, smod_53169[15:0]}) < $signed({1'h0, sel_53232}) ? smod_53169[15:0] : sel_53232;
  assign umul_53427 = umul22b_16b_x_6b(array_index_53365, 6'h35);
  assign add_53429 = {1'h0, umul_53233[21:7]} + 16'h007d;
  assign sel_53434 = $signed({1'h0, smod_53175[15:0]}) < $signed({1'h0, sel_53240}) ? smod_53175[15:0] : sel_53240;
  assign smod_53438 = $unsigned($signed({8'h00, add_53297, umul_53101[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53443 = $unsigned($signed({8'h00, add_53305, umul_53109[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53448 = $unsigned($signed({8'h00, add_53313, umul_53117[0]}) % $signed(32'h0000_3ffd));
  assign smod_53453 = $unsigned($signed({8'h00, add_53321, umul_53125[0]}) % $signed(32'h0000_3ffd));
  assign smod_53458 = $unsigned($signed({9'h000, add_53329, umul_53133[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53463 = $unsigned($signed({9'h000, add_53337, umul_53141[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53468 = $unsigned($signed({9'h000, add_53345, umul_53149[0]}) % $signed(32'h0000_3ffd));
  assign smod_53473 = $unsigned($signed({9'h000, add_53353, umul_53157[0]}) % $signed(32'h0000_3ffd));
  assign umul_53489 = umul23b_16b_x_7b(array_index_52783, 7'h49);
  assign add_53491 = {1'h0, umul_53295[22:3]} + 21'h00_07e9;
  assign sel_53496 = $signed({1'h0, smod_53244[15:0]}) < $signed({1'h0, sel_53302}) ? smod_53244[15:0] : sel_53302;
  assign umul_53497 = umul23b_16b_x_7b(array_index_52789, 7'h49);
  assign add_53499 = {1'h0, umul_53303[22:3]} + 21'h00_07e9;
  assign sel_53504 = $signed({1'h0, smod_53249[15:0]}) < $signed({1'h0, sel_53310}) ? smod_53249[15:0] : sel_53310;
  assign umul_53505 = umul23b_16b_x_7b(array_index_52969, 7'h47);
  assign add_53507 = {1'h0, umul_53311[22:1]} + 23'h00_1f8b;
  assign sel_53512 = $signed({1'h0, smod_53254[15:0]}) < $signed({1'h0, sel_53318}) ? smod_53254[15:0] : sel_53318;
  assign umul_53513 = umul23b_16b_x_7b(array_index_52975, 7'h47);
  assign add_53515 = {1'h0, umul_53319[22:1]} + 23'h00_1f8b;
  assign sel_53520 = $signed({1'h0, smod_53259[15:0]}) < $signed({1'h0, sel_53326}) ? smod_53259[15:0] : sel_53326;
  assign umul_53521 = umul22b_16b_x_6b(array_index_53165, 6'h3d);
  assign add_53523 = {1'h0, umul_53327[21:2]} + 21'h00_0fb9;
  assign sel_53528 = $signed({1'h0, smod_53264[15:0]}) < $signed({1'h0, sel_53334}) ? smod_53264[15:0] : sel_53334;
  assign umul_53529 = umul22b_16b_x_6b(array_index_53171, 6'h3d);
  assign add_53531 = {1'h0, umul_53335[21:2]} + 21'h00_0fb9;
  assign sel_53536 = $signed({1'h0, smod_53269[15:0]}) < $signed({1'h0, sel_53342}) ? smod_53269[15:0] : sel_53342;
  assign umul_53537 = umul22b_16b_x_6b(array_index_53359, 6'h3b);
  assign add_53539 = {1'h0, umul_53343[21:1]} + 22'h00_1f59;
  assign sel_53544 = $signed({1'h0, smod_53274[15:0]}) < $signed({1'h0, sel_53350}) ? smod_53274[15:0] : sel_53350;
  assign umul_53545 = umul22b_16b_x_6b(array_index_53365, 6'h3b);
  assign add_53547 = {1'h0, umul_53351[21:1]} + 22'h00_1f59;
  assign sel_53552 = $signed({1'h0, smod_53279[15:0]}) < $signed({1'h0, sel_53358}) ? smod_53279[15:0] : sel_53358;
  assign array_index_53553 = set1_unflattened[5'h09];
  assign smod_53557 = $unsigned($signed({9'h000, add_53421, umul_53225[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_53559 = set2_unflattened[5'h09];
  assign smod_53563 = $unsigned($signed({9'h000, add_53429, umul_53233[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_53613 = umul22b_16b_x_6b(array_index_53553, 6'h35);
  assign add_53615 = {1'h0, umul_53419[21:7]} + 16'h007d;
  assign sel_53620 = $signed({1'h0, smod_53363[15:0]}) < $signed({1'h0, sel_53426}) ? smod_53363[15:0] : sel_53426;
  assign umul_53621 = umul22b_16b_x_6b(array_index_53559, 6'h35);
  assign add_53623 = {1'h0, umul_53427[21:7]} + 16'h007d;
  assign sel_53628 = $signed({1'h0, smod_53369[15:0]}) < $signed({1'h0, sel_53434}) ? smod_53369[15:0] : sel_53434;
  assign smod_53632 = $unsigned($signed({8'h00, add_53491, umul_53295[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53637 = $unsigned($signed({8'h00, add_53499, umul_53303[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53642 = $unsigned($signed({8'h00, add_53507, umul_53311[0]}) % $signed(32'h0000_3ffd));
  assign smod_53647 = $unsigned($signed({8'h00, add_53515, umul_53319[0]}) % $signed(32'h0000_3ffd));
  assign smod_53652 = $unsigned($signed({9'h000, add_53523, umul_53327[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53657 = $unsigned($signed({9'h000, add_53531, umul_53335[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53662 = $unsigned($signed({9'h000, add_53539, umul_53343[0]}) % $signed(32'h0000_3ffd));
  assign smod_53667 = $unsigned($signed({9'h000, add_53547, umul_53351[0]}) % $signed(32'h0000_3ffd));
  assign umul_53683 = umul23b_16b_x_7b(array_index_52969, 7'h49);
  assign add_53685 = {1'h0, umul_53489[22:3]} + 21'h00_07e9;
  assign sel_53690 = $signed({1'h0, smod_53438[15:0]}) < $signed({1'h0, sel_53496}) ? smod_53438[15:0] : sel_53496;
  assign umul_53691 = umul23b_16b_x_7b(array_index_52975, 7'h49);
  assign add_53693 = {1'h0, umul_53497[22:3]} + 21'h00_07e9;
  assign sel_53698 = $signed({1'h0, smod_53443[15:0]}) < $signed({1'h0, sel_53504}) ? smod_53443[15:0] : sel_53504;
  assign umul_53699 = umul23b_16b_x_7b(array_index_53165, 7'h47);
  assign add_53701 = {1'h0, umul_53505[22:1]} + 23'h00_1f8b;
  assign sel_53706 = $signed({1'h0, smod_53448[15:0]}) < $signed({1'h0, sel_53512}) ? smod_53448[15:0] : sel_53512;
  assign umul_53707 = umul23b_16b_x_7b(array_index_53171, 7'h47);
  assign add_53709 = {1'h0, umul_53513[22:1]} + 23'h00_1f8b;
  assign sel_53714 = $signed({1'h0, smod_53453[15:0]}) < $signed({1'h0, sel_53520}) ? smod_53453[15:0] : sel_53520;
  assign umul_53715 = umul22b_16b_x_6b(array_index_53359, 6'h3d);
  assign add_53717 = {1'h0, umul_53521[21:2]} + 21'h00_0fb9;
  assign sel_53722 = $signed({1'h0, smod_53458[15:0]}) < $signed({1'h0, sel_53528}) ? smod_53458[15:0] : sel_53528;
  assign umul_53723 = umul22b_16b_x_6b(array_index_53365, 6'h3d);
  assign add_53725 = {1'h0, umul_53529[21:2]} + 21'h00_0fb9;
  assign sel_53730 = $signed({1'h0, smod_53463[15:0]}) < $signed({1'h0, sel_53536}) ? smod_53463[15:0] : sel_53536;
  assign umul_53731 = umul22b_16b_x_6b(array_index_53553, 6'h3b);
  assign add_53733 = {1'h0, umul_53537[21:1]} + 22'h00_1f59;
  assign sel_53738 = $signed({1'h0, smod_53468[15:0]}) < $signed({1'h0, sel_53544}) ? smod_53468[15:0] : sel_53544;
  assign umul_53739 = umul22b_16b_x_6b(array_index_53559, 6'h3b);
  assign add_53741 = {1'h0, umul_53545[21:1]} + 22'h00_1f59;
  assign sel_53746 = $signed({1'h0, smod_53473[15:0]}) < $signed({1'h0, sel_53552}) ? smod_53473[15:0] : sel_53552;
  assign array_index_53747 = set1_unflattened[5'h0a];
  assign smod_53751 = $unsigned($signed({9'h000, add_53615, umul_53419[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_53753 = set2_unflattened[5'h0a];
  assign smod_53757 = $unsigned($signed({9'h000, add_53623, umul_53427[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_53807 = umul22b_16b_x_6b(array_index_53747, 6'h35);
  assign add_53809 = {1'h0, umul_53613[21:7]} + 16'h007d;
  assign sel_53814 = $signed({1'h0, smod_53557[15:0]}) < $signed({1'h0, sel_53620}) ? smod_53557[15:0] : sel_53620;
  assign umul_53815 = umul22b_16b_x_6b(array_index_53753, 6'h35);
  assign add_53817 = {1'h0, umul_53621[21:7]} + 16'h007d;
  assign sel_53822 = $signed({1'h0, smod_53563[15:0]}) < $signed({1'h0, sel_53628}) ? smod_53563[15:0] : sel_53628;
  assign smod_53826 = $unsigned($signed({8'h00, add_53685, umul_53489[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53831 = $unsigned($signed({8'h00, add_53693, umul_53497[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_53836 = $unsigned($signed({8'h00, add_53701, umul_53505[0]}) % $signed(32'h0000_3ffd));
  assign smod_53841 = $unsigned($signed({8'h00, add_53709, umul_53513[0]}) % $signed(32'h0000_3ffd));
  assign smod_53846 = $unsigned($signed({9'h000, add_53717, umul_53521[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53851 = $unsigned($signed({9'h000, add_53725, umul_53529[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_53856 = $unsigned($signed({9'h000, add_53733, umul_53537[0]}) % $signed(32'h0000_3ffd));
  assign smod_53861 = $unsigned($signed({9'h000, add_53741, umul_53545[0]}) % $signed(32'h0000_3ffd));
  assign umul_53877 = umul23b_16b_x_7b(array_index_53165, 7'h49);
  assign add_53879 = {1'h0, umul_53683[22:3]} + 21'h00_07e9;
  assign sel_53884 = $signed({1'h0, smod_53632[15:0]}) < $signed({1'h0, sel_53690}) ? smod_53632[15:0] : sel_53690;
  assign umul_53885 = umul23b_16b_x_7b(array_index_53171, 7'h49);
  assign add_53887 = {1'h0, umul_53691[22:3]} + 21'h00_07e9;
  assign sel_53892 = $signed({1'h0, smod_53637[15:0]}) < $signed({1'h0, sel_53698}) ? smod_53637[15:0] : sel_53698;
  assign umul_53893 = umul23b_16b_x_7b(array_index_53359, 7'h47);
  assign add_53895 = {1'h0, umul_53699[22:1]} + 23'h00_1f8b;
  assign sel_53900 = $signed({1'h0, smod_53642[15:0]}) < $signed({1'h0, sel_53706}) ? smod_53642[15:0] : sel_53706;
  assign umul_53901 = umul23b_16b_x_7b(array_index_53365, 7'h47);
  assign add_53903 = {1'h0, umul_53707[22:1]} + 23'h00_1f8b;
  assign sel_53908 = $signed({1'h0, smod_53647[15:0]}) < $signed({1'h0, sel_53714}) ? smod_53647[15:0] : sel_53714;
  assign umul_53909 = umul22b_16b_x_6b(array_index_53553, 6'h3d);
  assign add_53911 = {1'h0, umul_53715[21:2]} + 21'h00_0fb9;
  assign sel_53916 = $signed({1'h0, smod_53652[15:0]}) < $signed({1'h0, sel_53722}) ? smod_53652[15:0] : sel_53722;
  assign umul_53917 = umul22b_16b_x_6b(array_index_53559, 6'h3d);
  assign add_53919 = {1'h0, umul_53723[21:2]} + 21'h00_0fb9;
  assign sel_53924 = $signed({1'h0, smod_53657[15:0]}) < $signed({1'h0, sel_53730}) ? smod_53657[15:0] : sel_53730;
  assign umul_53925 = umul22b_16b_x_6b(array_index_53747, 6'h3b);
  assign add_53927 = {1'h0, umul_53731[21:1]} + 22'h00_1f59;
  assign sel_53932 = $signed({1'h0, smod_53662[15:0]}) < $signed({1'h0, sel_53738}) ? smod_53662[15:0] : sel_53738;
  assign umul_53933 = umul22b_16b_x_6b(array_index_53753, 6'h3b);
  assign add_53935 = {1'h0, umul_53739[21:1]} + 22'h00_1f59;
  assign sel_53940 = $signed({1'h0, smod_53667[15:0]}) < $signed({1'h0, sel_53746}) ? smod_53667[15:0] : sel_53746;
  assign array_index_53941 = set1_unflattened[5'h0b];
  assign smod_53945 = $unsigned($signed({9'h000, add_53809, umul_53613[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_53947 = set2_unflattened[5'h0b];
  assign smod_53951 = $unsigned($signed({9'h000, add_53817, umul_53621[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_54001 = umul22b_16b_x_6b(array_index_53941, 6'h35);
  assign add_54003 = {1'h0, umul_53807[21:7]} + 16'h007d;
  assign sel_54008 = $signed({1'h0, smod_53751[15:0]}) < $signed({1'h0, sel_53814}) ? smod_53751[15:0] : sel_53814;
  assign umul_54009 = umul22b_16b_x_6b(array_index_53947, 6'h35);
  assign add_54011 = {1'h0, umul_53815[21:7]} + 16'h007d;
  assign sel_54016 = $signed({1'h0, smod_53757[15:0]}) < $signed({1'h0, sel_53822}) ? smod_53757[15:0] : sel_53822;
  assign smod_54020 = $unsigned($signed({8'h00, add_53879, umul_53683[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54025 = $unsigned($signed({8'h00, add_53887, umul_53691[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54030 = $unsigned($signed({8'h00, add_53895, umul_53699[0]}) % $signed(32'h0000_3ffd));
  assign smod_54035 = $unsigned($signed({8'h00, add_53903, umul_53707[0]}) % $signed(32'h0000_3ffd));
  assign smod_54040 = $unsigned($signed({9'h000, add_53911, umul_53715[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54045 = $unsigned($signed({9'h000, add_53919, umul_53723[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54050 = $unsigned($signed({9'h000, add_53927, umul_53731[0]}) % $signed(32'h0000_3ffd));
  assign smod_54055 = $unsigned($signed({9'h000, add_53935, umul_53739[0]}) % $signed(32'h0000_3ffd));
  assign umul_54071 = umul23b_16b_x_7b(array_index_53359, 7'h49);
  assign add_54073 = {1'h0, umul_53877[22:3]} + 21'h00_07e9;
  assign sel_54078 = $signed({1'h0, smod_53826[15:0]}) < $signed({1'h0, sel_53884}) ? smod_53826[15:0] : sel_53884;
  assign umul_54079 = umul23b_16b_x_7b(array_index_53365, 7'h49);
  assign add_54081 = {1'h0, umul_53885[22:3]} + 21'h00_07e9;
  assign sel_54086 = $signed({1'h0, smod_53831[15:0]}) < $signed({1'h0, sel_53892}) ? smod_53831[15:0] : sel_53892;
  assign umul_54087 = umul23b_16b_x_7b(array_index_53553, 7'h47);
  assign add_54089 = {1'h0, umul_53893[22:1]} + 23'h00_1f8b;
  assign sel_54094 = $signed({1'h0, smod_53836[15:0]}) < $signed({1'h0, sel_53900}) ? smod_53836[15:0] : sel_53900;
  assign umul_54095 = umul23b_16b_x_7b(array_index_53559, 7'h47);
  assign add_54097 = {1'h0, umul_53901[22:1]} + 23'h00_1f8b;
  assign sel_54102 = $signed({1'h0, smod_53841[15:0]}) < $signed({1'h0, sel_53908}) ? smod_53841[15:0] : sel_53908;
  assign umul_54103 = umul22b_16b_x_6b(array_index_53747, 6'h3d);
  assign add_54105 = {1'h0, umul_53909[21:2]} + 21'h00_0fb9;
  assign sel_54110 = $signed({1'h0, smod_53846[15:0]}) < $signed({1'h0, sel_53916}) ? smod_53846[15:0] : sel_53916;
  assign umul_54111 = umul22b_16b_x_6b(array_index_53753, 6'h3d);
  assign add_54113 = {1'h0, umul_53917[21:2]} + 21'h00_0fb9;
  assign sel_54118 = $signed({1'h0, smod_53851[15:0]}) < $signed({1'h0, sel_53924}) ? smod_53851[15:0] : sel_53924;
  assign umul_54119 = umul22b_16b_x_6b(array_index_53941, 6'h3b);
  assign add_54121 = {1'h0, umul_53925[21:1]} + 22'h00_1f59;
  assign sel_54126 = $signed({1'h0, smod_53856[15:0]}) < $signed({1'h0, sel_53932}) ? smod_53856[15:0] : sel_53932;
  assign umul_54127 = umul22b_16b_x_6b(array_index_53947, 6'h3b);
  assign add_54129 = {1'h0, umul_53933[21:1]} + 22'h00_1f59;
  assign sel_54134 = $signed({1'h0, smod_53861[15:0]}) < $signed({1'h0, sel_53940}) ? smod_53861[15:0] : sel_53940;
  assign array_index_54135 = set1_unflattened[5'h0c];
  assign smod_54139 = $unsigned($signed({9'h000, add_54003, umul_53807[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_54141 = set2_unflattened[5'h0c];
  assign smod_54145 = $unsigned($signed({9'h000, add_54011, umul_53815[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_54195 = umul22b_16b_x_6b(array_index_54135, 6'h35);
  assign add_54197 = {1'h0, umul_54001[21:7]} + 16'h007d;
  assign sel_54202 = $signed({1'h0, smod_53945[15:0]}) < $signed({1'h0, sel_54008}) ? smod_53945[15:0] : sel_54008;
  assign umul_54203 = umul22b_16b_x_6b(array_index_54141, 6'h35);
  assign add_54205 = {1'h0, umul_54009[21:7]} + 16'h007d;
  assign sel_54210 = $signed({1'h0, smod_53951[15:0]}) < $signed({1'h0, sel_54016}) ? smod_53951[15:0] : sel_54016;
  assign smod_54214 = $unsigned($signed({8'h00, add_54073, umul_53877[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54219 = $unsigned($signed({8'h00, add_54081, umul_53885[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54224 = $unsigned($signed({8'h00, add_54089, umul_53893[0]}) % $signed(32'h0000_3ffd));
  assign smod_54229 = $unsigned($signed({8'h00, add_54097, umul_53901[0]}) % $signed(32'h0000_3ffd));
  assign smod_54234 = $unsigned($signed({9'h000, add_54105, umul_53909[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54239 = $unsigned($signed({9'h000, add_54113, umul_53917[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54244 = $unsigned($signed({9'h000, add_54121, umul_53925[0]}) % $signed(32'h0000_3ffd));
  assign smod_54249 = $unsigned($signed({9'h000, add_54129, umul_53933[0]}) % $signed(32'h0000_3ffd));
  assign umul_54265 = umul23b_16b_x_7b(array_index_53553, 7'h49);
  assign add_54267 = {1'h0, umul_54071[22:3]} + 21'h00_07e9;
  assign sel_54272 = $signed({1'h0, smod_54020[15:0]}) < $signed({1'h0, sel_54078}) ? smod_54020[15:0] : sel_54078;
  assign umul_54273 = umul23b_16b_x_7b(array_index_53559, 7'h49);
  assign add_54275 = {1'h0, umul_54079[22:3]} + 21'h00_07e9;
  assign sel_54280 = $signed({1'h0, smod_54025[15:0]}) < $signed({1'h0, sel_54086}) ? smod_54025[15:0] : sel_54086;
  assign umul_54281 = umul23b_16b_x_7b(array_index_53747, 7'h47);
  assign add_54283 = {1'h0, umul_54087[22:1]} + 23'h00_1f8b;
  assign sel_54288 = $signed({1'h0, smod_54030[15:0]}) < $signed({1'h0, sel_54094}) ? smod_54030[15:0] : sel_54094;
  assign umul_54289 = umul23b_16b_x_7b(array_index_53753, 7'h47);
  assign add_54291 = {1'h0, umul_54095[22:1]} + 23'h00_1f8b;
  assign sel_54296 = $signed({1'h0, smod_54035[15:0]}) < $signed({1'h0, sel_54102}) ? smod_54035[15:0] : sel_54102;
  assign umul_54297 = umul22b_16b_x_6b(array_index_53941, 6'h3d);
  assign add_54299 = {1'h0, umul_54103[21:2]} + 21'h00_0fb9;
  assign sel_54304 = $signed({1'h0, smod_54040[15:0]}) < $signed({1'h0, sel_54110}) ? smod_54040[15:0] : sel_54110;
  assign umul_54305 = umul22b_16b_x_6b(array_index_53947, 6'h3d);
  assign add_54307 = {1'h0, umul_54111[21:2]} + 21'h00_0fb9;
  assign sel_54312 = $signed({1'h0, smod_54045[15:0]}) < $signed({1'h0, sel_54118}) ? smod_54045[15:0] : sel_54118;
  assign umul_54313 = umul22b_16b_x_6b(array_index_54135, 6'h3b);
  assign add_54315 = {1'h0, umul_54119[21:1]} + 22'h00_1f59;
  assign sel_54320 = $signed({1'h0, smod_54050[15:0]}) < $signed({1'h0, sel_54126}) ? smod_54050[15:0] : sel_54126;
  assign umul_54321 = umul22b_16b_x_6b(array_index_54141, 6'h3b);
  assign add_54323 = {1'h0, umul_54127[21:1]} + 22'h00_1f59;
  assign sel_54328 = $signed({1'h0, smod_54055[15:0]}) < $signed({1'h0, sel_54134}) ? smod_54055[15:0] : sel_54134;
  assign array_index_54329 = set1_unflattened[5'h0d];
  assign smod_54333 = $unsigned($signed({9'h000, add_54197, umul_54001[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_54335 = set2_unflattened[5'h0d];
  assign smod_54339 = $unsigned($signed({9'h000, add_54205, umul_54009[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_54389 = umul22b_16b_x_6b(array_index_54329, 6'h35);
  assign add_54391 = {1'h0, umul_54195[21:7]} + 16'h007d;
  assign sel_54396 = $signed({1'h0, smod_54139[15:0]}) < $signed({1'h0, sel_54202}) ? smod_54139[15:0] : sel_54202;
  assign umul_54397 = umul22b_16b_x_6b(array_index_54335, 6'h35);
  assign add_54399 = {1'h0, umul_54203[21:7]} + 16'h007d;
  assign sel_54404 = $signed({1'h0, smod_54145[15:0]}) < $signed({1'h0, sel_54210}) ? smod_54145[15:0] : sel_54210;
  assign smod_54408 = $unsigned($signed({8'h00, add_54267, umul_54071[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54413 = $unsigned($signed({8'h00, add_54275, umul_54079[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54418 = $unsigned($signed({8'h00, add_54283, umul_54087[0]}) % $signed(32'h0000_3ffd));
  assign smod_54423 = $unsigned($signed({8'h00, add_54291, umul_54095[0]}) % $signed(32'h0000_3ffd));
  assign smod_54428 = $unsigned($signed({9'h000, add_54299, umul_54103[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54433 = $unsigned($signed({9'h000, add_54307, umul_54111[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54438 = $unsigned($signed({9'h000, add_54315, umul_54119[0]}) % $signed(32'h0000_3ffd));
  assign smod_54443 = $unsigned($signed({9'h000, add_54323, umul_54127[0]}) % $signed(32'h0000_3ffd));
  assign umul_54459 = umul23b_16b_x_7b(array_index_53747, 7'h49);
  assign add_54461 = {1'h0, umul_54265[22:3]} + 21'h00_07e9;
  assign sel_54466 = $signed({1'h0, smod_54214[15:0]}) < $signed({1'h0, sel_54272}) ? smod_54214[15:0] : sel_54272;
  assign umul_54467 = umul23b_16b_x_7b(array_index_53753, 7'h49);
  assign add_54469 = {1'h0, umul_54273[22:3]} + 21'h00_07e9;
  assign sel_54474 = $signed({1'h0, smod_54219[15:0]}) < $signed({1'h0, sel_54280}) ? smod_54219[15:0] : sel_54280;
  assign umul_54475 = umul23b_16b_x_7b(array_index_53941, 7'h47);
  assign add_54477 = {1'h0, umul_54281[22:1]} + 23'h00_1f8b;
  assign sel_54482 = $signed({1'h0, smod_54224[15:0]}) < $signed({1'h0, sel_54288}) ? smod_54224[15:0] : sel_54288;
  assign umul_54483 = umul23b_16b_x_7b(array_index_53947, 7'h47);
  assign add_54485 = {1'h0, umul_54289[22:1]} + 23'h00_1f8b;
  assign sel_54490 = $signed({1'h0, smod_54229[15:0]}) < $signed({1'h0, sel_54296}) ? smod_54229[15:0] : sel_54296;
  assign umul_54491 = umul22b_16b_x_6b(array_index_54135, 6'h3d);
  assign add_54493 = {1'h0, umul_54297[21:2]} + 21'h00_0fb9;
  assign sel_54498 = $signed({1'h0, smod_54234[15:0]}) < $signed({1'h0, sel_54304}) ? smod_54234[15:0] : sel_54304;
  assign umul_54499 = umul22b_16b_x_6b(array_index_54141, 6'h3d);
  assign add_54501 = {1'h0, umul_54305[21:2]} + 21'h00_0fb9;
  assign sel_54506 = $signed({1'h0, smod_54239[15:0]}) < $signed({1'h0, sel_54312}) ? smod_54239[15:0] : sel_54312;
  assign umul_54507 = umul22b_16b_x_6b(array_index_54329, 6'h3b);
  assign add_54509 = {1'h0, umul_54313[21:1]} + 22'h00_1f59;
  assign sel_54514 = $signed({1'h0, smod_54244[15:0]}) < $signed({1'h0, sel_54320}) ? smod_54244[15:0] : sel_54320;
  assign umul_54515 = umul22b_16b_x_6b(array_index_54335, 6'h3b);
  assign add_54517 = {1'h0, umul_54321[21:1]} + 22'h00_1f59;
  assign sel_54522 = $signed({1'h0, smod_54249[15:0]}) < $signed({1'h0, sel_54328}) ? smod_54249[15:0] : sel_54328;
  assign array_index_54523 = set1_unflattened[5'h0e];
  assign smod_54527 = $unsigned($signed({9'h000, add_54391, umul_54195[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_54529 = set2_unflattened[5'h0e];
  assign smod_54533 = $unsigned($signed({9'h000, add_54399, umul_54203[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_54583 = umul22b_16b_x_6b(array_index_54523, 6'h35);
  assign add_54585 = {1'h0, umul_54389[21:7]} + 16'h007d;
  assign sel_54590 = $signed({1'h0, smod_54333[15:0]}) < $signed({1'h0, sel_54396}) ? smod_54333[15:0] : sel_54396;
  assign umul_54591 = umul22b_16b_x_6b(array_index_54529, 6'h35);
  assign add_54593 = {1'h0, umul_54397[21:7]} + 16'h007d;
  assign sel_54598 = $signed({1'h0, smod_54339[15:0]}) < $signed({1'h0, sel_54404}) ? smod_54339[15:0] : sel_54404;
  assign smod_54602 = $unsigned($signed({8'h00, add_54461, umul_54265[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54607 = $unsigned($signed({8'h00, add_54469, umul_54273[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54612 = $unsigned($signed({8'h00, add_54477, umul_54281[0]}) % $signed(32'h0000_3ffd));
  assign smod_54617 = $unsigned($signed({8'h00, add_54485, umul_54289[0]}) % $signed(32'h0000_3ffd));
  assign smod_54622 = $unsigned($signed({9'h000, add_54493, umul_54297[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54627 = $unsigned($signed({9'h000, add_54501, umul_54305[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54632 = $unsigned($signed({9'h000, add_54509, umul_54313[0]}) % $signed(32'h0000_3ffd));
  assign smod_54637 = $unsigned($signed({9'h000, add_54517, umul_54321[0]}) % $signed(32'h0000_3ffd));
  assign umul_54653 = umul23b_16b_x_7b(array_index_53941, 7'h49);
  assign add_54655 = {1'h0, umul_54459[22:3]} + 21'h00_07e9;
  assign sel_54660 = $signed({1'h0, smod_54408[15:0]}) < $signed({1'h0, sel_54466}) ? smod_54408[15:0] : sel_54466;
  assign umul_54661 = umul23b_16b_x_7b(array_index_53947, 7'h49);
  assign add_54663 = {1'h0, umul_54467[22:3]} + 21'h00_07e9;
  assign sel_54668 = $signed({1'h0, smod_54413[15:0]}) < $signed({1'h0, sel_54474}) ? smod_54413[15:0] : sel_54474;
  assign umul_54669 = umul23b_16b_x_7b(array_index_54135, 7'h47);
  assign add_54671 = {1'h0, umul_54475[22:1]} + 23'h00_1f8b;
  assign sel_54676 = $signed({1'h0, smod_54418[15:0]}) < $signed({1'h0, sel_54482}) ? smod_54418[15:0] : sel_54482;
  assign umul_54677 = umul23b_16b_x_7b(array_index_54141, 7'h47);
  assign add_54679 = {1'h0, umul_54483[22:1]} + 23'h00_1f8b;
  assign sel_54684 = $signed({1'h0, smod_54423[15:0]}) < $signed({1'h0, sel_54490}) ? smod_54423[15:0] : sel_54490;
  assign umul_54685 = umul22b_16b_x_6b(array_index_54329, 6'h3d);
  assign add_54687 = {1'h0, umul_54491[21:2]} + 21'h00_0fb9;
  assign sel_54692 = $signed({1'h0, smod_54428[15:0]}) < $signed({1'h0, sel_54498}) ? smod_54428[15:0] : sel_54498;
  assign umul_54693 = umul22b_16b_x_6b(array_index_54335, 6'h3d);
  assign add_54695 = {1'h0, umul_54499[21:2]} + 21'h00_0fb9;
  assign sel_54700 = $signed({1'h0, smod_54433[15:0]}) < $signed({1'h0, sel_54506}) ? smod_54433[15:0] : sel_54506;
  assign umul_54701 = umul22b_16b_x_6b(array_index_54523, 6'h3b);
  assign add_54703 = {1'h0, umul_54507[21:1]} + 22'h00_1f59;
  assign sel_54708 = $signed({1'h0, smod_54438[15:0]}) < $signed({1'h0, sel_54514}) ? smod_54438[15:0] : sel_54514;
  assign umul_54709 = umul22b_16b_x_6b(array_index_54529, 6'h3b);
  assign add_54711 = {1'h0, umul_54515[21:1]} + 22'h00_1f59;
  assign sel_54716 = $signed({1'h0, smod_54443[15:0]}) < $signed({1'h0, sel_54522}) ? smod_54443[15:0] : sel_54522;
  assign array_index_54717 = set1_unflattened[5'h0f];
  assign smod_54721 = $unsigned($signed({9'h000, add_54585, umul_54389[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_54723 = set2_unflattened[5'h0f];
  assign smod_54727 = $unsigned($signed({9'h000, add_54593, umul_54397[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_54777 = umul22b_16b_x_6b(array_index_54717, 6'h35);
  assign add_54779 = {1'h0, umul_54583[21:7]} + 16'h007d;
  assign sel_54784 = $signed({1'h0, smod_54527[15:0]}) < $signed({1'h0, sel_54590}) ? smod_54527[15:0] : sel_54590;
  assign umul_54785 = umul22b_16b_x_6b(array_index_54723, 6'h35);
  assign add_54787 = {1'h0, umul_54591[21:7]} + 16'h007d;
  assign sel_54792 = $signed({1'h0, smod_54533[15:0]}) < $signed({1'h0, sel_54598}) ? smod_54533[15:0] : sel_54598;
  assign smod_54796 = $unsigned($signed({8'h00, add_54655, umul_54459[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54801 = $unsigned($signed({8'h00, add_54663, umul_54467[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54806 = $unsigned($signed({8'h00, add_54671, umul_54475[0]}) % $signed(32'h0000_3ffd));
  assign smod_54811 = $unsigned($signed({8'h00, add_54679, umul_54483[0]}) % $signed(32'h0000_3ffd));
  assign smod_54816 = $unsigned($signed({9'h000, add_54687, umul_54491[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54821 = $unsigned($signed({9'h000, add_54695, umul_54499[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_54826 = $unsigned($signed({9'h000, add_54703, umul_54507[0]}) % $signed(32'h0000_3ffd));
  assign smod_54831 = $unsigned($signed({9'h000, add_54711, umul_54515[0]}) % $signed(32'h0000_3ffd));
  assign umul_54847 = umul23b_16b_x_7b(array_index_54135, 7'h49);
  assign add_54849 = {1'h0, umul_54653[22:3]} + 21'h00_07e9;
  assign sel_54854 = $signed({1'h0, smod_54602[15:0]}) < $signed({1'h0, sel_54660}) ? smod_54602[15:0] : sel_54660;
  assign umul_54855 = umul23b_16b_x_7b(array_index_54141, 7'h49);
  assign add_54857 = {1'h0, umul_54661[22:3]} + 21'h00_07e9;
  assign sel_54862 = $signed({1'h0, smod_54607[15:0]}) < $signed({1'h0, sel_54668}) ? smod_54607[15:0] : sel_54668;
  assign umul_54863 = umul23b_16b_x_7b(array_index_54329, 7'h47);
  assign add_54865 = {1'h0, umul_54669[22:1]} + 23'h00_1f8b;
  assign sel_54870 = $signed({1'h0, smod_54612[15:0]}) < $signed({1'h0, sel_54676}) ? smod_54612[15:0] : sel_54676;
  assign umul_54871 = umul23b_16b_x_7b(array_index_54335, 7'h47);
  assign add_54873 = {1'h0, umul_54677[22:1]} + 23'h00_1f8b;
  assign sel_54878 = $signed({1'h0, smod_54617[15:0]}) < $signed({1'h0, sel_54684}) ? smod_54617[15:0] : sel_54684;
  assign umul_54879 = umul22b_16b_x_6b(array_index_54523, 6'h3d);
  assign add_54881 = {1'h0, umul_54685[21:2]} + 21'h00_0fb9;
  assign sel_54886 = $signed({1'h0, smod_54622[15:0]}) < $signed({1'h0, sel_54692}) ? smod_54622[15:0] : sel_54692;
  assign umul_54887 = umul22b_16b_x_6b(array_index_54529, 6'h3d);
  assign add_54889 = {1'h0, umul_54693[21:2]} + 21'h00_0fb9;
  assign sel_54894 = $signed({1'h0, smod_54627[15:0]}) < $signed({1'h0, sel_54700}) ? smod_54627[15:0] : sel_54700;
  assign umul_54895 = umul22b_16b_x_6b(array_index_54717, 6'h3b);
  assign add_54897 = {1'h0, umul_54701[21:1]} + 22'h00_1f59;
  assign sel_54902 = $signed({1'h0, smod_54632[15:0]}) < $signed({1'h0, sel_54708}) ? smod_54632[15:0] : sel_54708;
  assign umul_54903 = umul22b_16b_x_6b(array_index_54723, 6'h3b);
  assign add_54905 = {1'h0, umul_54709[21:1]} + 22'h00_1f59;
  assign sel_54910 = $signed({1'h0, smod_54637[15:0]}) < $signed({1'h0, sel_54716}) ? smod_54637[15:0] : sel_54716;
  assign array_index_54911 = set1_unflattened[5'h10];
  assign smod_54915 = $unsigned($signed({9'h000, add_54779, umul_54583[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_54917 = set2_unflattened[5'h10];
  assign smod_54921 = $unsigned($signed({9'h000, add_54787, umul_54591[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_54971 = umul22b_16b_x_6b(array_index_54911, 6'h35);
  assign add_54973 = {1'h0, umul_54777[21:7]} + 16'h007d;
  assign sel_54978 = $signed({1'h0, smod_54721[15:0]}) < $signed({1'h0, sel_54784}) ? smod_54721[15:0] : sel_54784;
  assign umul_54979 = umul22b_16b_x_6b(array_index_54917, 6'h35);
  assign add_54981 = {1'h0, umul_54785[21:7]} + 16'h007d;
  assign sel_54986 = $signed({1'h0, smod_54727[15:0]}) < $signed({1'h0, sel_54792}) ? smod_54727[15:0] : sel_54792;
  assign smod_54990 = $unsigned($signed({8'h00, add_54849, umul_54653[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_54995 = $unsigned($signed({8'h00, add_54857, umul_54661[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55000 = $unsigned($signed({8'h00, add_54865, umul_54669[0]}) % $signed(32'h0000_3ffd));
  assign smod_55005 = $unsigned($signed({8'h00, add_54873, umul_54677[0]}) % $signed(32'h0000_3ffd));
  assign smod_55010 = $unsigned($signed({9'h000, add_54881, umul_54685[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55015 = $unsigned($signed({9'h000, add_54889, umul_54693[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55020 = $unsigned($signed({9'h000, add_54897, umul_54701[0]}) % $signed(32'h0000_3ffd));
  assign smod_55025 = $unsigned($signed({9'h000, add_54905, umul_54709[0]}) % $signed(32'h0000_3ffd));
  assign umul_55041 = umul23b_16b_x_7b(array_index_54329, 7'h49);
  assign add_55043 = {1'h0, umul_54847[22:3]} + 21'h00_07e9;
  assign sel_55048 = $signed({1'h0, smod_54796[15:0]}) < $signed({1'h0, sel_54854}) ? smod_54796[15:0] : sel_54854;
  assign umul_55049 = umul23b_16b_x_7b(array_index_54335, 7'h49);
  assign add_55051 = {1'h0, umul_54855[22:3]} + 21'h00_07e9;
  assign sel_55056 = $signed({1'h0, smod_54801[15:0]}) < $signed({1'h0, sel_54862}) ? smod_54801[15:0] : sel_54862;
  assign umul_55057 = umul23b_16b_x_7b(array_index_54523, 7'h47);
  assign add_55059 = {1'h0, umul_54863[22:1]} + 23'h00_1f8b;
  assign sel_55064 = $signed({1'h0, smod_54806[15:0]}) < $signed({1'h0, sel_54870}) ? smod_54806[15:0] : sel_54870;
  assign umul_55065 = umul23b_16b_x_7b(array_index_54529, 7'h47);
  assign add_55067 = {1'h0, umul_54871[22:1]} + 23'h00_1f8b;
  assign sel_55072 = $signed({1'h0, smod_54811[15:0]}) < $signed({1'h0, sel_54878}) ? smod_54811[15:0] : sel_54878;
  assign umul_55073 = umul22b_16b_x_6b(array_index_54717, 6'h3d);
  assign add_55075 = {1'h0, umul_54879[21:2]} + 21'h00_0fb9;
  assign sel_55080 = $signed({1'h0, smod_54816[15:0]}) < $signed({1'h0, sel_54886}) ? smod_54816[15:0] : sel_54886;
  assign umul_55081 = umul22b_16b_x_6b(array_index_54723, 6'h3d);
  assign add_55083 = {1'h0, umul_54887[21:2]} + 21'h00_0fb9;
  assign sel_55088 = $signed({1'h0, smod_54821[15:0]}) < $signed({1'h0, sel_54894}) ? smod_54821[15:0] : sel_54894;
  assign umul_55089 = umul22b_16b_x_6b(array_index_54911, 6'h3b);
  assign add_55091 = {1'h0, umul_54895[21:1]} + 22'h00_1f59;
  assign sel_55096 = $signed({1'h0, smod_54826[15:0]}) < $signed({1'h0, sel_54902}) ? smod_54826[15:0] : sel_54902;
  assign umul_55097 = umul22b_16b_x_6b(array_index_54917, 6'h3b);
  assign add_55099 = {1'h0, umul_54903[21:1]} + 22'h00_1f59;
  assign sel_55104 = $signed({1'h0, smod_54831[15:0]}) < $signed({1'h0, sel_54910}) ? smod_54831[15:0] : sel_54910;
  assign array_index_55105 = set1_unflattened[5'h11];
  assign smod_55109 = $unsigned($signed({9'h000, add_54973, umul_54777[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_55111 = set2_unflattened[5'h11];
  assign smod_55115 = $unsigned($signed({9'h000, add_54981, umul_54785[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_55165 = umul22b_16b_x_6b(array_index_55105, 6'h35);
  assign add_55167 = {1'h0, umul_54971[21:7]} + 16'h007d;
  assign sel_55172 = $signed({1'h0, smod_54915[15:0]}) < $signed({1'h0, sel_54978}) ? smod_54915[15:0] : sel_54978;
  assign umul_55173 = umul22b_16b_x_6b(array_index_55111, 6'h35);
  assign add_55175 = {1'h0, umul_54979[21:7]} + 16'h007d;
  assign sel_55180 = $signed({1'h0, smod_54921[15:0]}) < $signed({1'h0, sel_54986}) ? smod_54921[15:0] : sel_54986;
  assign smod_55184 = $unsigned($signed({8'h00, add_55043, umul_54847[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55189 = $unsigned($signed({8'h00, add_55051, umul_54855[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55194 = $unsigned($signed({8'h00, add_55059, umul_54863[0]}) % $signed(32'h0000_3ffd));
  assign smod_55199 = $unsigned($signed({8'h00, add_55067, umul_54871[0]}) % $signed(32'h0000_3ffd));
  assign smod_55204 = $unsigned($signed({9'h000, add_55075, umul_54879[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55209 = $unsigned($signed({9'h000, add_55083, umul_54887[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55214 = $unsigned($signed({9'h000, add_55091, umul_54895[0]}) % $signed(32'h0000_3ffd));
  assign smod_55219 = $unsigned($signed({9'h000, add_55099, umul_54903[0]}) % $signed(32'h0000_3ffd));
  assign umul_55235 = umul23b_16b_x_7b(array_index_54523, 7'h49);
  assign add_55237 = {1'h0, umul_55041[22:3]} + 21'h00_07e9;
  assign sel_55242 = $signed({1'h0, smod_54990[15:0]}) < $signed({1'h0, sel_55048}) ? smod_54990[15:0] : sel_55048;
  assign umul_55243 = umul23b_16b_x_7b(array_index_54529, 7'h49);
  assign add_55245 = {1'h0, umul_55049[22:3]} + 21'h00_07e9;
  assign sel_55250 = $signed({1'h0, smod_54995[15:0]}) < $signed({1'h0, sel_55056}) ? smod_54995[15:0] : sel_55056;
  assign umul_55251 = umul23b_16b_x_7b(array_index_54717, 7'h47);
  assign add_55253 = {1'h0, umul_55057[22:1]} + 23'h00_1f8b;
  assign sel_55258 = $signed({1'h0, smod_55000[15:0]}) < $signed({1'h0, sel_55064}) ? smod_55000[15:0] : sel_55064;
  assign umul_55259 = umul23b_16b_x_7b(array_index_54723, 7'h47);
  assign add_55261 = {1'h0, umul_55065[22:1]} + 23'h00_1f8b;
  assign sel_55266 = $signed({1'h0, smod_55005[15:0]}) < $signed({1'h0, sel_55072}) ? smod_55005[15:0] : sel_55072;
  assign umul_55267 = umul22b_16b_x_6b(array_index_54911, 6'h3d);
  assign add_55269 = {1'h0, umul_55073[21:2]} + 21'h00_0fb9;
  assign sel_55274 = $signed({1'h0, smod_55010[15:0]}) < $signed({1'h0, sel_55080}) ? smod_55010[15:0] : sel_55080;
  assign umul_55275 = umul22b_16b_x_6b(array_index_54917, 6'h3d);
  assign add_55277 = {1'h0, umul_55081[21:2]} + 21'h00_0fb9;
  assign sel_55282 = $signed({1'h0, smod_55015[15:0]}) < $signed({1'h0, sel_55088}) ? smod_55015[15:0] : sel_55088;
  assign umul_55283 = umul22b_16b_x_6b(array_index_55105, 6'h3b);
  assign add_55285 = {1'h0, umul_55089[21:1]} + 22'h00_1f59;
  assign sel_55290 = $signed({1'h0, smod_55020[15:0]}) < $signed({1'h0, sel_55096}) ? smod_55020[15:0] : sel_55096;
  assign umul_55291 = umul22b_16b_x_6b(array_index_55111, 6'h3b);
  assign add_55293 = {1'h0, umul_55097[21:1]} + 22'h00_1f59;
  assign sel_55298 = $signed({1'h0, smod_55025[15:0]}) < $signed({1'h0, sel_55104}) ? smod_55025[15:0] : sel_55104;
  assign array_index_55299 = set1_unflattened[5'h12];
  assign smod_55303 = $unsigned($signed({9'h000, add_55167, umul_54971[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_55305 = set2_unflattened[5'h12];
  assign smod_55309 = $unsigned($signed({9'h000, add_55175, umul_54979[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_55359 = umul22b_16b_x_6b(array_index_55299, 6'h35);
  assign add_55361 = {1'h0, umul_55165[21:7]} + 16'h007d;
  assign sel_55366 = $signed({1'h0, smod_55109[15:0]}) < $signed({1'h0, sel_55172}) ? smod_55109[15:0] : sel_55172;
  assign umul_55367 = umul22b_16b_x_6b(array_index_55305, 6'h35);
  assign add_55369 = {1'h0, umul_55173[21:7]} + 16'h007d;
  assign sel_55374 = $signed({1'h0, smod_55115[15:0]}) < $signed({1'h0, sel_55180}) ? smod_55115[15:0] : sel_55180;
  assign smod_55378 = $unsigned($signed({8'h00, add_55237, umul_55041[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55383 = $unsigned($signed({8'h00, add_55245, umul_55049[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55388 = $unsigned($signed({8'h00, add_55253, umul_55057[0]}) % $signed(32'h0000_3ffd));
  assign smod_55393 = $unsigned($signed({8'h00, add_55261, umul_55065[0]}) % $signed(32'h0000_3ffd));
  assign smod_55398 = $unsigned($signed({9'h000, add_55269, umul_55073[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55403 = $unsigned($signed({9'h000, add_55277, umul_55081[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55408 = $unsigned($signed({9'h000, add_55285, umul_55089[0]}) % $signed(32'h0000_3ffd));
  assign smod_55413 = $unsigned($signed({9'h000, add_55293, umul_55097[0]}) % $signed(32'h0000_3ffd));
  assign umul_55429 = umul23b_16b_x_7b(array_index_54717, 7'h49);
  assign add_55431 = {1'h0, umul_55235[22:3]} + 21'h00_07e9;
  assign sel_55436 = $signed({1'h0, smod_55184[15:0]}) < $signed({1'h0, sel_55242}) ? smod_55184[15:0] : sel_55242;
  assign umul_55437 = umul23b_16b_x_7b(array_index_54723, 7'h49);
  assign add_55439 = {1'h0, umul_55243[22:3]} + 21'h00_07e9;
  assign sel_55444 = $signed({1'h0, smod_55189[15:0]}) < $signed({1'h0, sel_55250}) ? smod_55189[15:0] : sel_55250;
  assign umul_55445 = umul23b_16b_x_7b(array_index_54911, 7'h47);
  assign add_55447 = {1'h0, umul_55251[22:1]} + 23'h00_1f8b;
  assign sel_55452 = $signed({1'h0, smod_55194[15:0]}) < $signed({1'h0, sel_55258}) ? smod_55194[15:0] : sel_55258;
  assign umul_55453 = umul23b_16b_x_7b(array_index_54917, 7'h47);
  assign add_55455 = {1'h0, umul_55259[22:1]} + 23'h00_1f8b;
  assign sel_55460 = $signed({1'h0, smod_55199[15:0]}) < $signed({1'h0, sel_55266}) ? smod_55199[15:0] : sel_55266;
  assign umul_55461 = umul22b_16b_x_6b(array_index_55105, 6'h3d);
  assign add_55463 = {1'h0, umul_55267[21:2]} + 21'h00_0fb9;
  assign sel_55468 = $signed({1'h0, smod_55204[15:0]}) < $signed({1'h0, sel_55274}) ? smod_55204[15:0] : sel_55274;
  assign umul_55469 = umul22b_16b_x_6b(array_index_55111, 6'h3d);
  assign add_55471 = {1'h0, umul_55275[21:2]} + 21'h00_0fb9;
  assign sel_55476 = $signed({1'h0, smod_55209[15:0]}) < $signed({1'h0, sel_55282}) ? smod_55209[15:0] : sel_55282;
  assign umul_55477 = umul22b_16b_x_6b(array_index_55299, 6'h3b);
  assign add_55479 = {1'h0, umul_55283[21:1]} + 22'h00_1f59;
  assign sel_55484 = $signed({1'h0, smod_55214[15:0]}) < $signed({1'h0, sel_55290}) ? smod_55214[15:0] : sel_55290;
  assign umul_55485 = umul22b_16b_x_6b(array_index_55305, 6'h3b);
  assign add_55487 = {1'h0, umul_55291[21:1]} + 22'h00_1f59;
  assign sel_55492 = $signed({1'h0, smod_55219[15:0]}) < $signed({1'h0, sel_55298}) ? smod_55219[15:0] : sel_55298;
  assign array_index_55493 = set1_unflattened[5'h13];
  assign smod_55497 = $unsigned($signed({9'h000, add_55361, umul_55165[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_55499 = set2_unflattened[5'h13];
  assign smod_55503 = $unsigned($signed({9'h000, add_55369, umul_55173[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_55553 = umul22b_16b_x_6b(array_index_55493, 6'h35);
  assign add_55555 = {1'h0, umul_55359[21:7]} + 16'h007d;
  assign sel_55560 = $signed({1'h0, smod_55303[15:0]}) < $signed({1'h0, sel_55366}) ? smod_55303[15:0] : sel_55366;
  assign umul_55561 = umul22b_16b_x_6b(array_index_55499, 6'h35);
  assign add_55563 = {1'h0, umul_55367[21:7]} + 16'h007d;
  assign sel_55568 = $signed({1'h0, smod_55309[15:0]}) < $signed({1'h0, sel_55374}) ? smod_55309[15:0] : sel_55374;
  assign smod_55572 = $unsigned($signed({8'h00, add_55431, umul_55235[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55577 = $unsigned($signed({8'h00, add_55439, umul_55243[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55582 = $unsigned($signed({8'h00, add_55447, umul_55251[0]}) % $signed(32'h0000_3ffd));
  assign smod_55587 = $unsigned($signed({8'h00, add_55455, umul_55259[0]}) % $signed(32'h0000_3ffd));
  assign smod_55592 = $unsigned($signed({9'h000, add_55463, umul_55267[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55597 = $unsigned($signed({9'h000, add_55471, umul_55275[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55602 = $unsigned($signed({9'h000, add_55479, umul_55283[0]}) % $signed(32'h0000_3ffd));
  assign smod_55607 = $unsigned($signed({9'h000, add_55487, umul_55291[0]}) % $signed(32'h0000_3ffd));
  assign umul_55623 = umul23b_16b_x_7b(array_index_54911, 7'h49);
  assign add_55625 = {1'h0, umul_55429[22:3]} + 21'h00_07e9;
  assign sel_55630 = $signed({1'h0, smod_55378[15:0]}) < $signed({1'h0, sel_55436}) ? smod_55378[15:0] : sel_55436;
  assign umul_55631 = umul23b_16b_x_7b(array_index_54917, 7'h49);
  assign add_55633 = {1'h0, umul_55437[22:3]} + 21'h00_07e9;
  assign sel_55638 = $signed({1'h0, smod_55383[15:0]}) < $signed({1'h0, sel_55444}) ? smod_55383[15:0] : sel_55444;
  assign umul_55639 = umul23b_16b_x_7b(array_index_55105, 7'h47);
  assign add_55641 = {1'h0, umul_55445[22:1]} + 23'h00_1f8b;
  assign sel_55646 = $signed({1'h0, smod_55388[15:0]}) < $signed({1'h0, sel_55452}) ? smod_55388[15:0] : sel_55452;
  assign umul_55647 = umul23b_16b_x_7b(array_index_55111, 7'h47);
  assign add_55649 = {1'h0, umul_55453[22:1]} + 23'h00_1f8b;
  assign sel_55654 = $signed({1'h0, smod_55393[15:0]}) < $signed({1'h0, sel_55460}) ? smod_55393[15:0] : sel_55460;
  assign umul_55655 = umul22b_16b_x_6b(array_index_55299, 6'h3d);
  assign add_55657 = {1'h0, umul_55461[21:2]} + 21'h00_0fb9;
  assign sel_55662 = $signed({1'h0, smod_55398[15:0]}) < $signed({1'h0, sel_55468}) ? smod_55398[15:0] : sel_55468;
  assign umul_55663 = umul22b_16b_x_6b(array_index_55305, 6'h3d);
  assign add_55665 = {1'h0, umul_55469[21:2]} + 21'h00_0fb9;
  assign sel_55670 = $signed({1'h0, smod_55403[15:0]}) < $signed({1'h0, sel_55476}) ? smod_55403[15:0] : sel_55476;
  assign umul_55671 = umul22b_16b_x_6b(array_index_55493, 6'h3b);
  assign add_55673 = {1'h0, umul_55477[21:1]} + 22'h00_1f59;
  assign sel_55678 = $signed({1'h0, smod_55408[15:0]}) < $signed({1'h0, sel_55484}) ? smod_55408[15:0] : sel_55484;
  assign umul_55679 = umul22b_16b_x_6b(array_index_55499, 6'h3b);
  assign add_55681 = {1'h0, umul_55485[21:1]} + 22'h00_1f59;
  assign sel_55686 = $signed({1'h0, smod_55413[15:0]}) < $signed({1'h0, sel_55492}) ? smod_55413[15:0] : sel_55492;
  assign array_index_55687 = set1_unflattened[5'h14];
  assign smod_55691 = $unsigned($signed({9'h000, add_55555, umul_55359[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_55693 = set2_unflattened[5'h14];
  assign smod_55697 = $unsigned($signed({9'h000, add_55563, umul_55367[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_55747 = umul22b_16b_x_6b(array_index_55687, 6'h35);
  assign add_55749 = {1'h0, umul_55553[21:7]} + 16'h007d;
  assign sel_55754 = $signed({1'h0, smod_55497[15:0]}) < $signed({1'h0, sel_55560}) ? smod_55497[15:0] : sel_55560;
  assign umul_55755 = umul22b_16b_x_6b(array_index_55693, 6'h35);
  assign add_55757 = {1'h0, umul_55561[21:7]} + 16'h007d;
  assign sel_55762 = $signed({1'h0, smod_55503[15:0]}) < $signed({1'h0, sel_55568}) ? smod_55503[15:0] : sel_55568;
  assign smod_55766 = $unsigned($signed({8'h00, add_55625, umul_55429[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55771 = $unsigned($signed({8'h00, add_55633, umul_55437[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55776 = $unsigned($signed({8'h00, add_55641, umul_55445[0]}) % $signed(32'h0000_3ffd));
  assign smod_55781 = $unsigned($signed({8'h00, add_55649, umul_55453[0]}) % $signed(32'h0000_3ffd));
  assign smod_55786 = $unsigned($signed({9'h000, add_55657, umul_55461[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55791 = $unsigned($signed({9'h000, add_55665, umul_55469[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55796 = $unsigned($signed({9'h000, add_55673, umul_55477[0]}) % $signed(32'h0000_3ffd));
  assign smod_55801 = $unsigned($signed({9'h000, add_55681, umul_55485[0]}) % $signed(32'h0000_3ffd));
  assign umul_55817 = umul23b_16b_x_7b(array_index_55105, 7'h49);
  assign add_55819 = {1'h0, umul_55623[22:3]} + 21'h00_07e9;
  assign sel_55824 = $signed({1'h0, smod_55572[15:0]}) < $signed({1'h0, sel_55630}) ? smod_55572[15:0] : sel_55630;
  assign umul_55825 = umul23b_16b_x_7b(array_index_55111, 7'h49);
  assign add_55827 = {1'h0, umul_55631[22:3]} + 21'h00_07e9;
  assign sel_55832 = $signed({1'h0, smod_55577[15:0]}) < $signed({1'h0, sel_55638}) ? smod_55577[15:0] : sel_55638;
  assign umul_55833 = umul23b_16b_x_7b(array_index_55299, 7'h47);
  assign add_55835 = {1'h0, umul_55639[22:1]} + 23'h00_1f8b;
  assign sel_55840 = $signed({1'h0, smod_55582[15:0]}) < $signed({1'h0, sel_55646}) ? smod_55582[15:0] : sel_55646;
  assign umul_55841 = umul23b_16b_x_7b(array_index_55305, 7'h47);
  assign add_55843 = {1'h0, umul_55647[22:1]} + 23'h00_1f8b;
  assign sel_55848 = $signed({1'h0, smod_55587[15:0]}) < $signed({1'h0, sel_55654}) ? smod_55587[15:0] : sel_55654;
  assign umul_55849 = umul22b_16b_x_6b(array_index_55493, 6'h3d);
  assign add_55851 = {1'h0, umul_55655[21:2]} + 21'h00_0fb9;
  assign sel_55856 = $signed({1'h0, smod_55592[15:0]}) < $signed({1'h0, sel_55662}) ? smod_55592[15:0] : sel_55662;
  assign umul_55857 = umul22b_16b_x_6b(array_index_55499, 6'h3d);
  assign add_55859 = {1'h0, umul_55663[21:2]} + 21'h00_0fb9;
  assign sel_55864 = $signed({1'h0, smod_55597[15:0]}) < $signed({1'h0, sel_55670}) ? smod_55597[15:0] : sel_55670;
  assign umul_55865 = umul22b_16b_x_6b(array_index_55687, 6'h3b);
  assign add_55867 = {1'h0, umul_55671[21:1]} + 22'h00_1f59;
  assign sel_55872 = $signed({1'h0, smod_55602[15:0]}) < $signed({1'h0, sel_55678}) ? smod_55602[15:0] : sel_55678;
  assign umul_55873 = umul22b_16b_x_6b(array_index_55693, 6'h3b);
  assign add_55875 = {1'h0, umul_55679[21:1]} + 22'h00_1f59;
  assign sel_55880 = $signed({1'h0, smod_55607[15:0]}) < $signed({1'h0, sel_55686}) ? smod_55607[15:0] : sel_55686;
  assign array_index_55881 = set1_unflattened[5'h15];
  assign smod_55885 = $unsigned($signed({9'h000, add_55749, umul_55553[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_55887 = set2_unflattened[5'h15];
  assign smod_55891 = $unsigned($signed({9'h000, add_55757, umul_55561[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_55941 = umul22b_16b_x_6b(array_index_55881, 6'h35);
  assign add_55943 = {1'h0, umul_55747[21:7]} + 16'h007d;
  assign sel_55948 = $signed({1'h0, smod_55691[15:0]}) < $signed({1'h0, sel_55754}) ? smod_55691[15:0] : sel_55754;
  assign umul_55949 = umul22b_16b_x_6b(array_index_55887, 6'h35);
  assign add_55951 = {1'h0, umul_55755[21:7]} + 16'h007d;
  assign sel_55956 = $signed({1'h0, smod_55697[15:0]}) < $signed({1'h0, sel_55762}) ? smod_55697[15:0] : sel_55762;
  assign smod_55960 = $unsigned($signed({8'h00, add_55819, umul_55623[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55965 = $unsigned($signed({8'h00, add_55827, umul_55631[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_55970 = $unsigned($signed({8'h00, add_55835, umul_55639[0]}) % $signed(32'h0000_3ffd));
  assign smod_55975 = $unsigned($signed({8'h00, add_55843, umul_55647[0]}) % $signed(32'h0000_3ffd));
  assign smod_55980 = $unsigned($signed({9'h000, add_55851, umul_55655[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55985 = $unsigned($signed({9'h000, add_55859, umul_55663[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_55990 = $unsigned($signed({9'h000, add_55867, umul_55671[0]}) % $signed(32'h0000_3ffd));
  assign smod_55995 = $unsigned($signed({9'h000, add_55875, umul_55679[0]}) % $signed(32'h0000_3ffd));
  assign umul_56011 = umul23b_16b_x_7b(array_index_55299, 7'h49);
  assign add_56013 = {1'h0, umul_55817[22:3]} + 21'h00_07e9;
  assign sel_56018 = $signed({1'h0, smod_55766[15:0]}) < $signed({1'h0, sel_55824}) ? smod_55766[15:0] : sel_55824;
  assign umul_56019 = umul23b_16b_x_7b(array_index_55305, 7'h49);
  assign add_56021 = {1'h0, umul_55825[22:3]} + 21'h00_07e9;
  assign sel_56026 = $signed({1'h0, smod_55771[15:0]}) < $signed({1'h0, sel_55832}) ? smod_55771[15:0] : sel_55832;
  assign umul_56027 = umul23b_16b_x_7b(array_index_55493, 7'h47);
  assign add_56029 = {1'h0, umul_55833[22:1]} + 23'h00_1f8b;
  assign sel_56034 = $signed({1'h0, smod_55776[15:0]}) < $signed({1'h0, sel_55840}) ? smod_55776[15:0] : sel_55840;
  assign umul_56035 = umul23b_16b_x_7b(array_index_55499, 7'h47);
  assign add_56037 = {1'h0, umul_55841[22:1]} + 23'h00_1f8b;
  assign sel_56042 = $signed({1'h0, smod_55781[15:0]}) < $signed({1'h0, sel_55848}) ? smod_55781[15:0] : sel_55848;
  assign umul_56043 = umul22b_16b_x_6b(array_index_55687, 6'h3d);
  assign add_56045 = {1'h0, umul_55849[21:2]} + 21'h00_0fb9;
  assign sel_56050 = $signed({1'h0, smod_55786[15:0]}) < $signed({1'h0, sel_55856}) ? smod_55786[15:0] : sel_55856;
  assign umul_56051 = umul22b_16b_x_6b(array_index_55693, 6'h3d);
  assign add_56053 = {1'h0, umul_55857[21:2]} + 21'h00_0fb9;
  assign sel_56058 = $signed({1'h0, smod_55791[15:0]}) < $signed({1'h0, sel_55864}) ? smod_55791[15:0] : sel_55864;
  assign umul_56059 = umul22b_16b_x_6b(array_index_55881, 6'h3b);
  assign add_56061 = {1'h0, umul_55865[21:1]} + 22'h00_1f59;
  assign sel_56066 = $signed({1'h0, smod_55796[15:0]}) < $signed({1'h0, sel_55872}) ? smod_55796[15:0] : sel_55872;
  assign umul_56067 = umul22b_16b_x_6b(array_index_55887, 6'h3b);
  assign add_56069 = {1'h0, umul_55873[21:1]} + 22'h00_1f59;
  assign sel_56074 = $signed({1'h0, smod_55801[15:0]}) < $signed({1'h0, sel_55880}) ? smod_55801[15:0] : sel_55880;
  assign array_index_56075 = set1_unflattened[5'h16];
  assign smod_56079 = $unsigned($signed({9'h000, add_55943, umul_55747[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_56081 = set2_unflattened[5'h16];
  assign smod_56085 = $unsigned($signed({9'h000, add_55951, umul_55755[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_56135 = umul22b_16b_x_6b(array_index_56075, 6'h35);
  assign add_56137 = {1'h0, umul_55941[21:7]} + 16'h007d;
  assign sel_56142 = $signed({1'h0, smod_55885[15:0]}) < $signed({1'h0, sel_55948}) ? smod_55885[15:0] : sel_55948;
  assign umul_56143 = umul22b_16b_x_6b(array_index_56081, 6'h35);
  assign add_56145 = {1'h0, umul_55949[21:7]} + 16'h007d;
  assign sel_56150 = $signed({1'h0, smod_55891[15:0]}) < $signed({1'h0, sel_55956}) ? smod_55891[15:0] : sel_55956;
  assign smod_56154 = $unsigned($signed({8'h00, add_56013, umul_55817[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56159 = $unsigned($signed({8'h00, add_56021, umul_55825[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56164 = $unsigned($signed({8'h00, add_56029, umul_55833[0]}) % $signed(32'h0000_3ffd));
  assign smod_56169 = $unsigned($signed({8'h00, add_56037, umul_55841[0]}) % $signed(32'h0000_3ffd));
  assign smod_56174 = $unsigned($signed({9'h000, add_56045, umul_55849[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56179 = $unsigned($signed({9'h000, add_56053, umul_55857[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56184 = $unsigned($signed({9'h000, add_56061, umul_55865[0]}) % $signed(32'h0000_3ffd));
  assign smod_56189 = $unsigned($signed({9'h000, add_56069, umul_55873[0]}) % $signed(32'h0000_3ffd));
  assign umul_56205 = umul23b_16b_x_7b(array_index_55493, 7'h49);
  assign add_56207 = {1'h0, umul_56011[22:3]} + 21'h00_07e9;
  assign sel_56212 = $signed({1'h0, smod_55960[15:0]}) < $signed({1'h0, sel_56018}) ? smod_55960[15:0] : sel_56018;
  assign umul_56213 = umul23b_16b_x_7b(array_index_55499, 7'h49);
  assign add_56215 = {1'h0, umul_56019[22:3]} + 21'h00_07e9;
  assign sel_56220 = $signed({1'h0, smod_55965[15:0]}) < $signed({1'h0, sel_56026}) ? smod_55965[15:0] : sel_56026;
  assign umul_56221 = umul23b_16b_x_7b(array_index_55687, 7'h47);
  assign add_56223 = {1'h0, umul_56027[22:1]} + 23'h00_1f8b;
  assign sel_56228 = $signed({1'h0, smod_55970[15:0]}) < $signed({1'h0, sel_56034}) ? smod_55970[15:0] : sel_56034;
  assign umul_56229 = umul23b_16b_x_7b(array_index_55693, 7'h47);
  assign add_56231 = {1'h0, umul_56035[22:1]} + 23'h00_1f8b;
  assign sel_56236 = $signed({1'h0, smod_55975[15:0]}) < $signed({1'h0, sel_56042}) ? smod_55975[15:0] : sel_56042;
  assign umul_56237 = umul22b_16b_x_6b(array_index_55881, 6'h3d);
  assign add_56239 = {1'h0, umul_56043[21:2]} + 21'h00_0fb9;
  assign sel_56244 = $signed({1'h0, smod_55980[15:0]}) < $signed({1'h0, sel_56050}) ? smod_55980[15:0] : sel_56050;
  assign umul_56245 = umul22b_16b_x_6b(array_index_55887, 6'h3d);
  assign add_56247 = {1'h0, umul_56051[21:2]} + 21'h00_0fb9;
  assign sel_56252 = $signed({1'h0, smod_55985[15:0]}) < $signed({1'h0, sel_56058}) ? smod_55985[15:0] : sel_56058;
  assign umul_56253 = umul22b_16b_x_6b(array_index_56075, 6'h3b);
  assign add_56255 = {1'h0, umul_56059[21:1]} + 22'h00_1f59;
  assign sel_56260 = $signed({1'h0, smod_55990[15:0]}) < $signed({1'h0, sel_56066}) ? smod_55990[15:0] : sel_56066;
  assign umul_56261 = umul22b_16b_x_6b(array_index_56081, 6'h3b);
  assign add_56263 = {1'h0, umul_56067[21:1]} + 22'h00_1f59;
  assign sel_56268 = $signed({1'h0, smod_55995[15:0]}) < $signed({1'h0, sel_56074}) ? smod_55995[15:0] : sel_56074;
  assign array_index_56269 = set1_unflattened[5'h17];
  assign smod_56273 = $unsigned($signed({9'h000, add_56137, umul_55941[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_56275 = set2_unflattened[5'h17];
  assign smod_56279 = $unsigned($signed({9'h000, add_56145, umul_55949[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_56329 = umul22b_16b_x_6b(array_index_56269, 6'h35);
  assign add_56331 = {1'h0, umul_56135[21:7]} + 16'h007d;
  assign sel_56336 = $signed({1'h0, smod_56079[15:0]}) < $signed({1'h0, sel_56142}) ? smod_56079[15:0] : sel_56142;
  assign umul_56337 = umul22b_16b_x_6b(array_index_56275, 6'h35);
  assign add_56339 = {1'h0, umul_56143[21:7]} + 16'h007d;
  assign sel_56344 = $signed({1'h0, smod_56085[15:0]}) < $signed({1'h0, sel_56150}) ? smod_56085[15:0] : sel_56150;
  assign smod_56348 = $unsigned($signed({8'h00, add_56207, umul_56011[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56353 = $unsigned($signed({8'h00, add_56215, umul_56019[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56358 = $unsigned($signed({8'h00, add_56223, umul_56027[0]}) % $signed(32'h0000_3ffd));
  assign smod_56363 = $unsigned($signed({8'h00, add_56231, umul_56035[0]}) % $signed(32'h0000_3ffd));
  assign smod_56368 = $unsigned($signed({9'h000, add_56239, umul_56043[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56373 = $unsigned($signed({9'h000, add_56247, umul_56051[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56378 = $unsigned($signed({9'h000, add_56255, umul_56059[0]}) % $signed(32'h0000_3ffd));
  assign smod_56383 = $unsigned($signed({9'h000, add_56263, umul_56067[0]}) % $signed(32'h0000_3ffd));
  assign umul_56399 = umul23b_16b_x_7b(array_index_55687, 7'h49);
  assign add_56401 = {1'h0, umul_56205[22:3]} + 21'h00_07e9;
  assign sel_56406 = $signed({1'h0, smod_56154[15:0]}) < $signed({1'h0, sel_56212}) ? smod_56154[15:0] : sel_56212;
  assign umul_56407 = umul23b_16b_x_7b(array_index_55693, 7'h49);
  assign add_56409 = {1'h0, umul_56213[22:3]} + 21'h00_07e9;
  assign sel_56414 = $signed({1'h0, smod_56159[15:0]}) < $signed({1'h0, sel_56220}) ? smod_56159[15:0] : sel_56220;
  assign umul_56415 = umul23b_16b_x_7b(array_index_55881, 7'h47);
  assign add_56417 = {1'h0, umul_56221[22:1]} + 23'h00_1f8b;
  assign sel_56422 = $signed({1'h0, smod_56164[15:0]}) < $signed({1'h0, sel_56228}) ? smod_56164[15:0] : sel_56228;
  assign umul_56423 = umul23b_16b_x_7b(array_index_55887, 7'h47);
  assign add_56425 = {1'h0, umul_56229[22:1]} + 23'h00_1f8b;
  assign sel_56430 = $signed({1'h0, smod_56169[15:0]}) < $signed({1'h0, sel_56236}) ? smod_56169[15:0] : sel_56236;
  assign umul_56431 = umul22b_16b_x_6b(array_index_56075, 6'h3d);
  assign add_56433 = {1'h0, umul_56237[21:2]} + 21'h00_0fb9;
  assign sel_56438 = $signed({1'h0, smod_56174[15:0]}) < $signed({1'h0, sel_56244}) ? smod_56174[15:0] : sel_56244;
  assign umul_56439 = umul22b_16b_x_6b(array_index_56081, 6'h3d);
  assign add_56441 = {1'h0, umul_56245[21:2]} + 21'h00_0fb9;
  assign sel_56446 = $signed({1'h0, smod_56179[15:0]}) < $signed({1'h0, sel_56252}) ? smod_56179[15:0] : sel_56252;
  assign umul_56447 = umul22b_16b_x_6b(array_index_56269, 6'h3b);
  assign add_56449 = {1'h0, umul_56253[21:1]} + 22'h00_1f59;
  assign sel_56454 = $signed({1'h0, smod_56184[15:0]}) < $signed({1'h0, sel_56260}) ? smod_56184[15:0] : sel_56260;
  assign umul_56455 = umul22b_16b_x_6b(array_index_56275, 6'h3b);
  assign add_56457 = {1'h0, umul_56261[21:1]} + 22'h00_1f59;
  assign sel_56462 = $signed({1'h0, smod_56189[15:0]}) < $signed({1'h0, sel_56268}) ? smod_56189[15:0] : sel_56268;
  assign array_index_56463 = set1_unflattened[5'h18];
  assign smod_56467 = $unsigned($signed({9'h000, add_56331, umul_56135[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_56469 = set2_unflattened[5'h18];
  assign smod_56473 = $unsigned($signed({9'h000, add_56339, umul_56143[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_56523 = umul22b_16b_x_6b(array_index_56463, 6'h35);
  assign add_56525 = {1'h0, umul_56329[21:7]} + 16'h007d;
  assign sel_56530 = $signed({1'h0, smod_56273[15:0]}) < $signed({1'h0, sel_56336}) ? smod_56273[15:0] : sel_56336;
  assign umul_56531 = umul22b_16b_x_6b(array_index_56469, 6'h35);
  assign add_56533 = {1'h0, umul_56337[21:7]} + 16'h007d;
  assign sel_56538 = $signed({1'h0, smod_56279[15:0]}) < $signed({1'h0, sel_56344}) ? smod_56279[15:0] : sel_56344;
  assign smod_56542 = $unsigned($signed({8'h00, add_56401, umul_56205[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56547 = $unsigned($signed({8'h00, add_56409, umul_56213[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56552 = $unsigned($signed({8'h00, add_56417, umul_56221[0]}) % $signed(32'h0000_3ffd));
  assign smod_56557 = $unsigned($signed({8'h00, add_56425, umul_56229[0]}) % $signed(32'h0000_3ffd));
  assign smod_56562 = $unsigned($signed({9'h000, add_56433, umul_56237[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56567 = $unsigned($signed({9'h000, add_56441, umul_56245[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56572 = $unsigned($signed({9'h000, add_56449, umul_56253[0]}) % $signed(32'h0000_3ffd));
  assign smod_56577 = $unsigned($signed({9'h000, add_56457, umul_56261[0]}) % $signed(32'h0000_3ffd));
  assign umul_56593 = umul23b_16b_x_7b(array_index_55881, 7'h49);
  assign add_56595 = {1'h0, umul_56399[22:3]} + 21'h00_07e9;
  assign sel_56600 = $signed({1'h0, smod_56348[15:0]}) < $signed({1'h0, sel_56406}) ? smod_56348[15:0] : sel_56406;
  assign umul_56601 = umul23b_16b_x_7b(array_index_55887, 7'h49);
  assign add_56603 = {1'h0, umul_56407[22:3]} + 21'h00_07e9;
  assign sel_56608 = $signed({1'h0, smod_56353[15:0]}) < $signed({1'h0, sel_56414}) ? smod_56353[15:0] : sel_56414;
  assign umul_56609 = umul23b_16b_x_7b(array_index_56075, 7'h47);
  assign add_56611 = {1'h0, umul_56415[22:1]} + 23'h00_1f8b;
  assign sel_56616 = $signed({1'h0, smod_56358[15:0]}) < $signed({1'h0, sel_56422}) ? smod_56358[15:0] : sel_56422;
  assign umul_56617 = umul23b_16b_x_7b(array_index_56081, 7'h47);
  assign add_56619 = {1'h0, umul_56423[22:1]} + 23'h00_1f8b;
  assign sel_56624 = $signed({1'h0, smod_56363[15:0]}) < $signed({1'h0, sel_56430}) ? smod_56363[15:0] : sel_56430;
  assign umul_56625 = umul22b_16b_x_6b(array_index_56269, 6'h3d);
  assign add_56627 = {1'h0, umul_56431[21:2]} + 21'h00_0fb9;
  assign sel_56632 = $signed({1'h0, smod_56368[15:0]}) < $signed({1'h0, sel_56438}) ? smod_56368[15:0] : sel_56438;
  assign umul_56633 = umul22b_16b_x_6b(array_index_56275, 6'h3d);
  assign add_56635 = {1'h0, umul_56439[21:2]} + 21'h00_0fb9;
  assign sel_56640 = $signed({1'h0, smod_56373[15:0]}) < $signed({1'h0, sel_56446}) ? smod_56373[15:0] : sel_56446;
  assign umul_56641 = umul22b_16b_x_6b(array_index_56463, 6'h3b);
  assign add_56643 = {1'h0, umul_56447[21:1]} + 22'h00_1f59;
  assign sel_56648 = $signed({1'h0, smod_56378[15:0]}) < $signed({1'h0, sel_56454}) ? smod_56378[15:0] : sel_56454;
  assign umul_56649 = umul22b_16b_x_6b(array_index_56469, 6'h3b);
  assign add_56651 = {1'h0, umul_56455[21:1]} + 22'h00_1f59;
  assign sel_56656 = $signed({1'h0, smod_56383[15:0]}) < $signed({1'h0, sel_56462}) ? smod_56383[15:0] : sel_56462;
  assign array_index_56657 = set1_unflattened[5'h19];
  assign smod_56661 = $unsigned($signed({9'h000, add_56525, umul_56329[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_56663 = set2_unflattened[5'h19];
  assign smod_56667 = $unsigned($signed({9'h000, add_56533, umul_56337[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_56717 = umul22b_16b_x_6b(array_index_56657, 6'h35);
  assign add_56719 = {1'h0, umul_56523[21:7]} + 16'h007d;
  assign sel_56724 = $signed({1'h0, smod_56467[15:0]}) < $signed({1'h0, sel_56530}) ? smod_56467[15:0] : sel_56530;
  assign umul_56725 = umul22b_16b_x_6b(array_index_56663, 6'h35);
  assign add_56727 = {1'h0, umul_56531[21:7]} + 16'h007d;
  assign sel_56732 = $signed({1'h0, smod_56473[15:0]}) < $signed({1'h0, sel_56538}) ? smod_56473[15:0] : sel_56538;
  assign smod_56736 = $unsigned($signed({8'h00, add_56595, umul_56399[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56741 = $unsigned($signed({8'h00, add_56603, umul_56407[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56746 = $unsigned($signed({8'h00, add_56611, umul_56415[0]}) % $signed(32'h0000_3ffd));
  assign smod_56751 = $unsigned($signed({8'h00, add_56619, umul_56423[0]}) % $signed(32'h0000_3ffd));
  assign smod_56756 = $unsigned($signed({9'h000, add_56627, umul_56431[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56761 = $unsigned($signed({9'h000, add_56635, umul_56439[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56766 = $unsigned($signed({9'h000, add_56643, umul_56447[0]}) % $signed(32'h0000_3ffd));
  assign smod_56771 = $unsigned($signed({9'h000, add_56651, umul_56455[0]}) % $signed(32'h0000_3ffd));
  assign umul_56787 = umul23b_16b_x_7b(array_index_56075, 7'h49);
  assign add_56789 = {1'h0, umul_56593[22:3]} + 21'h00_07e9;
  assign sel_56794 = $signed({1'h0, smod_56542[15:0]}) < $signed({1'h0, sel_56600}) ? smod_56542[15:0] : sel_56600;
  assign umul_56795 = umul23b_16b_x_7b(array_index_56081, 7'h49);
  assign add_56797 = {1'h0, umul_56601[22:3]} + 21'h00_07e9;
  assign sel_56802 = $signed({1'h0, smod_56547[15:0]}) < $signed({1'h0, sel_56608}) ? smod_56547[15:0] : sel_56608;
  assign umul_56803 = umul23b_16b_x_7b(array_index_56269, 7'h47);
  assign add_56805 = {1'h0, umul_56609[22:1]} + 23'h00_1f8b;
  assign sel_56810 = $signed({1'h0, smod_56552[15:0]}) < $signed({1'h0, sel_56616}) ? smod_56552[15:0] : sel_56616;
  assign umul_56811 = umul23b_16b_x_7b(array_index_56275, 7'h47);
  assign add_56813 = {1'h0, umul_56617[22:1]} + 23'h00_1f8b;
  assign sel_56818 = $signed({1'h0, smod_56557[15:0]}) < $signed({1'h0, sel_56624}) ? smod_56557[15:0] : sel_56624;
  assign umul_56819 = umul22b_16b_x_6b(array_index_56463, 6'h3d);
  assign add_56821 = {1'h0, umul_56625[21:2]} + 21'h00_0fb9;
  assign sel_56826 = $signed({1'h0, smod_56562[15:0]}) < $signed({1'h0, sel_56632}) ? smod_56562[15:0] : sel_56632;
  assign umul_56827 = umul22b_16b_x_6b(array_index_56469, 6'h3d);
  assign add_56829 = {1'h0, umul_56633[21:2]} + 21'h00_0fb9;
  assign sel_56834 = $signed({1'h0, smod_56567[15:0]}) < $signed({1'h0, sel_56640}) ? smod_56567[15:0] : sel_56640;
  assign umul_56835 = umul22b_16b_x_6b(array_index_56657, 6'h3b);
  assign add_56837 = {1'h0, umul_56641[21:1]} + 22'h00_1f59;
  assign sel_56842 = $signed({1'h0, smod_56572[15:0]}) < $signed({1'h0, sel_56648}) ? smod_56572[15:0] : sel_56648;
  assign umul_56843 = umul22b_16b_x_6b(array_index_56663, 6'h3b);
  assign add_56845 = {1'h0, umul_56649[21:1]} + 22'h00_1f59;
  assign sel_56850 = $signed({1'h0, smod_56577[15:0]}) < $signed({1'h0, sel_56656}) ? smod_56577[15:0] : sel_56656;
  assign array_index_56851 = set1_unflattened[5'h1a];
  assign smod_56855 = $unsigned($signed({9'h000, add_56719, umul_56523[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_56857 = set2_unflattened[5'h1a];
  assign smod_56861 = $unsigned($signed({9'h000, add_56727, umul_56531[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_56911 = umul22b_16b_x_6b(array_index_56851, 6'h35);
  assign add_56913 = {1'h0, umul_56717[21:7]} + 16'h007d;
  assign sel_56918 = $signed({1'h0, smod_56661[15:0]}) < $signed({1'h0, sel_56724}) ? smod_56661[15:0] : sel_56724;
  assign umul_56919 = umul22b_16b_x_6b(array_index_56857, 6'h35);
  assign add_56921 = {1'h0, umul_56725[21:7]} + 16'h007d;
  assign sel_56926 = $signed({1'h0, smod_56667[15:0]}) < $signed({1'h0, sel_56732}) ? smod_56667[15:0] : sel_56732;
  assign smod_56930 = $unsigned($signed({8'h00, add_56789, umul_56593[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56935 = $unsigned($signed({8'h00, add_56797, umul_56601[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_56940 = $unsigned($signed({8'h00, add_56805, umul_56609[0]}) % $signed(32'h0000_3ffd));
  assign smod_56945 = $unsigned($signed({8'h00, add_56813, umul_56617[0]}) % $signed(32'h0000_3ffd));
  assign smod_56950 = $unsigned($signed({9'h000, add_56821, umul_56625[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56955 = $unsigned($signed({9'h000, add_56829, umul_56633[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_56960 = $unsigned($signed({9'h000, add_56837, umul_56641[0]}) % $signed(32'h0000_3ffd));
  assign smod_56965 = $unsigned($signed({9'h000, add_56845, umul_56649[0]}) % $signed(32'h0000_3ffd));
  assign umul_56981 = umul23b_16b_x_7b(array_index_56269, 7'h49);
  assign add_56983 = {1'h0, umul_56787[22:3]} + 21'h00_07e9;
  assign sel_56988 = $signed({1'h0, smod_56736[15:0]}) < $signed({1'h0, sel_56794}) ? smod_56736[15:0] : sel_56794;
  assign umul_56989 = umul23b_16b_x_7b(array_index_56275, 7'h49);
  assign add_56991 = {1'h0, umul_56795[22:3]} + 21'h00_07e9;
  assign sel_56996 = $signed({1'h0, smod_56741[15:0]}) < $signed({1'h0, sel_56802}) ? smod_56741[15:0] : sel_56802;
  assign umul_56997 = umul23b_16b_x_7b(array_index_56463, 7'h47);
  assign add_56999 = {1'h0, umul_56803[22:1]} + 23'h00_1f8b;
  assign sel_57004 = $signed({1'h0, smod_56746[15:0]}) < $signed({1'h0, sel_56810}) ? smod_56746[15:0] : sel_56810;
  assign umul_57005 = umul23b_16b_x_7b(array_index_56469, 7'h47);
  assign add_57007 = {1'h0, umul_56811[22:1]} + 23'h00_1f8b;
  assign sel_57012 = $signed({1'h0, smod_56751[15:0]}) < $signed({1'h0, sel_56818}) ? smod_56751[15:0] : sel_56818;
  assign umul_57013 = umul22b_16b_x_6b(array_index_56657, 6'h3d);
  assign add_57015 = {1'h0, umul_56819[21:2]} + 21'h00_0fb9;
  assign sel_57020 = $signed({1'h0, smod_56756[15:0]}) < $signed({1'h0, sel_56826}) ? smod_56756[15:0] : sel_56826;
  assign umul_57021 = umul22b_16b_x_6b(array_index_56663, 6'h3d);
  assign add_57023 = {1'h0, umul_56827[21:2]} + 21'h00_0fb9;
  assign sel_57028 = $signed({1'h0, smod_56761[15:0]}) < $signed({1'h0, sel_56834}) ? smod_56761[15:0] : sel_56834;
  assign umul_57029 = umul22b_16b_x_6b(array_index_56851, 6'h3b);
  assign add_57031 = {1'h0, umul_56835[21:1]} + 22'h00_1f59;
  assign sel_57036 = $signed({1'h0, smod_56766[15:0]}) < $signed({1'h0, sel_56842}) ? smod_56766[15:0] : sel_56842;
  assign umul_57037 = umul22b_16b_x_6b(array_index_56857, 6'h3b);
  assign add_57039 = {1'h0, umul_56843[21:1]} + 22'h00_1f59;
  assign sel_57044 = $signed({1'h0, smod_56771[15:0]}) < $signed({1'h0, sel_56850}) ? smod_56771[15:0] : sel_56850;
  assign array_index_57045 = set1_unflattened[5'h1b];
  assign smod_57049 = $unsigned($signed({9'h000, add_56913, umul_56717[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_57051 = set2_unflattened[5'h1b];
  assign smod_57055 = $unsigned($signed({9'h000, add_56921, umul_56725[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_57105 = umul22b_16b_x_6b(array_index_57045, 6'h35);
  assign add_57107 = {1'h0, umul_56911[21:7]} + 16'h007d;
  assign sel_57112 = $signed({1'h0, smod_56855[15:0]}) < $signed({1'h0, sel_56918}) ? smod_56855[15:0] : sel_56918;
  assign umul_57113 = umul22b_16b_x_6b(array_index_57051, 6'h35);
  assign add_57115 = {1'h0, umul_56919[21:7]} + 16'h007d;
  assign sel_57120 = $signed({1'h0, smod_56861[15:0]}) < $signed({1'h0, sel_56926}) ? smod_56861[15:0] : sel_56926;
  assign smod_57124 = $unsigned($signed({8'h00, add_56983, umul_56787[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57129 = $unsigned($signed({8'h00, add_56991, umul_56795[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57134 = $unsigned($signed({8'h00, add_56999, umul_56803[0]}) % $signed(32'h0000_3ffd));
  assign smod_57139 = $unsigned($signed({8'h00, add_57007, umul_56811[0]}) % $signed(32'h0000_3ffd));
  assign smod_57144 = $unsigned($signed({9'h000, add_57015, umul_56819[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57149 = $unsigned($signed({9'h000, add_57023, umul_56827[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57154 = $unsigned($signed({9'h000, add_57031, umul_56835[0]}) % $signed(32'h0000_3ffd));
  assign smod_57159 = $unsigned($signed({9'h000, add_57039, umul_56843[0]}) % $signed(32'h0000_3ffd));
  assign umul_57175 = umul23b_16b_x_7b(array_index_56463, 7'h49);
  assign add_57177 = {1'h0, umul_56981[22:3]} + 21'h00_07e9;
  assign sel_57182 = $signed({1'h0, smod_56930[15:0]}) < $signed({1'h0, sel_56988}) ? smod_56930[15:0] : sel_56988;
  assign umul_57183 = umul23b_16b_x_7b(array_index_56469, 7'h49);
  assign add_57185 = {1'h0, umul_56989[22:3]} + 21'h00_07e9;
  assign sel_57190 = $signed({1'h0, smod_56935[15:0]}) < $signed({1'h0, sel_56996}) ? smod_56935[15:0] : sel_56996;
  assign umul_57191 = umul23b_16b_x_7b(array_index_56657, 7'h47);
  assign add_57193 = {1'h0, umul_56997[22:1]} + 23'h00_1f8b;
  assign sel_57198 = $signed({1'h0, smod_56940[15:0]}) < $signed({1'h0, sel_57004}) ? smod_56940[15:0] : sel_57004;
  assign umul_57199 = umul23b_16b_x_7b(array_index_56663, 7'h47);
  assign add_57201 = {1'h0, umul_57005[22:1]} + 23'h00_1f8b;
  assign sel_57206 = $signed({1'h0, smod_56945[15:0]}) < $signed({1'h0, sel_57012}) ? smod_56945[15:0] : sel_57012;
  assign umul_57207 = umul22b_16b_x_6b(array_index_56851, 6'h3d);
  assign add_57209 = {1'h0, umul_57013[21:2]} + 21'h00_0fb9;
  assign sel_57214 = $signed({1'h0, smod_56950[15:0]}) < $signed({1'h0, sel_57020}) ? smod_56950[15:0] : sel_57020;
  assign umul_57215 = umul22b_16b_x_6b(array_index_56857, 6'h3d);
  assign add_57217 = {1'h0, umul_57021[21:2]} + 21'h00_0fb9;
  assign sel_57222 = $signed({1'h0, smod_56955[15:0]}) < $signed({1'h0, sel_57028}) ? smod_56955[15:0] : sel_57028;
  assign umul_57223 = umul22b_16b_x_6b(array_index_57045, 6'h3b);
  assign add_57225 = {1'h0, umul_57029[21:1]} + 22'h00_1f59;
  assign sel_57230 = $signed({1'h0, smod_56960[15:0]}) < $signed({1'h0, sel_57036}) ? smod_56960[15:0] : sel_57036;
  assign umul_57231 = umul22b_16b_x_6b(array_index_57051, 6'h3b);
  assign add_57233 = {1'h0, umul_57037[21:1]} + 22'h00_1f59;
  assign sel_57238 = $signed({1'h0, smod_56965[15:0]}) < $signed({1'h0, sel_57044}) ? smod_56965[15:0] : sel_57044;
  assign array_index_57239 = set1_unflattened[5'h1c];
  assign smod_57243 = $unsigned($signed({9'h000, add_57107, umul_56911[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_57245 = set2_unflattened[5'h1c];
  assign smod_57249 = $unsigned($signed({9'h000, add_57115, umul_56919[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_57299 = umul22b_16b_x_6b(array_index_57239, 6'h35);
  assign add_57301 = {1'h0, umul_57105[21:7]} + 16'h007d;
  assign sel_57306 = $signed({1'h0, smod_57049[15:0]}) < $signed({1'h0, sel_57112}) ? smod_57049[15:0] : sel_57112;
  assign umul_57307 = umul22b_16b_x_6b(array_index_57245, 6'h35);
  assign add_57309 = {1'h0, umul_57113[21:7]} + 16'h007d;
  assign sel_57314 = $signed({1'h0, smod_57055[15:0]}) < $signed({1'h0, sel_57120}) ? smod_57055[15:0] : sel_57120;
  assign smod_57318 = $unsigned($signed({8'h00, add_57177, umul_56981[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57323 = $unsigned($signed({8'h00, add_57185, umul_56989[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57328 = $unsigned($signed({8'h00, add_57193, umul_56997[0]}) % $signed(32'h0000_3ffd));
  assign smod_57333 = $unsigned($signed({8'h00, add_57201, umul_57005[0]}) % $signed(32'h0000_3ffd));
  assign smod_57338 = $unsigned($signed({9'h000, add_57209, umul_57013[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57343 = $unsigned($signed({9'h000, add_57217, umul_57021[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57348 = $unsigned($signed({9'h000, add_57225, umul_57029[0]}) % $signed(32'h0000_3ffd));
  assign smod_57353 = $unsigned($signed({9'h000, add_57233, umul_57037[0]}) % $signed(32'h0000_3ffd));
  assign umul_57369 = umul23b_16b_x_7b(array_index_56657, 7'h49);
  assign add_57371 = {1'h0, umul_57175[22:3]} + 21'h00_07e9;
  assign sel_57376 = $signed({1'h0, smod_57124[15:0]}) < $signed({1'h0, sel_57182}) ? smod_57124[15:0] : sel_57182;
  assign umul_57377 = umul23b_16b_x_7b(array_index_56663, 7'h49);
  assign add_57379 = {1'h0, umul_57183[22:3]} + 21'h00_07e9;
  assign sel_57384 = $signed({1'h0, smod_57129[15:0]}) < $signed({1'h0, sel_57190}) ? smod_57129[15:0] : sel_57190;
  assign umul_57385 = umul23b_16b_x_7b(array_index_56851, 7'h47);
  assign add_57387 = {1'h0, umul_57191[22:1]} + 23'h00_1f8b;
  assign sel_57392 = $signed({1'h0, smod_57134[15:0]}) < $signed({1'h0, sel_57198}) ? smod_57134[15:0] : sel_57198;
  assign umul_57393 = umul23b_16b_x_7b(array_index_56857, 7'h47);
  assign add_57395 = {1'h0, umul_57199[22:1]} + 23'h00_1f8b;
  assign sel_57400 = $signed({1'h0, smod_57139[15:0]}) < $signed({1'h0, sel_57206}) ? smod_57139[15:0] : sel_57206;
  assign umul_57401 = umul22b_16b_x_6b(array_index_57045, 6'h3d);
  assign add_57403 = {1'h0, umul_57207[21:2]} + 21'h00_0fb9;
  assign sel_57408 = $signed({1'h0, smod_57144[15:0]}) < $signed({1'h0, sel_57214}) ? smod_57144[15:0] : sel_57214;
  assign umul_57409 = umul22b_16b_x_6b(array_index_57051, 6'h3d);
  assign add_57411 = {1'h0, umul_57215[21:2]} + 21'h00_0fb9;
  assign sel_57416 = $signed({1'h0, smod_57149[15:0]}) < $signed({1'h0, sel_57222}) ? smod_57149[15:0] : sel_57222;
  assign umul_57417 = umul22b_16b_x_6b(array_index_57239, 6'h3b);
  assign add_57419 = {1'h0, umul_57223[21:1]} + 22'h00_1f59;
  assign sel_57424 = $signed({1'h0, smod_57154[15:0]}) < $signed({1'h0, sel_57230}) ? smod_57154[15:0] : sel_57230;
  assign umul_57425 = umul22b_16b_x_6b(array_index_57245, 6'h3b);
  assign add_57427 = {1'h0, umul_57231[21:1]} + 22'h00_1f59;
  assign sel_57432 = $signed({1'h0, smod_57159[15:0]}) < $signed({1'h0, sel_57238}) ? smod_57159[15:0] : sel_57238;
  assign array_index_57433 = set1_unflattened[5'h1d];
  assign smod_57437 = $unsigned($signed({9'h000, add_57301, umul_57105[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_57439 = set2_unflattened[5'h1d];
  assign smod_57443 = $unsigned($signed({9'h000, add_57309, umul_57113[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_57493 = umul22b_16b_x_6b(array_index_57433, 6'h35);
  assign add_57495 = {1'h0, umul_57299[21:7]} + 16'h007d;
  assign sel_57500 = $signed({1'h0, smod_57243[15:0]}) < $signed({1'h0, sel_57306}) ? smod_57243[15:0] : sel_57306;
  assign umul_57501 = umul22b_16b_x_6b(array_index_57439, 6'h35);
  assign add_57503 = {1'h0, umul_57307[21:7]} + 16'h007d;
  assign sel_57508 = $signed({1'h0, smod_57249[15:0]}) < $signed({1'h0, sel_57314}) ? smod_57249[15:0] : sel_57314;
  assign smod_57512 = $unsigned($signed({8'h00, add_57371, umul_57175[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57517 = $unsigned($signed({8'h00, add_57379, umul_57183[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57522 = $unsigned($signed({8'h00, add_57387, umul_57191[0]}) % $signed(32'h0000_3ffd));
  assign smod_57527 = $unsigned($signed({8'h00, add_57395, umul_57199[0]}) % $signed(32'h0000_3ffd));
  assign smod_57532 = $unsigned($signed({9'h000, add_57403, umul_57207[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57537 = $unsigned($signed({9'h000, add_57411, umul_57215[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57542 = $unsigned($signed({9'h000, add_57419, umul_57223[0]}) % $signed(32'h0000_3ffd));
  assign smod_57547 = $unsigned($signed({9'h000, add_57427, umul_57231[0]}) % $signed(32'h0000_3ffd));
  assign umul_57561 = umul23b_16b_x_7b(array_index_56851, 7'h49);
  assign add_57563 = {1'h0, umul_57369[22:3]} + 21'h00_07e9;
  assign sel_57568 = $signed({1'h0, smod_57318[15:0]}) < $signed({1'h0, sel_57376}) ? smod_57318[15:0] : sel_57376;
  assign umul_57569 = umul23b_16b_x_7b(array_index_56857, 7'h49);
  assign add_57571 = {1'h0, umul_57377[22:3]} + 21'h00_07e9;
  assign sel_57576 = $signed({1'h0, smod_57323[15:0]}) < $signed({1'h0, sel_57384}) ? smod_57323[15:0] : sel_57384;
  assign umul_57577 = umul23b_16b_x_7b(array_index_57045, 7'h47);
  assign add_57579 = {1'h0, umul_57385[22:1]} + 23'h00_1f8b;
  assign sel_57584 = $signed({1'h0, smod_57328[15:0]}) < $signed({1'h0, sel_57392}) ? smod_57328[15:0] : sel_57392;
  assign umul_57585 = umul23b_16b_x_7b(array_index_57051, 7'h47);
  assign add_57587 = {1'h0, umul_57393[22:1]} + 23'h00_1f8b;
  assign sel_57592 = $signed({1'h0, smod_57333[15:0]}) < $signed({1'h0, sel_57400}) ? smod_57333[15:0] : sel_57400;
  assign umul_57593 = umul22b_16b_x_6b(array_index_57239, 6'h3d);
  assign add_57595 = {1'h0, umul_57401[21:2]} + 21'h00_0fb9;
  assign sel_57600 = $signed({1'h0, smod_57338[15:0]}) < $signed({1'h0, sel_57408}) ? smod_57338[15:0] : sel_57408;
  assign umul_57601 = umul22b_16b_x_6b(array_index_57245, 6'h3d);
  assign add_57603 = {1'h0, umul_57409[21:2]} + 21'h00_0fb9;
  assign sel_57608 = $signed({1'h0, smod_57343[15:0]}) < $signed({1'h0, sel_57416}) ? smod_57343[15:0] : sel_57416;
  assign umul_57609 = umul22b_16b_x_6b(array_index_57433, 6'h3b);
  assign add_57611 = {1'h0, umul_57417[21:1]} + 22'h00_1f59;
  assign sel_57616 = $signed({1'h0, smod_57348[15:0]}) < $signed({1'h0, sel_57424}) ? smod_57348[15:0] : sel_57424;
  assign umul_57617 = umul22b_16b_x_6b(array_index_57439, 6'h3b);
  assign add_57619 = {1'h0, umul_57425[21:1]} + 22'h00_1f59;
  assign sel_57624 = $signed({1'h0, smod_57353[15:0]}) < $signed({1'h0, sel_57432}) ? smod_57353[15:0] : sel_57432;
  assign smod_57627 = $unsigned($signed({9'h000, add_57495, umul_57299[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_57631 = $unsigned($signed({9'h000, add_57503, umul_57307[6:0]}) % $signed(32'h0000_3ffd));
  assign add_57682 = {1'h0, umul_57493[21:7]} + 16'h007d;
  assign sel_57687 = $signed({1'h0, smod_57437[15:0]}) < $signed({1'h0, sel_57500}) ? smod_57437[15:0] : sel_57500;
  assign add_57689 = {1'h0, umul_57501[21:7]} + 16'h007d;
  assign sel_57694 = $signed({1'h0, smod_57443[15:0]}) < $signed({1'h0, sel_57508}) ? smod_57443[15:0] : sel_57508;
  assign smod_57698 = $unsigned($signed({8'h00, add_57563, umul_57369[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57703 = $unsigned($signed({8'h00, add_57571, umul_57377[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57708 = $unsigned($signed({8'h00, add_57579, umul_57385[0]}) % $signed(32'h0000_3ffd));
  assign smod_57713 = $unsigned($signed({8'h00, add_57587, umul_57393[0]}) % $signed(32'h0000_3ffd));
  assign smod_57718 = $unsigned($signed({9'h000, add_57595, umul_57401[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57723 = $unsigned($signed({9'h000, add_57603, umul_57409[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57727 = $unsigned($signed({9'h000, add_57611, umul_57417[0]}) % $signed(32'h0000_3ffd));
  assign smod_57731 = $unsigned($signed({9'h000, add_57619, umul_57425[0]}) % $signed(32'h0000_3ffd));
  assign umul_57741 = umul23b_16b_x_7b(array_index_57045, 7'h49);
  assign add_57743 = {1'h0, umul_57561[22:3]} + 21'h00_07e9;
  assign sel_57748 = $signed({1'h0, smod_57512[15:0]}) < $signed({1'h0, sel_57568}) ? smod_57512[15:0] : sel_57568;
  assign umul_57749 = umul23b_16b_x_7b(array_index_57051, 7'h49);
  assign add_57751 = {1'h0, umul_57569[22:3]} + 21'h00_07e9;
  assign sel_57756 = $signed({1'h0, smod_57517[15:0]}) < $signed({1'h0, sel_57576}) ? smod_57517[15:0] : sel_57576;
  assign umul_57757 = umul23b_16b_x_7b(array_index_57239, 7'h47);
  assign add_57759 = {1'h0, umul_57577[22:1]} + 23'h00_1f8b;
  assign sel_57764 = $signed({1'h0, smod_57522[15:0]}) < $signed({1'h0, sel_57584}) ? smod_57522[15:0] : sel_57584;
  assign umul_57765 = umul23b_16b_x_7b(array_index_57245, 7'h47);
  assign add_57767 = {1'h0, umul_57585[22:1]} + 23'h00_1f8b;
  assign sel_57772 = $signed({1'h0, smod_57527[15:0]}) < $signed({1'h0, sel_57592}) ? smod_57527[15:0] : sel_57592;
  assign umul_57773 = umul22b_16b_x_6b(array_index_57433, 6'h3d);
  assign add_57775 = {1'h0, umul_57593[21:2]} + 21'h00_0fb9;
  assign sel_57780 = $signed({1'h0, smod_57532[15:0]}) < $signed({1'h0, sel_57600}) ? smod_57532[15:0] : sel_57600;
  assign umul_57781 = umul22b_16b_x_6b(array_index_57439, 6'h3d);
  assign add_57783 = {1'h0, umul_57601[21:2]} + 21'h00_0fb9;
  assign sel_57788 = $signed({1'h0, smod_57537[15:0]}) < $signed({1'h0, sel_57608}) ? smod_57537[15:0] : sel_57608;
  assign add_57790 = {1'h0, umul_57609[21:1]} + 22'h00_1f59;
  assign sel_57795 = $signed({1'h0, smod_57542[15:0]}) < $signed({1'h0, sel_57616}) ? smod_57542[15:0] : sel_57616;
  assign add_57797 = {1'h0, umul_57617[21:1]} + 22'h00_1f59;
  assign sel_57802 = $signed({1'h0, smod_57547[15:0]}) < $signed({1'h0, sel_57624}) ? smod_57547[15:0] : sel_57624;
  assign smod_57803 = $unsigned($signed({9'h000, add_57682, umul_57493[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_57805 = $unsigned($signed({9'h000, add_57689, umul_57501[6:0]}) % $signed(32'h0000_3ffd));
  assign sel_57854 = $signed({1'h0, smod_57627[15:0]}) < $signed({1'h0, sel_57687}) ? smod_57627[15:0] : sel_57687;
  assign sel_57858 = $signed({1'h0, smod_57631[15:0]}) < $signed({1'h0, sel_57694}) ? smod_57631[15:0] : sel_57694;
  assign smod_57862 = $unsigned($signed({8'h00, add_57743, umul_57561[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57867 = $unsigned($signed({8'h00, add_57751, umul_57569[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57872 = $unsigned($signed({8'h00, add_57759, umul_57577[0]}) % $signed(32'h0000_3ffd));
  assign smod_57877 = $unsigned($signed({8'h00, add_57767, umul_57585[0]}) % $signed(32'h0000_3ffd));
  assign smod_57881 = $unsigned($signed({9'h000, add_57775, umul_57593[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57885 = $unsigned($signed({9'h000, add_57783, umul_57601[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_57887 = $unsigned($signed({9'h000, add_57790, umul_57609[0]}) % $signed(32'h0000_3ffd));
  assign smod_57889 = $unsigned($signed({9'h000, add_57797, umul_57617[0]}) % $signed(32'h0000_3ffd));
  assign umul_57895 = umul23b_16b_x_7b(array_index_57239, 7'h49);
  assign add_57897 = {1'h0, umul_57741[22:3]} + 21'h00_07e9;
  assign sel_57902 = $signed({1'h0, smod_57698[15:0]}) < $signed({1'h0, sel_57748}) ? smod_57698[15:0] : sel_57748;
  assign umul_57903 = umul23b_16b_x_7b(array_index_57245, 7'h49);
  assign add_57905 = {1'h0, umul_57749[22:3]} + 21'h00_07e9;
  assign sel_57910 = $signed({1'h0, smod_57703[15:0]}) < $signed({1'h0, sel_57756}) ? smod_57703[15:0] : sel_57756;
  assign umul_57911 = umul23b_16b_x_7b(array_index_57433, 7'h47);
  assign add_57913 = {1'h0, umul_57757[22:1]} + 23'h00_1f8b;
  assign sel_57918 = $signed({1'h0, smod_57708[15:0]}) < $signed({1'h0, sel_57764}) ? smod_57708[15:0] : sel_57764;
  assign umul_57919 = umul23b_16b_x_7b(array_index_57439, 7'h47);
  assign add_57921 = {1'h0, umul_57765[22:1]} + 23'h00_1f8b;
  assign sel_57926 = $signed({1'h0, smod_57713[15:0]}) < $signed({1'h0, sel_57772}) ? smod_57713[15:0] : sel_57772;
  assign add_57928 = {1'h0, umul_57773[21:2]} + 21'h00_0fb9;
  assign sel_57933 = $signed({1'h0, smod_57718[15:0]}) < $signed({1'h0, sel_57780}) ? smod_57718[15:0] : sel_57780;
  assign add_57935 = {1'h0, umul_57781[21:2]} + 21'h00_0fb9;
  assign sel_57940 = $signed({1'h0, smod_57723[15:0]}) < $signed({1'h0, sel_57788}) ? smod_57723[15:0] : sel_57788;
  assign sel_57944 = $signed({1'h0, smod_57727[15:0]}) < $signed({1'h0, sel_57795}) ? smod_57727[15:0] : sel_57795;
  assign sel_57948 = $signed({1'h0, smod_57731[15:0]}) < $signed({1'h0, sel_57802}) ? smod_57731[15:0] : sel_57802;
  assign smod_57992 = $unsigned($signed({8'h00, add_57897, umul_57741[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_57997 = $unsigned($signed({8'h00, add_57905, umul_57749[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_58001 = $unsigned($signed({8'h00, add_57913, umul_57757[0]}) % $signed(32'h0000_3ffd));
  assign smod_58005 = $unsigned($signed({8'h00, add_57921, umul_57765[0]}) % $signed(32'h0000_3ffd));
  assign smod_58007 = $unsigned($signed({9'h000, add_57928, umul_57773[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_58009 = $unsigned($signed({9'h000, add_57935, umul_57781[1:0]}) % $signed(32'h0000_3ffd));
  assign umul_58015 = umul23b_16b_x_7b(array_index_57433, 7'h49);
  assign add_58017 = {1'h0, umul_57895[22:3]} + 21'h00_07e9;
  assign sel_58022 = $signed({1'h0, smod_57862[15:0]}) < $signed({1'h0, sel_57902}) ? smod_57862[15:0] : sel_57902;
  assign umul_58023 = umul23b_16b_x_7b(array_index_57439, 7'h49);
  assign add_58025 = {1'h0, umul_57903[22:3]} + 21'h00_07e9;
  assign sel_58030 = $signed({1'h0, smod_57867[15:0]}) < $signed({1'h0, sel_57910}) ? smod_57867[15:0] : sel_57910;
  assign add_58032 = {1'h0, umul_57911[22:1]} + 23'h00_1f8b;
  assign sel_58037 = $signed({1'h0, smod_57872[15:0]}) < $signed({1'h0, sel_57918}) ? smod_57872[15:0] : sel_57918;
  assign add_58039 = {1'h0, umul_57919[22:1]} + 23'h00_1f8b;
  assign sel_58044 = $signed({1'h0, smod_57877[15:0]}) < $signed({1'h0, sel_57926}) ? smod_57877[15:0] : sel_57926;
  assign sel_58048 = $signed({1'h0, smod_57881[15:0]}) < $signed({1'h0, sel_57933}) ? smod_57881[15:0] : sel_57933;
  assign sel_58052 = $signed({1'h0, smod_57885[15:0]}) < $signed({1'h0, sel_57940}) ? smod_57885[15:0] : sel_57940;
  assign concat_58055 = {1'h0, ($signed({1'h0, smod_57803[15:0]}) < $signed({1'h0, sel_57854}) ? smod_57803[15:0] : sel_57854) == ($signed({1'h0, smod_57805[15:0]}) < $signed({1'h0, sel_57858}) ? smod_57805[15:0] : sel_57858)};
  assign add_58082 = concat_58055 + 2'h1;
  assign smod_58085 = $unsigned($signed({8'h00, add_58017, umul_57895[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_58089 = $unsigned($signed({8'h00, add_58025, umul_57903[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_58091 = $unsigned($signed({8'h00, add_58032, umul_57911[0]}) % $signed(32'h0000_3ffd));
  assign smod_58093 = $unsigned($signed({8'h00, add_58039, umul_57919[0]}) % $signed(32'h0000_3ffd));
  assign add_58100 = {1'h0, umul_58015[22:3]} + 21'h00_07e9;
  assign sel_58105 = $signed({1'h0, smod_57992[15:0]}) < $signed({1'h0, sel_58022}) ? smod_57992[15:0] : sel_58022;
  assign add_58107 = {1'h0, umul_58023[22:3]} + 21'h00_07e9;
  assign sel_58112 = $signed({1'h0, smod_57997[15:0]}) < $signed({1'h0, sel_58030}) ? smod_57997[15:0] : sel_58030;
  assign sel_58116 = $signed({1'h0, smod_58001[15:0]}) < $signed({1'h0, sel_58037}) ? smod_58001[15:0] : sel_58037;
  assign sel_58120 = $signed({1'h0, smod_58005[15:0]}) < $signed({1'h0, sel_58044}) ? smod_58005[15:0] : sel_58044;
  assign concat_58123 = {1'h0, ($signed({1'h0, smod_57887[15:0]}) < $signed({1'h0, sel_57944}) ? smod_57887[15:0] : sel_57944) == ($signed({1'h0, smod_57889[15:0]}) < $signed({1'h0, sel_57948}) ? smod_57889[15:0] : sel_57948) ? add_58082 : concat_58055};
  assign add_58138 = concat_58123 + 3'h1;
  assign smod_58139 = $unsigned($signed({8'h00, add_58100, umul_58015[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_58141 = $unsigned($signed({8'h00, add_58107, umul_58023[2:0]}) % $signed(32'h0000_3ffd));
  assign sel_58150 = $signed({1'h0, smod_58085[15:0]}) < $signed({1'h0, sel_58105}) ? smod_58085[15:0] : sel_58105;
  assign sel_58154 = $signed({1'h0, smod_58089[15:0]}) < $signed({1'h0, sel_58112}) ? smod_58089[15:0] : sel_58112;
  assign concat_58157 = {1'h0, ($signed({1'h0, smod_58007[15:0]}) < $signed({1'h0, sel_58048}) ? smod_58007[15:0] : sel_58048) == ($signed({1'h0, smod_58009[15:0]}) < $signed({1'h0, sel_58052}) ? smod_58009[15:0] : sel_58052) ? add_58138 : concat_58123};
  assign add_58164 = concat_58157 + 4'h1;
  assign concat_58171 = {1'h0, ($signed({1'h0, smod_58091[15:0]}) < $signed({1'h0, sel_58116}) ? smod_58091[15:0] : sel_58116) == ($signed({1'h0, smod_58093[15:0]}) < $signed({1'h0, sel_58120}) ? smod_58093[15:0] : sel_58120) ? add_58164 : concat_58157};
  assign add_58174 = concat_58171 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, smod_58139[15:0]}) < $signed({1'h0, sel_58150}) ? smod_58139[15:0] : sel_58150) == ($signed({1'h0, smod_58141[15:0]}) < $signed({1'h0, sel_58154}) ? smod_58141[15:0] : sel_58154) ? add_58174 : concat_58171}, {set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
