module min_hash(set1, set2, out);
  wire _00000_, _00001_, _00002_, _00003_, _00004_, _00005_, _00006_, _00007_, _00008_, _00009_, _00010_, _00011_, _00012_, _00013_, _00014_, _00015_, _00016_, _00017_, _00018_, _00019_, _00020_, _00021_, _00022_, _00023_, _00024_, _00025_, _00026_, _00027_, _00028_, _00029_, _00030_, _00031_, _00032_, _00033_, _00034_, _00035_, _00036_, _00037_, _00038_, _00039_, _00040_, _00041_, _00042_, _00043_, _00044_, _00045_, _00046_, _00047_, _00048_, _00049_, _00050_, _00051_, _00052_, _00053_, _00054_, _00055_, _00056_, _00057_, _00058_, _00059_, _00060_, _00061_, _00062_, _00063_, _00064_, _00065_, _00066_, _00067_, _00068_, _00069_, _00070_, _00071_, _00072_, _00073_, _00074_, _00075_, _00076_, _00077_, _00078_, _00079_, _00080_, _00081_, _00082_, _00083_, _00084_, _00085_, _00086_, _00087_, _00088_, _00089_, _00090_, _00091_, _00092_, _00093_, _00094_, _00095_, _00096_, _00097_, _00098_, _00099_, _00100_, _00101_, _00102_, _00103_, _00104_, _00105_, _00106_, _00107_, _00108_, _00109_, _00110_, _00111_, _00112_, _00113_, _00114_, _00115_, _00116_, _00117_, _00118_, _00119_, _00120_, _00121_, _00122_, _00123_, _00124_, _00125_, _00126_, _00127_, _00128_, _00129_, _00130_, _00131_, _00132_, _00133_, _00134_, _00135_, _00136_, _00137_, _00138_, _00139_, _00140_, _00141_, _00142_, _00143_, _00144_, _00145_, _00146_, _00147_, _00148_, _00149_, _00150_, _00151_, _00152_, _00153_, _00154_, _00155_, _00156_, _00157_, _00158_, _00159_, _00160_, _00161_, _00162_, _00163_, _00164_, _00165_, _00166_, _00167_, _00168_, _00169_, _00170_, _00171_, _00172_, _00173_, _00174_, _00175_, _00176_, _00177_, _00178_, _00179_, _00180_, _00181_, _00182_, _00183_, _00184_, _00185_, _00186_, _00187_, _00188_, _00189_, _00190_, _00191_, _00192_, _00193_, _00194_, _00195_, _00196_, _00197_, _00198_, _00199_, _00200_, _00201_, _00202_, _00203_, _00204_, _00205_, _00206_, _00207_, _00208_, _00209_, _00210_, _00211_, _00212_, _00213_, _00214_, _00215_, _00216_, _00217_, _00218_, _00219_, _00220_, _00221_, _00222_, _00223_, _00224_, _00225_, _00226_, _00227_, _00228_, _00229_, _00230_, _00231_, _00232_, _00233_, _00234_, _00235_, _00236_, _00237_, _00238_, _00239_, _00240_, _00241_, _00242_, _00243_, _00244_, _00245_, _00246_, _00247_, _00248_, _00249_, _00250_, _00251_, _00252_, _00253_, _00254_, _00255_, _00256_, _00257_, _00258_, _00259_, _00260_, _00261_, _00262_, _00263_, _00264_, _00265_, _00266_, _00267_, _00268_, _00269_, _00270_, _00271_, _00272_, _00273_, _00274_, _00275_, _00276_, _00277_, _00278_, _00279_, _00280_, _00281_, _00282_, _00283_, _00284_, _00285_, _00286_, _00287_, _00288_, _00289_, _00290_, _00291_, _00292_, _00293_, _00294_, _00295_, _00296_, _00297_, _00298_, _00299_, _00300_, _00301_, _00302_, _00303_, _00304_, _00305_, _00306_, _00307_, _00308_, _00309_, _00310_, _00311_, _00312_, _00313_, _00314_, _00315_, _00316_, _00317_, _00318_, _00319_, _00320_, _00321_, _00322_, _00323_, _00324_, _00325_, _00326_, _00327_, _00328_, _00329_, _00330_, _00331_, _00332_, _00333_, _00334_, _00335_, _00336_, _00337_, _00338_, _00339_, _00340_, _00341_, _00342_, _00343_, _00344_, _00345_, _00346_, _00347_, _00348_, _00349_, _00350_, _00351_, _00352_, _00353_, _00354_, _00355_, _00356_, _00357_, _00358_, _00359_, _00360_, _00361_, _00362_, _00363_, _00364_, _00365_, _00366_, _00367_, _00368_, _00369_, _00370_, _00371_, _00372_, _00373_, _00374_, _00375_, _00376_, _00377_, _00378_, _00379_, _00380_, _00381_, _00382_, _00383_, _00384_, _00385_, _00386_, _00387_, _00388_, _00389_, _00390_, _00391_, _00392_, _00393_, _00394_, _00395_, _00396_, _00397_, _00398_, _00399_, _00400_, _00401_, _00402_, _00403_, _00404_, _00405_, _00406_, _00407_, _00408_, _00409_, _00410_, _00411_, _00412_, _00413_, _00414_, _00415_, _00416_, _00417_, _00418_, _00419_, _00420_, _00421_, _00422_, _00423_, _00424_, _00425_, _00426_, _00427_, _00428_, _00429_, _00430_, _00431_, _00432_, _00433_, _00434_, _00435_, _00436_, _00437_, _00438_, _00439_, _00440_, _00441_, _00442_, _00443_, _00444_, _00445_, _00446_, _00447_, _00448_, _00449_, _00450_, _00451_, _00452_, _00453_, _00454_, _00455_, _00456_, _00457_, _00458_, _00459_, _00460_, _00461_, _00462_, _00463_, _00464_, _00465_, _00466_, _00467_, _00468_, _00469_, _00470_, _00471_, _00472_, _00473_, _00474_, _00475_, _00476_, _00477_, _00478_, _00479_, _00480_, _00481_, _00482_, _00483_, _00484_, _00485_, _00486_, _00487_, _00488_, _00489_, _00490_, _00491_, _00492_, _00493_, _00494_, _00495_, _00496_, _00497_, _00498_, _00499_, _00500_, _00501_, _00502_, _00503_, _00504_, _00505_, _00506_, _00507_, _00508_, _00509_, _00510_, _00511_, _00512_, _00513_, _00514_, _00515_, _00516_, _00517_, _00518_, _00519_, _00520_, _00521_, _00522_, _00523_, _00524_, _00525_, _00526_, _00527_, _00528_, _00529_, _00530_, _00531_, _00532_, _00533_, _00534_, _00535_, _00536_, _00537_, _00538_, _00539_, _00540_, _00541_, _00542_, _00543_, _00544_, _00545_, _00546_, _00547_, _00548_, _00549_, _00550_, _00551_, _00552_, _00553_, _00554_, _00555_, _00556_, _00557_, _00558_, _00559_, _00560_, _00561_, _00562_, _00563_, _00564_, _00565_, _00566_, _00567_, _00568_, _00569_, _00570_, _00571_, _00572_, _00573_, _00574_, _00575_, _00576_, _00577_, _00578_, _00579_, _00580_, _00581_, _00582_, _00583_, _00584_, _00585_, _00586_, _00587_, _00588_, _00589_, _00590_, _00591_, _00592_, _00593_, _00594_, _00595_, _00596_, _00597_, _00598_, _00599_, _00600_, _00601_, _00602_, _00603_, _00604_, _00605_, _00606_, _00607_, _00608_, _00609_, _00610_, _00611_, _00612_, _00613_, _00614_, _00615_, _00616_, _00617_, _00618_, _00619_, _00620_, _00621_, _00622_, _00623_, _00624_, _00625_, _00626_, _00627_, _00628_, _00629_, _00630_, _00631_, _00632_, _00633_, _00634_, _00635_, _00636_, _00637_, _00638_, _00639_, _00640_, _00641_, _00642_, _00643_, _00644_, _00645_, _00646_, _00647_, _00648_, _00649_, _00650_, _00651_, _00652_, _00653_, _00654_, _00655_, _00656_, _00657_, _00658_, _00659_, _00660_, _00661_, _00662_, _00663_, _00664_, _00665_, _00666_, _00667_, _00668_, _00669_, _00670_, _00671_, _00672_, _00673_, _00674_, _00675_, _00676_, _00677_, _00678_, _00679_, _00680_, _00681_, _00682_, _00683_, _00684_, _00685_, _00686_, _00687_, _00688_, _00689_, _00690_, _00691_, _00692_, _00693_, _00694_, _00695_, _00696_, _00697_, _00698_, _00699_, _00700_, _00701_, _00702_, _00703_, _00704_, _00705_, _00706_, _00707_, _00708_, _00709_, _00710_, _00711_, _00712_, _00713_, _00714_, _00715_, _00716_, _00717_, _00718_, _00719_, _00720_, _00721_, _00722_, _00723_, _00724_, _00725_, _00726_, _00727_, _00728_, _00729_, _00730_, _00731_, _00732_, _00733_, _00734_, _00735_, _00736_, _00737_, _00738_, _00739_, _00740_, _00741_, _00742_, _00743_, _00744_, _00745_, _00746_, _00747_, _00748_, _00749_, _00750_, _00751_, _00752_, _00753_, _00754_, _00755_, _00756_, _00757_, _00758_, _00759_, _00760_, _00761_, _00762_, _00763_, _00764_, _00765_, _00766_, _00767_, _00768_, _00769_, _00770_, _00771_, _00772_, _00773_, _00774_, _00775_, _00776_, _00777_, _00778_, _00779_, _00780_, _00781_, _00782_, _00783_, _00784_, _00785_, _00786_, _00787_, _00788_, _00789_, _00790_, _00791_, _00792_, _00793_, _00794_, _00795_, _00796_, _00797_, _00798_, _00799_, _00800_, _00801_, _00802_, _00803_, _00804_, _00805_, _00806_, _00807_, _00808_, _00809_, _00810_, _00811_, _00812_, _00813_, _00814_, _00815_, _00816_, _00817_, _00818_, _00819_, _00820_, _00821_, _00822_, _00823_, _00824_, _00825_, _00826_, _00827_, _00828_, _00829_, _00830_, _00831_, _00832_, _00833_, _00834_, _00835_, _00836_, _00837_, _00838_, _00839_, _00840_, _00841_, _00842_, _00843_, _00844_, _00845_, _00846_, _00847_, _00848_, _00849_, _00850_, _00851_, _00852_, _00853_, _00854_, _00855_, _00856_, _00857_, _00858_, _00859_, _00860_, _00861_, _00862_, _00863_, _00864_, _00865_, _00866_, _00867_, _00868_, _00869_, _00870_, _00871_, _00872_, _00873_, _00874_, _00875_, _00876_, _00877_, _00878_, _00879_, _00880_, _00881_, _00882_, _00883_, _00884_, _00885_, _00886_, _00887_, _00888_, _00889_, _00890_, _00891_, _00892_, _00893_, _00894_, _00895_, _00896_, _00897_, _00898_, _00899_, _00900_, _00901_, _00902_, _00903_, _00904_, _00905_, _00906_, _00907_, _00908_, _00909_, _00910_, _00911_, _00912_, _00913_, _00914_, _00915_, _00916_, _00917_, _00918_, _00919_, _00920_, _00921_, _00922_, _00923_, _00924_, _00925_, _00926_, _00927_, _00928_, _00929_, _00930_, _00931_, _00932_, _00933_, _00934_, _00935_, _00936_, _00937_, _00938_, _00939_, _00940_, _00941_, _00942_, _00943_, _00944_, _00945_, _00946_, _00947_, _00948_, _00949_, _00950_, _00951_, _00952_, _00953_, _00954_, _00955_, _00956_, _00957_, _00958_, _00959_, _00960_, _00961_, _00962_, _00963_, _00964_, _00965_, _00966_, _00967_, _00968_, _00969_, _00970_, _00971_, _00972_, _00973_, _00974_, _00975_, _00976_, _00977_, _00978_, _00979_, _00980_, _00981_, _00982_, _00983_, _00984_, _00985_, _00986_, _00987_, _00988_, _00989_, _00990_, _00991_, _00992_, _00993_, _00994_, _00995_, _00996_, _00997_, _00998_, _00999_, _01000_, _01001_, _01002_, _01003_, _01004_, _01005_, _01006_, _01007_, _01008_, _01009_, _01010_, _01011_, _01012_, _01013_, _01014_, _01015_, _01016_, _01017_, _01018_, _01019_, _01020_, _01021_, _01022_, _01023_, _01024_, _01025_, _01026_, _01027_, _01028_, _01029_, _01030_, _01031_, _01032_, _01033_, _01034_, _01035_, _01036_, _01037_, _01038_, _01039_, _01040_, _01041_, _01042_, _01043_, _01044_, _01045_, _01046_, _01047_, _01048_, _01049_, _01050_, _01051_, _01052_, _01053_, _01054_, _01055_, _01056_, _01057_, _01058_, _01059_, _01060_, _01061_, _01062_, _01063_, _01064_, _01065_, _01066_, _01067_, _01068_, _01069_, _01070_, _01071_, _01072_, _01073_, _01074_, _01075_, _01076_, _01077_, _01078_, _01079_, _01080_, _01081_, _01082_, _01083_, _01084_, _01085_, _01086_, _01087_, _01088_, _01089_, _01090_, _01091_, _01092_, _01093_, _01094_, _01095_, _01096_, _01097_, _01098_, _01099_, _01100_, _01101_, _01102_, _01103_, _01104_, _01105_, _01106_, _01107_, _01108_, _01109_, _01110_, _01111_, _01112_, _01113_, _01114_, _01115_, _01116_, _01117_, _01118_, _01119_, _01120_, _01121_, _01122_, _01123_, _01124_, _01125_, _01126_, _01127_, _01128_, _01129_, _01130_, _01131_, _01132_, _01133_, _01134_, _01135_, _01136_, _01137_, _01138_, _01139_, _01140_, _01141_, _01142_, _01143_, _01144_, _01145_, _01146_, _01147_, _01148_, _01149_, _01150_, _01151_, _01152_, _01153_, _01154_, _01155_, _01156_, _01157_, _01158_, _01159_, _01160_, _01161_, _01162_, _01163_, _01164_, _01165_, _01166_, _01167_, _01168_, _01169_, _01170_, _01171_, _01172_, _01173_, _01174_, _01175_, _01176_, _01177_, _01178_, _01179_, _01180_, _01181_, _01182_, _01183_, _01184_, _01185_, _01186_, _01187_, _01188_, _01189_, _01190_, _01191_, _01192_, _01193_, _01194_, _01195_, _01196_, _01197_, _01198_, _01199_, _01200_, _01201_, _01202_, _01203_, _01204_, _01205_, _01206_, _01207_, _01208_, _01209_, _01210_, _01211_, _01212_, _01213_, _01214_, _01215_, _01216_, _01217_, _01218_, _01219_, _01220_, _01221_, _01222_, _01223_, _01224_, _01225_, _01226_, _01227_, _01228_, _01229_, _01230_, _01231_, _01232_, _01233_, _01234_, _01235_, _01236_, _01237_, _01238_, _01239_, _01240_, _01241_, _01242_, _01243_, _01244_, _01245_, _01246_, _01247_, _01248_, _01249_, _01250_, _01251_, _01252_, _01253_, _01254_, _01255_, _01256_, _01257_, _01258_, _01259_, _01260_, _01261_, _01262_, _01263_, _01264_, _01265_, _01266_, _01267_, _01268_, _01269_, _01270_, _01271_, _01272_, _01273_, _01274_, _01275_, _01276_, _01277_, _01278_, _01279_, _01280_, _01281_, _01282_, _01283_, _01284_, _01285_, _01286_, _01287_, _01288_, _01289_, _01290_, _01291_, _01292_, _01293_, _01294_, _01295_, _01296_, _01297_, _01298_, _01299_, _01300_, _01301_, _01302_, _01303_, _01304_, _01305_, _01306_, _01307_, _01308_, _01309_, _01310_, _01311_, _01312_, _01313_, _01314_, _01315_, _01316_, _01317_, _01318_, _01319_, _01320_, _01321_, _01322_, _01323_, _01324_, _01325_, _01326_, _01327_, _01328_, _01329_, _01330_, _01331_, _01332_, _01333_, _01334_, _01335_, _01336_, _01337_, _01338_, _01339_, _01340_, _01341_, _01342_, _01343_, _01344_, _01345_, _01346_, _01347_, _01348_, _01349_, _01350_, _01351_, _01352_, _01353_, _01354_, _01355_, _01356_, _01357_, _01358_, _01359_, _01360_, _01361_, _01362_, _01363_, _01364_, _01365_, _01366_, _01367_, _01368_, _01369_, _01370_, _01371_, _01372_, _01373_, _01374_, _01375_, _01376_, _01377_, _01378_, _01379_, _01380_, _01381_, _01382_, _01383_, _01384_, _01385_, _01386_, _01387_, _01388_, _01389_, _01390_, _01391_, _01392_, _01393_, _01394_, _01395_, _01396_, _01397_, _01398_, _01399_, _01400_, _01401_, _01402_, _01403_, _01404_, _01405_, _01406_, _01407_, _01408_, _01409_, _01410_, _01411_, _01412_, _01413_, _01414_, _01415_, _01416_, _01417_, _01418_, _01419_, _01420_, _01421_, _01422_, _01423_, _01424_, _01425_, _01426_, _01427_, _01428_, _01429_, _01430_, _01431_, _01432_, _01433_, _01434_, _01435_, _01436_, _01437_, _01438_, _01439_, _01440_, _01441_, _01442_, _01443_, _01444_, _01445_, _01446_, _01447_, _01448_, _01449_, _01450_, _01451_, _01452_, _01453_, _01454_, _01455_, _01456_, _01457_, _01458_, _01459_, _01460_, _01461_, _01462_, _01463_, _01464_, _01465_, _01466_, _01467_, _01468_, _01469_, _01470_, _01471_, _01472_, _01473_, _01474_, _01475_, _01476_, _01477_, _01478_, _01479_, _01480_, _01481_, _01482_, _01483_, _01484_, _01485_, _01486_, _01487_, _01488_, _01489_, _01490_, _01491_, _01492_, _01493_, _01494_, _01495_, _01496_, _01497_, _01498_, _01499_, _01500_, _01501_, _01502_, _01503_, _01504_, _01505_, _01506_, _01507_, _01508_, _01509_, _01510_, _01511_, _01512_, _01513_, _01514_, _01515_, _01516_, _01517_, _01518_, _01519_, _01520_, _01521_, _01522_, _01523_, _01524_, _01525_, _01526_, _01527_, _01528_, _01529_, _01530_, _01531_, _01532_, _01533_, _01534_, _01535_, _01536_, _01537_, _01538_, _01539_, _01540_, _01541_, _01542_, _01543_, _01544_, _01545_, _01546_, _01547_, _01548_, _01549_, _01550_, _01551_, _01552_, _01553_, _01554_, _01555_, _01556_, _01557_, _01558_, _01559_, _01560_, _01561_, _01562_, _01563_, _01564_, _01565_, _01566_, _01567_, _01568_, _01569_, _01570_, _01571_, _01572_, _01573_, _01574_, _01575_, _01576_, _01577_, _01578_, _01579_, _01580_, _01581_, _01582_, _01583_, _01584_, _01585_, _01586_, _01587_, _01588_, _01589_, _01590_, _01591_, _01592_, _01593_, _01594_, _01595_, _01596_, _01597_, _01598_, _01599_, _01600_, _01601_, _01602_, _01603_, _01604_, _01605_, _01606_, _01607_, _01608_, _01609_, _01610_, _01611_, _01612_, _01613_, _01614_, _01615_, _01616_, _01617_, _01618_, _01619_, _01620_, _01621_, _01622_, _01623_, _01624_, _01625_, _01626_, _01627_, _01628_, _01629_, _01630_, _01631_, _01632_, _01633_, _01634_, _01635_, _01636_, _01637_, _01638_, _01639_, _01640_, _01641_, _01642_, _01643_, _01644_, _01645_, _01646_, _01647_, _01648_, _01649_, _01650_, _01651_, _01652_, _01653_, _01654_, _01655_, _01656_, _01657_, _01658_, _01659_, _01660_, _01661_, _01662_, _01663_, _01664_, _01665_, _01666_, _01667_, _01668_, _01669_, _01670_, _01671_, _01672_, _01673_, _01674_, _01675_, _01676_, _01677_, _01678_, _01679_, _01680_, _01681_, _01682_, _01683_, _01684_, _01685_, _01686_, _01687_, _01688_, _01689_, _01690_, _01691_, _01692_, _01693_, _01694_, _01695_, _01696_, _01697_, _01698_, _01699_, _01700_, _01701_, _01702_, _01703_, _01704_, _01705_, _01706_, _01707_, _01708_, _01709_, _01710_, _01711_, _01712_, _01713_, _01714_, _01715_, _01716_, _01717_, _01718_, _01719_, _01720_, _01721_, _01722_, _01723_, _01724_, _01725_, _01726_, _01727_, _01728_, _01729_, _01730_, _01731_, _01732_, _01733_, _01734_, _01735_, _01736_, _01737_, _01738_, _01739_, _01740_, _01741_, _01742_, _01743_, _01744_, _01745_, _01746_, _01747_, _01748_, _01749_, _01750_, _01751_, _01752_, _01753_, _01754_, _01755_, _01756_, _01757_, _01758_, _01759_, _01760_, _01761_, _01762_, _01763_, _01764_, _01765_, _01766_, _01767_, _01768_, _01769_, _01770_, _01771_, _01772_, _01773_, _01774_, _01775_, _01776_, _01777_, _01778_, _01779_, _01780_, _01781_, _01782_, _01783_, _01784_, _01785_, _01786_, _01787_, _01788_, _01789_, _01790_, _01791_, _01792_, _01793_, _01794_, _01795_, _01796_, _01797_, _01798_, _01799_, _01800_, _01801_, _01802_, _01803_, _01804_, _01805_, _01806_, _01807_, _01808_, _01809_, _01810_, _01811_, _01812_, _01813_, _01814_, _01815_, _01816_, _01817_, _01818_, _01819_, _01820_, _01821_, _01822_, _01823_, _01824_, _01825_, _01826_, _01827_, _01828_, _01829_, _01830_, _01831_, _01832_, _01833_, _01834_, _01835_, _01836_, _01837_, _01838_, _01839_, _01840_, _01841_, _01842_, _01843_, _01844_, _01845_, _01846_, _01847_, _01848_, _01849_, _01850_, _01851_, _01852_, _01853_, _01854_, _01855_, _01856_, _01857_, _01858_, _01859_, _01860_, _01861_, _01862_, _01863_, _01864_, _01865_, _01866_, _01867_, _01868_, _01869_, _01870_, _01871_, _01872_, _01873_, _01874_, _01875_, _01876_, _01877_, _01878_, _01879_, _01880_, _01881_, _01882_, _01883_, _01884_, _01885_, _01886_, _01887_, _01888_, _01889_, _01890_, _01891_, _01892_, _01893_, _01894_, _01895_, _01896_, _01897_, _01898_, _01899_, _01900_, _01901_, _01902_, _01903_, _01904_, _01905_, _01906_, _01907_, _01908_, _01909_, _01910_, _01911_, _01912_, _01913_, _01914_, _01915_, _01916_, _01917_, _01918_, _01919_, _01920_, _01921_, _01922_, _01923_, _01924_, _01925_, _01926_, _01927_, _01928_, _01929_, _01930_, _01931_, _01932_, _01933_, _01934_, _01935_, _01936_, _01937_, _01938_, _01939_, _01940_, _01941_, _01942_, _01943_, _01944_, _01945_, _01946_, _01947_, _01948_, _01949_, _01950_, _01951_, _01952_, _01953_, _01954_, _01955_, _01956_, _01957_, _01958_, _01959_, _01960_, _01961_, _01962_, _01963_, _01964_, _01965_, _01966_, _01967_, _01968_, _01969_, _01970_, _01971_, _01972_, _01973_, _01974_, _01975_, _01976_, _01977_, _01978_, _01979_, _01980_, _01981_, _01982_, _01983_, _01984_, _01985_, _01986_, _01987_, _01988_, _01989_, _01990_, _01991_, _01992_, _01993_, _01994_, _01995_, _01996_, _01997_, _01998_, _01999_, _02000_, _02001_, _02002_, _02003_, _02004_, _02005_, _02006_, _02007_, _02008_, _02009_, _02010_, _02011_, _02012_, _02013_, _02014_, _02015_, _02016_, _02017_, _02018_, _02019_, _02020_, _02021_, _02022_, _02023_, _02024_, _02025_, _02026_, _02027_, _02028_, _02029_, _02030_, _02031_, _02032_, _02033_, _02034_, _02035_, _02036_, _02037_, _02038_, _02039_, _02040_, _02041_, _02042_, _02043_, _02044_, _02045_, _02046_, _02047_, _02048_, _02049_, _02050_, _02051_, _02052_, _02053_, _02054_, _02055_, _02056_, _02057_, _02058_, _02059_, _02060_, _02061_, _02062_, _02063_, _02064_, _02065_, _02066_, _02067_, _02068_, _02069_, _02070_, _02071_, _02072_, _02073_, _02074_, _02075_, _02076_, _02077_, _02078_, _02079_, _02080_, _02081_, _02082_, _02083_, _02084_, _02085_, _02086_, _02087_, _02088_, _02089_, _02090_, _02091_, _02092_, _02093_, _02094_, _02095_, _02096_, _02097_, _02098_, _02099_, _02100_, _02101_, _02102_, _02103_, _02104_, _02105_, _02106_, _02107_, _02108_, _02109_, _02110_, _02111_, _02112_, _02113_, _02114_, _02115_, _02116_, _02117_, _02118_, _02119_, _02120_, _02121_, _02122_, _02123_, _02124_, _02125_, _02126_, _02127_, _02128_, _02129_, _02130_, _02131_, _02132_, _02133_, _02134_, _02135_, _02136_, _02137_, _02138_, _02139_, _02140_, _02141_, _02142_, _02143_, _02144_, _02145_, _02146_, _02147_, _02148_, _02149_, _02150_, _02151_, _02152_, _02153_, _02154_, _02155_, _02156_, _02157_, _02158_, _02159_, _02160_, _02161_, _02162_, _02163_, _02164_, _02165_, _02166_, _02167_, _02168_, _02169_, _02170_, _02171_, _02172_, _02173_, _02174_, _02175_, _02176_, _02177_, _02178_, _02179_, _02180_, _02181_, _02182_, _02183_, _02184_, _02185_, _02186_, _02187_, _02188_, _02189_, _02190_, _02191_, _02192_, _02193_, _02194_, _02195_, _02196_, _02197_, _02198_, _02199_, _02200_, _02201_, _02202_, _02203_, _02204_, _02205_, _02206_, _02207_, _02208_, _02209_, _02210_, _02211_, _02212_, _02213_, _02214_, _02215_, _02216_, _02217_, _02218_, _02219_, _02220_, _02221_, _02222_, _02223_, _02224_, _02225_, _02226_, _02227_, _02228_, _02229_, _02230_, _02231_, _02232_, _02233_, _02234_, _02235_, _02236_, _02237_, _02238_, _02239_, _02240_, _02241_, _02242_, _02243_, _02244_, _02245_, _02246_, _02247_, _02248_, _02249_, _02250_, _02251_, _02252_, _02253_, _02254_, _02255_, _02256_, _02257_, _02258_, _02259_, _02260_, _02261_, _02262_, _02263_, _02264_, _02265_, _02266_, _02267_, _02268_, _02269_, _02270_, _02271_, _02272_, _02273_, _02274_, _02275_, _02276_, _02277_, _02278_, _02279_, _02280_, _02281_, _02282_, _02283_, _02284_, _02285_, _02286_, _02287_, _02288_, _02289_, _02290_, _02291_, _02292_, _02293_, _02294_, _02295_, _02296_, _02297_, _02298_, _02299_, _02300_, _02301_, _02302_, _02303_, _02304_, _02305_, _02306_, _02307_, _02308_, _02309_, _02310_, _02311_, _02312_, _02313_, _02314_, _02315_, _02316_, _02317_, _02318_, _02319_, _02320_, _02321_, _02322_, _02323_, _02324_, _02325_, _02326_, _02327_, _02328_, _02329_, _02330_, _02331_, _02332_, _02333_, _02334_, _02335_, _02336_, _02337_, _02338_, _02339_, _02340_, _02341_, _02342_, _02343_, _02344_, _02345_, _02346_, _02347_, _02348_, _02349_, _02350_, _02351_, _02352_, _02353_, _02354_, _02355_, _02356_, _02357_, _02358_, _02359_, _02360_, _02361_, _02362_, _02363_, _02364_, _02365_, _02366_, _02367_, _02368_, _02369_, _02370_, _02371_, _02372_, _02373_, _02374_, _02375_, _02376_, _02377_, _02378_, _02379_, _02380_, _02381_, _02382_, _02383_, _02384_, _02385_, _02386_, _02387_, _02388_, _02389_, _02390_, _02391_, _02392_, _02393_, _02394_, _02395_, _02396_, _02397_, _02398_, _02399_, _02400_, _02401_, _02402_, _02403_, _02404_, _02405_, _02406_, _02407_, _02408_, _02409_, _02410_, _02411_, _02412_, _02413_, _02414_, _02415_, _02416_, _02417_, _02418_, _02419_, _02420_, _02421_, _02422_, _02423_, _02424_, _02425_, _02426_, _02427_, _02428_, _02429_, _02430_, _02431_, _02432_, _02433_, _02434_, _02435_, _02436_, _02437_, _02438_, _02439_, _02440_, _02441_, _02442_, _02443_, _02444_, _02445_, _02446_, _02447_, _02448_, _02449_, _02450_, _02451_, _02452_, _02453_, _02454_, _02455_, _02456_, _02457_, _02458_, _02459_, _02460_, _02461_, _02462_, _02463_, _02464_, _02465_, _02466_, _02467_, _02468_, _02469_, _02470_, _02471_, _02472_, _02473_, _02474_, _02475_, _02476_, _02477_, _02478_, _02479_, _02480_, _02481_, _02482_, _02483_, _02484_, _02485_, _02486_, _02487_, _02488_, _02489_, _02490_, _02491_, _02492_, _02493_, _02494_, _02495_, _02496_, _02497_, _02498_, _02499_, _02500_, _02501_, _02502_, _02503_, _02504_, _02505_, _02506_, _02507_, _02508_, _02509_, _02510_, _02511_, _02512_, _02513_, _02514_, _02515_, _02516_, _02517_, _02518_, _02519_, _02520_, _02521_, _02522_, _02523_, _02524_, _02525_, _02526_, _02527_, _02528_, _02529_, _02530_, _02531_, _02532_, _02533_, _02534_, _02535_, _02536_, _02537_, _02538_, _02539_, _02540_, _02541_, _02542_, _02543_, _02544_, _02545_, _02546_, _02547_, _02548_, _02549_, _02550_, _02551_, _02552_, _02553_, _02554_, _02555_, _02556_, _02557_, _02558_, _02559_, _02560_, _02561_, _02562_, _02563_, _02564_, _02565_, _02566_, _02567_, _02568_, _02569_, _02570_, _02571_, _02572_, _02573_, _02574_, _02575_, _02576_, _02577_, _02578_, _02579_, _02580_, _02581_, _02582_, _02583_, _02584_, _02585_, _02586_, _02587_, _02588_, _02589_, _02590_, _02591_, _02592_, _02593_, _02594_, _02595_, _02596_, _02597_, _02598_, _02599_, _02600_, _02601_, _02602_, _02603_, _02604_, _02605_, _02606_, _02607_, _02608_, _02609_, _02610_, _02611_, _02612_, _02613_, _02614_, _02615_, _02616_, _02617_, _02618_, _02619_, _02620_, _02621_, _02622_, _02623_, _02624_, _02625_, _02626_, _02627_, _02628_, _02629_, _02630_, _02631_, _02632_, _02633_, _02634_, _02635_, _02636_, _02637_, _02638_, _02639_, _02640_, _02641_, _02642_, _02643_, _02644_, _02645_, _02646_, _02647_, _02648_, _02649_, _02650_, _02651_, _02652_, _02653_, _02654_, _02655_, _02656_, _02657_, _02658_, _02659_, _02660_, _02661_, _02662_, _02663_, _02664_, _02665_, _02666_, _02667_, _02668_, _02669_, _02670_, _02671_, _02672_, _02673_, _02674_, _02675_, _02676_, _02677_, _02678_, _02679_, _02680_, _02681_, _02682_, _02683_, _02684_, _02685_, _02686_, _02687_, _02688_, _02689_, _02690_, _02691_, _02692_, _02693_, _02694_, _02695_, _02696_, _02697_, _02698_, _02699_, _02700_, _02701_, _02702_, _02703_, _02704_, _02705_, _02706_, _02707_, _02708_, _02709_, _02710_, _02711_, _02712_, _02713_, _02714_, _02715_, _02716_, _02717_, _02718_, _02719_, _02720_, _02721_, _02722_, _02723_, _02724_, _02725_, _02726_, _02727_, _02728_, _02729_, _02730_, _02731_, _02732_, _02733_, _02734_, _02735_, _02736_, _02737_, _02738_, _02739_, _02740_, _02741_, _02742_, _02743_, _02744_, _02745_, _02746_, _02747_, _02748_, _02749_, _02750_, _02751_, _02752_, _02753_, _02754_, _02755_, _02756_, _02757_, _02758_, _02759_, _02760_, _02761_, _02762_, _02763_, _02764_, _02765_, _02766_, _02767_, _02768_, _02769_, _02770_, _02771_, _02772_, _02773_, _02774_, _02775_, _02776_, _02777_, _02778_, _02779_, _02780_, _02781_, _02782_, _02783_, _02784_, _02785_, _02786_, _02787_, _02788_, _02789_, _02790_, _02791_, _02792_, _02793_, _02794_, _02795_, _02796_, _02797_, _02798_, _02799_, _02800_, _02801_, _02802_, _02803_, _02804_, _02805_, _02806_, _02807_, _02808_, _02809_, _02810_, _02811_, _02812_, _02813_, _02814_, _02815_, _02816_, _02817_, _02818_, _02819_, _02820_, _02821_, _02822_, _02823_, _02824_, _02825_, _02826_, _02827_, _02828_, _02829_, _02830_, _02831_, _02832_, _02833_, _02834_, _02835_, _02836_, _02837_, _02838_, _02839_, _02840_, _02841_, _02842_, _02843_, _02844_, _02845_, _02846_, _02847_, _02848_, _02849_, _02850_, _02851_, _02852_, _02853_, _02854_, _02855_, _02856_, _02857_, _02858_, _02859_, _02860_, _02861_, _02862_, _02863_, _02864_, _02865_, _02866_, _02867_, _02868_, _02869_, _02870_, _02871_, _02872_, _02873_, _02874_, _02875_, _02876_, _02877_, _02878_, _02879_, _02880_, _02881_, _02882_, _02883_, _02884_, _02885_, _02886_, _02887_, _02888_, _02889_, _02890_, _02891_, _02892_, _02893_, _02894_, _02895_, _02896_, _02897_, _02898_, _02899_, _02900_, _02901_, _02902_, _02903_, _02904_, _02905_, _02906_, _02907_, _02908_, _02909_, _02910_, _02911_, _02912_, _02913_, _02914_, _02915_, _02916_, _02917_, _02918_, _02919_, _02920_, _02921_, _02922_, _02923_, _02924_, _02925_, _02926_, _02927_, _02928_, _02929_, _02930_, _02931_, _02932_, _02933_, _02934_, _02935_, _02936_, _02937_, _02938_, _02939_, _02940_, _02941_, _02942_, _02943_, _02944_, _02945_, _02946_, _02947_, _02948_, _02949_, _02950_, _02951_, _02952_, _02953_, _02954_, _02955_, _02956_, _02957_, _02958_, _02959_, _02960_, _02961_, _02962_, _02963_, _02964_, _02965_, _02966_, _02967_, _02968_, _02969_, _02970_, _02971_, _02972_, _02973_, _02974_, _02975_, _02976_, _02977_, _02978_, _02979_, _02980_, _02981_, _02982_, _02983_, _02984_, _02985_, _02986_, _02987_, _02988_, _02989_, _02990_, _02991_, _02992_, _02993_, _02994_, _02995_, _02996_, _02997_, _02998_, _02999_, _03000_, _03001_, _03002_, _03003_, _03004_, _03005_, _03006_, _03007_, _03008_, _03009_, _03010_, _03011_, _03012_, _03013_, _03014_, _03015_, _03016_, _03017_, _03018_, _03019_, _03020_, _03021_, _03022_, _03023_, _03024_, _03025_, _03026_, _03027_, _03028_, _03029_, _03030_, _03031_, _03032_, _03033_, _03034_, _03035_, _03036_, _03037_, _03038_, _03039_, _03040_, _03041_, _03042_, _03043_, _03044_, _03045_, _03046_, _03047_, _03048_, _03049_, _03050_, _03051_, _03052_, _03053_, _03054_, _03055_, _03056_, _03057_, _03058_, _03059_, _03060_, _03061_, _03062_, _03063_, _03064_, _03065_, _03066_, _03067_, _03068_, _03069_, _03070_, _03071_, _03072_, _03073_, _03074_, _03075_, _03076_, _03077_, _03078_, _03079_, _03080_, _03081_, _03082_, _03083_, _03084_, _03085_, _03086_, _03087_, _03088_, _03089_, _03090_, _03091_, _03092_, _03093_, _03094_, _03095_, _03096_, _03097_, _03098_, _03099_, _03100_, _03101_, _03102_, _03103_, _03104_, _03105_, _03106_, _03107_, _03108_, _03109_, _03110_, _03111_, _03112_, _03113_, _03114_, _03115_, _03116_, _03117_, _03118_, _03119_, _03120_, _03121_, _03122_, _03123_, _03124_, _03125_, _03126_, _03127_, _03128_, _03129_, _03130_, _03131_, _03132_, _03133_, _03134_, _03135_, _03136_, _03137_, _03138_, _03139_, _03140_, _03141_, _03142_, _03143_, _03144_, _03145_, _03146_, _03147_, _03148_, _03149_, _03150_, _03151_, _03152_, _03153_, _03154_, _03155_, _03156_, _03157_, _03158_, _03159_, _03160_, _03161_, _03162_, _03163_, _03164_, _03165_, _03166_, _03167_, _03168_, _03169_, _03170_, _03171_, _03172_, _03173_, _03174_, _03175_, _03176_, _03177_, _03178_, _03179_, _03180_, _03181_, _03182_, _03183_, _03184_, _03185_, _03186_, _03187_, _03188_, _03189_, _03190_, _03191_, _03192_, _03193_, _03194_, _03195_, _03196_, _03197_, _03198_, _03199_, _03200_, _03201_, _03202_, _03203_, _03204_, _03205_, _03206_, _03207_, _03208_, _03209_, _03210_, _03211_, _03212_, _03213_, _03214_, _03215_, _03216_, _03217_, _03218_, _03219_, _03220_, _03221_, _03222_, _03223_, _03224_, _03225_, _03226_, _03227_, _03228_, _03229_, _03230_, _03231_, _03232_, _03233_, _03234_, _03235_, _03236_, _03237_, _03238_, _03239_, _03240_, _03241_, _03242_, _03243_, _03244_, _03245_, _03246_, _03247_, _03248_, _03249_, _03250_, _03251_, _03252_, _03253_, _03254_, _03255_, _03256_, _03257_, _03258_, _03259_, _03260_, _03261_, _03262_, _03263_, _03264_, _03265_, _03266_, _03267_, _03268_, _03269_, _03270_, _03271_, _03272_, _03273_, _03274_, _03275_, _03276_, _03277_, _03278_, _03279_, _03280_, _03281_, _03282_, _03283_, _03284_, _03285_, _03286_, _03287_, _03288_, _03289_, _03290_, _03291_, _03292_, _03293_, _03294_, _03295_, _03296_, _03297_, _03298_, _03299_, _03300_, _03301_, _03302_, _03303_, _03304_, _03305_, _03306_, _03307_, _03308_, _03309_, _03310_, _03311_, _03312_, _03313_, _03314_, _03315_, _03316_, _03317_, _03318_, _03319_, _03320_, _03321_, _03322_, _03323_, _03324_, _03325_, _03326_, _03327_, _03328_, _03329_, _03330_, _03331_, _03332_, _03333_, _03334_, _03335_, _03336_, _03337_, _03338_, _03339_, _03340_, _03341_, _03342_, _03343_, _03344_, _03345_, _03346_, _03347_, _03348_, _03349_, _03350_, _03351_, _03352_, _03353_, _03354_, _03355_, _03356_, _03357_, _03358_, _03359_, _03360_, _03361_, _03362_, _03363_, _03364_, _03365_, _03366_, _03367_, _03368_, _03369_, _03370_, _03371_, _03372_, _03373_, _03374_, _03375_, _03376_, _03377_, _03378_, _03379_, _03380_, _03381_, _03382_, _03383_, _03384_, _03385_, _03386_, _03387_, _03388_, _03389_, _03390_, _03391_, _03392_, _03393_, _03394_, _03395_, _03396_, _03397_, _03398_, _03399_, _03400_, _03401_, _03402_, _03403_, _03404_, _03405_, _03406_, _03407_, _03408_, _03409_, _03410_, _03411_, _03412_, _03413_, _03414_, _03415_, _03416_, _03417_, _03418_, _03419_, _03420_, _03421_, _03422_, _03423_, _03424_, _03425_, _03426_, _03427_, _03428_, _03429_, _03430_, _03431_, _03432_, _03433_, _03434_, _03435_, _03436_, _03437_, _03438_, _03439_, _03440_, _03441_, _03442_, _03443_, _03444_, _03445_, _03446_, _03447_, _03448_, _03449_, _03450_, _03451_, _03452_, _03453_, _03454_, _03455_, _03456_, _03457_, _03458_, _03459_, _03460_, _03461_, _03462_, _03463_, _03464_, _03465_, _03466_, _03467_, _03468_, _03469_, _03470_, _03471_, _03472_, _03473_, _03474_, _03475_, _03476_, _03477_, _03478_, _03479_, _03480_, _03481_, _03482_, _03483_, _03484_, _03485_, _03486_, _03487_, _03488_, _03489_, _03490_, _03491_, _03492_, _03493_, _03494_, _03495_, _03496_, _03497_, _03498_, _03499_, _03500_, _03501_, _03502_, _03503_, _03504_, _03505_, _03506_, _03507_, _03508_, _03509_, _03510_, _03511_, _03512_, _03513_, _03514_, _03515_, _03516_, _03517_, _03518_, _03519_, _03520_, _03521_, _03522_, _03523_, _03524_, _03525_, _03526_, _03527_, _03528_, _03529_, _03530_, _03531_, _03532_, _03533_, _03534_, _03535_, _03536_, _03537_, _03538_, _03539_, _03540_, _03541_, _03542_, _03543_, _03544_, _03545_, _03546_, _03547_, _03548_, _03549_, _03550_, _03551_, _03552_, _03553_, _03554_, _03555_, _03556_, _03557_, _03558_, _03559_, _03560_, _03561_, _03562_, _03563_, _03564_, _03565_, _03566_, _03567_, _03568_, _03569_, _03570_, _03571_, _03572_, _03573_, _03574_, _03575_, _03576_, _03577_, _03578_, _03579_, _03580_, _03581_, _03582_, _03583_, _03584_, _03585_, _03586_, _03587_, _03588_, _03589_, _03590_, _03591_, _03592_, _03593_, _03594_, _03595_, _03596_, _03597_, _03598_, _03599_, _03600_, _03601_, _03602_, _03603_, _03604_, _03605_, _03606_, _03607_, _03608_, _03609_, _03610_, _03611_, _03612_, _03613_, _03614_, _03615_, _03616_, _03617_, _03618_, _03619_, _03620_, _03621_, _03622_, _03623_, _03624_, _03625_, _03626_, _03627_, _03628_, _03629_, _03630_, _03631_, _03632_, _03633_, _03634_, _03635_, _03636_, _03637_, _03638_, _03639_, _03640_, _03641_, _03642_, _03643_, _03644_, _03645_, _03646_, _03647_, _03648_, _03649_, _03650_, _03651_, _03652_, _03653_, _03654_, _03655_, _03656_, _03657_, _03658_, _03659_, _03660_, _03661_, _03662_, _03663_, _03664_, _03665_, _03666_, _03667_, _03668_, _03669_, _03670_, _03671_, _03672_, _03673_, _03674_, _03675_, _03676_, _03677_, _03678_, _03679_, _03680_, _03681_, _03682_, _03683_, _03684_, _03685_, _03686_, _03687_, _03688_, _03689_, _03690_, _03691_, _03692_, _03693_, _03694_, _03695_, _03696_, _03697_, _03698_, _03699_, _03700_, _03701_, _03702_, _03703_, _03704_, _03705_, _03706_, _03707_, _03708_, _03709_, _03710_, _03711_, _03712_, _03713_, _03714_, _03715_, _03716_, _03717_, _03718_, _03719_, _03720_, _03721_, _03722_, _03723_, _03724_, _03725_, _03726_, _03727_, _03728_, _03729_, _03730_, _03731_, _03732_, _03733_, _03734_, _03735_, _03736_, _03737_, _03738_, _03739_, _03740_, _03741_, _03742_, _03743_, _03744_, _03745_, _03746_, _03747_, _03748_, _03749_, _03750_, _03751_, _03752_, _03753_, _03754_, _03755_, _03756_, _03757_, _03758_, _03759_, _03760_, _03761_, _03762_, _03763_, _03764_, _03765_, _03766_, _03767_, _03768_, _03769_, _03770_, _03771_, _03772_, _03773_, _03774_, _03775_, _03776_, _03777_, _03778_, _03779_, _03780_, _03781_, _03782_, _03783_, _03784_, _03785_, _03786_, _03787_, _03788_, _03789_, _03790_, _03791_, _03792_, _03793_, _03794_, _03795_, _03796_, _03797_, _03798_, _03799_, _03800_, _03801_, _03802_, _03803_, _03804_, _03805_, _03806_, _03807_, _03808_, _03809_, _03810_, _03811_, _03812_, _03813_, _03814_, _03815_, _03816_, _03817_, _03818_, _03819_, _03820_, _03821_, _03822_, _03823_, _03824_, _03825_, _03826_, _03827_, _03828_, _03829_, _03830_, _03831_, _03832_, _03833_, _03834_, _03835_, _03836_, _03837_, _03838_, _03839_, _03840_, _03841_, _03842_, _03843_, _03844_, _03845_, _03846_, _03847_, _03848_, _03849_, _03850_, _03851_, _03852_, _03853_, _03854_, _03855_, _03856_, _03857_, _03858_, _03859_, _03860_, _03861_, _03862_, _03863_, _03864_, _03865_, _03866_, _03867_, _03868_, _03869_, _03870_, _03871_, _03872_, _03873_, _03874_, _03875_, _03876_, _03877_, _03878_, _03879_, _03880_, _03881_, _03882_, _03883_, _03884_, _03885_, _03886_, _03887_, _03888_, _03889_, _03890_, _03891_, _03892_, _03893_, _03894_, _03895_, _03896_, _03897_, _03898_, _03899_, _03900_, _03901_, _03902_, _03903_, _03904_, _03905_, _03906_, _03907_, _03908_, _03909_, _03910_, _03911_, _03912_, _03913_, _03914_, _03915_, _03916_, _03917_, _03918_, _03919_, _03920_, _03921_, _03922_, _03923_, _03924_, _03925_, _03926_, _03927_, _03928_, _03929_, _03930_, _03931_, _03932_, _03933_, _03934_, _03935_, _03936_, _03937_, _03938_, _03939_, _03940_, _03941_, _03942_, _03943_, _03944_, _03945_, _03946_, _03947_, _03948_, _03949_, _03950_, _03951_, _03952_, _03953_, _03954_, _03955_, _03956_, _03957_, _03958_, _03959_, _03960_, _03961_, _03962_, _03963_, _03964_, _03965_, _03966_, _03967_, _03968_, _03969_, _03970_, _03971_, _03972_, _03973_, _03974_, _03975_, _03976_, _03977_, _03978_, _03979_, _03980_, _03981_, _03982_, _03983_, _03984_, _03985_, _03986_, _03987_, _03988_, _03989_, _03990_, _03991_, _03992_, _03993_, _03994_, _03995_, _03996_, _03997_, _03998_, _03999_, _04000_, _04001_, _04002_, _04003_, _04004_, _04005_, _04006_, _04007_, _04008_, _04009_, _04010_, _04011_, _04012_, _04013_, _04014_, _04015_, _04016_, _04017_, _04018_, _04019_, _04020_, _04021_, _04022_, _04023_, _04024_, _04025_, _04026_, _04027_, _04028_, _04029_, _04030_, _04031_, _04032_, _04033_, _04034_, _04035_, _04036_, _04037_, _04038_, _04039_, _04040_, _04041_, _04042_, _04043_, _04044_, _04045_, _04046_, _04047_, _04048_, _04049_, _04050_, _04051_, _04052_, _04053_, _04054_, _04055_, _04056_, _04057_, _04058_, _04059_, _04060_, _04061_, _04062_, _04063_, _04064_, _04065_, _04066_, _04067_, _04068_, _04069_, _04070_, _04071_, _04072_, _04073_, _04074_, _04075_, _04076_, _04077_, _04078_, _04079_, _04080_, _04081_, _04082_, _04083_, _04084_, _04085_, _04086_, _04087_, _04088_, _04089_, _04090_, _04091_, _04092_, _04093_, _04094_, _04095_, _04096_, _04097_, _04098_, _04099_, _04100_, _04101_, _04102_, _04103_, _04104_, _04105_, _04106_, _04107_, _04108_, _04109_, _04110_, _04111_, _04112_, _04113_, _04114_, _04115_, _04116_, _04117_, _04118_, _04119_, _04120_, _04121_, _04122_, _04123_, _04124_, _04125_, _04126_, _04127_, _04128_, _04129_, _04130_, _04131_, _04132_, _04133_, _04134_, _04135_, _04136_, _04137_, _04138_, _04139_, _04140_, _04141_, _04142_, _04143_, _04144_, _04145_, _04146_, _04147_, _04148_, _04149_, _04150_, _04151_, _04152_, _04153_, _04154_, _04155_, _04156_, _04157_, _04158_, _04159_, _04160_, _04161_, _04162_, _04163_, _04164_, _04165_, _04166_, _04167_, _04168_, _04169_, _04170_, _04171_, _04172_, _04173_, _04174_, _04175_, _04176_, _04177_, _04178_, _04179_, _04180_, _04181_, _04182_, _04183_, _04184_, _04185_, _04186_, _04187_, _04188_, _04189_, _04190_, _04191_, _04192_, _04193_, _04194_, _04195_, _04196_, _04197_, _04198_, _04199_, _04200_, _04201_, _04202_, _04203_, _04204_, _04205_, _04206_, _04207_, _04208_, _04209_, _04210_, _04211_, _04212_, _04213_, _04214_, _04215_, _04216_, _04217_, _04218_, _04219_, _04220_, _04221_, _04222_, _04223_, _04224_, _04225_, _04226_, _04227_, _04228_, _04229_, _04230_, _04231_, _04232_, _04233_, _04234_, _04235_, _04236_, _04237_, _04238_, _04239_, _04240_, _04241_, _04242_, _04243_, _04244_, _04245_, _04246_, _04247_, _04248_, _04249_, _04250_, _04251_, _04252_, _04253_, _04254_, _04255_, _04256_, _04257_, _04258_, _04259_, _04260_, _04261_, _04262_, _04263_, _04264_, _04265_, _04266_, _04267_, _04268_, _04269_, _04270_, _04271_, _04272_, _04273_, _04274_, _04275_, _04276_, _04277_, _04278_, _04279_, _04280_, _04281_, _04282_, _04283_, _04284_, _04285_, _04286_, _04287_, _04288_, _04289_, _04290_, _04291_, _04292_, _04293_, _04294_, _04295_, _04296_, _04297_, _04298_, _04299_, _04300_, _04301_, _04302_, _04303_, _04304_, _04305_, _04306_, _04307_, _04308_, _04309_, _04310_, _04311_, _04312_, _04313_, _04314_, _04315_, _04316_, _04317_, _04318_, _04319_, _04320_, _04321_, _04322_, _04323_, _04324_, _04325_, _04326_, _04327_, _04328_, _04329_, _04330_, _04331_, _04332_, _04333_, _04334_, _04335_, _04336_, _04337_, _04338_, _04339_, _04340_, _04341_, _04342_, _04343_, _04344_, _04345_, _04346_, _04347_, _04348_, _04349_, _04350_, _04351_, _04352_, _04353_, _04354_, _04355_, _04356_, _04357_, _04358_, _04359_, _04360_, _04361_, _04362_, _04363_, _04364_, _04365_, _04366_, _04367_, _04368_, _04369_, _04370_, _04371_, _04372_, _04373_, _04374_, _04375_, _04376_, _04377_, _04378_, _04379_, _04380_, _04381_, _04382_, _04383_, _04384_, _04385_, _04386_, _04387_, _04388_, _04389_, _04390_, _04391_, _04392_, _04393_, _04394_, _04395_, _04396_, _04397_, _04398_, _04399_, _04400_, _04401_, _04402_, _04403_, _04404_, _04405_, _04406_, _04407_, _04408_, _04409_, _04410_, _04411_, _04412_, _04413_, _04414_, _04415_, _04416_, _04417_, _04418_, _04419_, _04420_, _04421_, _04422_, _04423_, _04424_, _04425_, _04426_, _04427_, _04428_, _04429_, _04430_, _04431_, _04432_, _04433_, _04434_, _04435_, _04436_, _04437_, _04438_, _04439_, _04440_, _04441_, _04442_, _04443_, _04444_, _04445_, _04446_, _04447_, _04448_, _04449_, _04450_, _04451_, _04452_, _04453_, _04454_, _04455_, _04456_, _04457_, _04458_, _04459_, _04460_, _04461_, _04462_, _04463_, _04464_, _04465_, _04466_, _04467_, _04468_, _04469_, _04470_, _04471_, _04472_, _04473_, _04474_, _04475_, _04476_, _04477_, _04478_, _04479_, _04480_, _04481_, _04482_, _04483_, _04484_, _04485_, _04486_, _04487_, _04488_, _04489_, _04490_, _04491_, _04492_, _04493_, _04494_, _04495_, _04496_, _04497_, _04498_, _04499_, _04500_, _04501_, _04502_, _04503_, _04504_, _04505_, _04506_, _04507_, _04508_, _04509_, _04510_, _04511_, _04512_, _04513_, _04514_, _04515_, _04516_, _04517_, _04518_, _04519_, _04520_, _04521_, _04522_, _04523_, _04524_, _04525_, _04526_, _04527_, _04528_, _04529_, _04530_, _04531_, _04532_, _04533_, _04534_, _04535_, _04536_, _04537_, _04538_, _04539_, _04540_, _04541_, _04542_, _04543_, _04544_, _04545_, _04546_, _04547_, _04548_, _04549_, _04550_, _04551_, _04552_, _04553_, _04554_, _04555_, _04556_, _04557_, _04558_, _04559_, _04560_, _04561_, _04562_, _04563_, _04564_, _04565_, _04566_, _04567_, _04568_, _04569_, _04570_, _04571_, _04572_, _04573_, _04574_, _04575_, _04576_, _04577_, _04578_, _04579_, _04580_, _04581_, _04582_, _04583_, _04584_, _04585_, _04586_, _04587_, _04588_, _04589_, _04590_, _04591_, _04592_, _04593_, _04594_, _04595_, _04596_, _04597_, _04598_, _04599_, _04600_, _04601_, _04602_, _04603_, _04604_, _04605_, _04606_, _04607_, _04608_, _04609_, _04610_, _04611_, _04612_, _04613_, _04614_, _04615_, _04616_, _04617_, _04618_, _04619_, _04620_, _04621_, _04622_, _04623_, _04624_, _04625_, _04626_, _04627_, _04628_, _04629_, _04630_, _04631_, _04632_, _04633_, _04634_, _04635_, _04636_, _04637_, _04638_, _04639_, _04640_, _04641_, _04642_, _04643_, _04644_, _04645_, _04646_, _04647_, _04648_, _04649_, _04650_, _04651_, _04652_, _04653_, _04654_, _04655_, _04656_, _04657_, _04658_, _04659_, _04660_, _04661_, _04662_, _04663_, _04664_, _04665_, _04666_, _04667_, _04668_, _04669_, _04670_, _04671_, _04672_, _04673_, _04674_, _04675_, _04676_, _04677_, _04678_, _04679_, _04680_, _04681_, _04682_, _04683_, _04684_, _04685_, _04686_, _04687_, _04688_, _04689_, _04690_, _04691_, _04692_, _04693_, _04694_, _04695_, _04696_, _04697_, _04698_, _04699_, _04700_, _04701_, _04702_, _04703_, _04704_, _04705_, _04706_, _04707_, _04708_, _04709_, _04710_, _04711_, _04712_, _04713_, _04714_, _04715_, _04716_, _04717_, _04718_, _04719_, _04720_, _04721_, _04722_, _04723_, _04724_, _04725_, _04726_, _04727_, _04728_, _04729_, _04730_, _04731_, _04732_, _04733_, _04734_, _04735_, _04736_, _04737_, _04738_, _04739_, _04740_, _04741_, _04742_, _04743_, _04744_, _04745_, _04746_, _04747_, _04748_, _04749_, _04750_, _04751_, _04752_, _04753_, _04754_, _04755_, _04756_, _04757_, _04758_, _04759_, _04760_, _04761_, _04762_, _04763_, _04764_, _04765_, _04766_, _04767_, _04768_, _04769_, _04770_, _04771_, _04772_, _04773_, _04774_, _04775_, _04776_, _04777_, _04778_, _04779_, _04780_, _04781_, _04782_, _04783_, _04784_, _04785_, _04786_, _04787_, _04788_, _04789_, _04790_, _04791_, _04792_, _04793_, _04794_, _04795_, _04796_, _04797_, _04798_, _04799_, _04800_, _04801_, _04802_, _04803_, _04804_, _04805_, _04806_, _04807_, _04808_, _04809_, _04810_, _04811_, _04812_, _04813_, _04814_, _04815_, _04816_, _04817_, _04818_, _04819_, _04820_, _04821_, _04822_, _04823_, _04824_, _04825_, _04826_, _04827_, _04828_, _04829_, _04830_, _04831_, _04832_, _04833_, _04834_, _04835_, _04836_, _04837_, _04838_, _04839_, _04840_, _04841_, _04842_, _04843_, _04844_, _04845_, _04846_, _04847_, _04848_, _04849_, _04850_, _04851_, _04852_, _04853_, _04854_, _04855_, _04856_, _04857_, _04858_, _04859_, _04860_, _04861_, _04862_, _04863_, _04864_, _04865_, _04866_, _04867_, _04868_, _04869_, _04870_, _04871_, _04872_, _04873_, _04874_, _04875_, _04876_, _04877_, _04878_, _04879_, _04880_, _04881_, _04882_, _04883_, _04884_, _04885_, _04886_, _04887_, _04888_, _04889_, _04890_, _04891_, _04892_, _04893_, _04894_, _04895_, _04896_, _04897_, _04898_, _04899_, _04900_, _04901_, _04902_, _04903_, _04904_, _04905_, _04906_, _04907_, _04908_, _04909_, _04910_, _04911_, _04912_, _04913_, _04914_, _04915_, _04916_, _04917_, _04918_, _04919_, _04920_, _04921_, _04922_, _04923_, _04924_, _04925_, _04926_, _04927_, _04928_, _04929_, _04930_, _04931_, _04932_, _04933_, _04934_, _04935_, _04936_, _04937_, _04938_, _04939_, _04940_, _04941_, _04942_, _04943_, _04944_, _04945_, _04946_, _04947_, _04948_, _04949_, _04950_, _04951_, _04952_, _04953_, _04954_, _04955_, _04956_, _04957_, _04958_, _04959_, _04960_, _04961_, _04962_, _04963_, _04964_, _04965_, _04966_, _04967_, _04968_, _04969_, _04970_, _04971_, _04972_, _04973_, _04974_, _04975_, _04976_, _04977_, _04978_, _04979_, _04980_, _04981_, _04982_, _04983_, _04984_, _04985_, _04986_, _04987_, _04988_, _04989_, _04990_, _04991_, _04992_, _04993_, _04994_, _04995_, _04996_, _04997_, _04998_, _04999_, _05000_, _05001_, _05002_, _05003_, _05004_, _05005_, _05006_, _05007_, _05008_, _05009_, _05010_, _05011_, _05012_, _05013_, _05014_, _05015_, _05016_, _05017_, _05018_, _05019_, _05020_, _05021_, _05022_, _05023_, _05024_, _05025_, _05026_, _05027_, _05028_, _05029_, _05030_, _05031_, _05032_, _05033_, _05034_, _05035_, _05036_, _05037_, _05038_, _05039_, _05040_, _05041_, _05042_, _05043_, _05044_, _05045_, _05046_, _05047_, _05048_, _05049_, _05050_, _05051_, _05052_, _05053_, _05054_, _05055_, _05056_, _05057_, _05058_, _05059_, _05060_, _05061_, _05062_, _05063_, _05064_, _05065_, _05066_, _05067_, _05068_, _05069_, _05070_, _05071_, _05072_, _05073_, _05074_, _05075_, _05076_, _05077_, _05078_, _05079_, _05080_, _05081_, _05082_, _05083_, _05084_, _05085_, _05086_, _05087_, _05088_, _05089_, _05090_, _05091_, _05092_, _05093_, _05094_, _05095_, _05096_, _05097_, _05098_, _05099_, _05100_, _05101_, _05102_, _05103_, _05104_, _05105_, _05106_, _05107_, _05108_, _05109_, _05110_, _05111_, _05112_, _05113_, _05114_, _05115_, _05116_, _05117_, _05118_, _05119_, _05120_, _05121_, _05122_, _05123_, _05124_, _05125_, _05126_, _05127_, _05128_, _05129_, _05130_, _05131_, _05132_, _05133_, _05134_, _05135_, _05136_, _05137_, _05138_, _05139_, _05140_, _05141_, _05142_, _05143_, _05144_, _05145_, _05146_, _05147_, _05148_, _05149_, _05150_, _05151_, _05152_, _05153_, _05154_, _05155_, _05156_, _05157_, _05158_, _05159_, _05160_, _05161_, _05162_, _05163_, _05164_, _05165_, _05166_, _05167_, _05168_, _05169_, _05170_, _05171_, _05172_, _05173_, _05174_, _05175_, _05176_, _05177_, _05178_, _05179_, _05180_, _05181_, _05182_, _05183_, _05184_, _05185_, _05186_, _05187_, _05188_, _05189_, _05190_, _05191_, _05192_, _05193_, _05194_, _05195_, _05196_, _05197_, _05198_, _05199_, _05200_, _05201_, _05202_, _05203_, _05204_, _05205_, _05206_, _05207_, _05208_, _05209_, _05210_, _05211_, _05212_, _05213_, _05214_, _05215_, _05216_, _05217_, _05218_, _05219_, _05220_, _05221_, _05222_, _05223_, _05224_, _05225_, _05226_, _05227_, _05228_, _05229_, _05230_, _05231_, _05232_, _05233_, _05234_, _05235_, _05236_, _05237_, _05238_, _05239_, _05240_, _05241_, _05242_, _05243_, _05244_, _05245_, _05246_, _05247_, _05248_, _05249_, _05250_, _05251_, _05252_, _05253_, _05254_, _05255_, _05256_, _05257_, _05258_, _05259_, _05260_, _05261_, _05262_, _05263_, _05264_, _05265_, _05266_, _05267_, _05268_, _05269_, _05270_, _05271_, _05272_, _05273_, _05274_, _05275_, _05276_, _05277_, _05278_, _05279_, _05280_, _05281_, _05282_, _05283_, _05284_, _05285_, _05286_, _05287_, _05288_, _05289_, _05290_, _05291_, _05292_, _05293_, _05294_, _05295_, _05296_, _05297_, _05298_, _05299_, _05300_, _05301_, _05302_, _05303_, _05304_, _05305_, _05306_, _05307_, _05308_, _05309_, _05310_, _05311_, _05312_, _05313_, _05314_, _05315_, _05316_, _05317_, _05318_, _05319_, _05320_, _05321_, _05322_, _05323_, _05324_, _05325_, _05326_, _05327_, _05328_, _05329_, _05330_, _05331_, _05332_, _05333_, _05334_, _05335_, _05336_, _05337_, _05338_, _05339_, _05340_, _05341_, _05342_, _05343_, _05344_, _05345_, _05346_, _05347_, _05348_, _05349_, _05350_, _05351_, _05352_, _05353_, _05354_, _05355_, _05356_, _05357_, _05358_, _05359_, _05360_, _05361_, _05362_, _05363_, _05364_, _05365_, _05366_, _05367_, _05368_, _05369_, _05370_, _05371_, _05372_, _05373_, _05374_, _05375_, _05376_, _05377_, _05378_, _05379_, _05380_, _05381_, _05382_, _05383_, _05384_, _05385_, _05386_, _05387_, _05388_, _05389_, _05390_, _05391_, _05392_, _05393_, _05394_, _05395_, _05396_, _05397_, _05398_, _05399_, _05400_, _05401_, _05402_, _05403_, _05404_, _05405_, _05406_, _05407_, _05408_, _05409_, _05410_, _05411_, _05412_, _05413_, _05414_, _05415_, _05416_, _05417_, _05418_, _05419_, _05420_, _05421_, _05422_, _05423_, _05424_, _05425_, _05426_, _05427_, _05428_, _05429_, _05430_, _05431_, _05432_, _05433_, _05434_, _05435_, _05436_, _05437_, _05438_, _05439_, _05440_, _05441_, _05442_, _05443_, _05444_, _05445_, _05446_, _05447_, _05448_, _05449_, _05450_, _05451_, _05452_, _05453_, _05454_, _05455_, _05456_, _05457_, _05458_, _05459_, _05460_, _05461_, _05462_, _05463_, _05464_, _05465_, _05466_, _05467_, _05468_, _05469_, _05470_, _05471_, _05472_, _05473_, _05474_, _05475_, _05476_, _05477_, _05478_, _05479_, _05480_, _05481_, _05482_, _05483_, _05484_, _05485_, _05486_, _05487_, _05488_, _05489_, _05490_, _05491_, _05492_, _05493_, _05494_, _05495_, _05496_, _05497_, _05498_, _05499_, _05500_, _05501_, _05502_, _05503_, _05504_, _05505_, _05506_, _05507_, _05508_, _05509_, _05510_, _05511_, _05512_, _05513_, _05514_, _05515_, _05516_, _05517_, _05518_, _05519_, _05520_, _05521_, _05522_, _05523_, _05524_, _05525_, _05526_, _05527_, _05528_, _05529_, _05530_, _05531_, _05532_, _05533_, _05534_, _05535_, _05536_, _05537_, _05538_, _05539_, _05540_, _05541_, _05542_, _05543_, _05544_, _05545_, _05546_, _05547_, _05548_, _05549_, _05550_, _05551_, _05552_, _05553_, _05554_, _05555_, _05556_, _05557_, _05558_, _05559_, _05560_, _05561_, _05562_, _05563_, _05564_, _05565_, _05566_, _05567_, _05568_, _05569_, _05570_, _05571_, _05572_, _05573_, _05574_, _05575_, _05576_, _05577_, _05578_, _05579_, _05580_, _05581_, _05582_, _05583_, _05584_, _05585_, _05586_, _05587_, _05588_, _05589_, _05590_, _05591_, _05592_, _05593_, _05594_, _05595_, _05596_, _05597_, _05598_, _05599_, _05600_, _05601_, _05602_, _05603_, _05604_, _05605_, _05606_, _05607_, _05608_, _05609_, _05610_, _05611_, _05612_, _05613_, _05614_, _05615_, _05616_, _05617_, _05618_, _05619_, _05620_, _05621_, _05622_, _05623_, _05624_, _05625_, _05626_, _05627_, _05628_, _05629_, _05630_, _05631_, _05632_, _05633_, _05634_, _05635_, _05636_, _05637_, _05638_, _05639_, _05640_, _05641_, _05642_, _05643_, _05644_, _05645_, _05646_, _05647_, _05648_, _05649_, _05650_, _05651_, _05652_, _05653_, _05654_, _05655_, _05656_, _05657_, _05658_, _05659_, _05660_, _05661_, _05662_, _05663_, _05664_, _05665_, _05666_, _05667_, _05668_, _05669_, _05670_, _05671_, _05672_, _05673_, _05674_, _05675_, _05676_, _05677_, _05678_, _05679_, _05680_, _05681_, _05682_, _05683_, _05684_, _05685_, _05686_, _05687_, _05688_, _05689_, _05690_, _05691_, _05692_, _05693_, _05694_, _05695_, _05696_, _05697_, _05698_, _05699_, _05700_, _05701_, _05702_, _05703_, _05704_, _05705_, _05706_, _05707_, _05708_, _05709_, _05710_, _05711_, _05712_, _05713_, _05714_, _05715_, _05716_, _05717_, _05718_, _05719_, _05720_, _05721_, _05722_, _05723_, _05724_, _05725_, _05726_, _05727_, _05728_, _05729_, _05730_, _05731_, _05732_, _05733_, _05734_, _05735_, _05736_, _05737_, _05738_, _05739_, _05740_, _05741_, _05742_, _05743_, _05744_, _05745_, _05746_, _05747_, _05748_, _05749_, _05750_, _05751_, _05752_, _05753_, _05754_, _05755_, _05756_, _05757_, _05758_, _05759_, _05760_, _05761_, _05762_, _05763_, _05764_, _05765_, _05766_, _05767_, _05768_, _05769_, _05770_, _05771_, _05772_, _05773_, _05774_, _05775_, _05776_, _05777_, _05778_, _05779_, _05780_, _05781_, _05782_, _05783_, _05784_, _05785_, _05786_, _05787_, _05788_, _05789_, _05790_, _05791_, _05792_, _05793_, _05794_, _05795_, _05796_, _05797_, _05798_, _05799_, _05800_, _05801_, _05802_, _05803_, _05804_, _05805_, _05806_, _05807_, _05808_, _05809_, _05810_, _05811_, _05812_, _05813_, _05814_, _05815_, _05816_, _05817_, _05818_, _05819_, _05820_, _05821_, _05822_, _05823_, _05824_, _05825_, _05826_, _05827_, _05828_, _05829_, _05830_, _05831_, _05832_, _05833_, _05834_, _05835_, _05836_, _05837_, _05838_, _05839_, _05840_, _05841_, _05842_, _05843_, _05844_, _05845_, _05846_, _05847_, _05848_, _05849_, _05850_, _05851_, _05852_, _05853_, _05854_, _05855_, _05856_, _05857_, _05858_, _05859_, _05860_, _05861_, _05862_, _05863_, _05864_, _05865_, _05866_, _05867_, _05868_, _05869_, _05870_, _05871_, _05872_, _05873_, _05874_, _05875_, _05876_, _05877_, _05878_, _05879_, _05880_, _05881_, _05882_, _05883_, _05884_, _05885_, _05886_, _05887_, _05888_, _05889_, _05890_, _05891_, _05892_, _05893_, _05894_, _05895_, _05896_, _05897_, _05898_, _05899_, _05900_, _05901_, _05902_, _05903_, _05904_, _05905_, _05906_, _05907_, _05908_, _05909_, _05910_, _05911_, _05912_, _05913_, _05914_, _05915_, _05916_, _05917_, _05918_, _05919_, _05920_, _05921_, _05922_, _05923_, _05924_, _05925_, _05926_, _05927_, _05928_, _05929_, _05930_, _05931_, _05932_, _05933_, _05934_, _05935_, _05936_, _05937_, _05938_, _05939_, _05940_, _05941_, _05942_, _05943_, _05944_, _05945_, _05946_, _05947_, _05948_, _05949_, _05950_, _05951_, _05952_, _05953_, _05954_, _05955_, _05956_, _05957_, _05958_, _05959_, _05960_, _05961_, _05962_, _05963_, _05964_, _05965_, _05966_, _05967_, _05968_, _05969_, _05970_, _05971_, _05972_, _05973_, _05974_, _05975_, _05976_, _05977_, _05978_, _05979_, _05980_, _05981_, _05982_, _05983_, _05984_, _05985_, _05986_, _05987_, _05988_, _05989_, _05990_, _05991_, _05992_, _05993_, _05994_, _05995_, _05996_, _05997_, _05998_, _05999_, _06000_, _06001_, _06002_, _06003_, _06004_, _06005_, _06006_, _06007_, _06008_, _06009_, _06010_, _06011_, _06012_, _06013_, _06014_, _06015_, _06016_, _06017_, _06018_, _06019_, _06020_, _06021_, _06022_, _06023_, _06024_, _06025_, _06026_, _06027_, _06028_, _06029_, _06030_, _06031_, _06032_, _06033_, _06034_, _06035_, _06036_, _06037_, _06038_, _06039_, _06040_, _06041_, _06042_, _06043_, _06044_, _06045_, _06046_, _06047_, _06048_, _06049_, _06050_, _06051_, _06052_, _06053_, _06054_, _06055_, _06056_, _06057_, _06058_, _06059_, _06060_, _06061_, _06062_, _06063_, _06064_, _06065_, _06066_, _06067_, _06068_, _06069_, _06070_, _06071_, _06072_, _06073_, _06074_, _06075_, _06076_, _06077_, _06078_, _06079_, _06080_, _06081_, _06082_, _06083_, _06084_, _06085_, _06086_, _06087_, _06088_, _06089_, _06090_, _06091_, _06092_, _06093_, _06094_, _06095_, _06096_, _06097_, _06098_, _06099_, _06100_, _06101_, _06102_, _06103_, _06104_, _06105_, _06106_, _06107_, _06108_, _06109_, _06110_, _06111_, _06112_, _06113_, _06114_, _06115_, _06116_, _06117_, _06118_, _06119_, _06120_, _06121_, _06122_, _06123_, _06124_, _06125_, _06126_, _06127_, _06128_, _06129_, _06130_, _06131_, _06132_, _06133_, _06134_, _06135_, _06136_, _06137_, _06138_, _06139_, _06140_, _06141_, _06142_, _06143_, _06144_, _06145_, _06146_, _06147_, _06148_, _06149_, _06150_, _06151_, _06152_, _06153_, _06154_, _06155_, _06156_, _06157_, _06158_, _06159_, _06160_, _06161_, _06162_, _06163_, _06164_, _06165_, _06166_, _06167_, _06168_, _06169_, _06170_, _06171_, _06172_, _06173_, _06174_, _06175_, _06176_, _06177_, _06178_, _06179_, _06180_, _06181_, _06182_, _06183_, _06184_, _06185_, _06186_, _06187_, _06188_, _06189_, _06190_, _06191_, _06192_, _06193_, _06194_, _06195_, _06196_, _06197_, _06198_, _06199_, _06200_, _06201_, _06202_, _06203_, _06204_, _06205_, _06206_, _06207_, _06208_, _06209_, _06210_, _06211_, _06212_, _06213_, _06214_, _06215_, _06216_, _06217_, _06218_, _06219_, _06220_, _06221_, _06222_, _06223_, _06224_, _06225_, _06226_, _06227_, _06228_, _06229_, _06230_, _06231_, _06232_, _06233_, _06234_, _06235_, _06236_, _06237_, _06238_, _06239_, _06240_, _06241_, _06242_, _06243_, _06244_, _06245_, _06246_, _06247_, _06248_, _06249_, _06250_, _06251_, _06252_, _06253_, _06254_, _06255_, _06256_, _06257_, _06258_, _06259_, _06260_, _06261_, _06262_, _06263_, _06264_, _06265_, _06266_, _06267_, _06268_, _06269_, _06270_, _06271_, _06272_, _06273_, _06274_, _06275_, _06276_, _06277_, _06278_, _06279_, _06280_, _06281_, _06282_, _06283_, _06284_, _06285_, _06286_, _06287_, _06288_, _06289_, _06290_, _06291_, _06292_, _06293_, _06294_, _06295_, _06296_, _06297_, _06298_, _06299_, _06300_, _06301_, _06302_, _06303_, _06304_, _06305_, _06306_, _06307_, _06308_, _06309_, _06310_, _06311_, _06312_, _06313_, _06314_, _06315_, _06316_, _06317_, _06318_, _06319_, _06320_, _06321_, _06322_, _06323_, _06324_, _06325_, _06326_, _06327_, _06328_, _06329_, _06330_, _06331_, _06332_, _06333_, _06334_, _06335_, _06336_, _06337_, _06338_, _06339_, _06340_, _06341_, _06342_, _06343_, _06344_, _06345_, _06346_, _06347_, _06348_, _06349_, _06350_, _06351_, _06352_, _06353_, _06354_, _06355_, _06356_, _06357_, _06358_, _06359_, _06360_, _06361_, _06362_, _06363_, _06364_, _06365_, _06366_, _06367_, _06368_, _06369_, _06370_, _06371_, _06372_, _06373_, _06374_, _06375_, _06376_, _06377_, _06378_, _06379_, _06380_, _06381_, _06382_, _06383_, _06384_, _06385_, _06386_, _06387_, _06388_, _06389_, _06390_, _06391_, _06392_, _06393_, _06394_, _06395_, _06396_, _06397_, _06398_, _06399_, _06400_, _06401_, _06402_, _06403_, _06404_, _06405_, _06406_, _06407_, _06408_, _06409_, _06410_, _06411_, _06412_, _06413_, _06414_, _06415_, _06416_, _06417_, _06418_, _06419_, _06420_, _06421_, _06422_, _06423_, _06424_, _06425_, _06426_, _06427_, _06428_, _06429_, _06430_, _06431_, _06432_, _06433_, _06434_, _06435_, _06436_, _06437_, _06438_, _06439_, _06440_, _06441_, _06442_, _06443_, _06444_, _06445_, _06446_, _06447_, _06448_, _06449_, _06450_, _06451_, _06452_, _06453_, _06454_, _06455_, _06456_, _06457_, _06458_, _06459_, _06460_, _06461_, _06462_, _06463_, _06464_, _06465_, _06466_, _06467_, _06468_, _06469_, _06470_, _06471_, _06472_, _06473_, _06474_, _06475_, _06476_, _06477_, _06478_, _06479_, _06480_, _06481_, _06482_, _06483_, _06484_, _06485_, _06486_, _06487_, _06488_, _06489_, _06490_, _06491_, _06492_, _06493_, _06494_, _06495_, _06496_, _06497_, _06498_, _06499_, _06500_, _06501_, _06502_, _06503_, _06504_, _06505_, _06506_, _06507_, _06508_, _06509_, _06510_, _06511_, _06512_, _06513_, _06514_, _06515_, _06516_, _06517_, _06518_, _06519_, _06520_, _06521_, _06522_, _06523_, _06524_, _06525_, _06526_, _06527_, _06528_, _06529_, _06530_, _06531_, _06532_, _06533_, _06534_, _06535_, _06536_, _06537_, _06538_, _06539_, _06540_, _06541_, _06542_, _06543_, _06544_, _06545_, _06546_, _06547_, _06548_, _06549_, _06550_, _06551_, _06552_, _06553_, _06554_, _06555_, _06556_, _06557_, _06558_, _06559_, _06560_, _06561_, _06562_, _06563_, _06564_, _06565_, _06566_, _06567_, _06568_, _06569_, _06570_, _06571_, _06572_, _06573_, _06574_, _06575_, _06576_, _06577_, _06578_, _06579_, _06580_, _06581_, _06582_, _06583_, _06584_, _06585_, _06586_, _06587_, _06588_, _06589_, _06590_, _06591_, _06592_, _06593_, _06594_, _06595_, _06596_, _06597_, _06598_, _06599_, _06600_, _06601_, _06602_, _06603_, _06604_, _06605_, _06606_, _06607_, _06608_, _06609_, _06610_, _06611_, _06612_, _06613_, _06614_, _06615_, _06616_, _06617_, _06618_, _06619_, _06620_, _06621_, _06622_, _06623_, _06624_, _06625_, _06626_, _06627_, _06628_, _06629_, _06630_, _06631_, _06632_, _06633_, _06634_, _06635_, _06636_, _06637_, _06638_, _06639_, _06640_, _06641_, _06642_, _06643_, _06644_, _06645_, _06646_, _06647_, _06648_, _06649_, _06650_, _06651_, _06652_, _06653_, _06654_, _06655_, _06656_, _06657_, _06658_, _06659_, _06660_, _06661_, _06662_, _06663_, _06664_, _06665_, _06666_, _06667_, _06668_, _06669_, _06670_, _06671_, _06672_, _06673_, _06674_, _06675_, _06676_, _06677_, _06678_, _06679_, _06680_, _06681_, _06682_, _06683_, _06684_, _06685_, _06686_, _06687_, _06688_, _06689_, _06690_, _06691_, _06692_, _06693_, _06694_, _06695_, _06696_, _06697_, _06698_, _06699_, _06700_, _06701_, _06702_, _06703_, _06704_, _06705_, _06706_, _06707_, _06708_, _06709_, _06710_, _06711_, _06712_, _06713_, _06714_, _06715_, _06716_, _06717_, _06718_, _06719_, _06720_, _06721_, _06722_, _06723_, _06724_, _06725_, _06726_, _06727_, _06728_, _06729_, _06730_, _06731_, _06732_, _06733_, _06734_, _06735_, _06736_, _06737_, _06738_, _06739_, _06740_, _06741_, _06742_, _06743_, _06744_, _06745_, _06746_, _06747_, _06748_, _06749_, _06750_, _06751_, _06752_, _06753_, _06754_, _06755_, _06756_, _06757_, _06758_, _06759_, _06760_, _06761_, _06762_, _06763_, _06764_, _06765_, _06766_, _06767_, _06768_, _06769_, _06770_, _06771_, _06772_, _06773_, _06774_, _06775_, _06776_, _06777_, _06778_, _06779_, _06780_, _06781_, _06782_, _06783_, _06784_, _06785_, _06786_, _06787_, _06788_, _06789_, _06790_, _06791_, _06792_, _06793_, _06794_, _06795_, _06796_, _06797_, _06798_, _06799_, _06800_, _06801_, _06802_, _06803_, _06804_, _06805_, _06806_, _06807_, _06808_, _06809_, _06810_, _06811_, _06812_, _06813_, _06814_, _06815_, _06816_, _06817_, _06818_, _06819_, _06820_, _06821_, _06822_, _06823_, _06824_, _06825_, _06826_, _06827_, _06828_, _06829_, _06830_, _06831_, _06832_, _06833_, _06834_, _06835_, _06836_, _06837_, _06838_, _06839_, _06840_, _06841_, _06842_, _06843_, _06844_, _06845_, _06846_, _06847_, _06848_, _06849_, _06850_, _06851_, _06852_, _06853_, _06854_, _06855_, _06856_, _06857_, _06858_, _06859_, _06860_, _06861_, _06862_, _06863_, _06864_, _06865_, _06866_, _06867_, _06868_, _06869_, _06870_, _06871_, _06872_, _06873_, _06874_, _06875_, _06876_, _06877_, _06878_, _06879_, _06880_, _06881_, _06882_, _06883_, _06884_, _06885_, _06886_, _06887_, _06888_, _06889_, _06890_, _06891_, _06892_, _06893_, _06894_, _06895_, _06896_, _06897_, _06898_, _06899_, _06900_, _06901_, _06902_, _06903_, _06904_, _06905_, _06906_, _06907_, _06908_, _06909_, _06910_, _06911_, _06912_, _06913_, _06914_, _06915_, _06916_, _06917_, _06918_, _06919_, _06920_, _06921_, _06922_, _06923_, _06924_, _06925_, _06926_, _06927_, _06928_, _06929_, _06930_, _06931_, _06932_, _06933_, _06934_, _06935_, _06936_, _06937_, _06938_, _06939_, _06940_, _06941_, _06942_, _06943_, _06944_, _06945_, _06946_, _06947_, _06948_, _06949_, _06950_, _06951_, _06952_, _06953_, _06954_, _06955_, _06956_, _06957_, _06958_, _06959_, _06960_, _06961_, _06962_, _06963_, _06964_, _06965_, _06966_, _06967_, _06968_, _06969_, _06970_, _06971_, _06972_, _06973_, _06974_, _06975_, _06976_, _06977_, _06978_, _06979_, _06980_, _06981_, _06982_, _06983_, _06984_, _06985_, _06986_, _06987_, _06988_, _06989_, _06990_, _06991_, _06992_, _06993_, _06994_, _06995_, _06996_, _06997_, _06998_, _06999_, _07000_, _07001_, _07002_, _07003_, _07004_, _07005_, _07006_, _07007_, _07008_, _07009_, _07010_, _07011_, _07012_, _07013_, _07014_, _07015_, _07016_, _07017_, _07018_, _07019_, _07020_, _07021_, _07022_, _07023_, _07024_, _07025_, _07026_, _07027_, _07028_, _07029_, _07030_, _07031_, _07032_, _07033_, _07034_, _07035_, _07036_, _07037_, _07038_, _07039_, _07040_, _07041_, _07042_, _07043_, _07044_, _07045_, _07046_, _07047_, _07048_, _07049_, _07050_, _07051_, _07052_, _07053_, _07054_, _07055_, _07056_, _07057_, _07058_, _07059_, _07060_, _07061_, _07062_, _07063_, _07064_, _07065_, _07066_, _07067_, _07068_, _07069_, _07070_, _07071_, _07072_, _07073_, _07074_, _07075_, _07076_, _07077_, _07078_, _07079_, _07080_, _07081_, _07082_, _07083_, _07084_, _07085_, _07086_, _07087_, _07088_, _07089_, _07090_, _07091_, _07092_, _07093_, _07094_, _07095_, _07096_, _07097_, _07098_, _07099_, _07100_, _07101_, _07102_, _07103_, _07104_, _07105_, _07106_, _07107_, _07108_, _07109_, _07110_, _07111_, _07112_, _07113_, _07114_, _07115_, _07116_, _07117_, _07118_, _07119_, _07120_, _07121_, _07122_, _07123_, _07124_, _07125_, _07126_, _07127_, _07128_, _07129_, _07130_, _07131_, _07132_, _07133_, _07134_, _07135_, _07136_, _07137_, _07138_, _07139_, _07140_, _07141_, _07142_, _07143_, _07144_, _07145_, _07146_, _07147_, _07148_, _07149_, _07150_, _07151_, _07152_, _07153_, _07154_, _07155_, _07156_, _07157_, _07158_, _07159_, _07160_, _07161_, _07162_, _07163_, _07164_, _07165_, _07166_, _07167_, _07168_, _07169_, _07170_, _07171_, _07172_, _07173_, _07174_, _07175_, _07176_, _07177_, _07178_, _07179_, _07180_, _07181_, _07182_, _07183_, _07184_, _07185_, _07186_, _07187_, _07188_, _07189_, _07190_, _07191_, _07192_, _07193_, _07194_, _07195_, _07196_, _07197_, _07198_, _07199_, _07200_, _07201_, _07202_, _07203_, _07204_, _07205_, _07206_, _07207_, _07208_, _07209_, _07210_, _07211_, _07212_, _07213_, _07214_, _07215_, _07216_, _07217_, _07218_, _07219_, _07220_, _07221_, _07222_, _07223_, _07224_, _07225_, _07226_, _07227_, _07228_, _07229_, _07230_, _07231_, _07232_, _07233_, _07234_, _07235_, _07236_, _07237_, _07238_, _07239_, _07240_, _07241_, _07242_, _07243_, _07244_, _07245_, _07246_, _07247_, _07248_, _07249_, _07250_, _07251_, _07252_, _07253_, _07254_, _07255_, _07256_, _07257_, _07258_, _07259_, _07260_, _07261_, _07262_, _07263_, _07264_, _07265_, _07266_, _07267_, _07268_, _07269_, _07270_, _07271_, _07272_, _07273_, _07274_, _07275_, _07276_, _07277_, _07278_, _07279_, _07280_, _07281_, _07282_, _07283_, _07284_, _07285_, _07286_, _07287_, _07288_, _07289_, _07290_, _07291_, _07292_, _07293_, _07294_, _07295_, _07296_, _07297_, _07298_, _07299_, _07300_, _07301_, _07302_, _07303_, _07304_, _07305_, _07306_, _07307_, _07308_, _07309_, _07310_, _07311_, _07312_, _07313_, _07314_, _07315_, _07316_, _07317_, _07318_, _07319_, _07320_, _07321_, _07322_, _07323_, _07324_, _07325_, _07326_, _07327_, _07328_, _07329_, _07330_, _07331_, _07332_, _07333_, _07334_, _07335_, _07336_, _07337_, _07338_, _07339_, _07340_, _07341_, _07342_, _07343_, _07344_, _07345_, _07346_, _07347_, _07348_, _07349_, _07350_, _07351_, _07352_, _07353_, _07354_, _07355_, _07356_, _07357_, _07358_, _07359_, _07360_, _07361_, _07362_, _07363_, _07364_, _07365_, _07366_, _07367_, _07368_, _07369_, _07370_, _07371_, _07372_, _07373_, _07374_, _07375_, _07376_, _07377_, _07378_, _07379_, _07380_, _07381_, _07382_, _07383_, _07384_, _07385_, _07386_, _07387_, _07388_, _07389_, _07390_, _07391_, _07392_, _07393_, _07394_, _07395_, _07396_, _07397_, _07398_, _07399_, _07400_, _07401_, _07402_, _07403_, _07404_, _07405_, _07406_, _07407_, _07408_, _07409_, _07410_, _07411_, _07412_, _07413_, _07414_, _07415_, _07416_, _07417_, _07418_, _07419_, _07420_, _07421_, _07422_, _07423_, _07424_, _07425_, _07426_, _07427_, _07428_, _07429_, _07430_, _07431_, _07432_, _07433_, _07434_, _07435_, _07436_, _07437_, _07438_, _07439_, _07440_, _07441_, _07442_, _07443_, _07444_, _07445_, _07446_, _07447_, _07448_, _07449_, _07450_, _07451_, _07452_, _07453_, _07454_, _07455_, _07456_, _07457_, _07458_, _07459_, _07460_, _07461_, _07462_, _07463_, _07464_, _07465_, _07466_, _07467_, _07468_, _07469_, _07470_, _07471_, _07472_, _07473_, _07474_, _07475_, _07476_, _07477_, _07478_, _07479_, _07480_, _07481_, _07482_, _07483_, _07484_, _07485_, _07486_, _07487_, _07488_, _07489_, _07490_, _07491_, _07492_, _07493_, _07494_, _07495_, _07496_, _07497_, _07498_, _07499_, _07500_, _07501_, _07502_, _07503_, _07504_, _07505_, _07506_, _07507_, _07508_, _07509_, _07510_, _07511_, _07512_, _07513_, _07514_, _07515_, _07516_, _07517_, _07518_, _07519_, _07520_, _07521_, _07522_, _07523_, _07524_, _07525_, _07526_, _07527_, _07528_, _07529_, _07530_, _07531_, _07532_, _07533_, _07534_, _07535_, _07536_, _07537_, _07538_, _07539_, _07540_, _07541_, _07542_, _07543_, _07544_, _07545_, _07546_, _07547_, _07548_, _07549_, _07550_, _07551_, _07552_, _07553_, _07554_, _07555_, _07556_, _07557_, _07558_, _07559_, _07560_, _07561_, _07562_, _07563_, _07564_, _07565_, _07566_, _07567_, _07568_, _07569_, _07570_, _07571_, _07572_, _07573_, _07574_, _07575_, _07576_, _07577_, _07578_, _07579_, _07580_, _07581_, _07582_, _07583_, _07584_, _07585_, _07586_, _07587_, _07588_, _07589_, _07590_, _07591_, _07592_, _07593_, _07594_, _07595_, _07596_, _07597_, _07598_, _07599_, _07600_, _07601_, _07602_, _07603_, _07604_, _07605_, _07606_, _07607_, _07608_, _07609_, _07610_, _07611_, _07612_, _07613_, _07614_, _07615_, _07616_, _07617_, _07618_, _07619_, _07620_, _07621_, _07622_, _07623_, _07624_, _07625_, _07626_, _07627_, _07628_, _07629_, _07630_, _07631_, _07632_, _07633_, _07634_, _07635_, _07636_, _07637_, _07638_, _07639_, _07640_, _07641_, _07642_, _07643_, _07644_, _07645_, _07646_, _07647_, _07648_, _07649_, _07650_, _07651_, _07652_, _07653_, _07654_, _07655_, _07656_, _07657_, _07658_, _07659_, _07660_, _07661_, _07662_, _07663_, _07664_, _07665_, _07666_, _07667_, _07668_, _07669_, _07670_, _07671_, _07672_, _07673_, _07674_, _07675_, _07676_, _07677_, _07678_, _07679_, _07680_, _07681_, _07682_, _07683_, _07684_, _07685_, _07686_, _07687_, _07688_, _07689_, _07690_, _07691_, _07692_, _07693_, _07694_, _07695_, _07696_, _07697_, _07698_, _07699_, _07700_, _07701_, _07702_, _07703_, _07704_, _07705_, _07706_, _07707_, _07708_, _07709_, _07710_, _07711_, _07712_, _07713_, _07714_, _07715_, _07716_, _07717_, _07718_, _07719_, _07720_, _07721_, _07722_, _07723_, _07724_, _07725_, _07726_, _07727_, _07728_, _07729_, _07730_, _07731_, _07732_, _07733_, _07734_, _07735_, _07736_, _07737_, _07738_, _07739_, _07740_, _07741_, _07742_, _07743_, _07744_, _07745_, _07746_, _07747_, _07748_, _07749_, _07750_, _07751_, _07752_, _07753_, _07754_, _07755_, _07756_, _07757_, _07758_, _07759_, _07760_, _07761_, _07762_, _07763_, _07764_, _07765_, _07766_, _07767_, _07768_, _07769_, _07770_, _07771_, _07772_, _07773_, _07774_, _07775_, _07776_, _07777_, _07778_, _07779_, _07780_, _07781_, _07782_, _07783_, _07784_, _07785_, _07786_, _07787_, _07788_, _07789_, _07790_, _07791_, _07792_, _07793_, _07794_, _07795_, _07796_, _07797_, _07798_, _07799_, _07800_, _07801_, _07802_, _07803_, _07804_, _07805_, _07806_, _07807_, _07808_, _07809_, _07810_, _07811_, _07812_, _07813_, _07814_, _07815_, _07816_, _07817_, _07818_, _07819_, _07820_, _07821_, _07822_, _07823_, _07824_, _07825_, _07826_, _07827_, _07828_, _07829_, _07830_, _07831_, _07832_, _07833_, _07834_, _07835_, _07836_, _07837_, _07838_, _07839_, _07840_, _07841_, _07842_, _07843_, _07844_, _07845_, _07846_, _07847_, _07848_, _07849_, _07850_, _07851_, _07852_, _07853_, _07854_, _07855_, _07856_, _07857_, _07858_, _07859_, _07860_, _07861_, _07862_, _07863_, _07864_, _07865_, _07866_, _07867_, _07868_, _07869_, _07870_, _07871_, _07872_, _07873_, _07874_, _07875_, _07876_, _07877_, _07878_, _07879_, _07880_, _07881_, _07882_, _07883_, _07884_, _07885_, _07886_, _07887_, _07888_, _07889_, _07890_, _07891_, _07892_, _07893_, _07894_, _07895_, _07896_, _07897_, _07898_, _07899_, _07900_, _07901_, _07902_, _07903_, _07904_, _07905_, _07906_, _07907_, _07908_, _07909_, _07910_, _07911_, _07912_, _07913_, _07914_, _07915_, _07916_, _07917_, _07918_, _07919_, _07920_, _07921_, _07922_, _07923_, _07924_, _07925_, _07926_, _07927_, _07928_, _07929_, _07930_, _07931_, _07932_, _07933_, _07934_, _07935_, _07936_, _07937_, _07938_, _07939_, _07940_, _07941_, _07942_, _07943_, _07944_, _07945_, _07946_, _07947_, _07948_, _07949_, _07950_, _07951_, _07952_, _07953_, _07954_, _07955_, _07956_, _07957_, _07958_, _07959_, _07960_, _07961_, _07962_, _07963_, _07964_, _07965_, _07966_, _07967_, _07968_, _07969_, _07970_, _07971_, _07972_, _07973_, _07974_, _07975_, _07976_, _07977_, _07978_, _07979_, _07980_, _07981_, _07982_, _07983_, _07984_, _07985_, _07986_, _07987_, _07988_, _07989_, _07990_, _07991_, _07992_, _07993_, _07994_, _07995_, _07996_, _07997_, _07998_, _07999_, _08000_, _08001_, _08002_, _08003_, _08004_, _08005_, _08006_, _08007_, _08008_, _08009_, _08010_, _08011_, _08012_, _08013_, _08014_, _08015_, _08016_, _08017_, _08018_, _08019_, _08020_, _08021_, _08022_, _08023_, _08024_, _08025_, _08026_, _08027_, _08028_, _08029_, _08030_, _08031_, _08032_, _08033_, _08034_, _08035_, _08036_, _08037_, _08038_, _08039_, _08040_, _08041_, _08042_, _08043_, _08044_, _08045_, _08046_, _08047_, _08048_, _08049_, _08050_, _08051_, _08052_, _08053_, _08054_, _08055_, _08056_, _08057_, _08058_, _08059_, _08060_, _08061_, _08062_, _08063_, _08064_, _08065_, _08066_, _08067_, _08068_, _08069_, _08070_, _08071_, _08072_, _08073_, _08074_, _08075_, _08076_, _08077_, _08078_, _08079_, _08080_, _08081_, _08082_, _08083_, _08084_, _08085_, _08086_, _08087_, _08088_, _08089_, _08090_, _08091_, _08092_, _08093_, _08094_, _08095_, _08096_, _08097_, _08098_, _08099_, _08100_, _08101_, _08102_, _08103_, _08104_, _08105_, _08106_, _08107_, _08108_, _08109_, _08110_, _08111_, _08112_, _08113_, _08114_, _08115_, _08116_, _08117_, _08118_, _08119_, _08120_, _08121_, _08122_, _08123_, _08124_, _08125_, _08126_, _08127_, _08128_, _08129_, _08130_, _08131_, _08132_, _08133_, _08134_, _08135_, _08136_, _08137_, _08138_, _08139_, _08140_, _08141_, _08142_, _08143_, _08144_, _08145_, _08146_, _08147_, _08148_, _08149_, _08150_, _08151_, _08152_, _08153_, _08154_, _08155_, _08156_, _08157_, _08158_, _08159_, _08160_, _08161_, _08162_, _08163_, _08164_, _08165_, _08166_, _08167_, _08168_, _08169_, _08170_, _08171_, _08172_, _08173_, _08174_, _08175_, _08176_, _08177_, _08178_, _08179_, _08180_, _08181_, _08182_, _08183_, _08184_, _08185_, _08186_, _08187_, _08188_, _08189_, _08190_, _08191_, _08192_, _08193_, _08194_, _08195_, _08196_, _08197_, _08198_, _08199_, _08200_, _08201_, _08202_, _08203_, _08204_, _08205_, _08206_, _08207_, _08208_, _08209_, _08210_, _08211_, _08212_, _08213_, _08214_, _08215_, _08216_, _08217_, _08218_, _08219_, _08220_, _08221_, _08222_, _08223_, _08224_, _08225_, _08226_, _08227_, _08228_, _08229_, _08230_, _08231_, _08232_, _08233_, _08234_, _08235_, _08236_, _08237_, _08238_, _08239_, _08240_, _08241_, _08242_, _08243_, _08244_, _08245_, _08246_, _08247_, _08248_, _08249_, _08250_, _08251_, _08252_, _08253_, _08254_, _08255_, _08256_, _08257_, _08258_, _08259_, _08260_, _08261_, _08262_, _08263_, _08264_, _08265_, _08266_, _08267_, _08268_, _08269_, _08270_, _08271_, _08272_, _08273_, _08274_, _08275_, _08276_, _08277_, _08278_, _08279_, _08280_, _08281_, _08282_, _08283_, _08284_, _08285_, _08286_, _08287_, _08288_, _08289_, _08290_, _08291_, _08292_, _08293_, _08294_, _08295_, _08296_, _08297_, _08298_, _08299_, _08300_, _08301_, _08302_, _08303_, _08304_, _08305_, _08306_, _08307_, _08308_, _08309_, _08310_, _08311_, _08312_, _08313_, _08314_, _08315_, _08316_, _08317_, _08318_, _08319_, _08320_, _08321_, _08322_, _08323_, _08324_, _08325_, _08326_, _08327_, _08328_, _08329_, _08330_, _08331_, _08332_, _08333_, _08334_, _08335_, _08336_, _08337_, _08338_, _08339_, _08340_, _08341_, _08342_, _08343_, _08344_, _08345_, _08346_, _08347_, _08348_, _08349_, _08350_, _08351_, _08352_, _08353_, _08354_, _08355_, _08356_, _08357_, _08358_, _08359_, _08360_, _08361_, _08362_, _08363_, _08364_, _08365_, _08366_, _08367_, _08368_, _08369_, _08370_, _08371_, _08372_, _08373_, _08374_, _08375_, _08376_, _08377_, _08378_, _08379_, _08380_, _08381_, _08382_, _08383_, _08384_, _08385_, _08386_, _08387_, _08388_, _08389_, _08390_, _08391_, _08392_, _08393_, _08394_, _08395_, _08396_, _08397_, _08398_, _08399_, _08400_, _08401_, _08402_, _08403_, _08404_, _08405_, _08406_, _08407_, _08408_, _08409_, _08410_, _08411_, _08412_, _08413_, _08414_, _08415_, _08416_, _08417_, _08418_, _08419_, _08420_, _08421_, _08422_, _08423_, _08424_, _08425_, _08426_, _08427_, _08428_, _08429_, _08430_, _08431_, _08432_, _08433_, _08434_, _08435_, _08436_, _08437_, _08438_, _08439_, _08440_, _08441_, _08442_, _08443_, _08444_, _08445_, _08446_, _08447_, _08448_, _08449_, _08450_, _08451_, _08452_, _08453_, _08454_, _08455_, _08456_, _08457_, _08458_, _08459_, _08460_, _08461_, _08462_, _08463_, _08464_, _08465_, _08466_, _08467_, _08468_, _08469_, _08470_, _08471_, _08472_, _08473_, _08474_, _08475_, _08476_, _08477_, _08478_, _08479_, _08480_, _08481_, _08482_, _08483_, _08484_, _08485_, _08486_, _08487_, _08488_, _08489_, _08490_, _08491_, _08492_, _08493_, _08494_, _08495_, _08496_, _08497_, _08498_, _08499_, _08500_, _08501_, _08502_, _08503_, _08504_, _08505_, _08506_, _08507_, _08508_, _08509_, _08510_, _08511_, _08512_, _08513_, _08514_, _08515_, _08516_, _08517_, _08518_, _08519_, _08520_, _08521_, _08522_, _08523_, _08524_, _08525_, _08526_, _08527_, _08528_, _08529_, _08530_, _08531_, _08532_, _08533_, _08534_, _08535_, _08536_, _08537_, _08538_, _08539_, _08540_, _08541_, _08542_, _08543_, _08544_, _08545_, _08546_, _08547_, _08548_, _08549_, _08550_, _08551_, _08552_, _08553_, _08554_, _08555_, _08556_, _08557_, _08558_, _08559_, _08560_, _08561_, _08562_, _08563_, _08564_, _08565_, _08566_, _08567_, _08568_, _08569_, _08570_, _08571_, _08572_, _08573_, _08574_, _08575_, _08576_, _08577_, _08578_, _08579_, _08580_, _08581_, _08582_, _08583_, _08584_, _08585_, _08586_, _08587_, _08588_, _08589_, _08590_, _08591_, _08592_, _08593_, _08594_, _08595_, _08596_, _08597_, _08598_, _08599_, _08600_, _08601_, _08602_, _08603_, _08604_, _08605_, _08606_, _08607_, _08608_, _08609_, _08610_, _08611_, _08612_, _08613_, _08614_, _08615_, _08616_, _08617_, _08618_, _08619_, _08620_, _08621_, _08622_, _08623_, _08624_, _08625_, _08626_, _08627_, _08628_, _08629_, _08630_, _08631_, _08632_, _08633_, _08634_, _08635_, _08636_, _08637_, _08638_, _08639_, _08640_, _08641_, _08642_, _08643_, _08644_, _08645_, _08646_, _08647_, _08648_, _08649_, _08650_, _08651_, _08652_, _08653_, _08654_, _08655_, _08656_, _08657_, _08658_, _08659_, _08660_, _08661_, _08662_, _08663_, _08664_, _08665_, _08666_, _08667_, _08668_, _08669_, _08670_, _08671_, _08672_, _08673_, _08674_, _08675_, _08676_, _08677_, _08678_, _08679_, _08680_, _08681_, _08682_, _08683_, _08684_, _08685_, _08686_, _08687_, _08688_, _08689_, _08690_, _08691_, _08692_, _08693_, _08694_, _08695_, _08696_, _08697_, _08698_, _08699_, _08700_, _08701_, _08702_, _08703_, _08704_, _08705_, _08706_, _08707_, _08708_, _08709_, _08710_, _08711_, _08712_, _08713_, _08714_, _08715_, _08716_, _08717_, _08718_, _08719_, _08720_, _08721_, _08722_, _08723_, _08724_, _08725_, _08726_, _08727_, _08728_, _08729_, _08730_, _08731_, _08732_, _08733_, _08734_, _08735_, _08736_, _08737_, _08738_, _08739_, _08740_, _08741_, _08742_, _08743_, _08744_, _08745_, _08746_, _08747_, _08748_, _08749_, _08750_, _08751_, _08752_, _08753_, _08754_, _08755_, _08756_, _08757_, _08758_, _08759_, _08760_, _08761_, _08762_, _08763_, _08764_, _08765_, _08766_, _08767_, _08768_, _08769_, _08770_, _08771_, _08772_, _08773_, _08774_, _08775_, _08776_, _08777_, _08778_, _08779_, _08780_, _08781_, _08782_, _08783_, _08784_, _08785_, _08786_, _08787_, _08788_, _08789_, _08790_, _08791_, _08792_, _08793_, _08794_, _08795_, _08796_, _08797_, _08798_, _08799_, _08800_, _08801_, _08802_, _08803_, _08804_, _08805_, _08806_, _08807_, _08808_, _08809_, _08810_, _08811_, _08812_, _08813_, _08814_, _08815_, _08816_, _08817_, _08818_, _08819_, _08820_, _08821_, _08822_, _08823_, _08824_, _08825_, _08826_, _08827_, _08828_, _08829_, _08830_, _08831_, _08832_, _08833_, _08834_, _08835_, _08836_, _08837_, _08838_, _08839_, _08840_, _08841_, _08842_, _08843_, _08844_, _08845_, _08846_, _08847_, _08848_, _08849_, _08850_, _08851_, _08852_, _08853_, _08854_, _08855_, _08856_, _08857_, _08858_, _08859_, _08860_, _08861_, _08862_, _08863_, _08864_, _08865_, _08866_, _08867_, _08868_, _08869_, _08870_, _08871_, _08872_, _08873_, _08874_, _08875_, _08876_, _08877_, _08878_, _08879_, _08880_, _08881_, _08882_, _08883_, _08884_, _08885_, _08886_, _08887_, _08888_, _08889_, _08890_, _08891_, _08892_, _08893_, _08894_, _08895_, _08896_, _08897_, _08898_, _08899_, _08900_, _08901_, _08902_, _08903_, _08904_, _08905_, _08906_, _08907_, _08908_, _08909_, _08910_, _08911_, _08912_, _08913_, _08914_, _08915_, _08916_, _08917_, _08918_, _08919_, _08920_, _08921_, _08922_, _08923_, _08924_, _08925_, _08926_, _08927_, _08928_, _08929_, _08930_, _08931_, _08932_, _08933_, _08934_, _08935_, _08936_, _08937_, _08938_, _08939_, _08940_, _08941_, _08942_, _08943_, _08944_, _08945_, _08946_, _08947_, _08948_, _08949_, _08950_, _08951_, _08952_, _08953_, _08954_, _08955_, _08956_, _08957_, _08958_, _08959_, _08960_, _08961_, _08962_, _08963_, _08964_, _08965_, _08966_, _08967_, _08968_, _08969_, _08970_, _08971_, _08972_, _08973_, _08974_, _08975_, _08976_, _08977_, _08978_, _08979_, _08980_, _08981_, _08982_, _08983_, _08984_, _08985_, _08986_, _08987_, _08988_, _08989_, _08990_, _08991_, _08992_, _08993_, _08994_, _08995_, _08996_, _08997_, _08998_, _08999_, _09000_, _09001_, _09002_, _09003_, _09004_, _09005_, _09006_, _09007_, _09008_, _09009_, _09010_, _09011_, _09012_, _09013_, _09014_, _09015_, _09016_, _09017_, _09018_, _09019_, _09020_, _09021_, _09022_, _09023_, _09024_, _09025_, _09026_, _09027_, _09028_, _09029_, _09030_, _09031_, _09032_, _09033_, _09034_, _09035_, _09036_, _09037_, _09038_, _09039_, _09040_, _09041_, _09042_, _09043_, _09044_, _09045_, _09046_, _09047_, _09048_, _09049_, _09050_, _09051_, _09052_, _09053_, _09054_, _09055_, _09056_, _09057_, _09058_, _09059_, _09060_, _09061_, _09062_, _09063_, _09064_, _09065_, _09066_, _09067_, _09068_, _09069_, _09070_, _09071_, _09072_, _09073_, _09074_, _09075_, _09076_, _09077_, _09078_, _09079_, _09080_, _09081_, _09082_, _09083_, _09084_, _09085_, _09086_, _09087_, _09088_, _09089_, _09090_, _09091_, _09092_, _09093_, _09094_, _09095_, _09096_, _09097_, _09098_, _09099_, _09100_, _09101_, _09102_, _09103_, _09104_, _09105_, _09106_, _09107_, _09108_, _09109_, _09110_, _09111_, _09112_, _09113_, _09114_, _09115_, _09116_, _09117_, _09118_, _09119_, _09120_, _09121_, _09122_, _09123_, _09124_, _09125_, _09126_, _09127_, _09128_, _09129_, _09130_, _09131_, _09132_, _09133_, _09134_, _09135_, _09136_, _09137_, _09138_, _09139_, _09140_, _09141_, _09142_, _09143_, _09144_, _09145_, _09146_, _09147_, _09148_, _09149_, _09150_, _09151_, _09152_, _09153_, _09154_, _09155_, _09156_, _09157_, _09158_, _09159_, _09160_, _09161_, _09162_, _09163_, _09164_, _09165_, _09166_, _09167_, _09168_, _09169_, _09170_, _09171_, _09172_, _09173_, _09174_, _09175_, _09176_, _09177_, _09178_, _09179_, _09180_, _09181_, _09182_, _09183_, _09184_, _09185_, _09186_, _09187_, _09188_, _09189_, _09190_, _09191_, _09192_, _09193_, _09194_, _09195_, _09196_, _09197_, _09198_, _09199_, _09200_, _09201_, _09202_, _09203_, _09204_, _09205_, _09206_, _09207_, _09208_, _09209_, _09210_, _09211_, _09212_, _09213_, _09214_, _09215_, _09216_, _09217_, _09218_, _09219_, _09220_, _09221_, _09222_, _09223_, _09224_, _09225_, _09226_, _09227_, _09228_, _09229_, _09230_, _09231_, _09232_, _09233_, _09234_, _09235_, _09236_, _09237_, _09238_, _09239_, _09240_, _09241_, _09242_, _09243_, _09244_, _09245_, _09246_, _09247_, _09248_, _09249_, _09250_, _09251_, _09252_, _09253_, _09254_, _09255_, _09256_, _09257_, _09258_, _09259_, _09260_, _09261_, _09262_, _09263_, _09264_, _09265_, _09266_, _09267_, _09268_, _09269_, _09270_, _09271_, _09272_, _09273_, _09274_, _09275_, _09276_, _09277_, _09278_, _09279_, _09280_, _09281_, _09282_, _09283_, _09284_, _09285_, _09286_, _09287_, _09288_, _09289_, _09290_, _09291_, _09292_, _09293_, _09294_, _09295_, _09296_, _09297_, _09298_, _09299_, _09300_, _09301_, _09302_, _09303_, _09304_, _09305_, _09306_, _09307_, _09308_, _09309_, _09310_, _09311_, _09312_, _09313_, _09314_, _09315_, _09316_, _09317_, _09318_, _09319_, _09320_, _09321_, _09322_, _09323_, _09324_, _09325_, _09326_, _09327_, _09328_, _09329_, _09330_, _09331_, _09332_, _09333_, _09334_, _09335_, _09336_, _09337_, _09338_, _09339_, _09340_, _09341_, _09342_, _09343_, _09344_, _09345_, _09346_, _09347_, _09348_, _09349_, _09350_, _09351_, _09352_, _09353_, _09354_, _09355_, _09356_, _09357_, _09358_, _09359_, _09360_, _09361_, _09362_, _09363_, _09364_, _09365_, _09366_, _09367_, _09368_, _09369_, _09370_, _09371_, _09372_, _09373_, _09374_, _09375_, _09376_, _09377_, _09378_, _09379_, _09380_, _09381_, _09382_, _09383_, _09384_, _09385_, _09386_, _09387_, _09388_, _09389_, _09390_, _09391_, _09392_, _09393_, _09394_, _09395_, _09396_, _09397_, _09398_, _09399_, _09400_, _09401_, _09402_, _09403_, _09404_, _09405_, _09406_, _09407_, _09408_, _09409_, _09410_, _09411_, _09412_, _09413_, _09414_, _09415_, _09416_, _09417_, _09418_, _09419_, _09420_, _09421_, _09422_, _09423_, _09424_, _09425_, _09426_, _09427_, _09428_, _09429_, _09430_, _09431_, _09432_, _09433_, _09434_, _09435_, _09436_, _09437_, _09438_, _09439_, _09440_, _09441_, _09442_, _09443_, _09444_, _09445_, _09446_, _09447_, _09448_, _09449_, _09450_, _09451_, _09452_, _09453_, _09454_, _09455_, _09456_, _09457_, _09458_, _09459_, _09460_, _09461_, _09462_, _09463_, _09464_, _09465_, _09466_, _09467_, _09468_, _09469_, _09470_, _09471_, _09472_, _09473_, _09474_, _09475_, _09476_, _09477_, _09478_, _09479_, _09480_, _09481_, _09482_, _09483_, _09484_, _09485_, _09486_, _09487_, _09488_, _09489_, _09490_, _09491_, _09492_, _09493_, _09494_, _09495_, _09496_, _09497_, _09498_, _09499_, _09500_, _09501_, _09502_, _09503_, _09504_, _09505_, _09506_, _09507_, _09508_, _09509_, _09510_, _09511_, _09512_, _09513_, _09514_, _09515_, _09516_, _09517_, _09518_, _09519_, _09520_, _09521_, _09522_, _09523_, _09524_, _09525_, _09526_, _09527_, _09528_, _09529_, _09530_, _09531_, _09532_, _09533_, _09534_, _09535_, _09536_, _09537_, _09538_, _09539_, _09540_, _09541_, _09542_, _09543_, _09544_, _09545_, _09546_, _09547_, _09548_, _09549_, _09550_, _09551_, _09552_, _09553_, _09554_, _09555_, _09556_, _09557_, _09558_, _09559_, _09560_, _09561_, _09562_, _09563_, _09564_, _09565_, _09566_, _09567_, _09568_, _09569_, _09570_, _09571_, _09572_, _09573_, _09574_, _09575_, _09576_, _09577_, _09578_, _09579_, _09580_, _09581_, _09582_, _09583_, _09584_, _09585_, _09586_, _09587_, _09588_, _09589_, _09590_, _09591_, _09592_, _09593_, _09594_, _09595_, _09596_, _09597_, _09598_, _09599_, _09600_, _09601_, _09602_, _09603_, _09604_, _09605_, _09606_, _09607_, _09608_, _09609_, _09610_, _09611_, _09612_, _09613_, _09614_, _09615_, _09616_, _09617_, _09618_, _09619_, _09620_, _09621_, _09622_, _09623_, _09624_, _09625_, _09626_, _09627_, _09628_, _09629_, _09630_, _09631_, _09632_, _09633_, _09634_, _09635_, _09636_, _09637_, _09638_, _09639_, _09640_, _09641_, _09642_, _09643_, _09644_, _09645_, _09646_, _09647_, _09648_, _09649_, _09650_, _09651_, _09652_, _09653_, _09654_, _09655_, _09656_, _09657_, _09658_, _09659_, _09660_, _09661_, _09662_, _09663_, _09664_, _09665_, _09666_, _09667_, _09668_, _09669_, _09670_, _09671_, _09672_, _09673_, _09674_, _09675_, _09676_, _09677_, _09678_, _09679_, _09680_, _09681_, _09682_, _09683_, _09684_, _09685_, _09686_, _09687_, _09688_, _09689_, _09690_, _09691_, _09692_, _09693_, _09694_, _09695_, _09696_, _09697_, _09698_, _09699_, _09700_, _09701_, _09702_, _09703_, _09704_, _09705_, _09706_, _09707_, _09708_, _09709_, _09710_, _09711_, _09712_, _09713_, _09714_, _09715_, _09716_, _09717_, _09718_, _09719_, _09720_, _09721_, _09722_, _09723_, _09724_, _09725_, _09726_, _09727_, _09728_, _09729_, _09730_, _09731_, _09732_, _09733_, _09734_, _09735_, _09736_, _09737_, _09738_, _09739_, _09740_, _09741_, _09742_, _09743_, _09744_, _09745_, _09746_, _09747_, _09748_, _09749_, _09750_, _09751_, _09752_, _09753_, _09754_, _09755_, _09756_, _09757_, _09758_, _09759_, _09760_, _09761_, _09762_, _09763_, _09764_, _09765_, _09766_, _09767_, _09768_, _09769_, _09770_, _09771_, _09772_, _09773_, _09774_, _09775_, _09776_, _09777_, _09778_, _09779_, _09780_, _09781_, _09782_, _09783_, _09784_, _09785_, _09786_, _09787_, _09788_, _09789_, _09790_, _09791_, _09792_, _09793_, _09794_, _09795_, _09796_, _09797_, _09798_, _09799_, _09800_, _09801_, _09802_, _09803_, _09804_, _09805_, _09806_, _09807_, _09808_, _09809_, _09810_, _09811_, _09812_, _09813_, _09814_, _09815_, _09816_, _09817_, _09818_, _09819_, _09820_, _09821_, _09822_, _09823_, _09824_, _09825_, _09826_, _09827_, _09828_, _09829_, _09830_, _09831_, _09832_, _09833_, _09834_, _09835_, _09836_, _09837_, _09838_, _09839_, _09840_, _09841_, _09842_, _09843_, _09844_, _09845_, _09846_, _09847_, _09848_, _09849_, _09850_, _09851_, _09852_, _09853_, _09854_, _09855_, _09856_, _09857_, _09858_, _09859_, _09860_, _09861_, _09862_, _09863_, _09864_, _09865_, _09866_, _09867_, _09868_, _09869_, _09870_, _09871_, _09872_, _09873_, _09874_, _09875_, _09876_, _09877_, _09878_, _09879_, _09880_, _09881_, _09882_, _09883_, _09884_, _09885_, _09886_, _09887_, _09888_, _09889_, _09890_, _09891_, _09892_, _09893_, _09894_, _09895_, _09896_, _09897_, _09898_, _09899_, _09900_, _09901_, _09902_, _09903_, _09904_, _09905_, _09906_, _09907_, _09908_, _09909_, _09910_, _09911_, _09912_, _09913_, _09914_, _09915_, _09916_, _09917_, _09918_, _09919_, _09920_, _09921_, _09922_, _09923_, _09924_, _09925_, _09926_, _09927_, _09928_, _09929_, _09930_, _09931_, _09932_, _09933_, _09934_, _09935_, _09936_, _09937_, _09938_, _09939_, _09940_, _09941_, _09942_, _09943_, _09944_, _09945_, _09946_, _09947_, _09948_, _09949_, _09950_, _09951_, _09952_, _09953_, _09954_, _09955_, _09956_, _09957_, _09958_, _09959_, _09960_, _09961_, _09962_, _09963_, _09964_, _09965_, _09966_, _09967_, _09968_, _09969_, _09970_, _09971_, _09972_, _09973_, _09974_, _09975_, _09976_, _09977_, _09978_, _09979_, _09980_, _09981_, _09982_, _09983_, _09984_, _09985_, _09986_, _09987_, _09988_, _09989_, _09990_, _09991_, _09992_, _09993_, _09994_, _09995_, _09996_, _09997_, _09998_, _09999_, _10000_, _10001_, _10002_, _10003_, _10004_, _10005_, _10006_, _10007_, _10008_, _10009_, _10010_, _10011_, _10012_, _10013_, _10014_, _10015_, _10016_, _10017_, _10018_, _10019_, _10020_, _10021_, _10022_, _10023_, _10024_, _10025_, _10026_, _10027_, _10028_, _10029_, _10030_, _10031_, _10032_, _10033_, _10034_, _10035_, _10036_, _10037_, _10038_, _10039_, _10040_, _10041_, _10042_, _10043_, _10044_, _10045_, _10046_, _10047_, _10048_, _10049_, _10050_, _10051_, _10052_, _10053_, _10054_, _10055_, _10056_, _10057_, _10058_, _10059_, _10060_, _10061_, _10062_, _10063_, _10064_, _10065_, _10066_, _10067_, _10068_, _10069_, _10070_, _10071_, _10072_, _10073_, _10074_, _10075_, _10076_, _10077_, _10078_, _10079_, _10080_, _10081_, _10082_, _10083_, _10084_, _10085_, _10086_, _10087_, _10088_, _10089_, _10090_, _10091_, _10092_, _10093_, _10094_, _10095_, _10096_, _10097_, _10098_, _10099_, _10100_, _10101_, _10102_, _10103_, _10104_, _10105_, _10106_, _10107_, _10108_, _10109_, _10110_, _10111_, _10112_, _10113_, _10114_, _10115_, _10116_, _10117_, _10118_, _10119_, _10120_, _10121_, _10122_, _10123_, _10124_, _10125_, _10126_, _10127_, _10128_, _10129_, _10130_, _10131_, _10132_, _10133_, _10134_, _10135_, _10136_, _10137_, _10138_, _10139_, _10140_, _10141_, _10142_, _10143_, _10144_, _10145_, _10146_, _10147_, _10148_, _10149_, _10150_, _10151_, _10152_, _10153_, _10154_, _10155_, _10156_, _10157_, _10158_, _10159_, _10160_, _10161_, _10162_, _10163_, _10164_, _10165_, _10166_, _10167_, _10168_, _10169_, _10170_, _10171_, _10172_, _10173_, _10174_, _10175_, _10176_, _10177_, _10178_, _10179_, _10180_, _10181_, _10182_, _10183_, _10184_, _10185_, _10186_, _10187_, _10188_, _10189_, _10190_, _10191_, _10192_, _10193_, _10194_, _10195_, _10196_, _10197_, _10198_, _10199_, _10200_, _10201_, _10202_, _10203_, _10204_, _10205_, _10206_, _10207_, _10208_, _10209_, _10210_, _10211_, _10212_, _10213_, _10214_, _10215_, _10216_, _10217_, _10218_, _10219_, _10220_, _10221_, _10222_, _10223_, _10224_, _10225_, _10226_, _10227_, _10228_, _10229_, _10230_, _10231_, _10232_, _10233_, _10234_, _10235_, _10236_, _10237_, _10238_, _10239_, _10240_, _10241_, _10242_, _10243_, _10244_, _10245_, _10246_, _10247_, _10248_, _10249_, _10250_, _10251_, _10252_, _10253_, _10254_, _10255_, _10256_, _10257_, _10258_, _10259_, _10260_, _10261_, _10262_, _10263_, _10264_, _10265_, _10266_, _10267_, _10268_, _10269_, _10270_, _10271_, _10272_, _10273_, _10274_, _10275_, _10276_, _10277_, _10278_, _10279_, _10280_, _10281_, _10282_, _10283_, _10284_, _10285_, _10286_, _10287_, _10288_, _10289_, _10290_, _10291_, _10292_, _10293_, _10294_, _10295_, _10296_, _10297_, _10298_, _10299_, _10300_, _10301_, _10302_, _10303_, _10304_, _10305_, _10306_, _10307_, _10308_, _10309_, _10310_, _10311_, _10312_, _10313_, _10314_, _10315_, _10316_, _10317_, _10318_, _10319_, _10320_, _10321_, _10322_, _10323_, _10324_, _10325_, _10326_, _10327_, _10328_, _10329_, _10330_, _10331_, _10332_, _10333_, _10334_, _10335_, _10336_, _10337_, _10338_, _10339_, _10340_, _10341_, _10342_, _10343_, _10344_, _10345_, _10346_, _10347_, _10348_, _10349_, _10350_, _10351_, _10352_, _10353_, _10354_, _10355_, _10356_, _10357_, _10358_, _10359_, _10360_, _10361_, _10362_, _10363_, _10364_, _10365_, _10366_, _10367_, _10368_, _10369_, _10370_, _10371_, _10372_, _10373_, _10374_, _10375_, _10376_, _10377_, _10378_, _10379_, _10380_, _10381_, _10382_, _10383_, _10384_, _10385_, _10386_, _10387_, _10388_, _10389_, _10390_, _10391_, _10392_, _10393_, _10394_, _10395_, _10396_, _10397_, _10398_, _10399_, _10400_, _10401_, _10402_, _10403_, _10404_, _10405_, _10406_, _10407_, _10408_, _10409_, _10410_, _10411_, _10412_, _10413_, _10414_, _10415_, _10416_, _10417_, _10418_, _10419_, _10420_, _10421_, _10422_, _10423_, _10424_, _10425_, _10426_, _10427_, _10428_, _10429_, _10430_, _10431_, _10432_, _10433_, _10434_, _10435_, _10436_, _10437_, _10438_, _10439_, _10440_, _10441_, _10442_, _10443_, _10444_, _10445_, _10446_, _10447_, _10448_, _10449_, _10450_, _10451_, _10452_, _10453_, _10454_, _10455_, _10456_, _10457_, _10458_, _10459_, _10460_, _10461_, _10462_, _10463_, _10464_, _10465_, _10466_, _10467_, _10468_, _10469_, _10470_, _10471_, _10472_, _10473_, _10474_, _10475_, _10476_, _10477_, _10478_, _10479_, _10480_, _10481_, _10482_, _10483_, _10484_, _10485_, _10486_, _10487_, _10488_, _10489_, _10490_, _10491_, _10492_, _10493_, _10494_, _10495_, _10496_, _10497_, _10498_, _10499_, _10500_, _10501_, _10502_, _10503_, _10504_, _10505_, _10506_, _10507_, _10508_, _10509_, _10510_, _10511_, _10512_, _10513_, _10514_, _10515_, _10516_, _10517_, _10518_, _10519_, _10520_, _10521_, _10522_, _10523_, _10524_, _10525_, _10526_, _10527_, _10528_, _10529_, _10530_, _10531_, _10532_, _10533_, _10534_, _10535_, _10536_, _10537_, _10538_, _10539_, _10540_, _10541_, _10542_, _10543_, _10544_, _10545_, _10546_, _10547_, _10548_, _10549_, _10550_, _10551_, _10552_, _10553_, _10554_, _10555_, _10556_, _10557_, _10558_, _10559_, _10560_, _10561_, _10562_, _10563_, _10564_, _10565_, _10566_, _10567_, _10568_, _10569_, _10570_, _10571_, _10572_, _10573_, _10574_, _10575_, _10576_, _10577_, _10578_, _10579_, _10580_, _10581_, _10582_, _10583_, _10584_, _10585_, _10586_, _10587_, _10588_, _10589_, _10590_, _10591_, _10592_, _10593_, _10594_, _10595_, _10596_, _10597_, _10598_, _10599_, _10600_, _10601_, _10602_, _10603_, _10604_, _10605_, _10606_, _10607_, _10608_, _10609_, _10610_, _10611_, _10612_, _10613_, _10614_, _10615_, _10616_, _10617_, _10618_, _10619_, _10620_, _10621_, _10622_, _10623_, _10624_, _10625_, _10626_, _10627_, _10628_, _10629_, _10630_, _10631_, _10632_, _10633_, _10634_, _10635_, _10636_, _10637_, _10638_, _10639_, _10640_, _10641_, _10642_, _10643_, _10644_, _10645_, _10646_, _10647_, _10648_, _10649_, _10650_, _10651_, _10652_, _10653_, _10654_, _10655_, _10656_, _10657_, _10658_, _10659_, _10660_, _10661_, _10662_, _10663_, _10664_, _10665_, _10666_, _10667_, _10668_, _10669_, _10670_, _10671_, _10672_, _10673_, _10674_, _10675_, _10676_, _10677_, _10678_, _10679_, _10680_, _10681_, _10682_, _10683_, _10684_, _10685_, _10686_, _10687_, _10688_, _10689_, _10690_, _10691_, _10692_, _10693_, _10694_, _10695_, _10696_, _10697_, _10698_, _10699_, _10700_, _10701_, _10702_, _10703_, _10704_, _10705_, _10706_, _10707_, _10708_, _10709_, _10710_, _10711_, _10712_, _10713_, _10714_, _10715_, _10716_, _10717_, _10718_, _10719_, _10720_, _10721_, _10722_, _10723_, _10724_, _10725_, _10726_, _10727_, _10728_, _10729_, _10730_, _10731_, _10732_, _10733_, _10734_, _10735_, _10736_, _10737_, _10738_, _10739_, _10740_, _10741_, _10742_, _10743_, _10744_, _10745_, _10746_, _10747_, _10748_, _10749_, _10750_, _10751_, _10752_, _10753_, _10754_, _10755_, _10756_, _10757_, _10758_, _10759_, _10760_, _10761_, _10762_, _10763_, _10764_, _10765_, _10766_, _10767_, _10768_, _10769_, _10770_, _10771_, _10772_, _10773_, _10774_, _10775_, _10776_, _10777_, _10778_, _10779_, _10780_, _10781_, _10782_, _10783_, _10784_, _10785_, _10786_, _10787_, _10788_, _10789_, _10790_, _10791_, _10792_, _10793_, _10794_, _10795_, _10796_, _10797_, _10798_, _10799_, _10800_, _10801_, _10802_, _10803_, _10804_, _10805_, _10806_, _10807_, _10808_, _10809_, _10810_, _10811_, _10812_, _10813_, _10814_, _10815_, _10816_, _10817_, _10818_, _10819_, _10820_, _10821_, _10822_, _10823_, _10824_, _10825_, _10826_, _10827_, _10828_, _10829_, _10830_, _10831_, _10832_, _10833_, _10834_, _10835_, _10836_, _10837_, _10838_, _10839_, _10840_, _10841_, _10842_, _10843_, _10844_, _10845_, _10846_, _10847_, _10848_, _10849_, _10850_, _10851_, _10852_, _10853_, _10854_, _10855_, _10856_, _10857_, _10858_, _10859_, _10860_, _10861_, _10862_, _10863_, _10864_, _10865_, _10866_, _10867_, _10868_, _10869_, _10870_, _10871_, _10872_, _10873_, _10874_, _10875_, _10876_, _10877_, _10878_, _10879_, _10880_, _10881_, _10882_, _10883_, _10884_, _10885_, _10886_, _10887_, _10888_, _10889_, _10890_, _10891_, _10892_, _10893_, _10894_, _10895_, _10896_, _10897_, _10898_, _10899_, _10900_, _10901_, _10902_, _10903_, _10904_, _10905_, _10906_, _10907_, _10908_, _10909_, _10910_, _10911_, _10912_, _10913_, _10914_, _10915_, _10916_, _10917_, _10918_, _10919_, _10920_, _10921_, _10922_, _10923_, _10924_, _10925_, _10926_, _10927_, _10928_, _10929_, _10930_, _10931_, _10932_, _10933_, _10934_, _10935_, _10936_, _10937_, _10938_, _10939_, _10940_, _10941_, _10942_, _10943_, _10944_, _10945_, _10946_, _10947_, _10948_, _10949_, _10950_, _10951_, _10952_, _10953_, _10954_, _10955_, _10956_, _10957_, _10958_, _10959_, _10960_, _10961_, _10962_, _10963_, _10964_, _10965_, _10966_, _10967_, _10968_, _10969_, _10970_, _10971_, _10972_, _10973_, _10974_, _10975_, _10976_, _10977_, _10978_, _10979_, _10980_, _10981_, _10982_, _10983_, _10984_, _10985_, _10986_, _10987_, _10988_, _10989_, _10990_, _10991_, _10992_, _10993_, _10994_, _10995_, _10996_, _10997_, _10998_, _10999_, _11000_, _11001_, _11002_, _11003_, _11004_, _11005_, _11006_, _11007_, _11008_, _11009_, _11010_, _11011_, _11012_, _11013_, _11014_, _11015_, _11016_, _11017_, _11018_, _11019_, _11020_, _11021_, _11022_, _11023_, _11024_, _11025_, _11026_, _11027_, _11028_, _11029_, _11030_, _11031_, _11032_, _11033_, _11034_, _11035_, _11036_, _11037_, _11038_, _11039_, _11040_, _11041_, _11042_, _11043_, _11044_, _11045_, _11046_, _11047_, _11048_, _11049_, _11050_, _11051_, _11052_, _11053_, _11054_, _11055_, _11056_, _11057_, _11058_, _11059_, _11060_, _11061_, _11062_, _11063_, _11064_, _11065_, _11066_, _11067_, _11068_, _11069_, _11070_, _11071_, _11072_, _11073_, _11074_, _11075_, _11076_, _11077_, _11078_, _11079_, _11080_, _11081_, _11082_, _11083_, _11084_, _11085_, _11086_, _11087_, _11088_, _11089_, _11090_, _11091_, _11092_, _11093_, _11094_, _11095_, _11096_, _11097_, _11098_, _11099_, _11100_, _11101_, _11102_, _11103_, _11104_, _11105_, _11106_, _11107_, _11108_, _11109_, _11110_, _11111_, _11112_, _11113_, _11114_, _11115_, _11116_, _11117_, _11118_, _11119_, _11120_, _11121_, _11122_, _11123_, _11124_, _11125_, _11126_, _11127_, _11128_, _11129_, _11130_, _11131_, _11132_, _11133_, _11134_, _11135_, _11136_, _11137_, _11138_, _11139_, _11140_, _11141_, _11142_, _11143_, _11144_, _11145_, _11146_, _11147_, _11148_, _11149_, _11150_, _11151_, _11152_, _11153_, _11154_, _11155_, _11156_, _11157_, _11158_, _11159_, _11160_, _11161_, _11162_, _11163_, _11164_, _11165_, _11166_, _11167_, _11168_, _11169_, _11170_, _11171_, _11172_, _11173_, _11174_, _11175_, _11176_, _11177_, _11178_, _11179_, _11180_, _11181_, _11182_, _11183_, _11184_, _11185_, _11186_, _11187_, _11188_, _11189_, _11190_, _11191_, _11192_, _11193_, _11194_, _11195_, _11196_, _11197_, _11198_, _11199_, _11200_, _11201_, _11202_, _11203_, _11204_, _11205_, _11206_, _11207_, _11208_, _11209_, _11210_, _11211_, _11212_, _11213_, _11214_, _11215_, _11216_, _11217_, _11218_, _11219_, _11220_, _11221_, _11222_, _11223_, _11224_, _11225_, _11226_, _11227_, _11228_, _11229_, _11230_, _11231_, _11232_, _11233_, _11234_, _11235_, _11236_, _11237_, _11238_, _11239_, _11240_, _11241_, _11242_, _11243_, _11244_, _11245_, _11246_, _11247_, _11248_, _11249_, _11250_, _11251_, _11252_, _11253_, _11254_, _11255_, _11256_, _11257_, _11258_, _11259_, _11260_, _11261_, _11262_, _11263_, _11264_, _11265_, _11266_, _11267_, _11268_, _11269_, _11270_, _11271_, _11272_, _11273_, _11274_, _11275_, _11276_, _11277_, _11278_, _11279_, _11280_, _11281_, _11282_, _11283_, _11284_, _11285_, _11286_, _11287_, _11288_, _11289_, _11290_, _11291_, _11292_, _11293_, _11294_, _11295_, _11296_, _11297_, _11298_, _11299_, _11300_, _11301_, _11302_, _11303_, _11304_, _11305_, _11306_, _11307_, _11308_, _11309_, _11310_, _11311_, _11312_, _11313_, _11314_, _11315_, _11316_, _11317_, _11318_, _11319_, _11320_, _11321_, _11322_, _11323_, _11324_, _11325_, _11326_, _11327_, _11328_, _11329_, _11330_, _11331_, _11332_, _11333_, _11334_, _11335_, _11336_, _11337_, _11338_, _11339_, _11340_, _11341_, _11342_, _11343_, _11344_, _11345_, _11346_, _11347_, _11348_, _11349_, _11350_, _11351_, _11352_, _11353_, _11354_, _11355_, _11356_, _11357_, _11358_, _11359_, _11360_, _11361_, _11362_, _11363_, _11364_, _11365_, _11366_, _11367_, _11368_, _11369_, _11370_, _11371_, _11372_, _11373_, _11374_, _11375_, _11376_, _11377_, _11378_, _11379_, _11380_, _11381_, _11382_, _11383_, _11384_, _11385_, _11386_, _11387_, _11388_, _11389_, _11390_, _11391_, _11392_, _11393_, _11394_, _11395_, _11396_, _11397_, _11398_, _11399_, _11400_, _11401_, _11402_, _11403_, _11404_, _11405_, _11406_, _11407_, _11408_, _11409_, _11410_, _11411_, _11412_, _11413_, _11414_, _11415_, _11416_, _11417_, _11418_, _11419_, _11420_, _11421_, _11422_, _11423_, _11424_, _11425_, _11426_, _11427_, _11428_, _11429_, _11430_, _11431_, _11432_, _11433_, _11434_, _11435_, _11436_, _11437_, _11438_, _11439_, _11440_, _11441_, _11442_, _11443_, _11444_, _11445_, _11446_, _11447_, _11448_, _11449_, _11450_, _11451_, _11452_, _11453_, _11454_, _11455_, _11456_, _11457_, _11458_, _11459_, _11460_, _11461_, _11462_, _11463_, _11464_, _11465_, _11466_, _11467_, _11468_, _11469_, _11470_, _11471_, _11472_, _11473_, _11474_, _11475_, _11476_, _11477_, _11478_, _11479_, _11480_, _11481_, _11482_, _11483_, _11484_, _11485_, _11486_, _11487_, _11488_, _11489_, _11490_, _11491_, _11492_, _11493_, _11494_, _11495_, _11496_, _11497_, _11498_, _11499_, _11500_, _11501_, _11502_, _11503_, _11504_, _11505_, _11506_, _11507_, _11508_, _11509_, _11510_, _11511_, _11512_, _11513_, _11514_, _11515_, _11516_, _11517_, _11518_, _11519_, _11520_, _11521_, _11522_, _11523_, _11524_, _11525_, _11526_, _11527_, _11528_, _11529_, _11530_, _11531_, _11532_, _11533_, _11534_, _11535_, _11536_, _11537_, _11538_, _11539_, _11540_, _11541_, _11542_, _11543_, _11544_, _11545_, _11546_, _11547_, _11548_, _11549_, _11550_, _11551_, _11552_, _11553_, _11554_, _11555_, _11556_, _11557_, _11558_, _11559_, _11560_, _11561_, _11562_, _11563_, _11564_, _11565_, _11566_, _11567_, _11568_, _11569_, _11570_, _11571_, _11572_, _11573_, _11574_, _11575_, _11576_, _11577_, _11578_, _11579_, _11580_, _11581_, _11582_, _11583_, _11584_, _11585_, _11586_, _11587_, _11588_, _11589_, _11590_, _11591_, _11592_, _11593_, _11594_, _11595_, _11596_, _11597_, _11598_, _11599_, _11600_, _11601_, _11602_, _11603_, _11604_, _11605_, _11606_, _11607_, _11608_, _11609_, _11610_, _11611_, _11612_, _11613_, _11614_, _11615_, _11616_, _11617_, _11618_, _11619_, _11620_, _11621_, _11622_, _11623_, _11624_, _11625_, _11626_, _11627_, _11628_, _11629_, _11630_, _11631_, _11632_, _11633_, _11634_, _11635_, _11636_, _11637_, _11638_, _11639_, _11640_, _11641_, _11642_, _11643_, _11644_, _11645_, _11646_, _11647_, _11648_, _11649_, _11650_, _11651_, _11652_, _11653_, _11654_, _11655_, _11656_, _11657_, _11658_, _11659_, _11660_, _11661_, _11662_, _11663_, _11664_, _11665_, _11666_, _11667_, _11668_, _11669_, _11670_, _11671_, _11672_, _11673_, _11674_, _11675_, _11676_, _11677_, _11678_, _11679_, _11680_, _11681_, _11682_, _11683_, _11684_, _11685_, _11686_, _11687_, _11688_, _11689_, _11690_, _11691_, _11692_, _11693_, _11694_, _11695_, _11696_, _11697_, _11698_, _11699_, _11700_, _11701_, _11702_, _11703_, _11704_, _11705_, _11706_, _11707_, _11708_, _11709_, _11710_, _11711_, _11712_, _11713_, _11714_, _11715_, _11716_, _11717_, _11718_, _11719_, _11720_, _11721_, _11722_, _11723_, _11724_, _11725_, _11726_, _11727_, _11728_, _11729_, _11730_, _11731_, _11732_, _11733_, _11734_, _11735_, _11736_, _11737_, _11738_, _11739_, _11740_, _11741_, _11742_, _11743_, _11744_, _11745_, _11746_, _11747_, _11748_, _11749_, _11750_, _11751_, _11752_, _11753_, _11754_, _11755_, _11756_, _11757_, _11758_, _11759_, _11760_, _11761_, _11762_, _11763_, _11764_, _11765_, _11766_, _11767_, _11768_, _11769_, _11770_, _11771_, _11772_, _11773_, _11774_, _11775_, _11776_, _11777_, _11778_, _11779_, _11780_, _11781_, _11782_, _11783_, _11784_, _11785_, _11786_, _11787_, _11788_, _11789_, _11790_, _11791_, _11792_, _11793_, _11794_, _11795_, _11796_, _11797_, _11798_, _11799_, _11800_, _11801_, _11802_, _11803_, _11804_, _11805_, _11806_, _11807_, _11808_, _11809_, _11810_, _11811_, _11812_, _11813_, _11814_, _11815_, _11816_, _11817_, _11818_, _11819_, _11820_, _11821_, _11822_, _11823_, _11824_, _11825_, _11826_, _11827_, _11828_, _11829_, _11830_, _11831_, _11832_, _11833_, _11834_, _11835_, _11836_, _11837_, _11838_, _11839_, _11840_, _11841_, _11842_, _11843_, _11844_, _11845_, _11846_, _11847_, _11848_, _11849_, _11850_, _11851_, _11852_, _11853_, _11854_, _11855_, _11856_, _11857_, _11858_, _11859_, _11860_, _11861_, _11862_, _11863_, _11864_, _11865_, _11866_, _11867_, _11868_, _11869_, _11870_, _11871_, _11872_, _11873_, _11874_, _11875_, _11876_, _11877_, _11878_, _11879_, _11880_, _11881_, _11882_, _11883_, _11884_, _11885_, _11886_, _11887_, _11888_, _11889_, _11890_, _11891_, _11892_, _11893_, _11894_, _11895_, _11896_, _11897_, _11898_, _11899_, _11900_, _11901_, _11902_, _11903_, _11904_, _11905_, _11906_, _11907_, _11908_, _11909_, _11910_, _11911_, _11912_, _11913_, _11914_, _11915_, _11916_, _11917_, _11918_, _11919_, _11920_, _11921_, _11922_, _11923_, _11924_, _11925_, _11926_, _11927_, _11928_, _11929_, _11930_, _11931_, _11932_, _11933_, _11934_, _11935_, _11936_, _11937_, _11938_, _11939_, _11940_, _11941_, _11942_, _11943_, _11944_, _11945_, _11946_, _11947_, _11948_, _11949_, _11950_, _11951_, _11952_, _11953_, _11954_, _11955_, _11956_, _11957_, _11958_, _11959_, _11960_, _11961_, _11962_, _11963_, _11964_, _11965_, _11966_, _11967_, _11968_, _11969_, _11970_, _11971_, _11972_, _11973_, _11974_, _11975_, _11976_, _11977_, _11978_, _11979_, _11980_, _11981_, _11982_, _11983_, _11984_, _11985_, _11986_, _11987_, _11988_, _11989_, _11990_, _11991_, _11992_, _11993_, _11994_, _11995_, _11996_, _11997_, _11998_, _11999_, _12000_, _12001_, _12002_, _12003_, _12004_, _12005_, _12006_, _12007_, _12008_, _12009_, _12010_, _12011_, _12012_, _12013_, _12014_, _12015_, _12016_, _12017_, _12018_, _12019_, _12020_, _12021_, _12022_, _12023_, _12024_, _12025_, _12026_, _12027_, _12028_, _12029_, _12030_, _12031_, _12032_, _12033_, _12034_, _12035_, _12036_, _12037_, _12038_, _12039_, _12040_, _12041_, _12042_, _12043_, _12044_, _12045_, _12046_, _12047_, _12048_, _12049_, _12050_, _12051_, _12052_, _12053_, _12054_, _12055_, _12056_, _12057_, _12058_, _12059_, _12060_, _12061_, _12062_, _12063_, _12064_, _12065_, _12066_, _12067_, _12068_, _12069_, _12070_, _12071_, _12072_, _12073_, _12074_, _12075_, _12076_, _12077_, _12078_, _12079_, _12080_, _12081_, _12082_, _12083_, _12084_, _12085_, _12086_, _12087_, _12088_, _12089_, _12090_, _12091_, _12092_, _12093_, _12094_, _12095_, _12096_, _12097_, _12098_, _12099_, _12100_, _12101_, _12102_, _12103_, _12104_, _12105_, _12106_, _12107_, _12108_, _12109_, _12110_, _12111_, _12112_, _12113_, _12114_, _12115_, _12116_, _12117_, _12118_, _12119_, _12120_, _12121_, _12122_, _12123_, _12124_, _12125_, _12126_, _12127_, _12128_, _12129_, _12130_, _12131_, _12132_, _12133_, _12134_, _12135_, _12136_, _12137_, _12138_, _12139_, _12140_, _12141_, _12142_, _12143_, _12144_, _12145_, _12146_, _12147_, _12148_, _12149_, _12150_, _12151_, _12152_, _12153_, _12154_, _12155_, _12156_, _12157_, _12158_, _12159_, _12160_, _12161_, _12162_, _12163_, _12164_, _12165_, _12166_, _12167_, _12168_, _12169_, _12170_, _12171_, _12172_, _12173_, _12174_, _12175_, _12176_, _12177_, _12178_, _12179_, _12180_, _12181_, _12182_, _12183_, _12184_, _12185_, _12186_, _12187_, _12188_, _12189_, _12190_, _12191_, _12192_, _12193_, _12194_, _12195_, _12196_, _12197_, _12198_, _12199_, _12200_, _12201_, _12202_, _12203_, _12204_, _12205_, _12206_, _12207_, _12208_, _12209_, _12210_, _12211_, _12212_, _12213_, _12214_, _12215_, _12216_, _12217_, _12218_, _12219_, _12220_, _12221_, _12222_, _12223_, _12224_, _12225_, _12226_, _12227_, _12228_, _12229_, _12230_, _12231_, _12232_, _12233_, _12234_, _12235_, _12236_, _12237_, _12238_, _12239_, _12240_, _12241_, _12242_, _12243_, _12244_, _12245_, _12246_, _12247_, _12248_, _12249_, _12250_, _12251_, _12252_, _12253_, _12254_, _12255_, _12256_, _12257_, _12258_, _12259_, _12260_, _12261_, _12262_, _12263_, _12264_, _12265_, _12266_, _12267_, _12268_, _12269_, _12270_, _12271_, _12272_, _12273_, _12274_, _12275_, _12276_, _12277_, _12278_, _12279_, _12280_, _12281_, _12282_, _12283_, _12284_, _12285_, _12286_, _12287_, _12288_, _12289_, _12290_, _12291_, _12292_, _12293_, _12294_, _12295_, _12296_, _12297_, _12298_, _12299_, _12300_, _12301_, _12302_, _12303_, _12304_, _12305_, _12306_, _12307_, _12308_, _12309_, _12310_, _12311_, _12312_, _12313_, _12314_, _12315_, _12316_, _12317_, _12318_, _12319_, _12320_, _12321_, _12322_, _12323_, _12324_, _12325_, _12326_, _12327_, _12328_, _12329_, _12330_, _12331_, _12332_, _12333_, _12334_, _12335_, _12336_, _12337_, _12338_, _12339_, _12340_, _12341_, _12342_, _12343_, _12344_, _12345_, _12346_, _12347_, _12348_, _12349_, _12350_, _12351_, _12352_, _12353_, _12354_, _12355_, _12356_, _12357_, _12358_, _12359_, _12360_, _12361_, _12362_, _12363_, _12364_, _12365_, _12366_, _12367_, _12368_, _12369_, _12370_, _12371_, _12372_, _12373_, _12374_, _12375_, _12376_, _12377_, _12378_, _12379_, _12380_, _12381_, _12382_, _12383_, _12384_, _12385_, _12386_, _12387_, _12388_, _12389_, _12390_, _12391_, _12392_, _12393_, _12394_, _12395_, _12396_, _12397_, _12398_, _12399_, _12400_, _12401_, _12402_, _12403_, _12404_, _12405_, _12406_, _12407_, _12408_, _12409_, _12410_, _12411_, _12412_, _12413_, _12414_, _12415_, _12416_, _12417_, _12418_, _12419_, _12420_, _12421_, _12422_, _12423_, _12424_, _12425_, _12426_, _12427_, _12428_, _12429_, _12430_, _12431_, _12432_, _12433_, _12434_, _12435_, _12436_, _12437_, _12438_, _12439_, _12440_, _12441_, _12442_, _12443_, _12444_, _12445_, _12446_, _12447_, _12448_, _12449_, _12450_, _12451_, _12452_, _12453_, _12454_, _12455_, _12456_, _12457_, _12458_, _12459_, _12460_, _12461_, _12462_, _12463_, _12464_, _12465_, _12466_, _12467_, _12468_, _12469_, _12470_, _12471_, _12472_, _12473_, _12474_, _12475_, _12476_, _12477_, _12478_, _12479_, _12480_, _12481_, _12482_, _12483_, _12484_, _12485_, _12486_, _12487_, _12488_, _12489_, _12490_, _12491_, _12492_, _12493_, _12494_, _12495_, _12496_, _12497_, _12498_, _12499_, _12500_, _12501_, _12502_, _12503_, _12504_, _12505_, _12506_, _12507_, _12508_, _12509_, _12510_, _12511_, _12512_, _12513_, _12514_, _12515_, _12516_, _12517_, _12518_, _12519_, _12520_, _12521_, _12522_, _12523_, _12524_, _12525_, _12526_, _12527_, _12528_, _12529_, _12530_, _12531_, _12532_, _12533_, _12534_, _12535_, _12536_, _12537_, _12538_, _12539_, _12540_, _12541_, _12542_, _12543_, _12544_, _12545_, _12546_, _12547_, _12548_, _12549_, _12550_, _12551_, _12552_, _12553_, _12554_, _12555_, _12556_, _12557_, _12558_, _12559_, _12560_, _12561_, _12562_, _12563_, _12564_, _12565_, _12566_, _12567_, _12568_, _12569_, _12570_, _12571_, _12572_, _12573_, _12574_, _12575_, _12576_, _12577_, _12578_, _12579_, _12580_, _12581_, _12582_, _12583_, _12584_, _12585_, _12586_, _12587_, _12588_, _12589_, _12590_, _12591_, _12592_, _12593_, _12594_, _12595_, _12596_, _12597_, _12598_, _12599_, _12600_, _12601_, _12602_, _12603_, _12604_, _12605_, _12606_, _12607_, _12608_, _12609_, _12610_, _12611_, _12612_, _12613_, _12614_, _12615_, _12616_, _12617_, _12618_, _12619_, _12620_, _12621_, _12622_, _12623_, _12624_, _12625_, _12626_, _12627_, _12628_, _12629_, _12630_, _12631_, _12632_, _12633_, _12634_, _12635_, _12636_, _12637_, _12638_, _12639_, _12640_, _12641_, _12642_, _12643_, _12644_, _12645_, _12646_, _12647_, _12648_, _12649_, _12650_, _12651_, _12652_, _12653_, _12654_, _12655_, _12656_, _12657_, _12658_, _12659_, _12660_, _12661_, _12662_, _12663_, _12664_, _12665_, _12666_, _12667_, _12668_, _12669_, _12670_, _12671_, _12672_, _12673_, _12674_, _12675_, _12676_, _12677_, _12678_, _12679_, _12680_, _12681_, _12682_, _12683_, _12684_, _12685_, _12686_, _12687_, _12688_, _12689_, _12690_, _12691_, _12692_, _12693_, _12694_, _12695_, _12696_, _12697_, _12698_, _12699_, _12700_, _12701_, _12702_, _12703_, _12704_, _12705_, _12706_, _12707_, _12708_, _12709_, _12710_, _12711_, _12712_, _12713_, _12714_, _12715_, _12716_, _12717_, _12718_, _12719_, _12720_, _12721_, _12722_, _12723_, _12724_, _12725_, _12726_, _12727_, _12728_, _12729_, _12730_, _12731_, _12732_, _12733_, _12734_, _12735_, _12736_, _12737_, _12738_, _12739_, _12740_, _12741_, _12742_, _12743_, _12744_, _12745_, _12746_, _12747_, _12748_, _12749_, _12750_, _12751_, _12752_, _12753_, _12754_, _12755_, _12756_, _12757_, _12758_, _12759_, _12760_, _12761_, _12762_, _12763_, _12764_, _12765_, _12766_, _12767_, _12768_, _12769_, _12770_, _12771_, _12772_, _12773_, _12774_, _12775_, _12776_, _12777_, _12778_, _12779_, _12780_, _12781_, _12782_, _12783_, _12784_, _12785_, _12786_, _12787_, _12788_, _12789_, _12790_, _12791_, _12792_, _12793_, _12794_, _12795_, _12796_, _12797_, _12798_, _12799_, _12800_, _12801_, _12802_, _12803_, _12804_, _12805_, _12806_, _12807_, _12808_, _12809_, _12810_, _12811_, _12812_, _12813_, _12814_, _12815_, _12816_, _12817_, _12818_, _12819_, _12820_, _12821_, _12822_, _12823_, _12824_, _12825_, _12826_, _12827_, _12828_, _12829_, _12830_, _12831_, _12832_, _12833_, _12834_, _12835_, _12836_, _12837_, _12838_, _12839_, _12840_, _12841_, _12842_, _12843_, _12844_, _12845_, _12846_, _12847_, _12848_, _12849_, _12850_, _12851_, _12852_, _12853_, _12854_, _12855_, _12856_, _12857_, _12858_, _12859_, _12860_, _12861_, _12862_, _12863_, _12864_, _12865_, _12866_, _12867_, _12868_, _12869_, _12870_, _12871_, _12872_, _12873_, _12874_, _12875_, _12876_, _12877_, _12878_, _12879_, _12880_, _12881_, _12882_, _12883_, _12884_, _12885_, _12886_, _12887_, _12888_, _12889_, _12890_, _12891_, _12892_, _12893_, _12894_, _12895_, _12896_, _12897_, _12898_, _12899_, _12900_, _12901_, _12902_, _12903_, _12904_, _12905_, _12906_, _12907_, _12908_, _12909_, _12910_, _12911_, _12912_, _12913_, _12914_, _12915_, _12916_, _12917_, _12918_, _12919_, _12920_, _12921_, _12922_, _12923_, _12924_, _12925_, _12926_, _12927_, _12928_, _12929_, _12930_, _12931_, _12932_, _12933_, _12934_, _12935_, _12936_, _12937_, _12938_, _12939_, _12940_, _12941_, _12942_, _12943_, _12944_, _12945_, _12946_, _12947_, _12948_, _12949_, _12950_, _12951_, _12952_, _12953_, _12954_, _12955_, _12956_, _12957_, _12958_, _12959_, _12960_, _12961_, _12962_, _12963_, _12964_, _12965_, _12966_, _12967_, _12968_, _12969_, _12970_, _12971_, _12972_, _12973_, _12974_, _12975_, _12976_, _12977_, _12978_, _12979_, _12980_, _12981_, _12982_, _12983_, _12984_, _12985_, _12986_, _12987_, _12988_, _12989_, _12990_, _12991_, _12992_, _12993_, _12994_, _12995_, _12996_, _12997_, _12998_, _12999_, _13000_, _13001_, _13002_, _13003_, _13004_, _13005_, _13006_, _13007_, _13008_, _13009_, _13010_, _13011_, _13012_, _13013_, _13014_, _13015_, _13016_, _13017_, _13018_, _13019_, _13020_, _13021_, _13022_, _13023_, _13024_, _13025_, _13026_, _13027_, _13028_, _13029_, _13030_, _13031_, _13032_, _13033_, _13034_, _13035_, _13036_, _13037_, _13038_, _13039_, _13040_, _13041_, _13042_, _13043_, _13044_, _13045_, _13046_, _13047_, _13048_, _13049_, _13050_, _13051_, _13052_, _13053_, _13054_, _13055_, _13056_, _13057_, _13058_, _13059_, _13060_, _13061_, _13062_, _13063_, _13064_, _13065_, _13066_, _13067_, _13068_, _13069_, _13070_, _13071_, _13072_, _13073_, _13074_, _13075_, _13076_, _13077_, _13078_, _13079_, _13080_, _13081_, _13082_, _13083_, _13084_, _13085_, _13086_, _13087_, _13088_, _13089_, _13090_, _13091_, _13092_, _13093_, _13094_, _13095_, _13096_, _13097_, _13098_, _13099_, _13100_, _13101_, _13102_, _13103_, _13104_, _13105_, _13106_, _13107_, _13108_, _13109_, _13110_, _13111_, _13112_, _13113_, _13114_, _13115_, _13116_, _13117_, _13118_, _13119_, _13120_, _13121_, _13122_, _13123_, _13124_, _13125_, _13126_, _13127_, _13128_, _13129_, _13130_, _13131_, _13132_, _13133_, _13134_, _13135_, _13136_, _13137_, _13138_, _13139_, _13140_, _13141_, _13142_, _13143_, _13144_, _13145_, _13146_, _13147_, _13148_, _13149_, _13150_, _13151_, _13152_, _13153_, _13154_, _13155_, _13156_, _13157_, _13158_, _13159_, _13160_, _13161_, _13162_, _13163_, _13164_, _13165_, _13166_, _13167_, _13168_, _13169_, _13170_, _13171_, _13172_, _13173_, _13174_, _13175_, _13176_, _13177_, _13178_, _13179_, _13180_, _13181_, _13182_, _13183_, _13184_, _13185_, _13186_, _13187_, _13188_, _13189_, _13190_, _13191_, _13192_, _13193_, _13194_, _13195_, _13196_, _13197_, _13198_, _13199_, _13200_, _13201_, _13202_, _13203_, _13204_, _13205_, _13206_, _13207_, _13208_, _13209_, _13210_, _13211_, _13212_, _13213_, _13214_, _13215_, _13216_, _13217_, _13218_, _13219_, _13220_, _13221_, _13222_, _13223_, _13224_, _13225_, _13226_, _13227_, _13228_, _13229_, _13230_, _13231_, _13232_, _13233_, _13234_, _13235_, _13236_, _13237_, _13238_, _13239_, _13240_, _13241_, _13242_, _13243_, _13244_, _13245_, _13246_, _13247_, _13248_, _13249_, _13250_, _13251_, _13252_, _13253_, _13254_, _13255_, _13256_, _13257_, _13258_, _13259_, _13260_, _13261_, _13262_, _13263_, _13264_, _13265_, _13266_, _13267_, _13268_, _13269_, _13270_, _13271_, _13272_, _13273_, _13274_, _13275_, _13276_, _13277_, _13278_, _13279_, _13280_, _13281_, _13282_, _13283_, _13284_, _13285_, _13286_, _13287_, _13288_, _13289_, _13290_, _13291_, _13292_, _13293_, _13294_, _13295_, _13296_, _13297_, _13298_, _13299_, _13300_, _13301_, _13302_, _13303_, _13304_, _13305_, _13306_, _13307_, _13308_, _13309_, _13310_, _13311_, _13312_, _13313_, _13314_, _13315_, _13316_, _13317_, _13318_, _13319_, _13320_, _13321_, _13322_, _13323_, _13324_, _13325_, _13326_, _13327_, _13328_, _13329_, _13330_, _13331_, _13332_, _13333_, _13334_, _13335_, _13336_, _13337_, _13338_, _13339_, _13340_, _13341_, _13342_, _13343_, _13344_, _13345_, _13346_, _13347_, _13348_, _13349_, _13350_, _13351_, _13352_, _13353_, _13354_, _13355_, _13356_, _13357_, _13358_, _13359_, _13360_, _13361_, _13362_, _13363_, _13364_, _13365_, _13366_, _13367_, _13368_, _13369_, _13370_, _13371_, _13372_, _13373_, _13374_, _13375_, _13376_, _13377_, _13378_, _13379_, _13380_, _13381_, _13382_, _13383_, _13384_, _13385_, _13386_, _13387_, _13388_, _13389_, _13390_, _13391_, _13392_, _13393_, _13394_, _13395_, _13396_, _13397_, _13398_, _13399_, _13400_, _13401_, _13402_, _13403_, _13404_, _13405_, _13406_, _13407_, _13408_, _13409_, _13410_, _13411_, _13412_, _13413_, _13414_, _13415_, _13416_, _13417_, _13418_, _13419_, _13420_, _13421_, _13422_, _13423_, _13424_, _13425_, _13426_, _13427_, _13428_, _13429_, _13430_, _13431_, _13432_, _13433_, _13434_, _13435_, _13436_, _13437_, _13438_, _13439_, _13440_, _13441_, _13442_, _13443_, _13444_, _13445_, _13446_, _13447_, _13448_, _13449_, _13450_, _13451_, _13452_, _13453_, _13454_, _13455_, _13456_, _13457_, _13458_, _13459_, _13460_, _13461_, _13462_, _13463_, _13464_, _13465_, _13466_, _13467_, _13468_, _13469_, _13470_, _13471_, _13472_, _13473_, _13474_, _13475_, _13476_, _13477_, _13478_, _13479_, _13480_, _13481_, _13482_, _13483_, _13484_, _13485_, _13486_, _13487_, _13488_, _13489_, _13490_, _13491_, _13492_, _13493_, _13494_, _13495_, _13496_, _13497_, _13498_, _13499_, _13500_, _13501_, _13502_, _13503_, _13504_, _13505_, _13506_, _13507_, _13508_, _13509_, _13510_, _13511_, _13512_, _13513_, _13514_, _13515_, _13516_, _13517_, _13518_, _13519_, _13520_, _13521_, _13522_, _13523_, _13524_, _13525_, _13526_, _13527_, _13528_, _13529_, _13530_, _13531_, _13532_, _13533_, _13534_, _13535_, _13536_, _13537_, _13538_, _13539_, _13540_, _13541_, _13542_, _13543_, _13544_, _13545_, _13546_, _13547_, _13548_, _13549_, _13550_, _13551_, _13552_, _13553_, _13554_, _13555_, _13556_, _13557_, _13558_, _13559_, _13560_, _13561_, _13562_, _13563_, _13564_, _13565_, _13566_, _13567_, _13568_, _13569_, _13570_, _13571_, _13572_, _13573_, _13574_, _13575_, _13576_, _13577_, _13578_, _13579_, _13580_, _13581_, _13582_, _13583_, _13584_, _13585_, _13586_, _13587_, _13588_, _13589_, _13590_, _13591_, _13592_, _13593_, _13594_, _13595_, _13596_, _13597_, _13598_, _13599_, _13600_, _13601_, _13602_, _13603_, _13604_, _13605_, _13606_, _13607_, _13608_, _13609_, _13610_, _13611_, _13612_, _13613_, _13614_, _13615_, _13616_, _13617_, _13618_, _13619_, _13620_, _13621_, _13622_, _13623_, _13624_, _13625_, _13626_, _13627_, _13628_, _13629_, _13630_, _13631_, _13632_, _13633_, _13634_, _13635_, _13636_, _13637_, _13638_, _13639_, _13640_, _13641_, _13642_, _13643_, _13644_, _13645_, _13646_, _13647_, _13648_, _13649_, _13650_, _13651_, _13652_, _13653_, _13654_, _13655_, _13656_, _13657_, _13658_, _13659_, _13660_, _13661_, _13662_, _13663_, _13664_, _13665_, _13666_, _13667_, _13668_, _13669_, _13670_, _13671_, _13672_, _13673_, _13674_, _13675_, _13676_, _13677_, _13678_, _13679_, _13680_, _13681_, _13682_, _13683_, _13684_, _13685_, _13686_, _13687_, _13688_, _13689_, _13690_, _13691_, _13692_, _13693_, _13694_, _13695_, _13696_, _13697_, _13698_, _13699_, _13700_, _13701_, _13702_, _13703_, _13704_, _13705_, _13706_, _13707_, _13708_, _13709_, _13710_, _13711_, _13712_, _13713_, _13714_, _13715_, _13716_, _13717_, _13718_, _13719_, _13720_, _13721_, _13722_, _13723_, _13724_, _13725_, _13726_, _13727_, _13728_, _13729_, _13730_, _13731_, _13732_, _13733_, _13734_, _13735_, _13736_, _13737_, _13738_, _13739_, _13740_, _13741_, _13742_, _13743_, _13744_, _13745_, _13746_, _13747_, _13748_, _13749_, _13750_, _13751_, _13752_, _13753_, _13754_, _13755_, _13756_, _13757_, _13758_, _13759_, _13760_, _13761_, _13762_, _13763_, _13764_, _13765_, _13766_, _13767_, _13768_, _13769_, _13770_, _13771_, _13772_, _13773_, _13774_, _13775_, _13776_, _13777_, _13778_, _13779_, _13780_, _13781_, _13782_, _13783_, _13784_, _13785_, _13786_, _13787_, _13788_, _13789_, _13790_, _13791_, _13792_, _13793_, _13794_, _13795_, _13796_, _13797_, _13798_, _13799_, _13800_, _13801_, _13802_, _13803_, _13804_, _13805_, _13806_, _13807_, _13808_, _13809_, _13810_, _13811_, _13812_, _13813_, _13814_, _13815_, _13816_, _13817_, _13818_, _13819_, _13820_, _13821_, _13822_, _13823_, _13824_, _13825_, _13826_, _13827_, _13828_, _13829_, _13830_, _13831_, _13832_, _13833_, _13834_, _13835_, _13836_, _13837_, _13838_, _13839_, _13840_, _13841_, _13842_, _13843_, _13844_, _13845_, _13846_, _13847_, _13848_, _13849_, _13850_, _13851_, _13852_, _13853_, _13854_, _13855_, _13856_, _13857_, _13858_, _13859_, _13860_, _13861_, _13862_, _13863_, _13864_, _13865_, _13866_, _13867_, _13868_, _13869_, _13870_, _13871_, _13872_, _13873_, _13874_, _13875_, _13876_, _13877_, _13878_, _13879_, _13880_, _13881_, _13882_, _13883_, _13884_, _13885_, _13886_, _13887_, _13888_, _13889_, _13890_, _13891_, _13892_, _13893_, _13894_, _13895_, _13896_, _13897_, _13898_, _13899_, _13900_, _13901_, _13902_, _13903_, _13904_, _13905_, _13906_, _13907_, _13908_, _13909_, _13910_, _13911_, _13912_, _13913_, _13914_, _13915_, _13916_, _13917_, _13918_, _13919_, _13920_, _13921_, _13922_, _13923_, _13924_, _13925_, _13926_, _13927_, _13928_, _13929_, _13930_, _13931_, _13932_, _13933_, _13934_, _13935_, _13936_, _13937_, _13938_, _13939_, _13940_, _13941_, _13942_, _13943_, _13944_, _13945_, _13946_, _13947_, _13948_, _13949_, _13950_, _13951_, _13952_, _13953_, _13954_, _13955_, _13956_, _13957_, _13958_, _13959_, _13960_, _13961_, _13962_, _13963_, _13964_, _13965_, _13966_, _13967_, _13968_, _13969_, _13970_, _13971_, _13972_, _13973_, _13974_, _13975_, _13976_, _13977_, _13978_, _13979_, _13980_, _13981_, _13982_, _13983_, _13984_, _13985_, _13986_, _13987_, _13988_, _13989_, _13990_, _13991_, _13992_, _13993_, _13994_, _13995_, _13996_, _13997_, _13998_, _13999_, _14000_, _14001_, _14002_, _14003_, _14004_, _14005_, _14006_, _14007_, _14008_, _14009_, _14010_, _14011_, _14012_, _14013_, _14014_, _14015_, _14016_, _14017_, _14018_, _14019_, _14020_, _14021_, _14022_, _14023_, _14024_, _14025_, _14026_, _14027_, _14028_, _14029_, _14030_, _14031_, _14032_, _14033_, _14034_, _14035_, _14036_, _14037_, _14038_, _14039_, _14040_, _14041_, _14042_, _14043_, _14044_, _14045_, _14046_, _14047_, _14048_, _14049_, _14050_, _14051_, _14052_, _14053_, _14054_, _14055_, _14056_, _14057_, _14058_, _14059_, _14060_, _14061_, _14062_, _14063_, _14064_, _14065_, _14066_, _14067_, _14068_, _14069_, _14070_, _14071_, _14072_, _14073_, _14074_, _14075_, _14076_, _14077_, _14078_, _14079_, _14080_, _14081_, _14082_, _14083_, _14084_, _14085_, _14086_, _14087_, _14088_, _14089_, _14090_, _14091_, _14092_, _14093_, _14094_, _14095_, _14096_, _14097_, _14098_, _14099_, _14100_, _14101_, _14102_, _14103_, _14104_, _14105_, _14106_, _14107_, _14108_, _14109_, _14110_, _14111_, _14112_, _14113_, _14114_, _14115_, _14116_, _14117_, _14118_, _14119_, _14120_, _14121_, _14122_, _14123_, _14124_, _14125_, _14126_, _14127_, _14128_, _14129_, _14130_, _14131_, _14132_, _14133_, _14134_, _14135_, _14136_, _14137_, _14138_, _14139_, _14140_, _14141_, _14142_, _14143_, _14144_, _14145_, _14146_, _14147_, _14148_, _14149_, _14150_, _14151_, _14152_, _14153_, _14154_, _14155_, _14156_, _14157_, _14158_, _14159_, _14160_, _14161_, _14162_, _14163_, _14164_, _14165_, _14166_, _14167_, _14168_, _14169_, _14170_, _14171_, _14172_, _14173_, _14174_, _14175_, _14176_, _14177_, _14178_, _14179_, _14180_, _14181_, _14182_, _14183_, _14184_, _14185_, _14186_, _14187_, _14188_, _14189_, _14190_, _14191_, _14192_, _14193_, _14194_, _14195_, _14196_, _14197_, _14198_, _14199_, _14200_, _14201_, _14202_, _14203_, _14204_, _14205_, _14206_, _14207_, _14208_, _14209_, _14210_, _14211_, _14212_, _14213_, _14214_, _14215_, _14216_, _14217_, _14218_, _14219_, _14220_, _14221_, _14222_, _14223_, _14224_, _14225_, _14226_, _14227_, _14228_, _14229_, _14230_, _14231_, _14232_, _14233_, _14234_, _14235_, _14236_, _14237_, _14238_, _14239_, _14240_, _14241_, _14242_, _14243_, _14244_, _14245_, _14246_, _14247_, _14248_, _14249_, _14250_, _14251_, _14252_, _14253_, _14254_, _14255_, _14256_, _14257_, _14258_, _14259_, _14260_, _14261_, _14262_, _14263_, _14264_, _14265_, _14266_, _14267_, _14268_, _14269_, _14270_, _14271_, _14272_, _14273_, _14274_, _14275_, _14276_, _14277_, _14278_, _14279_, _14280_, _14281_, _14282_, _14283_, _14284_, _14285_, _14286_, _14287_, _14288_, _14289_, _14290_, _14291_, _14292_, _14293_, _14294_, _14295_, _14296_, _14297_, _14298_, _14299_, _14300_, _14301_, _14302_, _14303_, _14304_, _14305_, _14306_, _14307_, _14308_, _14309_, _14310_, _14311_, _14312_, _14313_, _14314_, _14315_, _14316_, _14317_, _14318_, _14319_, _14320_, _14321_, _14322_, _14323_, _14324_, _14325_, _14326_, _14327_, _14328_, _14329_, _14330_, _14331_, _14332_, _14333_, _14334_, _14335_, _14336_, _14337_, _14338_, _14339_, _14340_, _14341_, _14342_, _14343_, _14344_, _14345_, _14346_, _14347_, _14348_, _14349_, _14350_, _14351_, _14352_, _14353_, _14354_, _14355_, _14356_, _14357_, _14358_, _14359_, _14360_, _14361_, _14362_, _14363_, _14364_, _14365_, _14366_, _14367_, _14368_, _14369_, _14370_, _14371_, _14372_, _14373_, _14374_, _14375_, _14376_, _14377_, _14378_, _14379_, _14380_, _14381_, _14382_, _14383_, _14384_, _14385_, _14386_, _14387_, _14388_, _14389_, _14390_, _14391_, _14392_, _14393_, _14394_, _14395_, _14396_, _14397_, _14398_, _14399_, _14400_, _14401_, _14402_, _14403_, _14404_, _14405_, _14406_, _14407_, _14408_, _14409_, _14410_, _14411_, _14412_, _14413_, _14414_, _14415_, _14416_, _14417_, _14418_, _14419_, _14420_, _14421_, _14422_, _14423_, _14424_, _14425_, _14426_, _14427_, _14428_, _14429_, _14430_, _14431_, _14432_, _14433_, _14434_, _14435_, _14436_, _14437_, _14438_, _14439_, _14440_, _14441_, _14442_, _14443_, _14444_, _14445_, _14446_, _14447_, _14448_, _14449_, _14450_, _14451_, _14452_, _14453_, _14454_, _14455_, _14456_, _14457_, _14458_, _14459_, _14460_, _14461_, _14462_, _14463_, _14464_, _14465_, _14466_, _14467_, _14468_, _14469_, _14470_, _14471_, _14472_, _14473_, _14474_, _14475_, _14476_, _14477_, _14478_, _14479_, _14480_, _14481_, _14482_, _14483_, _14484_, _14485_, _14486_, _14487_, _14488_, _14489_, _14490_, _14491_, _14492_, _14493_, _14494_, _14495_, _14496_, _14497_, _14498_, _14499_, _14500_, _14501_, _14502_, _14503_, _14504_, _14505_, _14506_, _14507_, _14508_, _14509_, _14510_, _14511_, _14512_, _14513_, _14514_, _14515_, _14516_, _14517_, _14518_, _14519_, _14520_, _14521_, _14522_, _14523_, _14524_, _14525_, _14526_, _14527_, _14528_, _14529_, _14530_, _14531_, _14532_, _14533_, _14534_, _14535_, _14536_, _14537_, _14538_, _14539_, _14540_, _14541_, _14542_, _14543_, _14544_, _14545_, _14546_, _14547_, _14548_, _14549_, _14550_, _14551_, _14552_, _14553_, _14554_, _14555_, _14556_, _14557_, _14558_, _14559_, _14560_, _14561_, _14562_, _14563_, _14564_, _14565_, _14566_, _14567_, _14568_, _14569_, _14570_, _14571_, _14572_, _14573_, _14574_, _14575_, _14576_, _14577_, _14578_, _14579_, _14580_, _14581_, _14582_, _14583_, _14584_, _14585_, _14586_, _14587_, _14588_, _14589_, _14590_, _14591_, _14592_, _14593_, _14594_, _14595_, _14596_, _14597_, _14598_, _14599_, _14600_, _14601_, _14602_, _14603_, _14604_, _14605_, _14606_, _14607_, _14608_, _14609_, _14610_, _14611_, _14612_, _14613_, _14614_, _14615_, _14616_, _14617_, _14618_, _14619_, _14620_, _14621_, _14622_, _14623_, _14624_, _14625_, _14626_, _14627_, _14628_, _14629_, _14630_, _14631_, _14632_, _14633_, _14634_, _14635_, _14636_, _14637_, _14638_, _14639_, _14640_, _14641_, _14642_, _14643_, _14644_, _14645_, _14646_, _14647_, _14648_, _14649_, _14650_, _14651_, _14652_, _14653_, _14654_, _14655_, _14656_, _14657_, _14658_, _14659_, _14660_, _14661_, _14662_, _14663_, _14664_, _14665_, _14666_, _14667_, _14668_, _14669_, _14670_, _14671_, _14672_, _14673_, _14674_, _14675_, _14676_, _14677_, _14678_, _14679_, _14680_, _14681_, _14682_, _14683_, _14684_, _14685_, _14686_, _14687_, _14688_, _14689_, _14690_, _14691_, _14692_, _14693_, _14694_, _14695_, _14696_, _14697_, _14698_, _14699_, _14700_, _14701_, _14702_, _14703_, _14704_, _14705_, _14706_, _14707_, _14708_, _14709_, _14710_, _14711_, _14712_, _14713_, _14714_, _14715_, _14716_, _14717_, _14718_, _14719_, _14720_, _14721_, _14722_, _14723_, _14724_, _14725_, _14726_, _14727_, _14728_, _14729_, _14730_, _14731_, _14732_, _14733_, _14734_, _14735_, _14736_, _14737_, _14738_, _14739_, _14740_, _14741_, _14742_, _14743_, _14744_, _14745_, _14746_, _14747_, _14748_, _14749_, _14750_, _14751_, _14752_, _14753_, _14754_, _14755_, _14756_, _14757_, _14758_, _14759_, _14760_, _14761_, _14762_, _14763_, _14764_, _14765_, _14766_, _14767_, _14768_, _14769_, _14770_, _14771_, _14772_, _14773_, _14774_, _14775_, _14776_, _14777_, _14778_, _14779_, _14780_, _14781_, _14782_, _14783_, _14784_, _14785_, _14786_, _14787_, _14788_, _14789_, _14790_, _14791_, _14792_, _14793_, _14794_, _14795_, _14796_, _14797_, _14798_, _14799_, _14800_, _14801_, _14802_, _14803_, _14804_, _14805_, _14806_, _14807_, _14808_, _14809_, _14810_, _14811_, _14812_, _14813_, _14814_, _14815_, _14816_, _14817_, _14818_, _14819_, _14820_, _14821_, _14822_, _14823_, _14824_, _14825_, _14826_, _14827_, _14828_, _14829_, _14830_, _14831_, _14832_, _14833_, _14834_, _14835_, _14836_, _14837_, _14838_, _14839_, _14840_, _14841_, _14842_, _14843_, _14844_, _14845_, _14846_, _14847_, _14848_, _14849_, _14850_, _14851_, _14852_, _14853_, _14854_, _14855_, _14856_, _14857_, _14858_, _14859_, _14860_, _14861_, _14862_, _14863_, _14864_, _14865_, _14866_, _14867_, _14868_, _14869_, _14870_, _14871_, _14872_, _14873_, _14874_, _14875_, _14876_, _14877_, _14878_, _14879_, _14880_, _14881_, _14882_, _14883_, _14884_, _14885_, _14886_, _14887_, _14888_, _14889_, _14890_, _14891_, _14892_, _14893_, _14894_, _14895_, _14896_, _14897_, _14898_, _14899_, _14900_, _14901_, _14902_, _14903_, _14904_, _14905_, _14906_, _14907_, _14908_, _14909_, _14910_, _14911_, _14912_, _14913_, _14914_, _14915_, _14916_, _14917_, _14918_, _14919_, _14920_, _14921_, _14922_, _14923_, _14924_, _14925_, _14926_, _14927_, _14928_, _14929_, _14930_, _14931_, _14932_, _14933_, _14934_, _14935_, _14936_, _14937_, _14938_, _14939_, _14940_, _14941_, _14942_, _14943_, _14944_, _14945_, _14946_, _14947_, _14948_, _14949_, _14950_, _14951_, _14952_, _14953_, _14954_, _14955_, _14956_, _14957_, _14958_, _14959_, _14960_, _14961_, _14962_, _14963_, _14964_, _14965_, _14966_, _14967_, _14968_, _14969_, _14970_, _14971_, _14972_, _14973_, _14974_, _14975_, _14976_, _14977_, _14978_, _14979_, _14980_, _14981_, _14982_, _14983_, _14984_, _14985_, _14986_, _14987_, _14988_, _14989_, _14990_, _14991_, _14992_, _14993_, _14994_, _14995_, _14996_, _14997_, _14998_, _14999_, _15000_, _15001_, _15002_, _15003_, _15004_, _15005_, _15006_, _15007_, _15008_, _15009_, _15010_, _15011_, _15012_, _15013_, _15014_, _15015_, _15016_, _15017_, _15018_, _15019_, _15020_, _15021_, _15022_, _15023_, _15024_, _15025_, _15026_, _15027_, _15028_, _15029_, _15030_, _15031_, _15032_, _15033_, _15034_, _15035_, _15036_, _15037_, _15038_, _15039_, _15040_, _15041_, _15042_, _15043_, _15044_, _15045_, _15046_, _15047_, _15048_, _15049_, _15050_, _15051_, _15052_, _15053_, _15054_, _15055_, _15056_, _15057_, _15058_, _15059_, _15060_, _15061_, _15062_, _15063_, _15064_, _15065_, _15066_, _15067_, _15068_, _15069_, _15070_, _15071_, _15072_, _15073_, _15074_, _15075_, _15076_, _15077_, _15078_, _15079_, _15080_, _15081_, _15082_, _15083_, _15084_, _15085_, _15086_, _15087_, _15088_, _15089_, _15090_, _15091_, _15092_, _15093_, _15094_, _15095_, _15096_, _15097_, _15098_, _15099_, _15100_, _15101_, _15102_, _15103_, _15104_, _15105_, _15106_, _15107_, _15108_, _15109_, _15110_, _15111_, _15112_, _15113_, _15114_, _15115_, _15116_, _15117_, _15118_, _15119_, _15120_, _15121_, _15122_, _15123_, _15124_, _15125_, _15126_, _15127_, _15128_, _15129_, _15130_, _15131_, _15132_, _15133_, _15134_, _15135_, _15136_, _15137_, _15138_, _15139_, _15140_, _15141_, _15142_, _15143_, _15144_, _15145_, _15146_, _15147_, _15148_, _15149_, _15150_, _15151_, _15152_, _15153_, _15154_, _15155_, _15156_, _15157_, _15158_, _15159_, _15160_, _15161_, _15162_, _15163_, _15164_, _15165_, _15166_, _15167_, _15168_, _15169_, _15170_, _15171_, _15172_, _15173_, _15174_, _15175_, _15176_, _15177_, _15178_, _15179_, _15180_, _15181_, _15182_, _15183_, _15184_, _15185_, _15186_, _15187_, _15188_, _15189_, _15190_, _15191_, _15192_, _15193_, _15194_, _15195_, _15196_, _15197_, _15198_, _15199_, _15200_, _15201_, _15202_, _15203_, _15204_, _15205_, _15206_, _15207_, _15208_, _15209_, _15210_, _15211_, _15212_, _15213_, _15214_, _15215_, _15216_, _15217_, _15218_, _15219_, _15220_, _15221_, _15222_, _15223_, _15224_, _15225_, _15226_, _15227_, _15228_, _15229_, _15230_, _15231_, _15232_, _15233_, _15234_, _15235_, _15236_, _15237_, _15238_, _15239_, _15240_, _15241_, _15242_, _15243_, _15244_, _15245_, _15246_, _15247_, _15248_, _15249_, _15250_, _15251_, _15252_, _15253_, _15254_, _15255_, _15256_, _15257_, _15258_, _15259_, _15260_, _15261_, _15262_, _15263_, _15264_, _15265_, _15266_, _15267_, _15268_, _15269_, _15270_, _15271_, _15272_, _15273_, _15274_, _15275_, _15276_, _15277_, _15278_, _15279_, _15280_, _15281_, _15282_, _15283_, _15284_, _15285_, _15286_, _15287_, _15288_, _15289_, _15290_, _15291_, _15292_, _15293_, _15294_, _15295_, _15296_, _15297_, _15298_, _15299_, _15300_, _15301_, _15302_, _15303_, _15304_, _15305_, _15306_, _15307_, _15308_, _15309_, _15310_, _15311_, _15312_, _15313_, _15314_, _15315_, _15316_, _15317_, _15318_, _15319_, _15320_, _15321_, _15322_, _15323_, _15324_, _15325_, _15326_, _15327_, _15328_, _15329_, _15330_, _15331_, _15332_, _15333_, _15334_, _15335_, _15336_, _15337_, _15338_, _15339_, _15340_, _15341_, _15342_, _15343_, _15344_, _15345_, _15346_, _15347_, _15348_, _15349_, _15350_, _15351_, _15352_, _15353_, _15354_, _15355_, _15356_, _15357_, _15358_, _15359_, _15360_, _15361_, _15362_, _15363_, _15364_, _15365_, _15366_, _15367_, _15368_, _15369_, _15370_, _15371_, _15372_, _15373_, _15374_, _15375_, _15376_, _15377_, _15378_, _15379_, _15380_, _15381_, _15382_, _15383_, _15384_, _15385_, _15386_, _15387_, _15388_, _15389_, _15390_, _15391_, _15392_, _15393_, _15394_, _15395_, _15396_, _15397_, _15398_, _15399_, _15400_, _15401_, _15402_, _15403_, _15404_, _15405_, _15406_, _15407_, _15408_, _15409_, _15410_, _15411_, _15412_, _15413_, _15414_, _15415_, _15416_, _15417_, _15418_, _15419_, _15420_, _15421_, _15422_, _15423_, _15424_, _15425_, _15426_, _15427_, _15428_, _15429_, _15430_, _15431_, _15432_, _15433_, _15434_, _15435_, _15436_, _15437_, _15438_, _15439_, _15440_, _15441_, _15442_, _15443_, _15444_, _15445_, _15446_, _15447_, _15448_, _15449_, _15450_, _15451_, _15452_, _15453_, _15454_, _15455_, _15456_, _15457_, _15458_, _15459_, _15460_, _15461_, _15462_, _15463_, _15464_, _15465_, _15466_, _15467_, _15468_, _15469_, _15470_, _15471_, _15472_, _15473_, _15474_, _15475_, _15476_, _15477_, _15478_, _15479_, _15480_, _15481_, _15482_, _15483_, _15484_, _15485_, _15486_, _15487_, _15488_, _15489_, _15490_, _15491_, _15492_, _15493_, _15494_, _15495_, _15496_, _15497_, _15498_, _15499_, _15500_, _15501_, _15502_, _15503_, _15504_, _15505_, _15506_, _15507_, _15508_, _15509_, _15510_, _15511_, _15512_, _15513_, _15514_, _15515_, _15516_, _15517_, _15518_, _15519_, _15520_, _15521_, _15522_, _15523_, _15524_, _15525_, _15526_, _15527_, _15528_, _15529_, _15530_, _15531_, _15532_, _15533_, _15534_, _15535_, _15536_, _15537_, _15538_, _15539_, _15540_, _15541_, _15542_, _15543_, _15544_, _15545_, _15546_, _15547_, _15548_, _15549_, _15550_, _15551_, _15552_, _15553_, _15554_, _15555_, _15556_, _15557_, _15558_, _15559_, _15560_, _15561_, _15562_, _15563_, _15564_, _15565_, _15566_, _15567_, _15568_, _15569_, _15570_, _15571_, _15572_, _15573_, _15574_, _15575_, _15576_, _15577_, _15578_, _15579_, _15580_, _15581_, _15582_, _15583_, _15584_, _15585_, _15586_, _15587_, _15588_, _15589_, _15590_, _15591_, _15592_, _15593_, _15594_, _15595_, _15596_, _15597_, _15598_, _15599_, _15600_, _15601_, _15602_, _15603_, _15604_, _15605_, _15606_, _15607_, _15608_, _15609_, _15610_, _15611_, _15612_, _15613_, _15614_, _15615_, _15616_, _15617_, _15618_, _15619_, _15620_, _15621_, _15622_, _15623_, _15624_, _15625_, _15626_, _15627_, _15628_, _15629_, _15630_, _15631_, _15632_, _15633_, _15634_, _15635_, _15636_, _15637_, _15638_, _15639_, _15640_, _15641_, _15642_, _15643_, _15644_, _15645_, _15646_, _15647_, _15648_, _15649_, _15650_, _15651_, _15652_, _15653_, _15654_, _15655_, _15656_, _15657_, _15658_, _15659_, _15660_, _15661_, _15662_, _15663_, _15664_, _15665_, _15666_, _15667_, _15668_, _15669_, _15670_, _15671_, _15672_, _15673_, _15674_, _15675_, _15676_, _15677_, _15678_, _15679_, _15680_, _15681_, _15682_, _15683_, _15684_, _15685_, _15686_, _15687_, _15688_, _15689_, _15690_, _15691_, _15692_, _15693_, _15694_, _15695_, _15696_, _15697_, _15698_, _15699_, _15700_, _15701_, _15702_, _15703_, _15704_, _15705_, _15706_, _15707_, _15708_, _15709_, _15710_, _15711_, _15712_, _15713_, _15714_, _15715_, _15716_, _15717_, _15718_, _15719_, _15720_, _15721_, _15722_, _15723_, _15724_, _15725_, _15726_, _15727_, _15728_, _15729_, _15730_, _15731_, _15732_, _15733_, _15734_, _15735_, _15736_, _15737_, _15738_, _15739_, _15740_, _15741_, _15742_, _15743_, _15744_, _15745_, _15746_, _15747_, _15748_, _15749_, _15750_, _15751_, _15752_, _15753_, _15754_, _15755_, _15756_, _15757_, _15758_, _15759_, _15760_, _15761_, _15762_, _15763_, _15764_, _15765_, _15766_, _15767_, _15768_, _15769_, _15770_, _15771_, _15772_, _15773_, _15774_, _15775_, _15776_, _15777_, _15778_, _15779_, _15780_, _15781_, _15782_, _15783_, _15784_, _15785_, _15786_, _15787_, _15788_, _15789_, _15790_, _15791_, _15792_, _15793_, _15794_, _15795_, _15796_, _15797_, _15798_, _15799_, _15800_, _15801_, _15802_, _15803_, _15804_, _15805_, _15806_, _15807_, _15808_, _15809_, _15810_, _15811_, _15812_, _15813_, _15814_, _15815_, _15816_, _15817_, _15818_, _15819_, _15820_, _15821_, _15822_, _15823_, _15824_, _15825_, _15826_, _15827_, _15828_, _15829_, _15830_, _15831_, _15832_, _15833_, _15834_, _15835_, _15836_, _15837_, _15838_, _15839_, _15840_, _15841_, _15842_, _15843_, _15844_, _15845_, _15846_, _15847_, _15848_, _15849_, _15850_, _15851_, _15852_, _15853_, _15854_, _15855_, _15856_, _15857_, _15858_, _15859_, _15860_, _15861_, _15862_, _15863_, _15864_, _15865_, _15866_, _15867_, _15868_, _15869_, _15870_, _15871_, _15872_, _15873_, _15874_, _15875_, _15876_, _15877_, _15878_, _15879_, _15880_, _15881_, _15882_, _15883_, _15884_, _15885_, _15886_, _15887_, _15888_, _15889_, _15890_, _15891_, _15892_, _15893_, _15894_, _15895_, _15896_, _15897_, _15898_, _15899_, _15900_, _15901_, _15902_, _15903_, _15904_, _15905_, _15906_, _15907_, _15908_, _15909_, _15910_, _15911_, _15912_, _15913_, _15914_, _15915_, _15916_, _15917_, _15918_, _15919_, _15920_, _15921_, _15922_, _15923_, _15924_, _15925_, _15926_, _15927_, _15928_, _15929_, _15930_, _15931_, _15932_, _15933_, _15934_, _15935_, _15936_, _15937_, _15938_, _15939_, _15940_, _15941_, _15942_, _15943_, _15944_, _15945_, _15946_, _15947_, _15948_, _15949_, _15950_, _15951_, _15952_, _15953_, _15954_, _15955_, _15956_, _15957_, _15958_, _15959_, _15960_, _15961_, _15962_, _15963_, _15964_, _15965_, _15966_, _15967_, _15968_, _15969_, _15970_, _15971_, _15972_, _15973_, _15974_, _15975_, _15976_, _15977_, _15978_, _15979_, _15980_, _15981_, _15982_, _15983_, _15984_, _15985_, _15986_, _15987_, _15988_, _15989_, _15990_, _15991_, _15992_, _15993_, _15994_, _15995_, _15996_, _15997_, _15998_, _15999_, _16000_, _16001_, _16002_, _16003_, _16004_, _16005_, _16006_, _16007_, _16008_, _16009_, _16010_, _16011_, _16012_, _16013_, _16014_, _16015_, _16016_, _16017_, _16018_, _16019_, _16020_, _16021_, _16022_, _16023_, _16024_, _16025_, _16026_, _16027_, _16028_, _16029_, _16030_, _16031_, _16032_, _16033_, _16034_, _16035_, _16036_, _16037_, _16038_, _16039_, _16040_, _16041_, _16042_, _16043_, _16044_, _16045_, _16046_, _16047_, _16048_, _16049_, _16050_, _16051_, _16052_, _16053_, _16054_, _16055_, _16056_, _16057_, _16058_, _16059_, _16060_, _16061_, _16062_, _16063_, _16064_, _16065_, _16066_, _16067_, _16068_, _16069_, _16070_, _16071_, _16072_, _16073_, _16074_, _16075_, _16076_, _16077_, _16078_, _16079_, _16080_, _16081_, _16082_, _16083_, _16084_, _16085_, _16086_, _16087_, _16088_, _16089_, _16090_, _16091_, _16092_, _16093_, _16094_, _16095_, _16096_, _16097_, _16098_, _16099_, _16100_, _16101_, _16102_, _16103_, _16104_, _16105_, _16106_, _16107_, _16108_, _16109_, _16110_, _16111_, _16112_, _16113_, _16114_, _16115_, _16116_, _16117_, _16118_, _16119_, _16120_, _16121_, _16122_, _16123_, _16124_, _16125_, _16126_, _16127_, _16128_, _16129_, _16130_, _16131_, _16132_, _16133_, _16134_, _16135_, _16136_, _16137_, _16138_, _16139_, _16140_, _16141_, _16142_, _16143_, _16144_, _16145_, _16146_, _16147_, _16148_, _16149_, _16150_, _16151_, _16152_, _16153_, _16154_, _16155_, _16156_, _16157_, _16158_, _16159_, _16160_, _16161_, _16162_, _16163_, _16164_, _16165_, _16166_, _16167_, _16168_, _16169_, _16170_, _16171_, _16172_, _16173_, _16174_, _16175_, _16176_, _16177_, _16178_, _16179_, _16180_, _16181_, _16182_, _16183_, _16184_, _16185_, _16186_, _16187_, _16188_, _16189_, _16190_, _16191_, _16192_, _16193_, _16194_, _16195_, _16196_, _16197_, _16198_, _16199_, _16200_, _16201_, _16202_, _16203_, _16204_, _16205_, _16206_, _16207_, _16208_, _16209_, _16210_, _16211_, _16212_, _16213_, _16214_, _16215_, _16216_, _16217_, _16218_, _16219_, _16220_, _16221_, _16222_, _16223_, _16224_, _16225_, _16226_, _16227_, _16228_, _16229_, _16230_, _16231_, _16232_, _16233_, _16234_, _16235_, _16236_, _16237_, _16238_, _16239_, _16240_, _16241_, _16242_, _16243_, _16244_, _16245_, _16246_, _16247_, _16248_, _16249_, _16250_, _16251_, _16252_, _16253_, _16254_, _16255_, _16256_, _16257_, _16258_, _16259_, _16260_, _16261_, _16262_, _16263_, _16264_, _16265_, _16266_, _16267_, _16268_, _16269_, _16270_, _16271_, _16272_, _16273_, _16274_, _16275_, _16276_, _16277_, _16278_, _16279_, _16280_, _16281_, _16282_, _16283_, _16284_, _16285_, _16286_, _16287_, _16288_, _16289_, _16290_, _16291_, _16292_, _16293_, _16294_, _16295_, _16296_, _16297_, _16298_, _16299_, _16300_, _16301_, _16302_, _16303_, _16304_, _16305_, _16306_, _16307_, _16308_, _16309_, _16310_, _16311_, _16312_, _16313_, _16314_, _16315_, _16316_, _16317_, _16318_, _16319_, _16320_, _16321_, _16322_, _16323_, _16324_, _16325_, _16326_, _16327_, _16328_, _16329_, _16330_, _16331_, _16332_, _16333_, _16334_, _16335_, _16336_, _16337_, _16338_, _16339_, _16340_, _16341_, _16342_, _16343_, _16344_, _16345_, _16346_, _16347_, _16348_, _16349_, _16350_, _16351_, _16352_, _16353_, _16354_, _16355_, _16356_, _16357_, _16358_, _16359_, _16360_, _16361_, _16362_, _16363_, _16364_, _16365_, _16366_, _16367_, _16368_, _16369_, _16370_, _16371_, _16372_, _16373_, _16374_, _16375_, _16376_, _16377_, _16378_, _16379_, _16380_, _16381_, _16382_, _16383_, _16384_, _16385_, _16386_, _16387_, _16388_, _16389_, _16390_, _16391_, _16392_, _16393_, _16394_, _16395_, _16396_, _16397_, _16398_, _16399_, _16400_, _16401_, _16402_, _16403_, _16404_, _16405_, _16406_, _16407_, _16408_, _16409_, _16410_, _16411_, _16412_, _16413_, _16414_, _16415_, _16416_, _16417_, _16418_, _16419_, _16420_, _16421_, _16422_, _16423_, _16424_, _16425_, _16426_, _16427_, _16428_, _16429_, _16430_, _16431_, _16432_, _16433_, _16434_, _16435_, _16436_, _16437_, _16438_, _16439_, _16440_, _16441_, _16442_, _16443_, _16444_, _16445_, _16446_, _16447_, _16448_, _16449_, _16450_, _16451_, _16452_, _16453_, _16454_, _16455_, _16456_, _16457_, _16458_, _16459_, _16460_, _16461_, _16462_, _16463_, _16464_, _16465_, _16466_, _16467_, _16468_, _16469_, _16470_, _16471_, _16472_, _16473_, _16474_, _16475_, _16476_, _16477_, _16478_, _16479_, _16480_, _16481_, _16482_, _16483_, _16484_, _16485_, _16486_, _16487_, _16488_, _16489_, _16490_, _16491_, _16492_, _16493_, _16494_, _16495_, _16496_, _16497_, _16498_, _16499_, _16500_, _16501_, _16502_, _16503_, _16504_, _16505_, _16506_, _16507_, _16508_, _16509_, _16510_, _16511_, _16512_, _16513_, _16514_, _16515_, _16516_, _16517_, _16518_, _16519_, _16520_, _16521_, _16522_, _16523_, _16524_, _16525_, _16526_, _16527_, _16528_, _16529_, _16530_, _16531_, _16532_, _16533_, _16534_, _16535_, _16536_, _16537_, _16538_, _16539_, _16540_, _16541_, _16542_, _16543_, _16544_, _16545_, _16546_, _16547_, _16548_, _16549_, _16550_, _16551_, _16552_, _16553_, _16554_, _16555_, _16556_, _16557_, _16558_, _16559_, _16560_, _16561_, _16562_, _16563_, _16564_, _16565_, _16566_, _16567_, _16568_, _16569_, _16570_, _16571_, _16572_, _16573_, _16574_, _16575_, _16576_, _16577_, _16578_, _16579_, _16580_, _16581_, _16582_, _16583_, _16584_, _16585_, _16586_, _16587_, _16588_, _16589_, _16590_, _16591_, _16592_, _16593_, _16594_, _16595_, _16596_, _16597_, _16598_, _16599_, _16600_, _16601_, _16602_, _16603_, _16604_, _16605_, _16606_, _16607_, _16608_, _16609_, _16610_, _16611_, _16612_, _16613_, _16614_, _16615_, _16616_, _16617_, _16618_, _16619_, _16620_, _16621_, _16622_, _16623_, _16624_, _16625_, _16626_, _16627_, _16628_, _16629_, _16630_, _16631_, _16632_, _16633_, _16634_, _16635_, _16636_, _16637_, _16638_, _16639_, _16640_, _16641_, _16642_, _16643_, _16644_, _16645_, _16646_, _16647_, _16648_, _16649_, _16650_, _16651_, _16652_, _16653_, _16654_, _16655_, _16656_, _16657_, _16658_, _16659_, _16660_, _16661_, _16662_, _16663_, _16664_, _16665_, _16666_, _16667_, _16668_, _16669_, _16670_, _16671_, _16672_, _16673_, _16674_, _16675_, _16676_, _16677_, _16678_, _16679_, _16680_, _16681_, _16682_, _16683_, _16684_, _16685_, _16686_, _16687_, _16688_, _16689_, _16690_, _16691_, _16692_, _16693_, _16694_, _16695_, _16696_, _16697_, _16698_, _16699_, _16700_, _16701_, _16702_, _16703_, _16704_, _16705_, _16706_, _16707_, _16708_, _16709_, _16710_, _16711_, _16712_, _16713_, _16714_, _16715_, _16716_, _16717_, _16718_, _16719_, _16720_, _16721_, _16722_, _16723_, _16724_, _16725_, _16726_, _16727_, _16728_, _16729_, _16730_, _16731_, _16732_, _16733_, _16734_, _16735_, _16736_, _16737_, _16738_, _16739_, _16740_, _16741_, _16742_, _16743_, _16744_, _16745_, _16746_, _16747_, _16748_, _16749_, _16750_, _16751_, _16752_, _16753_, _16754_, _16755_, _16756_, _16757_, _16758_, _16759_, _16760_, _16761_, _16762_, _16763_, _16764_, _16765_, _16766_, _16767_, _16768_, _16769_, _16770_, _16771_, _16772_, _16773_, _16774_, _16775_, _16776_, _16777_, _16778_, _16779_, _16780_, _16781_, _16782_, _16783_, _16784_, _16785_, _16786_, _16787_, _16788_, _16789_, _16790_, _16791_, _16792_, _16793_, _16794_, _16795_, _16796_, _16797_, _16798_, _16799_, _16800_, _16801_, _16802_, _16803_, _16804_, _16805_, _16806_, _16807_, _16808_, _16809_, _16810_, _16811_, _16812_, _16813_, _16814_, _16815_, _16816_, _16817_, _16818_, _16819_, _16820_, _16821_, _16822_, _16823_, _16824_, _16825_, _16826_, _16827_, _16828_, _16829_, _16830_, _16831_, _16832_, _16833_, _16834_, _16835_, _16836_, _16837_, _16838_, _16839_, _16840_, _16841_, _16842_, _16843_, _16844_, _16845_, _16846_, _16847_, _16848_, _16849_, _16850_, _16851_, _16852_, _16853_, _16854_, _16855_, _16856_, _16857_, _16858_, _16859_, _16860_, _16861_, _16862_, _16863_, _16864_, _16865_, _16866_, _16867_, _16868_, _16869_, _16870_, _16871_, _16872_, _16873_, _16874_, _16875_, _16876_, _16877_, _16878_, _16879_, _16880_, _16881_, _16882_, _16883_, _16884_, _16885_, _16886_, _16887_, _16888_, _16889_, _16890_, _16891_, _16892_, _16893_, _16894_, _16895_, _16896_, _16897_, _16898_, _16899_, _16900_, _16901_, _16902_, _16903_, _16904_, _16905_, _16906_, _16907_, _16908_, _16909_, _16910_, _16911_, _16912_, _16913_, _16914_, _16915_, _16916_, _16917_, _16918_, _16919_, _16920_, _16921_, _16922_, _16923_, _16924_, _16925_, _16926_, _16927_, _16928_, _16929_, _16930_, _16931_, _16932_, _16933_, _16934_, _16935_, _16936_, _16937_, _16938_, _16939_, _16940_, _16941_, _16942_, _16943_, _16944_, _16945_, _16946_, _16947_, _16948_, _16949_, _16950_, _16951_, _16952_, _16953_, _16954_, _16955_, _16956_, _16957_, _16958_, _16959_, _16960_, _16961_, _16962_, _16963_, _16964_, _16965_, _16966_, _16967_, _16968_, _16969_, _16970_, _16971_, _16972_, _16973_, _16974_, _16975_, _16976_, _16977_, _16978_, _16979_, _16980_, _16981_, _16982_, _16983_, _16984_, _16985_, _16986_, _16987_, _16988_, _16989_, _16990_, _16991_, _16992_, _16993_, _16994_, _16995_, _16996_, _16997_, _16998_, _16999_, _17000_, _17001_, _17002_, _17003_, _17004_, _17005_, _17006_, _17007_, _17008_, _17009_, _17010_, _17011_, _17012_, _17013_, _17014_, _17015_, _17016_, _17017_, _17018_, _17019_, _17020_, _17021_, _17022_, _17023_, _17024_, _17025_, _17026_, _17027_, _17028_, _17029_, _17030_, _17031_, _17032_, _17033_, _17034_, _17035_, _17036_, _17037_, _17038_, _17039_, _17040_, _17041_, _17042_, _17043_, _17044_, _17045_, _17046_, _17047_, _17048_, _17049_, _17050_, _17051_, _17052_, _17053_, _17054_, _17055_, _17056_, _17057_, _17058_, _17059_, _17060_, _17061_, _17062_, _17063_, _17064_, _17065_, _17066_, _17067_, _17068_, _17069_, _17070_, _17071_, _17072_, _17073_, _17074_, _17075_, _17076_, _17077_, _17078_, _17079_, _17080_, _17081_, _17082_, _17083_, _17084_, _17085_, _17086_, _17087_, _17088_, _17089_, _17090_, _17091_, _17092_, _17093_, _17094_, _17095_, _17096_, _17097_, _17098_, _17099_, _17100_, _17101_, _17102_, _17103_, _17104_, _17105_, _17106_, _17107_, _17108_, _17109_, _17110_, _17111_, _17112_, _17113_, _17114_, _17115_, _17116_, _17117_, _17118_, _17119_, _17120_, _17121_, _17122_, _17123_, _17124_, _17125_, _17126_, _17127_, _17128_, _17129_, _17130_, _17131_, _17132_, _17133_, _17134_, _17135_, _17136_, _17137_, _17138_, _17139_, _17140_, _17141_, _17142_, _17143_, _17144_, _17145_, _17146_, _17147_, _17148_, _17149_, _17150_, _17151_, _17152_, _17153_, _17154_, _17155_, _17156_, _17157_, _17158_, _17159_, _17160_, _17161_, _17162_, _17163_, _17164_, _17165_, _17166_, _17167_, _17168_, _17169_, _17170_, _17171_, _17172_, _17173_, _17174_, _17175_, _17176_, _17177_, _17178_, _17179_, _17180_, _17181_, _17182_, _17183_, _17184_, _17185_, _17186_, _17187_, _17188_, _17189_, _17190_, _17191_, _17192_, _17193_, _17194_, _17195_, _17196_, _17197_, _17198_, _17199_, _17200_, _17201_, _17202_, _17203_, _17204_, _17205_, _17206_, _17207_, _17208_, _17209_, _17210_, _17211_, _17212_, _17213_, _17214_, _17215_, _17216_, _17217_, _17218_, _17219_, _17220_, _17221_, _17222_, _17223_, _17224_, _17225_, _17226_, _17227_, _17228_, _17229_, _17230_, _17231_, _17232_, _17233_, _17234_, _17235_, _17236_, _17237_, _17238_, _17239_, _17240_, _17241_, _17242_, _17243_, _17244_, _17245_, _17246_, _17247_, _17248_, _17249_, _17250_, _17251_, _17252_, _17253_, _17254_, _17255_, _17256_, _17257_, _17258_, _17259_, _17260_, _17261_, _17262_, _17263_, _17264_, _17265_, _17266_, _17267_, _17268_, _17269_, _17270_, _17271_, _17272_, _17273_, _17274_, _17275_, _17276_, _17277_, _17278_, _17279_, _17280_, _17281_, _17282_, _17283_, _17284_, _17285_, _17286_, _17287_, _17288_, _17289_, _17290_, _17291_, _17292_, _17293_, _17294_, _17295_, _17296_, _17297_, _17298_, _17299_, _17300_, _17301_, _17302_, _17303_, _17304_, _17305_, _17306_, _17307_, _17308_, _17309_, _17310_, _17311_, _17312_, _17313_, _17314_, _17315_, _17316_, _17317_, _17318_, _17319_, _17320_, _17321_, _17322_, _17323_, _17324_, _17325_, _17326_, _17327_, _17328_, _17329_, _17330_, _17331_, _17332_, _17333_, _17334_, _17335_, _17336_, _17337_, _17338_, _17339_, _17340_, _17341_, _17342_, _17343_, _17344_, _17345_, _17346_, _17347_, _17348_, _17349_, _17350_, _17351_, _17352_, _17353_, _17354_, _17355_, _17356_, _17357_, _17358_, _17359_, _17360_, _17361_, _17362_, _17363_, _17364_, _17365_, _17366_, _17367_, _17368_, _17369_, _17370_, _17371_, _17372_, _17373_, _17374_, _17375_, _17376_, _17377_, _17378_, _17379_, _17380_, _17381_, _17382_, _17383_, _17384_, _17385_, _17386_, _17387_, _17388_, _17389_, _17390_, _17391_, _17392_, _17393_, _17394_, _17395_, _17396_, _17397_, _17398_, _17399_, _17400_, _17401_, _17402_, _17403_, _17404_, _17405_, _17406_, _17407_, _17408_, _17409_, _17410_, _17411_, _17412_, _17413_, _17414_, _17415_, _17416_, _17417_, _17418_, _17419_, _17420_, _17421_, _17422_, _17423_, _17424_, _17425_, _17426_, _17427_, _17428_, _17429_, _17430_, _17431_, _17432_, _17433_, _17434_, _17435_, _17436_, _17437_, _17438_, _17439_, _17440_, _17441_, _17442_, _17443_, _17444_, _17445_, _17446_, _17447_, _17448_, _17449_, _17450_, _17451_, _17452_, _17453_, _17454_, _17455_, _17456_, _17457_, _17458_, _17459_, _17460_, _17461_, _17462_, _17463_, _17464_, _17465_, _17466_, _17467_, _17468_, _17469_, _17470_, _17471_, _17472_, _17473_, _17474_, _17475_, _17476_, _17477_, _17478_, _17479_, _17480_, _17481_, _17482_, _17483_, _17484_, _17485_, _17486_, _17487_, _17488_, _17489_, _17490_, _17491_, _17492_, _17493_, _17494_, _17495_, _17496_, _17497_, _17498_, _17499_, _17500_, _17501_, _17502_, _17503_, _17504_, _17505_, _17506_, _17507_, _17508_, _17509_, _17510_, _17511_, _17512_, _17513_, _17514_, _17515_, _17516_, _17517_, _17518_, _17519_, _17520_, _17521_, _17522_, _17523_, _17524_, _17525_, _17526_, _17527_, _17528_, _17529_, _17530_, _17531_, _17532_, _17533_, _17534_, _17535_, _17536_, _17537_, _17538_, _17539_, _17540_, _17541_, _17542_, _17543_, _17544_, _17545_, _17546_, _17547_, _17548_, _17549_, _17550_, _17551_, _17552_, _17553_, _17554_, _17555_, _17556_, _17557_, _17558_, _17559_, _17560_, _17561_, _17562_, _17563_, _17564_, _17565_, _17566_, _17567_, _17568_, _17569_, _17570_, _17571_, _17572_, _17573_, _17574_, _17575_, _17576_, _17577_, _17578_, _17579_, _17580_, _17581_, _17582_, _17583_, _17584_, _17585_, _17586_, _17587_, _17588_, _17589_, _17590_, _17591_, _17592_, _17593_, _17594_, _17595_, _17596_, _17597_, _17598_, _17599_, _17600_, _17601_, _17602_, _17603_, _17604_, _17605_, _17606_, _17607_, _17608_, _17609_, _17610_, _17611_, _17612_, _17613_, _17614_, _17615_, _17616_, _17617_, _17618_, _17619_, _17620_, _17621_, _17622_, _17623_, _17624_, _17625_, _17626_, _17627_, _17628_, _17629_, _17630_, _17631_, _17632_, _17633_, _17634_, _17635_, _17636_, _17637_, _17638_, _17639_, _17640_, _17641_, _17642_, _17643_, _17644_, _17645_, _17646_, _17647_, _17648_, _17649_, _17650_, _17651_, _17652_, _17653_, _17654_, _17655_, _17656_, _17657_, _17658_, _17659_, _17660_, _17661_, _17662_, _17663_, _17664_, _17665_, _17666_, _17667_, _17668_, _17669_, _17670_, _17671_, _17672_, _17673_, _17674_, _17675_, _17676_, _17677_, _17678_, _17679_, _17680_, _17681_, _17682_, _17683_, _17684_, _17685_, _17686_, _17687_, _17688_, _17689_, _17690_, _17691_, _17692_, _17693_, _17694_, _17695_, _17696_, _17697_, _17698_, _17699_, _17700_, _17701_, _17702_, _17703_, _17704_, _17705_, _17706_, _17707_, _17708_, _17709_, _17710_, _17711_, _17712_, _17713_, _17714_, _17715_, _17716_, _17717_, _17718_, _17719_, _17720_, _17721_, _17722_, _17723_, _17724_, _17725_, _17726_, _17727_, _17728_, _17729_, _17730_, _17731_, _17732_, _17733_, _17734_, _17735_, _17736_, _17737_, _17738_, _17739_, _17740_, _17741_, _17742_, _17743_, _17744_, _17745_, _17746_, _17747_, _17748_, _17749_, _17750_, _17751_, _17752_, _17753_, _17754_, _17755_, _17756_, _17757_, _17758_, _17759_, _17760_, _17761_, _17762_, _17763_, _17764_, _17765_, _17766_, _17767_, _17768_, _17769_, _17770_, _17771_, _17772_, _17773_, _17774_, _17775_, _17776_, _17777_, _17778_, _17779_, _17780_, _17781_, _17782_, _17783_, _17784_, _17785_, _17786_, _17787_, _17788_, _17789_, _17790_, _17791_, _17792_, _17793_, _17794_, _17795_, _17796_, _17797_, _17798_, _17799_, _17800_, _17801_, _17802_, _17803_, _17804_, _17805_, _17806_, _17807_, _17808_, _17809_, _17810_, _17811_, _17812_, _17813_, _17814_, _17815_, _17816_, _17817_, _17818_, _17819_, _17820_, _17821_, _17822_, _17823_, _17824_, _17825_, _17826_, _17827_, _17828_, _17829_, _17830_, _17831_, _17832_, _17833_, _17834_, _17835_, _17836_, _17837_, _17838_, _17839_, _17840_, _17841_, _17842_, _17843_, _17844_, _17845_, _17846_, _17847_, _17848_, _17849_, _17850_, _17851_, _17852_, _17853_, _17854_, _17855_, _17856_, _17857_, _17858_, _17859_, _17860_, _17861_, _17862_, _17863_, _17864_, _17865_, _17866_, _17867_, _17868_, _17869_, _17870_, _17871_, _17872_, _17873_, _17874_, _17875_, _17876_, _17877_, _17878_, _17879_, _17880_, _17881_, _17882_, _17883_, _17884_, _17885_, _17886_, _17887_, _17888_, _17889_, _17890_, _17891_, _17892_, _17893_, _17894_, _17895_, _17896_, _17897_, _17898_, _17899_, _17900_, _17901_, _17902_, _17903_, _17904_, _17905_, _17906_, _17907_, _17908_, _17909_, _17910_, _17911_, _17912_, _17913_, _17914_, _17915_, _17916_, _17917_, _17918_, _17919_, _17920_, _17921_, _17922_, _17923_, _17924_, _17925_, _17926_, _17927_, _17928_, _17929_, _17930_, _17931_, _17932_, _17933_, _17934_, _17935_, _17936_, _17937_, _17938_, _17939_, _17940_, _17941_, _17942_, _17943_, _17944_, _17945_, _17946_, _17947_, _17948_, _17949_, _17950_, _17951_, _17952_, _17953_, _17954_, _17955_, _17956_, _17957_, _17958_, _17959_, _17960_, _17961_, _17962_, _17963_, _17964_, _17965_, _17966_, _17967_, _17968_, _17969_, _17970_, _17971_, _17972_, _17973_, _17974_, _17975_, _17976_, _17977_, _17978_, _17979_, _17980_, _17981_, _17982_, _17983_, _17984_, _17985_, _17986_, _17987_, _17988_, _17989_, _17990_, _17991_, _17992_, _17993_, _17994_, _17995_, _17996_, _17997_, _17998_, _17999_, _18000_, _18001_, _18002_, _18003_, _18004_, _18005_, _18006_, _18007_, _18008_, _18009_, _18010_, _18011_, _18012_, _18013_, _18014_, _18015_, _18016_, _18017_, _18018_, _18019_, _18020_, _18021_, _18022_, _18023_, _18024_, _18025_, _18026_, _18027_, _18028_, _18029_, _18030_, _18031_, _18032_, _18033_, _18034_, _18035_, _18036_, _18037_, _18038_, _18039_, _18040_, _18041_, _18042_, _18043_, _18044_, _18045_, _18046_, _18047_, _18048_, _18049_, _18050_, _18051_, _18052_, _18053_, _18054_, _18055_, _18056_, _18057_, _18058_, _18059_, _18060_, _18061_, _18062_, _18063_, _18064_, _18065_, _18066_, _18067_, _18068_, _18069_, _18070_, _18071_, _18072_, _18073_, _18074_, _18075_, _18076_, _18077_, _18078_, _18079_, _18080_, _18081_, _18082_, _18083_, _18084_, _18085_, _18086_, _18087_, _18088_, _18089_, _18090_, _18091_, _18092_, _18093_, _18094_, _18095_, _18096_, _18097_, _18098_, _18099_, _18100_, _18101_, _18102_, _18103_, _18104_, _18105_, _18106_, _18107_, _18108_, _18109_, _18110_, _18111_, _18112_, _18113_, _18114_, _18115_, _18116_, _18117_, _18118_, _18119_, _18120_, _18121_, _18122_, _18123_, _18124_, _18125_, _18126_, _18127_, _18128_, _18129_, _18130_, _18131_, _18132_, _18133_, _18134_, _18135_, _18136_, _18137_, _18138_, _18139_, _18140_, _18141_, _18142_, _18143_, _18144_, _18145_, _18146_, _18147_, _18148_, _18149_, _18150_, _18151_, _18152_, _18153_, _18154_, _18155_, _18156_, _18157_, _18158_, _18159_, _18160_, _18161_, _18162_, _18163_, _18164_, _18165_, _18166_, _18167_, _18168_, _18169_, _18170_, _18171_, _18172_, _18173_, _18174_, _18175_, _18176_, _18177_, _18178_, _18179_, _18180_, _18181_, _18182_, _18183_, _18184_, _18185_, _18186_, _18187_, _18188_, _18189_, _18190_, _18191_, _18192_, _18193_, _18194_, _18195_, _18196_, _18197_, _18198_, _18199_, _18200_, _18201_, _18202_, _18203_, _18204_, _18205_, _18206_, _18207_, _18208_, _18209_, _18210_, _18211_, _18212_, _18213_, _18214_, _18215_, _18216_, _18217_, _18218_, _18219_, _18220_, _18221_, _18222_, _18223_, _18224_, _18225_, _18226_, _18227_, _18228_, _18229_, _18230_, _18231_, _18232_, _18233_, _18234_, _18235_, _18236_, _18237_, _18238_, _18239_, _18240_, _18241_, _18242_, _18243_, _18244_, _18245_, _18246_, _18247_, _18248_, _18249_, _18250_, _18251_, _18252_, _18253_, _18254_, _18255_, _18256_, _18257_, _18258_, _18259_, _18260_, _18261_, _18262_, _18263_, _18264_, _18265_, _18266_, _18267_, _18268_, _18269_, _18270_, _18271_, _18272_, _18273_, _18274_, _18275_, _18276_, _18277_, _18278_, _18279_, _18280_, _18281_, _18282_, _18283_, _18284_, _18285_, _18286_, _18287_, _18288_, _18289_, _18290_, _18291_, _18292_, _18293_, _18294_, _18295_, _18296_, _18297_, _18298_, _18299_, _18300_, _18301_, _18302_, _18303_, _18304_, _18305_, _18306_, _18307_, _18308_, _18309_, _18310_, _18311_, _18312_, _18313_, _18314_, _18315_, _18316_, _18317_, _18318_, _18319_, _18320_, _18321_, _18322_, _18323_, _18324_, _18325_, _18326_, _18327_, _18328_, _18329_, _18330_, _18331_, _18332_, _18333_, _18334_, _18335_, _18336_, _18337_, _18338_, _18339_, _18340_, _18341_, _18342_, _18343_, _18344_, _18345_, _18346_, _18347_, _18348_, _18349_, _18350_, _18351_, _18352_, _18353_, _18354_, _18355_, _18356_, _18357_, _18358_, _18359_, _18360_, _18361_, _18362_, _18363_, _18364_, _18365_, _18366_, _18367_, _18368_, _18369_, _18370_, _18371_, _18372_, _18373_, _18374_, _18375_, _18376_, _18377_, _18378_, _18379_, _18380_, _18381_, _18382_, _18383_, _18384_, _18385_, _18386_, _18387_, _18388_, _18389_, _18390_, _18391_, _18392_, _18393_, _18394_, _18395_, _18396_, _18397_, _18398_, _18399_, _18400_, _18401_, _18402_, _18403_, _18404_, _18405_, _18406_, _18407_, _18408_, _18409_, _18410_, _18411_, _18412_, _18413_, _18414_, _18415_, _18416_, _18417_, _18418_, _18419_, _18420_, _18421_, _18422_, _18423_, _18424_, _18425_, _18426_, _18427_, _18428_, _18429_, _18430_, _18431_, _18432_, _18433_, _18434_, _18435_, _18436_, _18437_, _18438_, _18439_, _18440_, _18441_, _18442_, _18443_, _18444_, _18445_, _18446_, _18447_, _18448_, _18449_, _18450_, _18451_, _18452_, _18453_, _18454_, _18455_, _18456_, _18457_, _18458_, _18459_, _18460_, _18461_, _18462_, _18463_, _18464_, _18465_, _18466_, _18467_, _18468_, _18469_, _18470_, _18471_, _18472_, _18473_, _18474_, _18475_, _18476_, _18477_, _18478_, _18479_, _18480_, _18481_, _18482_, _18483_, _18484_, _18485_, _18486_, _18487_, _18488_, _18489_, _18490_, _18491_, _18492_, _18493_, _18494_, _18495_, _18496_, _18497_, _18498_, _18499_, _18500_, _18501_, _18502_, _18503_, _18504_, _18505_, _18506_, _18507_, _18508_, _18509_, _18510_, _18511_, _18512_, _18513_, _18514_, _18515_, _18516_, _18517_, _18518_, _18519_, _18520_, _18521_, _18522_, _18523_, _18524_, _18525_, _18526_, _18527_, _18528_, _18529_, _18530_, _18531_, _18532_, _18533_, _18534_, _18535_, _18536_, _18537_, _18538_, _18539_, _18540_, _18541_, _18542_, _18543_, _18544_, _18545_, _18546_, _18547_, _18548_, _18549_, _18550_, _18551_, _18552_, _18553_, _18554_, _18555_, _18556_, _18557_, _18558_, _18559_, _18560_, _18561_, _18562_, _18563_, _18564_, _18565_, _18566_, _18567_, _18568_, _18569_, _18570_, _18571_, _18572_, _18573_, _18574_, _18575_, _18576_, _18577_, _18578_, _18579_, _18580_, _18581_, _18582_, _18583_, _18584_, _18585_, _18586_, _18587_, _18588_, _18589_, _18590_, _18591_, _18592_, _18593_, _18594_, _18595_, _18596_, _18597_, _18598_, _18599_, _18600_, _18601_, _18602_, _18603_, _18604_, _18605_, _18606_, _18607_, _18608_, _18609_, _18610_, _18611_, _18612_, _18613_, _18614_, _18615_, _18616_, _18617_, _18618_, _18619_, _18620_, _18621_, _18622_, _18623_, _18624_, _18625_, _18626_, _18627_, _18628_, _18629_, _18630_, _18631_, _18632_, _18633_, _18634_, _18635_, _18636_, _18637_, _18638_, _18639_, _18640_, _18641_, _18642_, _18643_, _18644_, _18645_, _18646_, _18647_, _18648_, _18649_, _18650_, _18651_, _18652_, _18653_, _18654_, _18655_, _18656_, _18657_, _18658_, _18659_, _18660_, _18661_, _18662_, _18663_, _18664_, _18665_, _18666_, _18667_, _18668_, _18669_, _18670_, _18671_, _18672_, _18673_, _18674_, _18675_, _18676_, _18677_, _18678_, _18679_, _18680_, _18681_, _18682_, _18683_, _18684_, _18685_, _18686_, _18687_, _18688_, _18689_, _18690_, _18691_, _18692_, _18693_, _18694_, _18695_, _18696_, _18697_, _18698_, _18699_, _18700_, _18701_, _18702_, _18703_, _18704_, _18705_, _18706_, _18707_, _18708_, _18709_, _18710_, _18711_, _18712_, _18713_, _18714_, _18715_, _18716_, _18717_, _18718_, _18719_, _18720_, _18721_, _18722_, _18723_, _18724_, _18725_, _18726_, _18727_, _18728_, _18729_, _18730_, _18731_, _18732_, _18733_, _18734_, _18735_, _18736_, _18737_, _18738_, _18739_, _18740_, _18741_, _18742_, _18743_, _18744_, _18745_, _18746_, _18747_, _18748_, _18749_, _18750_, _18751_, _18752_, _18753_, _18754_, _18755_, _18756_, _18757_, _18758_, _18759_, _18760_, _18761_, _18762_, _18763_, _18764_, _18765_, _18766_, _18767_, _18768_, _18769_, _18770_, _18771_, _18772_, _18773_, _18774_, _18775_, _18776_, _18777_, _18778_, _18779_, _18780_, _18781_, _18782_, _18783_, _18784_, _18785_, _18786_, _18787_, _18788_, _18789_, _18790_, _18791_, _18792_, _18793_, _18794_, _18795_, _18796_, _18797_, _18798_, _18799_, _18800_, _18801_, _18802_, _18803_, _18804_, _18805_, _18806_, _18807_, _18808_, _18809_, _18810_, _18811_, _18812_, _18813_, _18814_, _18815_, _18816_, _18817_, _18818_, _18819_, _18820_, _18821_, _18822_, _18823_, _18824_, _18825_, _18826_, _18827_, _18828_, _18829_, _18830_, _18831_, _18832_, _18833_, _18834_, _18835_, _18836_, _18837_, _18838_, _18839_, _18840_, _18841_, _18842_, _18843_, _18844_, _18845_, _18846_, _18847_, _18848_, _18849_, _18850_, _18851_, _18852_, _18853_, _18854_, _18855_, _18856_, _18857_, _18858_, _18859_, _18860_, _18861_, _18862_, _18863_, _18864_, _18865_, _18866_, _18867_, _18868_, _18869_, _18870_, _18871_, _18872_, _18873_, _18874_, _18875_, _18876_, _18877_, _18878_, _18879_, _18880_, _18881_, _18882_, _18883_, _18884_, _18885_, _18886_, _18887_, _18888_, _18889_, _18890_, _18891_, _18892_, _18893_, _18894_, _18895_, _18896_, _18897_, _18898_, _18899_, _18900_, _18901_, _18902_, _18903_, _18904_, _18905_, _18906_, _18907_, _18908_, _18909_, _18910_, _18911_, _18912_, _18913_, _18914_, _18915_, _18916_, _18917_, _18918_, _18919_, _18920_, _18921_, _18922_, _18923_, _18924_, _18925_, _18926_, _18927_, _18928_, _18929_, _18930_, _18931_, _18932_, _18933_, _18934_, _18935_, _18936_, _18937_, _18938_, _18939_, _18940_, _18941_, _18942_, _18943_, _18944_, _18945_, _18946_, _18947_, _18948_, _18949_, _18950_, _18951_, _18952_, _18953_, _18954_, _18955_, _18956_, _18957_, _18958_, _18959_, _18960_, _18961_, _18962_, _18963_, _18964_, _18965_, _18966_, _18967_, _18968_, _18969_, _18970_, _18971_, _18972_, _18973_, _18974_, _18975_, _18976_, _18977_, _18978_, _18979_, _18980_, _18981_, _18982_, _18983_, _18984_, _18985_, _18986_, _18987_, _18988_, _18989_, _18990_, _18991_, _18992_, _18993_, _18994_, _18995_, _18996_, _18997_, _18998_, _18999_, _19000_, _19001_, _19002_, _19003_, _19004_, _19005_, _19006_, _19007_, _19008_, _19009_, _19010_, _19011_, _19012_, _19013_, _19014_, _19015_, _19016_, _19017_, _19018_, _19019_, _19020_, _19021_, _19022_, _19023_, _19024_, _19025_, _19026_, _19027_, _19028_, _19029_, _19030_, _19031_, _19032_, _19033_, _19034_, _19035_, _19036_, _19037_, _19038_, _19039_, _19040_, _19041_, _19042_, _19043_, _19044_, _19045_, _19046_, _19047_, _19048_, _19049_, _19050_, _19051_, _19052_, _19053_, _19054_, _19055_, _19056_, _19057_, _19058_, _19059_, _19060_, _19061_, _19062_, _19063_, _19064_, _19065_, _19066_, _19067_, _19068_, _19069_, _19070_, _19071_, _19072_, _19073_, _19074_, _19075_, _19076_, _19077_, _19078_, _19079_, _19080_, _19081_, _19082_, _19083_, _19084_, _19085_, _19086_, _19087_, _19088_, _19089_, _19090_, _19091_, _19092_, _19093_, _19094_, _19095_, _19096_, _19097_, _19098_, _19099_, _19100_, _19101_, _19102_, _19103_, _19104_, _19105_, _19106_, _19107_, _19108_, _19109_, _19110_, _19111_, _19112_, _19113_, _19114_, _19115_, _19116_, _19117_, _19118_, _19119_, _19120_, _19121_, _19122_, _19123_, _19124_, _19125_, _19126_, _19127_, _19128_, _19129_, _19130_, _19131_, _19132_, _19133_, _19134_, _19135_, _19136_, _19137_, _19138_, _19139_, _19140_, _19141_, _19142_, _19143_, _19144_, _19145_, _19146_, _19147_, _19148_, _19149_, _19150_, _19151_, _19152_, _19153_, _19154_, _19155_, _19156_, _19157_, _19158_, _19159_, _19160_, _19161_, _19162_, _19163_, _19164_, _19165_, _19166_, _19167_, _19168_, _19169_, _19170_, _19171_, _19172_, _19173_, _19174_, _19175_, _19176_, _19177_, _19178_, _19179_, _19180_, _19181_, _19182_, _19183_, _19184_, _19185_, _19186_, _19187_, _19188_, _19189_, _19190_, _19191_, _19192_, _19193_, _19194_, _19195_, _19196_, _19197_, _19198_, _19199_, _19200_, _19201_, _19202_, _19203_, _19204_, _19205_, _19206_, _19207_, _19208_, _19209_, _19210_, _19211_, _19212_, _19213_, _19214_, _19215_, _19216_, _19217_, _19218_, _19219_, _19220_, _19221_, _19222_, _19223_, _19224_, _19225_, _19226_, _19227_, _19228_, _19229_, _19230_, _19231_, _19232_, _19233_, _19234_, _19235_, _19236_, _19237_, _19238_, _19239_, _19240_, _19241_, _19242_, _19243_, _19244_, _19245_, _19246_, _19247_, _19248_, _19249_, _19250_, _19251_, _19252_, _19253_, _19254_, _19255_, _19256_, _19257_, _19258_, _19259_, _19260_, _19261_, _19262_, _19263_, _19264_, _19265_, _19266_, _19267_, _19268_, _19269_, _19270_, _19271_, _19272_, _19273_, _19274_, _19275_, _19276_, _19277_, _19278_, _19279_, _19280_, _19281_, _19282_, _19283_, _19284_, _19285_, _19286_, _19287_, _19288_, _19289_, _19290_, _19291_, _19292_, _19293_, _19294_, _19295_, _19296_, _19297_, _19298_, _19299_, _19300_, _19301_, _19302_, _19303_, _19304_, _19305_, _19306_, _19307_, _19308_, _19309_, _19310_, _19311_, _19312_, _19313_, _19314_, _19315_, _19316_, _19317_, _19318_, _19319_, _19320_, _19321_, _19322_, _19323_, _19324_, _19325_, _19326_, _19327_, _19328_, _19329_, _19330_, _19331_, _19332_, _19333_, _19334_, _19335_, _19336_, _19337_, _19338_, _19339_, _19340_, _19341_, _19342_, _19343_, _19344_, _19345_, _19346_, _19347_, _19348_, _19349_, _19350_, _19351_, _19352_, _19353_, _19354_, _19355_, _19356_, _19357_, _19358_, _19359_, _19360_, _19361_, _19362_, _19363_, _19364_, _19365_, _19366_, _19367_, _19368_, _19369_, _19370_, _19371_, _19372_, _19373_, _19374_, _19375_, _19376_, _19377_, _19378_, _19379_, _19380_, _19381_, _19382_, _19383_, _19384_, _19385_, _19386_, _19387_, _19388_, _19389_, _19390_, _19391_, _19392_, _19393_, _19394_, _19395_, _19396_, _19397_, _19398_, _19399_, _19400_, _19401_, _19402_, _19403_, _19404_, _19405_, _19406_, _19407_, _19408_, _19409_, _19410_, _19411_, _19412_, _19413_, _19414_, _19415_, _19416_, _19417_, _19418_, _19419_, _19420_, _19421_, _19422_, _19423_, _19424_, _19425_, _19426_, _19427_, _19428_, _19429_, _19430_, _19431_, _19432_, _19433_, _19434_, _19435_, _19436_, _19437_, _19438_, _19439_, _19440_, _19441_, _19442_, _19443_, _19444_, _19445_, _19446_, _19447_, _19448_, _19449_, _19450_, _19451_, _19452_, _19453_, _19454_, _19455_, _19456_, _19457_, _19458_, _19459_, _19460_, _19461_, _19462_, _19463_, _19464_, _19465_, _19466_, _19467_, _19468_, _19469_, _19470_, _19471_, _19472_, _19473_, _19474_, _19475_, _19476_, _19477_, _19478_, _19479_, _19480_, _19481_, _19482_, _19483_, _19484_, _19485_, _19486_, _19487_, _19488_, _19489_, _19490_, _19491_, _19492_, _19493_, _19494_, _19495_, _19496_, _19497_, _19498_, _19499_, _19500_, _19501_, _19502_, _19503_, _19504_, _19505_, _19506_, _19507_, _19508_, _19509_, _19510_, _19511_, _19512_, _19513_, _19514_, _19515_, _19516_, _19517_, _19518_, _19519_, _19520_, _19521_, _19522_, _19523_, _19524_, _19525_, _19526_, _19527_, _19528_, _19529_, _19530_, _19531_, _19532_, _19533_, _19534_, _19535_, _19536_, _19537_, _19538_, _19539_, _19540_, _19541_, _19542_, _19543_, _19544_, _19545_, _19546_, _19547_, _19548_, _19549_, _19550_, _19551_, _19552_, _19553_, _19554_, _19555_, _19556_, _19557_, _19558_, _19559_, _19560_, _19561_, _19562_, _19563_, _19564_, _19565_, _19566_, _19567_, _19568_, _19569_, _19570_, _19571_, _19572_, _19573_, _19574_, _19575_, _19576_, _19577_, _19578_, _19579_, _19580_, _19581_, _19582_, _19583_, _19584_, _19585_, _19586_, _19587_, _19588_, _19589_, _19590_, _19591_, _19592_, _19593_, _19594_, _19595_, _19596_, _19597_, _19598_, _19599_, _19600_, _19601_, _19602_, _19603_, _19604_, _19605_, _19606_, _19607_, _19608_, _19609_, _19610_, _19611_, _19612_, _19613_, _19614_, _19615_, _19616_, _19617_, _19618_, _19619_, _19620_, _19621_, _19622_, _19623_, _19624_, _19625_, _19626_, _19627_, _19628_, _19629_, _19630_, _19631_, _19632_, _19633_, _19634_, _19635_, _19636_, _19637_, _19638_, _19639_, _19640_, _19641_, _19642_, _19643_, _19644_, _19645_, _19646_, _19647_, _19648_, _19649_, _19650_, _19651_, _19652_, _19653_, _19654_, _19655_, _19656_, _19657_, _19658_, _19659_, _19660_, _19661_, _19662_, _19663_, _19664_, _19665_, _19666_, _19667_, _19668_, _19669_, _19670_, _19671_, _19672_, _19673_, _19674_, _19675_, _19676_, _19677_, _19678_, _19679_, _19680_, _19681_, _19682_, _19683_, _19684_, _19685_, _19686_, _19687_, _19688_, _19689_, _19690_, _19691_, _19692_, _19693_, _19694_, _19695_, _19696_, _19697_, _19698_, _19699_, _19700_, _19701_, _19702_, _19703_, _19704_, _19705_, _19706_, _19707_, _19708_, _19709_, _19710_, _19711_, _19712_, _19713_, _19714_, _19715_, _19716_, _19717_, _19718_, _19719_, _19720_, _19721_, _19722_, _19723_, _19724_, _19725_, _19726_, _19727_, _19728_, _19729_, _19730_, _19731_, _19732_, _19733_, _19734_, _19735_, _19736_, _19737_, _19738_, _19739_, _19740_, _19741_, _19742_, _19743_, _19744_, _19745_, _19746_, _19747_, _19748_, _19749_, _19750_, _19751_, _19752_, _19753_, _19754_, _19755_, _19756_, _19757_, _19758_, _19759_, _19760_, _19761_, _19762_, _19763_, _19764_, _19765_, _19766_, _19767_, _19768_, _19769_, _19770_, _19771_, _19772_, _19773_, _19774_, _19775_, _19776_, _19777_, _19778_, _19779_, _19780_, _19781_, _19782_, _19783_, _19784_, _19785_, _19786_, _19787_, _19788_, _19789_, _19790_, _19791_, _19792_, _19793_, _19794_, _19795_, _19796_, _19797_, _19798_, _19799_, _19800_, _19801_, _19802_, _19803_, _19804_, _19805_, _19806_, _19807_, _19808_, _19809_, _19810_, _19811_, _19812_, _19813_, _19814_, _19815_, _19816_, _19817_, _19818_, _19819_, _19820_, _19821_, _19822_, _19823_, _19824_, _19825_, _19826_, _19827_, _19828_, _19829_, _19830_, _19831_, _19832_, _19833_, _19834_, _19835_, _19836_, _19837_, _19838_, _19839_, _19840_, _19841_, _19842_, _19843_, _19844_, _19845_, _19846_, _19847_, _19848_, _19849_, _19850_, _19851_, _19852_, _19853_, _19854_, _19855_, _19856_, _19857_, _19858_, _19859_, _19860_, _19861_, _19862_, _19863_, _19864_, _19865_, _19866_, _19867_, _19868_, _19869_, _19870_, _19871_, _19872_, _19873_, _19874_, _19875_, _19876_, _19877_, _19878_, _19879_, _19880_, _19881_, _19882_, _19883_, _19884_, _19885_, _19886_, _19887_, _19888_, _19889_, _19890_, _19891_, _19892_, _19893_, _19894_, _19895_, _19896_, _19897_, _19898_, _19899_, _19900_, _19901_, _19902_, _19903_, _19904_, _19905_, _19906_, _19907_, _19908_, _19909_, _19910_, _19911_, _19912_, _19913_, _19914_, _19915_, _19916_, _19917_, _19918_, _19919_, _19920_, _19921_, _19922_, _19923_, _19924_, _19925_, _19926_, _19927_, _19928_, _19929_, _19930_, _19931_, _19932_, _19933_, _19934_, _19935_, _19936_, _19937_, _19938_, _19939_, _19940_, _19941_, _19942_, _19943_, _19944_, _19945_, _19946_, _19947_, _19948_, _19949_, _19950_, _19951_, _19952_, _19953_, _19954_, _19955_, _19956_, _19957_, _19958_, _19959_, _19960_, _19961_, _19962_, _19963_, _19964_, _19965_, _19966_, _19967_, _19968_, _19969_, _19970_, _19971_, _19972_, _19973_, _19974_, _19975_, _19976_, _19977_, _19978_, _19979_, _19980_, _19981_, _19982_, _19983_, _19984_, _19985_, _19986_, _19987_, _19988_, _19989_, _19990_, _19991_, _19992_, _19993_, _19994_, _19995_, _19996_, _19997_, _19998_, _19999_, _20000_, _20001_, _20002_, _20003_, _20004_, _20005_, _20006_, _20007_, _20008_, _20009_, _20010_, _20011_, _20012_, _20013_, _20014_, _20015_, _20016_, _20017_, _20018_, _20019_, _20020_, _20021_, _20022_, _20023_, _20024_, _20025_, _20026_, _20027_, _20028_, _20029_, _20030_, _20031_, _20032_, _20033_, _20034_, _20035_, _20036_, _20037_, _20038_, _20039_, _20040_, _20041_, _20042_, _20043_, _20044_, _20045_, _20046_, _20047_, _20048_, _20049_, _20050_, _20051_, _20052_, _20053_, _20054_, _20055_, _20056_, _20057_, _20058_, _20059_, _20060_, _20061_, _20062_, _20063_, _20064_, _20065_, _20066_, _20067_, _20068_, _20069_, _20070_, _20071_, _20072_, _20073_, _20074_, _20075_, _20076_, _20077_, _20078_, _20079_, _20080_, _20081_, _20082_, _20083_, _20084_, _20085_, _20086_, _20087_, _20088_, _20089_, _20090_, _20091_, _20092_, _20093_, _20094_, _20095_, _20096_, _20097_, _20098_, _20099_, _20100_, _20101_, _20102_, _20103_, _20104_, _20105_, _20106_, _20107_, _20108_, _20109_, _20110_, _20111_, _20112_, _20113_, _20114_, _20115_, _20116_, _20117_, _20118_, _20119_, _20120_, _20121_, _20122_, _20123_, _20124_, _20125_, _20126_, _20127_, _20128_, _20129_, _20130_, _20131_, _20132_, _20133_, _20134_, _20135_, _20136_, _20137_, _20138_, _20139_, _20140_, _20141_, _20142_, _20143_, _20144_, _20145_, _20146_, _20147_, _20148_, _20149_, _20150_, _20151_, _20152_, _20153_, _20154_, _20155_, _20156_, _20157_, _20158_, _20159_, _20160_, _20161_, _20162_, _20163_, _20164_, _20165_, _20166_, _20167_, _20168_, _20169_, _20170_, _20171_, _20172_, _20173_, _20174_, _20175_, _20176_, _20177_, _20178_, _20179_, _20180_, _20181_, _20182_, _20183_, _20184_, _20185_, _20186_, _20187_, _20188_, _20189_, _20190_, _20191_, _20192_, _20193_, _20194_, _20195_, _20196_, _20197_, _20198_, _20199_, _20200_, _20201_, _20202_, _20203_, _20204_, _20205_, _20206_, _20207_, _20208_, _20209_, _20210_, _20211_, _20212_, _20213_, _20214_, _20215_, _20216_, _20217_, _20218_, _20219_, _20220_, _20221_, _20222_, _20223_, _20224_, _20225_, _20226_, _20227_, _20228_, _20229_, _20230_, _20231_, _20232_, _20233_, _20234_, _20235_, _20236_, _20237_, _20238_, _20239_, _20240_, _20241_, _20242_, _20243_, _20244_, _20245_, _20246_, _20247_, _20248_, _20249_, _20250_, _20251_, _20252_, _20253_, _20254_, _20255_, _20256_, _20257_, _20258_, _20259_, _20260_, _20261_, _20262_, _20263_, _20264_, _20265_, _20266_, _20267_, _20268_, _20269_, _20270_, _20271_, _20272_, _20273_, _20274_, _20275_, _20276_, _20277_, _20278_, _20279_, _20280_, _20281_, _20282_, _20283_, _20284_, _20285_, _20286_, _20287_, _20288_, _20289_, _20290_, _20291_, _20292_, _20293_, _20294_, _20295_, _20296_, _20297_, _20298_, _20299_, _20300_, _20301_, _20302_, _20303_, _20304_, _20305_, _20306_, _20307_, _20308_, _20309_, _20310_, _20311_, _20312_, _20313_, _20314_, _20315_, _20316_, _20317_, _20318_, _20319_, _20320_, _20321_, _20322_, _20323_, _20324_, _20325_, _20326_, _20327_, _20328_, _20329_, _20330_, _20331_, _20332_, _20333_, _20334_, _20335_, _20336_, _20337_, _20338_, _20339_, _20340_, _20341_, _20342_, _20343_, _20344_, _20345_, _20346_, _20347_, _20348_, _20349_, _20350_, _20351_, _20352_, _20353_, _20354_, _20355_, _20356_, _20357_, _20358_, _20359_, _20360_, _20361_, _20362_, _20363_, _20364_, _20365_, _20366_, _20367_, _20368_, _20369_, _20370_, _20371_, _20372_, _20373_, _20374_, _20375_, _20376_, _20377_, _20378_, _20379_, _20380_, _20381_, _20382_, _20383_, _20384_, _20385_, _20386_, _20387_, _20388_, _20389_, _20390_, _20391_, _20392_, _20393_, _20394_, _20395_, _20396_, _20397_, _20398_, _20399_, _20400_, _20401_, _20402_, _20403_, _20404_, _20405_, _20406_, _20407_, _20408_, _20409_, _20410_, _20411_, _20412_, _20413_, _20414_, _20415_, _20416_, _20417_, _20418_, _20419_, _20420_, _20421_, _20422_, _20423_, _20424_, _20425_, _20426_, _20427_, _20428_, _20429_, _20430_, _20431_, _20432_, _20433_, _20434_, _20435_, _20436_, _20437_, _20438_, _20439_, _20440_, _20441_, _20442_, _20443_, _20444_, _20445_, _20446_, _20447_, _20448_, _20449_, _20450_, _20451_, _20452_, _20453_, _20454_, _20455_, _20456_, _20457_, _20458_, _20459_, _20460_, _20461_, _20462_, _20463_, _20464_, _20465_, _20466_, _20467_, _20468_, _20469_, _20470_, _20471_, _20472_, _20473_, _20474_, _20475_, _20476_, _20477_, _20478_, _20479_, _20480_, _20481_, _20482_, _20483_, _20484_, _20485_, _20486_, _20487_, _20488_, _20489_, _20490_, _20491_, _20492_, _20493_, _20494_, _20495_, _20496_, _20497_, _20498_, _20499_, _20500_, _20501_, _20502_, _20503_, _20504_, _20505_, _20506_, _20507_, _20508_, _20509_, _20510_, _20511_, _20512_, _20513_, _20514_, _20515_, _20516_, _20517_, _20518_, _20519_, _20520_, _20521_, _20522_, _20523_, _20524_, _20525_, _20526_, _20527_, _20528_, _20529_, _20530_, _20531_, _20532_, _20533_, _20534_, _20535_, _20536_, _20537_, _20538_, _20539_, _20540_, _20541_, _20542_, _20543_, _20544_, _20545_, _20546_, _20547_, _20548_, _20549_, _20550_, _20551_, _20552_, _20553_, _20554_, _20555_, _20556_, _20557_, _20558_, _20559_, _20560_, _20561_, _20562_, _20563_, _20564_, _20565_, _20566_, _20567_, _20568_, _20569_, _20570_, _20571_, _20572_, _20573_, _20574_, _20575_, _20576_, _20577_, _20578_, _20579_, _20580_, _20581_, _20582_, _20583_, _20584_, _20585_, _20586_, _20587_, _20588_, _20589_, _20590_, _20591_, _20592_, _20593_, _20594_, _20595_, _20596_, _20597_, _20598_, _20599_, _20600_, _20601_, _20602_, _20603_, _20604_, _20605_, _20606_, _20607_, _20608_, _20609_, _20610_, _20611_, _20612_, _20613_, _20614_, _20615_, _20616_, _20617_, _20618_, _20619_, _20620_, _20621_, _20622_, _20623_, _20624_, _20625_, _20626_, _20627_, _20628_, _20629_, _20630_, _20631_, _20632_, _20633_, _20634_, _20635_, _20636_, _20637_, _20638_, _20639_, _20640_, _20641_, _20642_, _20643_, _20644_, _20645_, _20646_, _20647_, _20648_, _20649_, _20650_, _20651_, _20652_, _20653_, _20654_, _20655_, _20656_, _20657_, _20658_, _20659_, _20660_, _20661_, _20662_, _20663_, _20664_, _20665_, _20666_, _20667_, _20668_, _20669_, _20670_, _20671_, _20672_, _20673_, _20674_, _20675_, _20676_, _20677_, _20678_, _20679_, _20680_, _20681_, _20682_, _20683_, _20684_, _20685_, _20686_, _20687_, _20688_, _20689_, _20690_, _20691_, _20692_, _20693_, _20694_, _20695_, _20696_, _20697_, _20698_, _20699_, _20700_, _20701_, _20702_, _20703_, _20704_, _20705_, _20706_, _20707_, _20708_, _20709_, _20710_, _20711_, _20712_, _20713_, _20714_, _20715_, _20716_, _20717_, _20718_, _20719_, _20720_, _20721_, _20722_, _20723_, _20724_, _20725_, _20726_, _20727_, _20728_, _20729_, _20730_, _20731_, _20732_, _20733_, _20734_, _20735_, _20736_, _20737_, _20738_, _20739_, _20740_, _20741_, _20742_, _20743_, _20744_, _20745_, _20746_, _20747_, _20748_, _20749_, _20750_, _20751_, _20752_, _20753_, _20754_, _20755_, _20756_, _20757_, _20758_, _20759_, _20760_, _20761_, _20762_, _20763_, _20764_, _20765_, _20766_, _20767_, _20768_, _20769_, _20770_, _20771_, _20772_, _20773_, _20774_, _20775_, _20776_, _20777_, _20778_, _20779_, _20780_, _20781_, _20782_, _20783_, _20784_, _20785_, _20786_, _20787_, _20788_, _20789_, _20790_, _20791_, _20792_, _20793_, _20794_, _20795_, _20796_, _20797_, _20798_, _20799_, _20800_, _20801_, _20802_, _20803_, _20804_, _20805_, _20806_, _20807_, _20808_, _20809_, _20810_, _20811_, _20812_, _20813_, _20814_, _20815_, _20816_, _20817_, _20818_, _20819_, _20820_, _20821_, _20822_, _20823_, _20824_, _20825_, _20826_, _20827_, _20828_, _20829_, _20830_, _20831_, _20832_, _20833_, _20834_, _20835_, _20836_, _20837_, _20838_, _20839_, _20840_, _20841_, _20842_, _20843_, _20844_, _20845_, _20846_, _20847_, _20848_, _20849_, _20850_, _20851_, _20852_, _20853_, _20854_, _20855_, _20856_, _20857_, _20858_, _20859_, _20860_, _20861_, _20862_, _20863_, _20864_, _20865_, _20866_, _20867_, _20868_, _20869_, _20870_, _20871_, _20872_, _20873_, _20874_, _20875_, _20876_, _20877_, _20878_, _20879_, _20880_, _20881_, _20882_, _20883_, _20884_, _20885_, _20886_, _20887_, _20888_, _20889_, _20890_, _20891_, _20892_, _20893_, _20894_, _20895_, _20896_, _20897_, _20898_, _20899_, _20900_, _20901_, _20902_, _20903_, _20904_, _20905_, _20906_, _20907_, _20908_, _20909_, _20910_, _20911_, _20912_, _20913_, _20914_, _20915_, _20916_, _20917_, _20918_, _20919_, _20920_, _20921_, _20922_, _20923_, _20924_, _20925_, _20926_, _20927_, _20928_, _20929_, _20930_, _20931_, _20932_, _20933_, _20934_, _20935_, _20936_, _20937_, _20938_, _20939_, _20940_, _20941_, _20942_, _20943_, _20944_, _20945_, _20946_, _20947_, _20948_, _20949_, _20950_, _20951_, _20952_, _20953_, _20954_, _20955_, _20956_, _20957_, _20958_, _20959_, _20960_, _20961_, _20962_, _20963_, _20964_, _20965_, _20966_, _20967_, _20968_, _20969_, _20970_, _20971_, _20972_, _20973_, _20974_, _20975_, _20976_, _20977_, _20978_, _20979_, _20980_, _20981_, _20982_, _20983_, _20984_, _20985_, _20986_, _20987_, _20988_, _20989_, _20990_, _20991_, _20992_, _20993_, _20994_, _20995_, _20996_, _20997_, _20998_, _20999_, _21000_, _21001_, _21002_, _21003_, _21004_, _21005_, _21006_, _21007_, _21008_, _21009_, _21010_, _21011_, _21012_, _21013_, _21014_, _21015_, _21016_, _21017_, _21018_, _21019_, _21020_, _21021_, _21022_, _21023_, _21024_, _21025_, _21026_, _21027_, _21028_, _21029_, _21030_, _21031_, _21032_, _21033_, _21034_, _21035_, _21036_, _21037_, _21038_, _21039_, _21040_, _21041_, _21042_, _21043_, _21044_, _21045_, _21046_, _21047_, _21048_, _21049_, _21050_, _21051_, _21052_, _21053_, _21054_, _21055_, _21056_, _21057_, _21058_, _21059_, _21060_, _21061_, _21062_, _21063_, _21064_, _21065_, _21066_, _21067_, _21068_, _21069_, _21070_, _21071_, _21072_, _21073_, _21074_, _21075_, _21076_, _21077_, _21078_, _21079_, _21080_, _21081_, _21082_, _21083_, _21084_, _21085_, _21086_, _21087_, _21088_, _21089_, _21090_, _21091_, _21092_, _21093_, _21094_, _21095_, _21096_, _21097_, _21098_, _21099_, _21100_, _21101_, _21102_, _21103_, _21104_, _21105_, _21106_, _21107_, _21108_, _21109_, _21110_, _21111_, _21112_, _21113_, _21114_, _21115_, _21116_, _21117_, _21118_, _21119_, _21120_, _21121_, _21122_, _21123_, _21124_, _21125_, _21126_, _21127_, _21128_, _21129_, _21130_, _21131_, _21132_, _21133_, _21134_, _21135_, _21136_, _21137_, _21138_, _21139_, _21140_, _21141_, _21142_, _21143_, _21144_, _21145_, _21146_, _21147_, _21148_, _21149_, _21150_, _21151_, _21152_, _21153_, _21154_, _21155_, _21156_, _21157_, _21158_, _21159_, _21160_, _21161_, _21162_, _21163_, _21164_, _21165_, _21166_, _21167_, _21168_, _21169_, _21170_, _21171_, _21172_, _21173_, _21174_, _21175_, _21176_, _21177_, _21178_, _21179_, _21180_, _21181_, _21182_, _21183_, _21184_, _21185_, _21186_, _21187_, _21188_, _21189_, _21190_, _21191_, _21192_, _21193_, _21194_, _21195_, _21196_, _21197_, _21198_, _21199_, _21200_, _21201_, _21202_, _21203_, _21204_, _21205_, _21206_, _21207_, _21208_, _21209_, _21210_, _21211_, _21212_, _21213_, _21214_, _21215_, _21216_, _21217_, _21218_, _21219_, _21220_, _21221_, _21222_, _21223_, _21224_, _21225_, _21226_, _21227_, _21228_, _21229_, _21230_, _21231_, _21232_, _21233_, _21234_, _21235_, _21236_, _21237_, _21238_, _21239_, _21240_, _21241_, _21242_, _21243_, _21244_, _21245_, _21246_, _21247_, _21248_, _21249_, _21250_, _21251_, _21252_, _21253_, _21254_, _21255_, _21256_, _21257_, _21258_, _21259_, _21260_, _21261_, _21262_, _21263_, _21264_, _21265_, _21266_, _21267_, _21268_, _21269_, _21270_, _21271_, _21272_, _21273_, _21274_, _21275_, _21276_, _21277_, _21278_, _21279_, _21280_, _21281_, _21282_, _21283_, _21284_, _21285_, _21286_, _21287_, _21288_, _21289_, _21290_, _21291_, _21292_, _21293_, _21294_, _21295_, _21296_, _21297_, _21298_, _21299_, _21300_, _21301_, _21302_, _21303_, _21304_, _21305_, _21306_, _21307_, _21308_, _21309_, _21310_, _21311_, _21312_, _21313_, _21314_, _21315_, _21316_, _21317_, _21318_, _21319_, _21320_, _21321_, _21322_, _21323_, _21324_, _21325_, _21326_, _21327_, _21328_, _21329_, _21330_, _21331_, _21332_, _21333_, _21334_, _21335_, _21336_, _21337_, _21338_, _21339_, _21340_, _21341_, _21342_, _21343_, _21344_, _21345_, _21346_, _21347_, _21348_, _21349_, _21350_, _21351_, _21352_, _21353_, _21354_, _21355_, _21356_, _21357_, _21358_, _21359_, _21360_, _21361_, _21362_, _21363_, _21364_, _21365_, _21366_, _21367_, _21368_, _21369_, _21370_, _21371_, _21372_, _21373_, _21374_, _21375_, _21376_, _21377_, _21378_, _21379_, _21380_, _21381_, _21382_, _21383_, _21384_, _21385_, _21386_, _21387_, _21388_, _21389_, _21390_, _21391_, _21392_, _21393_, _21394_, _21395_, _21396_, _21397_, _21398_, _21399_, _21400_, _21401_, _21402_, _21403_, _21404_, _21405_, _21406_, _21407_, _21408_, _21409_, _21410_, _21411_, _21412_, _21413_, _21414_, _21415_, _21416_, _21417_, _21418_, _21419_, _21420_, _21421_, _21422_, _21423_, _21424_, _21425_, _21426_, _21427_, _21428_, _21429_, _21430_, _21431_, _21432_, _21433_, _21434_, _21435_, _21436_, _21437_, _21438_, _21439_, _21440_, _21441_, _21442_, _21443_, _21444_, _21445_, _21446_, _21447_, _21448_, _21449_, _21450_, _21451_, _21452_, _21453_, _21454_, _21455_, _21456_, _21457_, _21458_, _21459_, _21460_, _21461_, _21462_, _21463_, _21464_, _21465_, _21466_, _21467_, _21468_, _21469_, _21470_, _21471_, _21472_, _21473_, _21474_, _21475_, _21476_, _21477_, _21478_, _21479_, _21480_, _21481_, _21482_, _21483_, _21484_, _21485_, _21486_, _21487_, _21488_, _21489_, _21490_, _21491_, _21492_, _21493_, _21494_, _21495_, _21496_, _21497_, _21498_, _21499_, _21500_, _21501_, _21502_, _21503_, _21504_, _21505_, _21506_, _21507_, _21508_, _21509_, _21510_, _21511_, _21512_, _21513_, _21514_, _21515_, _21516_, _21517_, _21518_, _21519_, _21520_, _21521_, _21522_, _21523_, _21524_, _21525_, _21526_, _21527_, _21528_, _21529_, _21530_, _21531_, _21532_, _21533_, _21534_, _21535_, _21536_, _21537_, _21538_, _21539_, _21540_, _21541_, _21542_, _21543_, _21544_, _21545_, _21546_, _21547_, _21548_, _21549_, _21550_, _21551_, _21552_, _21553_, _21554_, _21555_, _21556_, _21557_, _21558_, _21559_, _21560_, _21561_, _21562_, _21563_, _21564_, _21565_, _21566_, _21567_, _21568_, _21569_, _21570_, _21571_, _21572_, _21573_, _21574_, _21575_, _21576_, _21577_, _21578_, _21579_, _21580_, _21581_, _21582_, _21583_, _21584_, _21585_, _21586_, _21587_, _21588_, _21589_, _21590_, _21591_, _21592_, _21593_, _21594_, _21595_, _21596_, _21597_, _21598_, _21599_, _21600_, _21601_, _21602_, _21603_, _21604_, _21605_, _21606_, _21607_, _21608_, _21609_, _21610_, _21611_, _21612_, _21613_, _21614_, _21615_, _21616_, _21617_, _21618_, _21619_, _21620_, _21621_, _21622_, _21623_, _21624_, _21625_, _21626_, _21627_, _21628_, _21629_, _21630_, _21631_, _21632_, _21633_, _21634_, _21635_, _21636_, _21637_, _21638_, _21639_, _21640_, _21641_, _21642_, _21643_, _21644_, _21645_, _21646_, _21647_, _21648_, _21649_, _21650_, _21651_, _21652_, _21653_, _21654_, _21655_, _21656_, _21657_, _21658_, _21659_, _21660_, _21661_, _21662_, _21663_, _21664_, _21665_, _21666_, _21667_, _21668_, _21669_, _21670_, _21671_, _21672_, _21673_, _21674_, _21675_, _21676_, _21677_, _21678_, _21679_, _21680_, _21681_, _21682_, _21683_, _21684_, _21685_, _21686_, _21687_, _21688_, _21689_, _21690_, _21691_, _21692_, _21693_, _21694_, _21695_, _21696_, _21697_, _21698_, _21699_, _21700_, _21701_, _21702_, _21703_, _21704_, _21705_, _21706_, _21707_, _21708_, _21709_, _21710_, _21711_, _21712_, _21713_, _21714_, _21715_, _21716_, _21717_, _21718_, _21719_, _21720_, _21721_, _21722_, _21723_, _21724_, _21725_, _21726_, _21727_, _21728_, _21729_, _21730_, _21731_, _21732_, _21733_, _21734_, _21735_, _21736_, _21737_, _21738_, _21739_, _21740_, _21741_, _21742_, _21743_, _21744_, _21745_, _21746_, _21747_, _21748_, _21749_, _21750_, _21751_, _21752_, _21753_, _21754_, _21755_, _21756_, _21757_, _21758_, _21759_, _21760_, _21761_, _21762_, _21763_, _21764_, _21765_, _21766_, _21767_, _21768_, _21769_, _21770_, _21771_, _21772_, _21773_, _21774_, _21775_, _21776_, _21777_, _21778_, _21779_, _21780_, _21781_, _21782_, _21783_, _21784_, _21785_, _21786_, _21787_, _21788_, _21789_, _21790_, _21791_, _21792_, _21793_, _21794_, _21795_, _21796_, _21797_, _21798_, _21799_, _21800_, _21801_, _21802_, _21803_, _21804_, _21805_, _21806_, _21807_, _21808_, _21809_, _21810_, _21811_, _21812_, _21813_, _21814_, _21815_, _21816_, _21817_, _21818_, _21819_, _21820_, _21821_, _21822_, _21823_, _21824_, _21825_, _21826_, _21827_, _21828_, _21829_, _21830_, _21831_, _21832_, _21833_, _21834_, _21835_, _21836_, _21837_, _21838_, _21839_, _21840_, _21841_, _21842_, _21843_, _21844_, _21845_, _21846_, _21847_, _21848_, _21849_, _21850_, _21851_, _21852_, _21853_, _21854_, _21855_, _21856_, _21857_, _21858_, _21859_, _21860_, _21861_, _21862_, _21863_, _21864_, _21865_, _21866_, _21867_, _21868_, _21869_, _21870_, _21871_, _21872_, _21873_, _21874_, _21875_, _21876_, _21877_, _21878_, _21879_, _21880_, _21881_, _21882_, _21883_, _21884_, _21885_, _21886_, _21887_, _21888_, _21889_, _21890_, _21891_, _21892_, _21893_, _21894_, _21895_, _21896_, _21897_, _21898_, _21899_, _21900_, _21901_, _21902_, _21903_, _21904_, _21905_, _21906_, _21907_, _21908_, _21909_, _21910_, _21911_, _21912_, _21913_, _21914_, _21915_, _21916_, _21917_, _21918_, _21919_, _21920_, _21921_, _21922_, _21923_, _21924_, _21925_, _21926_, _21927_, _21928_, _21929_, _21930_, _21931_, _21932_, _21933_, _21934_, _21935_, _21936_, _21937_, _21938_, _21939_, _21940_, _21941_, _21942_, _21943_, _21944_, _21945_, _21946_, _21947_, _21948_, _21949_, _21950_, _21951_, _21952_, _21953_, _21954_, _21955_, _21956_, _21957_, _21958_, _21959_, _21960_, _21961_, _21962_, _21963_, _21964_, _21965_, _21966_, _21967_, _21968_, _21969_, _21970_, _21971_, _21972_, _21973_, _21974_, _21975_, _21976_, _21977_, _21978_, _21979_, _21980_, _21981_, _21982_, _21983_, _21984_, _21985_, _21986_, _21987_, _21988_, _21989_, _21990_, _21991_, _21992_, _21993_, _21994_, _21995_, _21996_, _21997_, _21998_, _21999_, _22000_, _22001_, _22002_, _22003_, _22004_, _22005_, _22006_, _22007_, _22008_, _22009_, _22010_, _22011_, _22012_, _22013_, _22014_, _22015_, _22016_, _22017_, _22018_, _22019_, _22020_, _22021_, _22022_, _22023_, _22024_, _22025_, _22026_, _22027_, _22028_, _22029_, _22030_, _22031_, _22032_, _22033_, _22034_, _22035_, _22036_, _22037_, _22038_, _22039_, _22040_, _22041_, _22042_, _22043_, _22044_, _22045_, _22046_, _22047_, _22048_, _22049_, _22050_, _22051_, _22052_, _22053_, _22054_, _22055_, _22056_, _22057_, _22058_, _22059_, _22060_, _22061_, _22062_, _22063_, _22064_, _22065_, _22066_, _22067_, _22068_, _22069_, _22070_, _22071_, _22072_, _22073_, _22074_, _22075_, _22076_, _22077_, _22078_, _22079_, _22080_, _22081_, _22082_, _22083_, _22084_, _22085_, _22086_, _22087_, _22088_, _22089_, _22090_, _22091_, _22092_, _22093_, _22094_, _22095_, _22096_, _22097_, _22098_, _22099_, _22100_, _22101_, _22102_, _22103_, _22104_, _22105_, _22106_, _22107_, _22108_, _22109_, _22110_, _22111_, _22112_, _22113_, _22114_, _22115_, _22116_, _22117_, _22118_, _22119_, _22120_, _22121_, _22122_, _22123_, _22124_, _22125_, _22126_, _22127_, _22128_, _22129_, _22130_, _22131_, _22132_, _22133_, _22134_, _22135_, _22136_, _22137_, _22138_, _22139_, _22140_, _22141_, _22142_, _22143_, _22144_, _22145_, _22146_, _22147_, _22148_, _22149_, _22150_, _22151_, _22152_, _22153_, _22154_, _22155_, _22156_, _22157_, _22158_, _22159_, _22160_, _22161_, _22162_, _22163_, _22164_, _22165_, _22166_, _22167_, _22168_, _22169_, _22170_, _22171_, _22172_, _22173_, _22174_, _22175_, _22176_, _22177_, _22178_, _22179_, _22180_, _22181_, _22182_, _22183_, _22184_, _22185_, _22186_, _22187_, _22188_, _22189_, _22190_, _22191_, _22192_, _22193_, _22194_, _22195_, _22196_, _22197_, _22198_, _22199_, _22200_, _22201_, _22202_, _22203_, _22204_, _22205_, _22206_, _22207_, _22208_, _22209_, _22210_, _22211_, _22212_, _22213_, _22214_, _22215_, _22216_, _22217_, _22218_, _22219_, _22220_, _22221_, _22222_, _22223_, _22224_, _22225_, _22226_, _22227_, _22228_, _22229_, _22230_, _22231_, _22232_, _22233_, _22234_, _22235_, _22236_, _22237_, _22238_, _22239_, _22240_, _22241_, _22242_, _22243_, _22244_, _22245_, _22246_, _22247_, _22248_, _22249_, _22250_, _22251_, _22252_, _22253_, _22254_, _22255_, _22256_, _22257_, _22258_, _22259_, _22260_, _22261_, _22262_, _22263_, _22264_, _22265_, _22266_, _22267_, _22268_, _22269_, _22270_, _22271_, _22272_, _22273_, _22274_, _22275_, _22276_, _22277_, _22278_, _22279_, _22280_, _22281_, _22282_, _22283_, _22284_, _22285_, _22286_, _22287_, _22288_, _22289_, _22290_, _22291_, _22292_, _22293_, _22294_, _22295_, _22296_, _22297_, _22298_, _22299_, _22300_, _22301_, _22302_, _22303_, _22304_, _22305_, _22306_, _22307_, _22308_, _22309_, _22310_, _22311_, _22312_, _22313_, _22314_, _22315_, _22316_, _22317_, _22318_, _22319_, _22320_, _22321_, _22322_, _22323_, _22324_, _22325_, _22326_, _22327_, _22328_, _22329_, _22330_, _22331_, _22332_, _22333_, _22334_, _22335_, _22336_, _22337_, _22338_, _22339_, _22340_, _22341_, _22342_, _22343_, _22344_, _22345_, _22346_, _22347_, _22348_, _22349_, _22350_, _22351_, _22352_, _22353_, _22354_, _22355_, _22356_, _22357_, _22358_, _22359_, _22360_, _22361_, _22362_, _22363_, _22364_, _22365_, _22366_, _22367_, _22368_, _22369_, _22370_, _22371_, _22372_, _22373_, _22374_, _22375_, _22376_, _22377_, _22378_, _22379_, _22380_, _22381_, _22382_, _22383_, _22384_, _22385_, _22386_, _22387_, _22388_, _22389_, _22390_, _22391_, _22392_, _22393_, _22394_, _22395_, _22396_, _22397_, _22398_, _22399_, _22400_, _22401_, _22402_, _22403_, _22404_, _22405_, _22406_, _22407_, _22408_, _22409_, _22410_, _22411_, _22412_, _22413_, _22414_, _22415_, _22416_, _22417_, _22418_, _22419_, _22420_, _22421_, _22422_, _22423_, _22424_, _22425_, _22426_, _22427_, _22428_, _22429_, _22430_, _22431_, _22432_, _22433_, _22434_, _22435_, _22436_, _22437_, _22438_, _22439_, _22440_, _22441_, _22442_, _22443_, _22444_, _22445_, _22446_, _22447_, _22448_, _22449_, _22450_, _22451_, _22452_, _22453_, _22454_, _22455_, _22456_, _22457_, _22458_, _22459_, _22460_, _22461_, _22462_, _22463_, _22464_, _22465_, _22466_, _22467_, _22468_, _22469_, _22470_, _22471_, _22472_, _22473_, _22474_, _22475_, _22476_, _22477_, _22478_, _22479_, _22480_, _22481_, _22482_, _22483_, _22484_, _22485_, _22486_, _22487_, _22488_, _22489_, _22490_, _22491_, _22492_, _22493_, _22494_, _22495_, _22496_, _22497_, _22498_, _22499_, _22500_, _22501_, _22502_, _22503_, _22504_, _22505_, _22506_, _22507_, _22508_, _22509_, _22510_, _22511_, _22512_, _22513_, _22514_, _22515_, _22516_, _22517_, _22518_, _22519_, _22520_, _22521_, _22522_, _22523_, _22524_, _22525_, _22526_, _22527_, _22528_, _22529_, _22530_, _22531_, _22532_, _22533_, _22534_, _22535_, _22536_, _22537_, _22538_, _22539_, _22540_, _22541_, _22542_, _22543_, _22544_, _22545_, _22546_, _22547_, _22548_, _22549_, _22550_, _22551_, _22552_, _22553_, _22554_, _22555_, _22556_, _22557_, _22558_, _22559_, _22560_, _22561_, _22562_, _22563_, _22564_, _22565_, _22566_, _22567_, _22568_, _22569_, _22570_, _22571_, _22572_, _22573_, _22574_, _22575_, _22576_, _22577_, _22578_, _22579_, _22580_, _22581_, _22582_, _22583_, _22584_, _22585_, _22586_, _22587_, _22588_, _22589_, _22590_, _22591_, _22592_, _22593_, _22594_, _22595_, _22596_, _22597_, _22598_, _22599_, _22600_, _22601_, _22602_, _22603_, _22604_, _22605_, _22606_, _22607_, _22608_, _22609_, _22610_, _22611_, _22612_, _22613_, _22614_, _22615_, _22616_, _22617_, _22618_, _22619_, _22620_, _22621_, _22622_, _22623_, _22624_, _22625_, _22626_, _22627_, _22628_, _22629_, _22630_, _22631_, _22632_, _22633_, _22634_, _22635_, _22636_, _22637_, _22638_, _22639_, _22640_, _22641_, _22642_, _22643_, _22644_, _22645_, _22646_, _22647_, _22648_, _22649_, _22650_, _22651_, _22652_, _22653_, _22654_, _22655_, _22656_, _22657_, _22658_, _22659_, _22660_, _22661_, _22662_, _22663_, _22664_, _22665_, _22666_, _22667_, _22668_, _22669_, _22670_, _22671_, _22672_, _22673_, _22674_, _22675_, _22676_, _22677_, _22678_, _22679_, _22680_, _22681_, _22682_, _22683_, _22684_, _22685_, _22686_, _22687_, _22688_, _22689_, _22690_, _22691_, _22692_, _22693_, _22694_, _22695_, _22696_, _22697_, _22698_, _22699_, _22700_, _22701_, _22702_, _22703_, _22704_, _22705_, _22706_, _22707_, _22708_, _22709_, _22710_, _22711_, _22712_, _22713_, _22714_, _22715_, _22716_, _22717_, _22718_, _22719_, _22720_, _22721_, _22722_, _22723_, _22724_, _22725_, _22726_, _22727_, _22728_, _22729_, _22730_, _22731_, _22732_, _22733_, _22734_, _22735_, _22736_, _22737_, _22738_, _22739_, _22740_, _22741_, _22742_, _22743_, _22744_, _22745_, _22746_, _22747_, _22748_, _22749_, _22750_, _22751_, _22752_, _22753_, _22754_, _22755_, _22756_, _22757_, _22758_, _22759_, _22760_, _22761_, _22762_, _22763_, _22764_, _22765_, _22766_, _22767_, _22768_, _22769_, _22770_, _22771_, _22772_, _22773_, _22774_, _22775_, _22776_, _22777_, _22778_, _22779_, _22780_, _22781_, _22782_, _22783_, _22784_, _22785_, _22786_, _22787_, _22788_, _22789_, _22790_, _22791_, _22792_, _22793_, _22794_, _22795_, _22796_, _22797_, _22798_, _22799_, _22800_, _22801_, _22802_, _22803_, _22804_, _22805_, _22806_, _22807_, _22808_, _22809_, _22810_, _22811_, _22812_, _22813_, _22814_, _22815_, _22816_, _22817_, _22818_, _22819_, _22820_, _22821_, _22822_, _22823_, _22824_, _22825_, _22826_, _22827_, _22828_, _22829_, _22830_, _22831_, _22832_, _22833_, _22834_, _22835_, _22836_, _22837_, _22838_, _22839_, _22840_, _22841_, _22842_, _22843_, _22844_, _22845_, _22846_, _22847_, _22848_, _22849_, _22850_, _22851_, _22852_, _22853_, _22854_, _22855_, _22856_, _22857_, _22858_, _22859_, _22860_, _22861_, _22862_, _22863_, _22864_, _22865_, _22866_, _22867_, _22868_, _22869_, _22870_, _22871_, _22872_, _22873_, _22874_, _22875_, _22876_, _22877_, _22878_, _22879_, _22880_, _22881_, _22882_, _22883_, _22884_, _22885_, _22886_, _22887_, _22888_, _22889_, _22890_, _22891_, _22892_, _22893_, _22894_, _22895_, _22896_, _22897_, _22898_, _22899_, _22900_, _22901_, _22902_, _22903_, _22904_, _22905_, _22906_, _22907_, _22908_, _22909_, _22910_, _22911_, _22912_, _22913_, _22914_, _22915_, _22916_, _22917_, _22918_, _22919_, _22920_, _22921_, _22922_, _22923_, _22924_, _22925_, _22926_, _22927_, _22928_, _22929_, _22930_, _22931_, _22932_, _22933_, _22934_, _22935_, _22936_, _22937_, _22938_, _22939_, _22940_, _22941_, _22942_, _22943_, _22944_, _22945_, _22946_, _22947_, _22948_, _22949_, _22950_, _22951_, _22952_, _22953_, _22954_, _22955_, _22956_, _22957_, _22958_, _22959_, _22960_, _22961_, _22962_, _22963_, _22964_, _22965_, _22966_, _22967_, _22968_, _22969_, _22970_, _22971_, _22972_, _22973_, _22974_, _22975_, _22976_, _22977_, _22978_, _22979_, _22980_, _22981_, _22982_, _22983_, _22984_, _22985_, _22986_, _22987_, _22988_, _22989_, _22990_, _22991_, _22992_, _22993_, _22994_, _22995_, _22996_, _22997_, _22998_, _22999_, _23000_, _23001_, _23002_, _23003_, _23004_, _23005_, _23006_, _23007_, _23008_, _23009_, _23010_, _23011_, _23012_, _23013_, _23014_, _23015_, _23016_, _23017_, _23018_, _23019_, _23020_, _23021_, _23022_, _23023_, _23024_, _23025_, _23026_, _23027_, _23028_, _23029_, _23030_, _23031_, _23032_, _23033_, _23034_, _23035_, _23036_, _23037_, _23038_, _23039_, _23040_, _23041_, _23042_, _23043_, _23044_, _23045_, _23046_, _23047_, _23048_, _23049_, _23050_, _23051_, _23052_, _23053_, _23054_, _23055_, _23056_, _23057_, _23058_, _23059_, _23060_, _23061_, _23062_, _23063_, _23064_, _23065_, _23066_, _23067_, _23068_, _23069_, _23070_, _23071_, _23072_, _23073_, _23074_, _23075_, _23076_, _23077_, _23078_, _23079_, _23080_, _23081_, _23082_, _23083_, _23084_, _23085_, _23086_, _23087_, _23088_, _23089_, _23090_, _23091_, _23092_, _23093_, _23094_, _23095_, _23096_, _23097_, _23098_, _23099_, _23100_, _23101_, _23102_, _23103_, _23104_, _23105_, _23106_, _23107_, _23108_, _23109_, _23110_, _23111_, _23112_, _23113_, _23114_, _23115_, _23116_, _23117_, _23118_, _23119_, _23120_, _23121_, _23122_, _23123_, _23124_, _23125_, _23126_, _23127_, _23128_, _23129_, _23130_, _23131_, _23132_, _23133_, _23134_, _23135_, _23136_, _23137_, _23138_, _23139_, _23140_, _23141_, _23142_, _23143_, _23144_, _23145_, _23146_, _23147_, _23148_, _23149_, _23150_, _23151_, _23152_, _23153_, _23154_, _23155_, _23156_, _23157_, _23158_, _23159_, _23160_, _23161_, _23162_, _23163_, _23164_, _23165_, _23166_, _23167_, _23168_, _23169_, _23170_, _23171_, _23172_, _23173_, _23174_, _23175_, _23176_, _23177_, _23178_, _23179_, _23180_, _23181_, _23182_, _23183_, _23184_, _23185_, _23186_, _23187_, _23188_, _23189_, _23190_, _23191_, _23192_, _23193_, _23194_, _23195_, _23196_, _23197_, _23198_, _23199_, _23200_, _23201_, _23202_, _23203_, _23204_, _23205_, _23206_, _23207_, _23208_, _23209_, _23210_, _23211_, _23212_, _23213_, _23214_, _23215_, _23216_, _23217_, _23218_, _23219_, _23220_, _23221_, _23222_, _23223_, _23224_, _23225_, _23226_, _23227_, _23228_, _23229_, _23230_, _23231_, _23232_, _23233_, _23234_, _23235_, _23236_, _23237_, _23238_, _23239_, _23240_, _23241_, _23242_, _23243_, _23244_, _23245_, _23246_, _23247_, _23248_, _23249_, _23250_, _23251_, _23252_, _23253_, _23254_, _23255_, _23256_, _23257_, _23258_, _23259_, _23260_, _23261_, _23262_, _23263_, _23264_, _23265_, _23266_, _23267_, _23268_, _23269_, _23270_, _23271_, _23272_, _23273_, _23274_, _23275_, _23276_, _23277_, _23278_, _23279_, _23280_, _23281_, _23282_, _23283_, _23284_, _23285_, _23286_, _23287_, _23288_, _23289_, _23290_, _23291_, _23292_, _23293_, _23294_, _23295_, _23296_, _23297_, _23298_, _23299_, _23300_, _23301_, _23302_, _23303_, _23304_, _23305_, _23306_, _23307_, _23308_, _23309_, _23310_, _23311_, _23312_, _23313_, _23314_, _23315_, _23316_, _23317_, _23318_, _23319_, _23320_, _23321_, _23322_, _23323_, _23324_, _23325_, _23326_, _23327_, _23328_, _23329_, _23330_, _23331_, _23332_, _23333_, _23334_, _23335_, _23336_, _23337_, _23338_, _23339_, _23340_, _23341_, _23342_, _23343_, _23344_, _23345_, _23346_, _23347_, _23348_, _23349_, _23350_, _23351_, _23352_, _23353_, _23354_, _23355_, _23356_, _23357_, _23358_, _23359_, _23360_, _23361_, _23362_, _23363_, _23364_, _23365_, _23366_, _23367_, _23368_, _23369_, _23370_, _23371_, _23372_, _23373_, _23374_, _23375_, _23376_, _23377_, _23378_, _23379_, _23380_, _23381_, _23382_, _23383_, _23384_, _23385_, _23386_, _23387_, _23388_, _23389_, _23390_, _23391_, _23392_, _23393_, _23394_, _23395_, _23396_, _23397_, _23398_, _23399_, _23400_, _23401_, _23402_, _23403_, _23404_, _23405_, _23406_, _23407_, _23408_, _23409_, _23410_, _23411_, _23412_, _23413_, _23414_, _23415_, _23416_, _23417_, _23418_, _23419_, _23420_, _23421_, _23422_, _23423_, _23424_, _23425_, _23426_, _23427_, _23428_, _23429_, _23430_, _23431_, _23432_, _23433_, _23434_, _23435_, _23436_, _23437_, _23438_, _23439_, _23440_, _23441_, _23442_, _23443_, _23444_, _23445_, _23446_, _23447_, _23448_, _23449_, _23450_, _23451_, _23452_, _23453_, _23454_, _23455_, _23456_, _23457_, _23458_, _23459_, _23460_, _23461_, _23462_, _23463_, _23464_, _23465_, _23466_, _23467_, _23468_, _23469_, _23470_, _23471_, _23472_, _23473_, _23474_, _23475_, _23476_, _23477_, _23478_, _23479_, _23480_, _23481_, _23482_, _23483_, _23484_, _23485_, _23486_, _23487_, _23488_, _23489_, _23490_, _23491_, _23492_, _23493_, _23494_, _23495_, _23496_, _23497_, _23498_, _23499_, _23500_, _23501_, _23502_, _23503_, _23504_, _23505_, _23506_, _23507_, _23508_, _23509_, _23510_, _23511_, _23512_, _23513_, _23514_, _23515_, _23516_, _23517_, _23518_, _23519_, _23520_, _23521_, _23522_, _23523_, _23524_, _23525_, _23526_, _23527_, _23528_, _23529_, _23530_, _23531_, _23532_, _23533_, _23534_, _23535_, _23536_, _23537_, _23538_, _23539_, _23540_, _23541_, _23542_, _23543_, _23544_, _23545_, _23546_, _23547_, _23548_, _23549_, _23550_, _23551_, _23552_, _23553_, _23554_, _23555_, _23556_, _23557_, _23558_, _23559_, _23560_, _23561_, _23562_, _23563_, _23564_, _23565_, _23566_, _23567_, _23568_, _23569_, _23570_, _23571_, _23572_, _23573_, _23574_, _23575_, _23576_, _23577_, _23578_, _23579_, _23580_, _23581_, _23582_, _23583_, _23584_, _23585_, _23586_, _23587_, _23588_, _23589_, _23590_, _23591_, _23592_, _23593_, _23594_, _23595_, _23596_, _23597_, _23598_, _23599_, _23600_, _23601_, _23602_, _23603_, _23604_, _23605_, _23606_, _23607_, _23608_, _23609_, _23610_, _23611_, _23612_, _23613_, _23614_, _23615_, _23616_, _23617_, _23618_, _23619_, _23620_, _23621_, _23622_, _23623_, _23624_, _23625_, _23626_, _23627_, _23628_, _23629_, _23630_, _23631_, _23632_, _23633_, _23634_, _23635_, _23636_, _23637_, _23638_, _23639_, _23640_, _23641_, _23642_, _23643_, _23644_, _23645_, _23646_, _23647_, _23648_, _23649_, _23650_, _23651_, _23652_, _23653_, _23654_, _23655_, _23656_, _23657_, _23658_, _23659_, _23660_, _23661_, _23662_, _23663_, _23664_, _23665_, _23666_, _23667_, _23668_, _23669_, _23670_, _23671_, _23672_, _23673_, _23674_, _23675_, _23676_, _23677_, _23678_, _23679_, _23680_, _23681_, _23682_, _23683_, _23684_, _23685_, _23686_, _23687_, _23688_, _23689_, _23690_, _23691_, _23692_, _23693_, _23694_, _23695_, _23696_, _23697_, _23698_, _23699_, _23700_, _23701_, _23702_, _23703_, _23704_, _23705_, _23706_, _23707_, _23708_, _23709_, _23710_, _23711_, _23712_, _23713_, _23714_, _23715_, _23716_, _23717_, _23718_, _23719_, _23720_, _23721_, _23722_, _23723_, _23724_, _23725_, _23726_, _23727_, _23728_, _23729_, _23730_, _23731_, _23732_, _23733_, _23734_, _23735_, _23736_, _23737_, _23738_, _23739_, _23740_, _23741_, _23742_, _23743_, _23744_, _23745_, _23746_, _23747_, _23748_, _23749_, _23750_, _23751_, _23752_, _23753_, _23754_, _23755_, _23756_, _23757_, _23758_, _23759_, _23760_, _23761_, _23762_, _23763_, _23764_, _23765_, _23766_, _23767_, _23768_, _23769_, _23770_, _23771_, _23772_, _23773_, _23774_, _23775_, _23776_, _23777_, _23778_, _23779_, _23780_, _23781_, _23782_, _23783_, _23784_, _23785_, _23786_, _23787_, _23788_, _23789_, _23790_, _23791_, _23792_, _23793_, _23794_, _23795_, _23796_, _23797_, _23798_, _23799_, _23800_, _23801_, _23802_, _23803_, _23804_, _23805_, _23806_, _23807_, _23808_, _23809_, _23810_, _23811_, _23812_, _23813_, _23814_, _23815_, _23816_, _23817_, _23818_, _23819_, _23820_, _23821_, _23822_, _23823_, _23824_, _23825_, _23826_, _23827_, _23828_, _23829_, _23830_, _23831_, _23832_, _23833_, _23834_, _23835_, _23836_, _23837_, _23838_, _23839_, _23840_, _23841_, _23842_, _23843_, _23844_, _23845_, _23846_, _23847_, _23848_, _23849_, _23850_, _23851_, _23852_, _23853_, _23854_, _23855_, _23856_, _23857_, _23858_, _23859_, _23860_, _23861_, _23862_, _23863_, _23864_, _23865_, _23866_, _23867_, _23868_, _23869_, _23870_, _23871_, _23872_, _23873_, _23874_, _23875_, _23876_, _23877_, _23878_, _23879_, _23880_, _23881_, _23882_, _23883_, _23884_, _23885_, _23886_, _23887_, _23888_, _23889_, _23890_, _23891_, _23892_, _23893_, _23894_, _23895_, _23896_, _23897_, _23898_, _23899_, _23900_, _23901_, _23902_, _23903_, _23904_, _23905_, _23906_, _23907_, _23908_, _23909_, _23910_, _23911_, _23912_, _23913_, _23914_, _23915_, _23916_, _23917_, _23918_, _23919_, _23920_, _23921_, _23922_, _23923_, _23924_, _23925_, _23926_, _23927_, _23928_, _23929_, _23930_, _23931_, _23932_, _23933_, _23934_, _23935_, _23936_, _23937_, _23938_, _23939_, _23940_, _23941_, _23942_, _23943_, _23944_, _23945_, _23946_, _23947_, _23948_, _23949_, _23950_, _23951_, _23952_, _23953_, _23954_, _23955_, _23956_, _23957_, _23958_, _23959_, _23960_, _23961_, _23962_, _23963_, _23964_, _23965_, _23966_, _23967_, _23968_, _23969_, _23970_, _23971_, _23972_, _23973_, _23974_, _23975_, _23976_, _23977_, _23978_, _23979_, _23980_, _23981_, _23982_, _23983_, _23984_, _23985_, _23986_, _23987_, _23988_, _23989_, _23990_, _23991_, _23992_, _23993_, _23994_, _23995_, _23996_, _23997_, _23998_, _23999_, _24000_, _24001_, _24002_, _24003_, _24004_, _24005_, _24006_, _24007_, _24008_, _24009_, _24010_, _24011_, _24012_, _24013_, _24014_, _24015_, _24016_, _24017_, _24018_, _24019_, _24020_, _24021_, _24022_, _24023_, _24024_, _24025_, _24026_, _24027_, _24028_, _24029_, _24030_, _24031_, _24032_, _24033_, _24034_, _24035_, _24036_, _24037_, _24038_, _24039_, _24040_, _24041_, _24042_, _24043_, _24044_, _24045_, _24046_, _24047_, _24048_, _24049_, _24050_, _24051_, _24052_, _24053_, _24054_, _24055_, _24056_, _24057_, _24058_, _24059_, _24060_, _24061_, _24062_, _24063_, _24064_, _24065_, _24066_, _24067_, _24068_, _24069_, _24070_, _24071_, _24072_, _24073_, _24074_, _24075_, _24076_, _24077_, _24078_, _24079_, _24080_, _24081_, _24082_, _24083_, _24084_, _24085_, _24086_, _24087_, _24088_, _24089_, _24090_, _24091_, _24092_, _24093_, _24094_, _24095_, _24096_, _24097_, _24098_, _24099_, _24100_, _24101_, _24102_, _24103_, _24104_, _24105_, _24106_, _24107_, _24108_, _24109_, _24110_, _24111_, _24112_, _24113_, _24114_, _24115_, _24116_, _24117_, _24118_, _24119_, _24120_, _24121_, _24122_, _24123_, _24124_, _24125_, _24126_, _24127_, _24128_, _24129_, _24130_, _24131_, _24132_, _24133_, _24134_, _24135_, _24136_, _24137_, _24138_, _24139_, _24140_, _24141_, _24142_, _24143_, _24144_, _24145_, _24146_, _24147_, _24148_, _24149_, _24150_, _24151_, _24152_, _24153_, _24154_, _24155_, _24156_, _24157_, _24158_, _24159_, _24160_, _24161_, _24162_, _24163_, _24164_, _24165_, _24166_, _24167_, _24168_, _24169_, _24170_, _24171_, _24172_, _24173_, _24174_, _24175_, _24176_, _24177_, _24178_, _24179_, _24180_, _24181_, _24182_, _24183_, _24184_, _24185_, _24186_, _24187_, _24188_, _24189_, _24190_, _24191_, _24192_, _24193_, _24194_, _24195_, _24196_, _24197_, _24198_, _24199_, _24200_, _24201_, _24202_, _24203_, _24204_, _24205_, _24206_, _24207_, _24208_, _24209_, _24210_, _24211_, _24212_, _24213_, _24214_, _24215_, _24216_, _24217_, _24218_, _24219_, _24220_, _24221_, _24222_, _24223_, _24224_, _24225_, _24226_, _24227_, _24228_, _24229_, _24230_, _24231_, _24232_, _24233_, _24234_, _24235_, _24236_, _24237_, _24238_, _24239_, _24240_, _24241_, _24242_, _24243_, _24244_, _24245_, _24246_, _24247_, _24248_, _24249_, _24250_, _24251_, _24252_, _24253_, _24254_, _24255_, _24256_, _24257_, _24258_, _24259_, _24260_, _24261_, _24262_, _24263_, _24264_, _24265_, _24266_, _24267_, _24268_, _24269_, _24270_, _24271_, _24272_, _24273_, _24274_, _24275_, _24276_, _24277_, _24278_, _24279_, _24280_, _24281_, _24282_, _24283_, _24284_, _24285_, _24286_, _24287_, _24288_, _24289_, _24290_, _24291_, _24292_, _24293_, _24294_, _24295_, _24296_, _24297_, _24298_, _24299_, _24300_, _24301_, _24302_, _24303_, _24304_, _24305_, _24306_, _24307_, _24308_, _24309_, _24310_, _24311_, _24312_, _24313_, _24314_, _24315_, _24316_, _24317_, _24318_, _24319_, _24320_, _24321_, _24322_, _24323_, _24324_, _24325_, _24326_, _24327_, _24328_, _24329_, _24330_, _24331_, _24332_, _24333_, _24334_, _24335_, _24336_, _24337_, _24338_, _24339_, _24340_, _24341_, _24342_, _24343_, _24344_, _24345_, _24346_, _24347_, _24348_, _24349_, _24350_, _24351_, _24352_, _24353_, _24354_, _24355_, _24356_, _24357_, _24358_, _24359_, _24360_, _24361_, _24362_, _24363_, _24364_, _24365_, _24366_, _24367_, _24368_, _24369_, _24370_, _24371_, _24372_, _24373_, _24374_, _24375_, _24376_, _24377_, _24378_, _24379_, _24380_, _24381_, _24382_, _24383_, _24384_, _24385_, _24386_, _24387_, _24388_, _24389_, _24390_, _24391_, _24392_, _24393_, _24394_, _24395_, _24396_, _24397_, _24398_, _24399_, _24400_, _24401_, _24402_, _24403_, _24404_, _24405_, _24406_, _24407_, _24408_, _24409_, _24410_, _24411_, _24412_, _24413_, _24414_, _24415_, _24416_, _24417_, _24418_, _24419_, _24420_, _24421_, _24422_, _24423_, _24424_, _24425_, _24426_, _24427_, _24428_, _24429_, _24430_, _24431_, _24432_, _24433_, _24434_, _24435_, _24436_, _24437_, _24438_, _24439_, _24440_, _24441_, _24442_, _24443_, _24444_, _24445_, _24446_, _24447_, _24448_, _24449_, _24450_, _24451_, _24452_, _24453_, _24454_, _24455_, _24456_, _24457_, _24458_, _24459_, _24460_, _24461_, _24462_, _24463_, _24464_, _24465_, _24466_, _24467_, _24468_, _24469_, _24470_, _24471_, _24472_, _24473_, _24474_, _24475_, _24476_, _24477_, _24478_, _24479_, _24480_, _24481_, _24482_, _24483_, _24484_, _24485_, _24486_, _24487_, _24488_, _24489_, _24490_, _24491_, _24492_, _24493_, _24494_, _24495_, _24496_, _24497_, _24498_, _24499_, _24500_, _24501_, _24502_, _24503_, _24504_, _24505_, _24506_, _24507_, _24508_, _24509_, _24510_, _24511_, _24512_, _24513_, _24514_, _24515_, _24516_, _24517_, _24518_, _24519_, _24520_, _24521_, _24522_, _24523_, _24524_, _24525_, _24526_, _24527_, _24528_, _24529_, _24530_, _24531_, _24532_, _24533_, _24534_, _24535_, _24536_, _24537_, _24538_, _24539_, _24540_, _24541_, _24542_, _24543_, _24544_, _24545_, _24546_, _24547_, _24548_, _24549_, _24550_, _24551_, _24552_, _24553_, _24554_, _24555_, _24556_, _24557_, _24558_, _24559_, _24560_, _24561_, _24562_, _24563_, _24564_, _24565_, _24566_, _24567_, _24568_, _24569_, _24570_, _24571_, _24572_, _24573_, _24574_, _24575_, _24576_, _24577_, _24578_, _24579_, _24580_, _24581_, _24582_, _24583_, _24584_, _24585_, _24586_, _24587_, _24588_, _24589_, _24590_, _24591_, _24592_, _24593_, _24594_, _24595_, _24596_, _24597_, _24598_, _24599_, _24600_, _24601_, _24602_, _24603_, _24604_, _24605_, _24606_, _24607_, _24608_, _24609_, _24610_, _24611_, _24612_, _24613_, _24614_, _24615_, _24616_, _24617_, _24618_, _24619_, _24620_, _24621_, _24622_, _24623_, _24624_, _24625_, _24626_, _24627_, _24628_, _24629_, _24630_, _24631_, _24632_, _24633_, _24634_, _24635_, _24636_, _24637_, _24638_, _24639_, _24640_, _24641_, _24642_, _24643_, _24644_, _24645_, _24646_, _24647_, _24648_, _24649_, _24650_, _24651_, _24652_, _24653_, _24654_, _24655_, _24656_, _24657_, _24658_, _24659_, _24660_, _24661_, _24662_, _24663_, _24664_, _24665_, _24666_, _24667_, _24668_, _24669_, _24670_, _24671_, _24672_, _24673_, _24674_, _24675_, _24676_, _24677_, _24678_, _24679_, _24680_, _24681_, _24682_, _24683_, _24684_, _24685_, _24686_, _24687_, _24688_, _24689_, _24690_, _24691_, _24692_, _24693_, _24694_, _24695_, _24696_, _24697_, _24698_, _24699_, _24700_, _24701_, _24702_, _24703_, _24704_, _24705_, _24706_, _24707_, _24708_, _24709_, _24710_, _24711_, _24712_, _24713_, _24714_, _24715_, _24716_, _24717_, _24718_, _24719_, _24720_, _24721_, _24722_, _24723_, _24724_, _24725_, _24726_, _24727_, _24728_, _24729_, _24730_, _24731_, _24732_, _24733_, _24734_, _24735_, _24736_, _24737_, _24738_, _24739_, _24740_, _24741_, _24742_, _24743_, _24744_, _24745_, _24746_, _24747_, _24748_, _24749_, _24750_, _24751_, _24752_, _24753_, _24754_, _24755_, _24756_, _24757_, _24758_, _24759_, _24760_, _24761_, _24762_, _24763_, _24764_, _24765_, _24766_, _24767_, _24768_, _24769_, _24770_, _24771_, _24772_, _24773_, _24774_, _24775_, _24776_, _24777_, _24778_, _24779_, _24780_, _24781_, _24782_, _24783_, _24784_, _24785_, _24786_, _24787_, _24788_, _24789_, _24790_, _24791_, _24792_, _24793_, _24794_, _24795_, _24796_, _24797_, _24798_, _24799_, _24800_, _24801_, _24802_, _24803_, _24804_, _24805_, _24806_, _24807_, _24808_, _24809_, _24810_, _24811_, _24812_, _24813_, _24814_, _24815_, _24816_, _24817_, _24818_, _24819_, _24820_, _24821_, _24822_, _24823_, _24824_, _24825_, _24826_, _24827_, _24828_, _24829_, _24830_, _24831_, _24832_, _24833_, _24834_, _24835_, _24836_, _24837_, _24838_, _24839_, _24840_, _24841_, _24842_, _24843_, _24844_, _24845_, _24846_, _24847_, _24848_, _24849_, _24850_, _24851_, _24852_, _24853_, _24854_, _24855_, _24856_, _24857_, _24858_, _24859_, _24860_, _24861_, _24862_, _24863_, _24864_, _24865_, _24866_, _24867_, _24868_, _24869_, _24870_, _24871_, _24872_, _24873_, _24874_, _24875_, _24876_, _24877_, _24878_, _24879_, _24880_, _24881_, _24882_, _24883_, _24884_, _24885_, _24886_, _24887_, _24888_, _24889_, _24890_, _24891_, _24892_, _24893_, _24894_, _24895_, _24896_, _24897_, _24898_, _24899_, _24900_, _24901_, _24902_, _24903_, _24904_, _24905_, _24906_, _24907_, _24908_, _24909_, _24910_, _24911_, _24912_, _24913_, _24914_, _24915_, _24916_, _24917_, _24918_, _24919_, _24920_, _24921_, _24922_, _24923_, _24924_, _24925_, _24926_, _24927_, _24928_, _24929_, _24930_, _24931_, _24932_, _24933_, _24934_, _24935_, _24936_, _24937_, _24938_, _24939_, _24940_, _24941_, _24942_, _24943_, _24944_, _24945_, _24946_, _24947_, _24948_, _24949_, _24950_, _24951_, _24952_, _24953_, _24954_, _24955_, _24956_, _24957_, _24958_, _24959_, _24960_, _24961_, _24962_, _24963_, _24964_, _24965_, _24966_, _24967_, _24968_, _24969_, _24970_, _24971_, _24972_, _24973_, _24974_, _24975_, _24976_, _24977_, _24978_, _24979_, _24980_, _24981_, _24982_, _24983_, _24984_, _24985_, _24986_, _24987_, _24988_, _24989_, _24990_, _24991_, _24992_, _24993_, _24994_, _24995_, _24996_, _24997_, _24998_, _24999_, _25000_, _25001_, _25002_, _25003_, _25004_, _25005_, _25006_, _25007_, _25008_, _25009_, _25010_, _25011_, _25012_, _25013_, _25014_, _25015_, _25016_, _25017_, _25018_, _25019_, _25020_, _25021_, _25022_, _25023_, _25024_, _25025_, _25026_, _25027_, _25028_, _25029_, _25030_, _25031_, _25032_, _25033_, _25034_, _25035_, _25036_, _25037_, _25038_, _25039_, _25040_, _25041_, _25042_, _25043_, _25044_, _25045_, _25046_, _25047_, _25048_, _25049_, _25050_, _25051_, _25052_, _25053_, _25054_, _25055_, _25056_, _25057_, _25058_, _25059_, _25060_, _25061_, _25062_, _25063_, _25064_, _25065_, _25066_, _25067_, _25068_, _25069_, _25070_, _25071_, _25072_, _25073_, _25074_, _25075_, _25076_, _25077_, _25078_, _25079_, _25080_, _25081_, _25082_, _25083_, _25084_, _25085_, _25086_, _25087_, _25088_, _25089_, _25090_, _25091_, _25092_, _25093_, _25094_, _25095_, _25096_, _25097_, _25098_, _25099_, _25100_, _25101_, _25102_, _25103_, _25104_, _25105_, _25106_, _25107_, _25108_, _25109_, _25110_, _25111_, _25112_, _25113_, _25114_, _25115_, _25116_, _25117_, _25118_, _25119_, _25120_, _25121_, _25122_, _25123_, _25124_, _25125_, _25126_, _25127_, _25128_, _25129_, _25130_, _25131_, _25132_, _25133_, _25134_, _25135_, _25136_, _25137_, _25138_, _25139_, _25140_, _25141_, _25142_, _25143_, _25144_, _25145_, _25146_, _25147_, _25148_, _25149_, _25150_, _25151_, _25152_, _25153_, _25154_, _25155_, _25156_, _25157_, _25158_, _25159_, _25160_, _25161_, _25162_, _25163_, _25164_, _25165_, _25166_, _25167_, _25168_, _25169_, _25170_, _25171_, _25172_, _25173_, _25174_, _25175_, _25176_, _25177_, _25178_, _25179_, _25180_, _25181_, _25182_, _25183_, _25184_, _25185_, _25186_, _25187_, _25188_, _25189_, _25190_, _25191_, _25192_, _25193_, _25194_, _25195_, _25196_, _25197_, _25198_, _25199_, _25200_, _25201_, _25202_, _25203_, _25204_, _25205_, _25206_, _25207_, _25208_, _25209_, _25210_, _25211_, _25212_, _25213_, _25214_, _25215_, _25216_, _25217_, _25218_, _25219_, _25220_, _25221_, _25222_, _25223_, _25224_, _25225_, _25226_, _25227_, _25228_, _25229_, _25230_, _25231_, _25232_, _25233_, _25234_, _25235_, _25236_, _25237_, _25238_, _25239_, _25240_, _25241_, _25242_, _25243_, _25244_, _25245_, _25246_, _25247_, _25248_, _25249_, _25250_, _25251_, _25252_, _25253_, _25254_, _25255_, _25256_, _25257_, _25258_, _25259_, _25260_, _25261_, _25262_, _25263_, _25264_, _25265_, _25266_, _25267_, _25268_, _25269_, _25270_, _25271_, _25272_, _25273_, _25274_, _25275_, _25276_, _25277_, _25278_, _25279_, _25280_, _25281_, _25282_, _25283_, _25284_, _25285_, _25286_, _25287_, _25288_, _25289_, _25290_, _25291_, _25292_, _25293_, _25294_, _25295_, _25296_, _25297_, _25298_, _25299_, _25300_, _25301_, _25302_, _25303_, _25304_, _25305_, _25306_, _25307_, _25308_, _25309_, _25310_, _25311_, _25312_, _25313_, _25314_, _25315_, _25316_, _25317_, _25318_, _25319_, _25320_, _25321_, _25322_, _25323_, _25324_, _25325_, _25326_, _25327_, _25328_, _25329_, _25330_, _25331_, _25332_, _25333_, _25334_, _25335_, _25336_, _25337_, _25338_, _25339_, _25340_, _25341_, _25342_, _25343_, _25344_, _25345_, _25346_, _25347_, _25348_, _25349_, _25350_, _25351_, _25352_, _25353_, _25354_, _25355_, _25356_, _25357_, _25358_, _25359_, _25360_, _25361_, _25362_, _25363_, _25364_, _25365_, _25366_, _25367_, _25368_, _25369_, _25370_, _25371_, _25372_, _25373_, _25374_, _25375_, _25376_, _25377_, _25378_, _25379_, _25380_, _25381_, _25382_, _25383_, _25384_, _25385_, _25386_, _25387_, _25388_, _25389_, _25390_, _25391_, _25392_, _25393_, _25394_, _25395_, _25396_, _25397_, _25398_, _25399_, _25400_, _25401_, _25402_, _25403_, _25404_, _25405_, _25406_, _25407_, _25408_, _25409_, _25410_, _25411_, _25412_, _25413_, _25414_, _25415_, _25416_, _25417_, _25418_, _25419_, _25420_, _25421_, _25422_, _25423_, _25424_, _25425_, _25426_, _25427_, _25428_, _25429_, _25430_, _25431_, _25432_, _25433_, _25434_, _25435_, _25436_, _25437_, _25438_, _25439_, _25440_, _25441_, _25442_, _25443_, _25444_, _25445_, _25446_, _25447_, _25448_, _25449_, _25450_, _25451_, _25452_, _25453_, _25454_, _25455_, _25456_, _25457_, _25458_, _25459_, _25460_, _25461_, _25462_, _25463_, _25464_, _25465_, _25466_, _25467_, _25468_, _25469_, _25470_, _25471_, _25472_, _25473_, _25474_, _25475_, _25476_, _25477_, _25478_, _25479_, _25480_, _25481_, _25482_, _25483_, _25484_, _25485_, _25486_, _25487_, _25488_, _25489_, _25490_, _25491_, _25492_, _25493_, _25494_, _25495_, _25496_, _25497_, _25498_, _25499_, _25500_, _25501_, _25502_, _25503_, _25504_, _25505_, _25506_, _25507_, _25508_, _25509_, _25510_, _25511_, _25512_, _25513_, _25514_, _25515_, _25516_, _25517_, _25518_, _25519_, _25520_, _25521_, _25522_, _25523_, _25524_, _25525_, _25526_, _25527_, _25528_, _25529_, _25530_, _25531_, _25532_, _25533_, _25534_, _25535_, _25536_, _25537_, _25538_, _25539_, _25540_, _25541_, _25542_, _25543_, _25544_, _25545_, _25546_, _25547_, _25548_, _25549_, _25550_, _25551_, _25552_, _25553_, _25554_, _25555_, _25556_, _25557_, _25558_, _25559_, _25560_, _25561_, _25562_, _25563_, _25564_, _25565_, _25566_, _25567_, _25568_, _25569_, _25570_, _25571_, _25572_, _25573_, _25574_, _25575_, _25576_, _25577_, _25578_, _25579_, _25580_, _25581_, _25582_, _25583_, _25584_, _25585_, _25586_, _25587_, _25588_, _25589_, _25590_, _25591_, _25592_, _25593_, _25594_, _25595_, _25596_, _25597_, _25598_, _25599_, _25600_, _25601_, _25602_, _25603_, _25604_, _25605_, _25606_, _25607_, _25608_, _25609_, _25610_, _25611_, _25612_, _25613_, _25614_, _25615_, _25616_, _25617_, _25618_, _25619_, _25620_, _25621_, _25622_, _25623_, _25624_, _25625_, _25626_, _25627_, _25628_, _25629_, _25630_, _25631_, _25632_, _25633_, _25634_, _25635_, _25636_, _25637_, _25638_, _25639_, _25640_, _25641_, _25642_, _25643_, _25644_, _25645_, _25646_, _25647_, _25648_, _25649_, _25650_, _25651_, _25652_, _25653_, _25654_, _25655_, _25656_, _25657_, _25658_, _25659_, _25660_, _25661_, _25662_, _25663_, _25664_, _25665_, _25666_, _25667_, _25668_, _25669_, _25670_, _25671_, _25672_, _25673_, _25674_, _25675_, _25676_, _25677_, _25678_, _25679_, _25680_, _25681_, _25682_, _25683_, _25684_, _25685_, _25686_, _25687_, _25688_, _25689_, _25690_, _25691_, _25692_, _25693_, _25694_, _25695_, _25696_, _25697_, _25698_, _25699_, _25700_, _25701_, _25702_, _25703_, _25704_, _25705_, _25706_, _25707_, _25708_, _25709_, _25710_, _25711_, _25712_, _25713_, _25714_, _25715_, _25716_, _25717_, _25718_, _25719_, _25720_, _25721_, _25722_, _25723_, _25724_, _25725_, _25726_, _25727_, _25728_, _25729_, _25730_, _25731_, _25732_, _25733_, _25734_, _25735_, _25736_, _25737_, _25738_, _25739_, _25740_, _25741_, _25742_, _25743_, _25744_, _25745_, _25746_, _25747_, _25748_, _25749_, _25750_, _25751_, _25752_, _25753_, _25754_, _25755_, _25756_, _25757_, _25758_, _25759_, _25760_, _25761_, _25762_, _25763_, _25764_, _25765_, _25766_, _25767_, _25768_, _25769_, _25770_, _25771_, _25772_, _25773_, _25774_, _25775_, _25776_, _25777_, _25778_, _25779_, _25780_, _25781_, _25782_, _25783_, _25784_, _25785_, _25786_, _25787_, _25788_, _25789_, _25790_, _25791_, _25792_, _25793_, _25794_, _25795_, _25796_, _25797_, _25798_, _25799_, _25800_, _25801_, _25802_, _25803_, _25804_, _25805_, _25806_, _25807_, _25808_, _25809_, _25810_, _25811_, _25812_, _25813_, _25814_, _25815_, _25816_, _25817_, _25818_, _25819_, _25820_, _25821_, _25822_, _25823_, _25824_, _25825_, _25826_, _25827_, _25828_, _25829_, _25830_, _25831_, _25832_, _25833_, _25834_, _25835_, _25836_, _25837_, _25838_, _25839_, _25840_, _25841_, _25842_, _25843_, _25844_, _25845_, _25846_, _25847_, _25848_, _25849_, _25850_, _25851_, _25852_, _25853_, _25854_, _25855_, _25856_, _25857_, _25858_, _25859_, _25860_, _25861_, _25862_, _25863_, _25864_, _25865_, _25866_, _25867_, _25868_, _25869_, _25870_, _25871_, _25872_, _25873_, _25874_, _25875_, _25876_, _25877_, _25878_, _25879_, _25880_, _25881_, _25882_, _25883_, _25884_, _25885_, _25886_, _25887_, _25888_, _25889_, _25890_, _25891_, _25892_, _25893_, _25894_, _25895_, _25896_, _25897_, _25898_, _25899_, _25900_, _25901_, _25902_, _25903_, _25904_, _25905_, _25906_, _25907_, _25908_, _25909_, _25910_, _25911_, _25912_, _25913_, _25914_, _25915_, _25916_, _25917_, _25918_, _25919_, _25920_, _25921_, _25922_, _25923_, _25924_, _25925_, _25926_, _25927_, _25928_, _25929_, _25930_, _25931_, _25932_, _25933_, _25934_, _25935_, _25936_, _25937_, _25938_, _25939_, _25940_, _25941_, _25942_, _25943_, _25944_, _25945_, _25946_, _25947_, _25948_, _25949_, _25950_, _25951_, _25952_, _25953_, _25954_, _25955_, _25956_, _25957_, _25958_, _25959_, _25960_, _25961_, _25962_, _25963_, _25964_, _25965_, _25966_, _25967_, _25968_, _25969_, _25970_, _25971_, _25972_, _25973_, _25974_, _25975_, _25976_, _25977_, _25978_, _25979_, _25980_, _25981_, _25982_, _25983_, _25984_, _25985_, _25986_, _25987_, _25988_, _25989_, _25990_, _25991_, _25992_, _25993_, _25994_, _25995_, _25996_, _25997_, _25998_, _25999_, _26000_, _26001_, _26002_, _26003_, _26004_, _26005_, _26006_, _26007_, _26008_, _26009_, _26010_, _26011_, _26012_, _26013_, _26014_, _26015_, _26016_, _26017_, _26018_, _26019_, _26020_, _26021_, _26022_, _26023_, _26024_, _26025_, _26026_, _26027_, _26028_, _26029_, _26030_, _26031_, _26032_, _26033_, _26034_, _26035_, _26036_, _26037_, _26038_, _26039_, _26040_, _26041_, _26042_, _26043_, _26044_, _26045_, _26046_, _26047_, _26048_, _26049_, _26050_, _26051_, _26052_, _26053_, _26054_, _26055_, _26056_, _26057_, _26058_, _26059_, _26060_, _26061_, _26062_, _26063_, _26064_, _26065_, _26066_, _26067_, _26068_, _26069_, _26070_, _26071_, _26072_, _26073_, _26074_, _26075_, _26076_, _26077_, _26078_, _26079_, _26080_, _26081_, _26082_, _26083_, _26084_, _26085_, _26086_, _26087_, _26088_, _26089_, _26090_, _26091_, _26092_, _26093_, _26094_, _26095_, _26096_, _26097_, _26098_, _26099_, _26100_, _26101_, _26102_, _26103_, _26104_, _26105_, _26106_, _26107_, _26108_, _26109_, _26110_, _26111_, _26112_, _26113_, _26114_, _26115_, _26116_, _26117_, _26118_, _26119_, _26120_, _26121_, _26122_, _26123_, _26124_, _26125_, _26126_, _26127_, _26128_, _26129_, _26130_, _26131_, _26132_, _26133_, _26134_, _26135_, _26136_, _26137_, _26138_, _26139_, _26140_, _26141_, _26142_, _26143_, _26144_, _26145_, _26146_, _26147_, _26148_, _26149_, _26150_, _26151_, _26152_, _26153_, _26154_, _26155_, _26156_, _26157_, _26158_, _26159_, _26160_, _26161_, _26162_, _26163_, _26164_, _26165_, _26166_, _26167_, _26168_, _26169_, _26170_, _26171_, _26172_, _26173_, _26174_, _26175_, _26176_, _26177_, _26178_, _26179_, _26180_, _26181_, _26182_, _26183_, _26184_, _26185_, _26186_, _26187_, _26188_, _26189_, _26190_, _26191_, _26192_, _26193_, _26194_, _26195_, _26196_, _26197_, _26198_, _26199_, _26200_, _26201_, _26202_, _26203_, _26204_, _26205_, _26206_, _26207_, _26208_, _26209_, _26210_, _26211_, _26212_, _26213_, _26214_, _26215_, _26216_, _26217_, _26218_, _26219_, _26220_, _26221_, _26222_, _26223_, _26224_, _26225_, _26226_, _26227_, _26228_, _26229_, _26230_, _26231_, _26232_, _26233_, _26234_, _26235_, _26236_, _26237_, _26238_, _26239_, _26240_, _26241_, _26242_, _26243_, _26244_, _26245_, _26246_, _26247_, _26248_, _26249_, _26250_, _26251_, _26252_, _26253_, _26254_, _26255_, _26256_, _26257_, _26258_, _26259_, _26260_, _26261_, _26262_, _26263_, _26264_, _26265_, _26266_, _26267_, _26268_, _26269_, _26270_, _26271_, _26272_, _26273_, _26274_, _26275_, _26276_, _26277_, _26278_, _26279_, _26280_, _26281_, _26282_, _26283_, _26284_, _26285_, _26286_, _26287_, _26288_, _26289_, _26290_, _26291_, _26292_, _26293_, _26294_, _26295_, _26296_, _26297_, _26298_, _26299_, _26300_, _26301_, _26302_, _26303_, _26304_, _26305_, _26306_, _26307_, _26308_, _26309_, _26310_, _26311_, _26312_, _26313_, _26314_, _26315_, _26316_, _26317_, _26318_, _26319_, _26320_, _26321_, _26322_, _26323_, _26324_, _26325_, _26326_, _26327_, _26328_, _26329_, _26330_, _26331_, _26332_, _26333_, _26334_, _26335_, _26336_, _26337_, _26338_, _26339_, _26340_, _26341_, _26342_, _26343_, _26344_, _26345_, _26346_, _26347_, _26348_, _26349_, _26350_, _26351_, _26352_, _26353_, _26354_, _26355_, _26356_, _26357_, _26358_, _26359_, _26360_, _26361_, _26362_, _26363_, _26364_, _26365_, _26366_, _26367_, _26368_, _26369_, _26370_, _26371_, _26372_, _26373_, _26374_, _26375_, _26376_, _26377_, _26378_, _26379_, _26380_, _26381_, _26382_, _26383_, _26384_, _26385_, _26386_, _26387_, _26388_, _26389_, _26390_, _26391_, _26392_, _26393_, _26394_, _26395_, _26396_, _26397_, _26398_, _26399_, _26400_, _26401_, _26402_, _26403_, _26404_, _26405_, _26406_, _26407_, _26408_, _26409_, _26410_, _26411_, _26412_, _26413_, _26414_, _26415_, _26416_, _26417_, _26418_, _26419_, _26420_, _26421_, _26422_, _26423_, _26424_, _26425_, _26426_, _26427_, _26428_, _26429_, _26430_, _26431_, _26432_, _26433_, _26434_, _26435_, _26436_, _26437_, _26438_, _26439_, _26440_, _26441_, _26442_, _26443_, _26444_, _26445_, _26446_, _26447_, _26448_, _26449_, _26450_, _26451_, _26452_, _26453_, _26454_, _26455_, _26456_, _26457_, _26458_, _26459_, _26460_, _26461_, _26462_, _26463_, _26464_, _26465_, _26466_, _26467_, _26468_, _26469_, _26470_, _26471_, _26472_, _26473_, _26474_, _26475_, _26476_, _26477_, _26478_, _26479_, _26480_, _26481_, _26482_, _26483_, _26484_, _26485_, _26486_, _26487_, _26488_, _26489_, _26490_, _26491_, _26492_, _26493_, _26494_, _26495_, _26496_, _26497_, _26498_, _26499_, _26500_, _26501_, _26502_, _26503_, _26504_, _26505_, _26506_, _26507_, _26508_, _26509_, _26510_, _26511_, _26512_, _26513_, _26514_, _26515_, _26516_, _26517_, _26518_, _26519_, _26520_, _26521_, _26522_, _26523_, _26524_, _26525_, _26526_, _26527_, _26528_, _26529_, _26530_, _26531_, _26532_, _26533_, _26534_, _26535_, _26536_, _26537_, _26538_, _26539_, _26540_, _26541_, _26542_, _26543_, _26544_, _26545_, _26546_, _26547_, _26548_, _26549_, _26550_, _26551_, _26552_, _26553_, _26554_, _26555_, _26556_, _26557_, _26558_, _26559_, _26560_, _26561_, _26562_, _26563_, _26564_, _26565_, _26566_, _26567_, _26568_, _26569_, _26570_, _26571_, _26572_, _26573_, _26574_, _26575_, _26576_, _26577_, _26578_, _26579_, _26580_, _26581_, _26582_, _26583_, _26584_, _26585_, _26586_, _26587_, _26588_, _26589_, _26590_, _26591_, _26592_, _26593_, _26594_, _26595_, _26596_, _26597_, _26598_, _26599_, _26600_, _26601_, _26602_, _26603_, _26604_, _26605_, _26606_, _26607_, _26608_, _26609_, _26610_, _26611_, _26612_, _26613_, _26614_, _26615_, _26616_, _26617_, _26618_, _26619_, _26620_, _26621_, _26622_, _26623_, _26624_, _26625_, _26626_, _26627_, _26628_, _26629_, _26630_, _26631_, _26632_, _26633_, _26634_, _26635_, _26636_, _26637_, _26638_, _26639_, _26640_, _26641_, _26642_, _26643_, _26644_, _26645_, _26646_, _26647_, _26648_, _26649_, _26650_, _26651_, _26652_, _26653_, _26654_, _26655_, _26656_, _26657_, _26658_, _26659_, _26660_, _26661_, _26662_, _26663_, _26664_, _26665_, _26666_, _26667_, _26668_, _26669_, _26670_, _26671_, _26672_, _26673_, _26674_, _26675_, _26676_, _26677_, _26678_, _26679_, _26680_, _26681_, _26682_, _26683_, _26684_, _26685_, _26686_, _26687_, _26688_, _26689_, _26690_, _26691_, _26692_, _26693_, _26694_, _26695_, _26696_, _26697_, _26698_, _26699_, _26700_, _26701_, _26702_, _26703_, _26704_, _26705_, _26706_, _26707_, _26708_, _26709_, _26710_, _26711_, _26712_, _26713_, _26714_, _26715_, _26716_, _26717_, _26718_, _26719_, _26720_, _26721_, _26722_, _26723_, _26724_, _26725_, _26726_, _26727_, _26728_, _26729_, _26730_, _26731_, _26732_, _26733_, _26734_, _26735_, _26736_, _26737_, _26738_, _26739_, _26740_, _26741_, _26742_, _26743_, _26744_, _26745_, _26746_, _26747_, _26748_, _26749_, _26750_, _26751_, _26752_, _26753_, _26754_, _26755_, _26756_, _26757_, _26758_, _26759_, _26760_, _26761_, _26762_, _26763_, _26764_, _26765_, _26766_, _26767_, _26768_, _26769_, _26770_, _26771_, _26772_, _26773_, _26774_, _26775_, _26776_, _26777_, _26778_, _26779_, _26780_, _26781_, _26782_, _26783_, _26784_, _26785_, _26786_, _26787_, _26788_, _26789_, _26790_, _26791_, _26792_, _26793_, _26794_, _26795_, _26796_, _26797_, _26798_, _26799_, _26800_, _26801_, _26802_, _26803_, _26804_, _26805_, _26806_, _26807_, _26808_, _26809_, _26810_, _26811_, _26812_, _26813_, _26814_, _26815_, _26816_, _26817_, _26818_, _26819_, _26820_, _26821_, _26822_, _26823_, _26824_, _26825_, _26826_, _26827_, _26828_, _26829_, _26830_, _26831_, _26832_, _26833_, _26834_, _26835_, _26836_, _26837_, _26838_, _26839_, _26840_, _26841_, _26842_, _26843_, _26844_, _26845_, _26846_, _26847_, _26848_, _26849_, _26850_, _26851_, _26852_, _26853_, _26854_, _26855_, _26856_, _26857_, _26858_, _26859_, _26860_, _26861_, _26862_, _26863_, _26864_, _26865_, _26866_, _26867_, _26868_, _26869_, _26870_, _26871_, _26872_, _26873_, _26874_, _26875_, _26876_, _26877_, _26878_, _26879_, _26880_, _26881_, _26882_, _26883_, _26884_, _26885_, _26886_, _26887_, _26888_, _26889_, _26890_, _26891_, _26892_, _26893_, _26894_, _26895_, _26896_, _26897_, _26898_, _26899_, _26900_, _26901_, _26902_, _26903_, _26904_, _26905_, _26906_, _26907_, _26908_, _26909_, _26910_, _26911_, _26912_, _26913_, _26914_, _26915_, _26916_, _26917_, _26918_, _26919_, _26920_, _26921_, _26922_, _26923_, _26924_, _26925_, _26926_, _26927_, _26928_, _26929_, _26930_, _26931_, _26932_, _26933_, _26934_, _26935_, _26936_, _26937_, _26938_, _26939_, _26940_, _26941_, _26942_, _26943_, _26944_, _26945_, _26946_, _26947_, _26948_, _26949_, _26950_, _26951_, _26952_, _26953_, _26954_, _26955_, _26956_, _26957_, _26958_, _26959_, _26960_, _26961_, _26962_, _26963_, _26964_, _26965_, _26966_, _26967_, _26968_, _26969_, _26970_, _26971_, _26972_, _26973_, _26974_, _26975_, _26976_, _26977_, _26978_, _26979_, _26980_, _26981_, _26982_, _26983_, _26984_, _26985_, _26986_, _26987_, _26988_, _26989_, _26990_, _26991_, _26992_, _26993_, _26994_, _26995_, _26996_, _26997_, _26998_, _26999_, _27000_, _27001_, _27002_, _27003_, _27004_, _27005_, _27006_, _27007_, _27008_, _27009_, _27010_, _27011_, _27012_, _27013_, _27014_, _27015_, _27016_, _27017_, _27018_, _27019_, _27020_, _27021_, _27022_, _27023_, _27024_, _27025_, _27026_, _27027_, _27028_, _27029_, _27030_, _27031_, _27032_, _27033_, _27034_, _27035_, _27036_, _27037_, _27038_, _27039_, _27040_, _27041_, _27042_, _27043_, _27044_, _27045_, _27046_, _27047_, _27048_, _27049_, _27050_, _27051_, _27052_, _27053_, _27054_, _27055_, _27056_, _27057_, _27058_, _27059_, _27060_, _27061_, _27062_, _27063_, _27064_, _27065_, _27066_, _27067_, _27068_, _27069_, _27070_, _27071_, _27072_, _27073_, _27074_, _27075_, _27076_, _27077_, _27078_, _27079_, , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , ;
  input [159:0] set1;
  input [159:0] set2;
  input set1[0], set1[1], set1[2], set1[3], set1[4], set1[5], set1[6], set1[7], set1[8], set1[9], set1[10], set1[11], set1[12], set1[13], set1[14], set1[15], set1[16], set1[17], set1[18], set1[19], set1[20], set1[21], set1[22], set1[23], set1[24], set1[25], set1[26], set1[27], set1[28], set1[29], set1[30], set1[31], set1[32], set1[33], set1[34], set1[35], set1[36], set1[37], set1[38], set1[39], set1[40], set1[41], set1[42], set1[43], set1[44], set1[45], set1[46], set1[47], set1[48], set1[49], set1[50], set1[51], set1[52], set1[53], set1[54], set1[55], set1[56], set1[57], set1[58], set1[59], set1[60], set1[61], set1[62], set1[63], set1[64], set1[65], set1[66], set1[67], set1[68], set1[69], set1[70], set1[71], set1[72], set1[73], set1[74], set1[75], set1[76], set1[77], set1[78], set1[79], set1[80], set1[81], set1[82], set1[83], set1[84], set1[85], set1[86], set1[87], set1[88], set1[89], set1[90], set1[91], set1[92], set1[93], set1[94], set1[95], set1[96], set1[97], set1[98], set1[99], set1[100], set1[101], set1[102], set1[103], set1[104], set1[105], set1[106], set1[107], set1[108], set1[109], set1[110], set1[111], set1[112], set1[113], set1[114], set1[115], set1[116], set1[117], set1[118], set1[119], set1[120], set1[121], set1[122], set1[123], set1[124], set1[125], set1[126], set1[127], set1[128], set1[129], set1[130], set1[131], set1[132], set1[133], set1[134], set1[135], set1[136], set1[137], set1[138], set1[139], set1[140], set1[141], set1[142], set1[143], set1[144], set1[145], set1[146], set1[147], set1[148], set1[149], set1[150], set1[151], set1[152], set1[153], set1[154], set1[155], set1[156], set1[157], set1[158], set1[159], set2[0], set2[1], set2[2], set2[3], set2[4], set2[5], set2[6], set2[7], set2[8], set2[9], set2[10], set2[11], set2[12], set2[13], set2[14], set2[15], set2[16], set2[17], set2[18], set2[19], set2[20], set2[21], set2[22], set2[23], set2[24], set2[25], set2[26], set2[27], set2[28], set2[29], set2[30], set2[31], set2[32], set2[33], set2[34], set2[35], set2[36], set2[37], set2[38], set2[39], set2[40], set2[41], set2[42], set2[43], set2[44], set2[45], set2[46], set2[47], set2[48], set2[49], set2[50], set2[51], set2[52], set2[53], set2[54], set2[55], set2[56], set2[57], set2[58], set2[59], set2[60], set2[61], set2[62], set2[63], set2[64], set2[65], set2[66], set2[67], set2[68], set2[69], set2[70], set2[71], set2[72], set2[73], set2[74], set2[75], set2[76], set2[77], set2[78], set2[79], set2[80], set2[81], set2[82], set2[83], set2[84], set2[85], set2[86], set2[87], set2[88], set2[89], set2[90], set2[91], set2[92], set2[93], set2[94], set2[95], set2[96], set2[97], set2[98], set2[99], set2[100], set2[101], set2[102], set2[103], set2[104], set2[105], set2[106], set2[107], set2[108], set2[109], set2[110], set2[111], set2[112], set2[113], set2[114], set2[115], set2[116], set2[117], set2[118], set2[119], set2[120], set2[121], set2[122], set2[123], set2[124], set2[125], set2[126], set2[127], set2[128], set2[129], set2[130], set2[131], set2[132], set2[133], set2[134], set2[135], set2[136], set2[137], set2[138], set2[139], set2[140], set2[141], set2[142], set2[143], set2[144], set2[145], set2[146], set2[147], set2[148], set2[149], set2[150], set2[151], set2[152], set2[153], set2[154], set2[155], set2[156], set2[157], set2[158], set2[159];
  output out[0], out[1], out[2], out[3], out[4], out[5], out[6], out[7], out[8], out[9], out[10], out[11], out[12], out[13], out[14], out[15], out[16], out[17], out[18], out[19], out[20], out[21], out[22], out[23], out[24], out[25], out[26], out[27], out[28], out[29], out[30], out[31], out[32], out[33], out[34], out[35], out[36], out[37], out[38], out[39], out[40], out[41], out[42], out[43], out[44], out[45], out[46], out[47], out[48], out[49], out[50], out[51], out[52], out[53], out[54], out[55], out[56], out[57], out[58], out[59], out[60], out[61], out[62], out[63], out[64], out[65], out[66], out[67], out[68], out[69], out[70], out[71], out[72], out[73], out[74], out[75], out[76], out[77], out[78], out[79], out[80], out[81], out[82], out[83], out[84], out[85], out[86], out[87], out[88], out[89], out[90], out[91], out[92], out[93], out[94], out[95], out[96], out[97], out[98], out[99], out[100], out[101], out[102], out[103], out[104], out[105], out[106], out[107], out[108], out[109], out[110], out[111], out[112], out[113], out[114], out[115], out[116], out[117], out[118], out[119], out[120], out[121], out[122], out[123], out[124], out[125], out[126], out[127], out[128], out[129], out[130], out[131], out[132], out[133], out[134], out[135], out[136], out[137], out[138], out[139], out[140], out[141], out[142], out[143], out[144], out[145], out[146], out[147], out[148], out[149], out[150], out[151], out[152], out[153], out[154], out[155], out[156], out[157], out[158], out[159], out[160], out[161], out[162], out[163], out[164], out[165], out[166], out[167], out[168], out[169], out[170], out[171], out[172], out[173], out[174], out[175], out[176], out[177], out[178], out[179], out[180], out[181], out[182], out[183], out[184], out[185], out[186], out[187], out[188], out[189], out[190], out[191], out[192], out[193], out[194], out[195], out[196], out[197], out[198], out[199], out[200], out[201], out[202], out[203], out[204], out[205], out[206], out[207], out[208], out[209], out[210], out[211], out[212], out[213], out[214], out[215], out[216], out[217], out[218], out[219], out[220], out[221], out[222], out[223], out[224], out[225], out[226], out[227], out[228], out[229], out[230], out[231], out[232], out[233], out[234], out[235], out[236], out[237], out[238], out[239], out[240], out[241], out[242], out[243], out[244], out[245], out[246], out[247], out[248], out[249], out[250], out[251], out[252], out[253], out[254], out[255], out[256], out[257], out[258], out[259], out[260], out[261], out[262], out[263], out[264], out[265], out[266], out[267], out[268], out[269], out[270], out[271], out[272], out[273], out[274], out[275], out[276], out[277], out[278], out[279], out[280], out[281], out[282], out[283], out[284], out[285], out[286], out[287], out[288], out[289], out[290], out[291], out[292], out[293], out[294], out[295], out[296], out[297], out[298], out[299], out[300], out[301], out[302], out[303], out[304], out[305], out[306], out[307], out[308], out[309], out[310], out[311], out[312], out[313], out[314], out[315], out[316], out[317], out[318], out[319], out[320], out[321], out[322], out[323], out[324], out[325], out[326], out[327], out[328], out[329], out[330], out[331], out[332], out[333], out[334], out[335];
  not g_27080_(out[304], _18562_);
  not g_27081_(out[288], _18573_);
  not g_27082_(out[160], _18584_);
  not g_27083_(out[171], _18595_);
  not g_27084_(out[167], _18606_);
  not g_27085_(out[166], _18617_);
  not g_27086_(out[165], _18628_);
  not g_27087_(out[164], _18639_);
  not g_27088_(out[161], _18650_);
  not g_27089_(out[162], _18661_);
  not g_27090_(out[163], _18672_);
  not g_27091_(out[168], _18683_);
  not g_27092_(out[169], _18694_);
  not g_27093_(out[170], _18705_);
  not g_27094_(out[187], _18716_);
  not g_27095_(out[183], _18727_);
  not g_27096_(out[182], _18738_);
  not g_27097_(out[181], _18749_);
  not g_27098_(out[180], _18760_);
  not g_27099_(out[177], _18771_);
  not g_27100_(out[176], _18782_);
  not g_27101_(out[178], _18793_);
  not g_27102_(out[179], _18804_);
  not g_27103_(out[184], _18815_);
  not g_27104_(out[185], _18826_);
  not g_27105_(out[186], _18837_);
  not g_27106_(out[203], _18848_);
  not g_27107_(out[199], _18859_);
  not g_27108_(out[198], _18870_);
  not g_27109_(out[197], _18881_);
  not g_27110_(out[196], _18892_);
  not g_27111_(out[193], _18903_);
  not g_27112_(out[192], _18914_);
  not g_27113_(out[194], _18925_);
  not g_27114_(out[195], _18936_);
  not g_27115_(out[200], _18947_);
  not g_27116_(out[219], _18958_);
  not g_27117_(out[215], _18969_);
  not g_27118_(out[214], _18980_);
  not g_27119_(out[213], _18991_);
  not g_27120_(out[212], _19002_);
  not g_27121_(out[209], _19013_);
  not g_27122_(out[208], _19024_);
  not g_27123_(out[210], _19035_);
  not g_27124_(out[211], _19046_);
  not g_27125_(out[216], _19057_);
  not g_27126_(out[217], _19068_);
  not g_27127_(out[218], _19079_);
  not g_27128_(out[235], _19090_);
  not g_27129_(out[231], _19101_);
  not g_27130_(out[230], _19112_);
  not g_27131_(out[229], _19123_);
  not g_27132_(out[228], _19134_);
  not g_27133_(out[225], _19145_);
  not g_27134_(out[224], _19156_);
  not g_27135_(out[226], _19167_);
  not g_27136_(out[227], _19178_);
  not g_27137_(out[232], _19189_);
  not g_27138_(out[233], _19200_);
  not g_27139_(out[234], _19211_);
  not g_27140_(out[251], _19222_);
  not g_27141_(out[247], _19233_);
  not g_27142_(out[246], _19244_);
  not g_27143_(out[245], _19255_);
  not g_27144_(out[244], _19266_);
  not g_27145_(out[241], _19277_);
  not g_27146_(out[240], _19288_);
  not g_27147_(out[242], _19299_);
  not g_27148_(out[243], _19310_);
  not g_27149_(out[248], _19321_);
  not g_27150_(out[249], _19332_);
  not g_27151_(out[250], _19343_);
  not g_27152_(out[267], _19354_);
  not g_27153_(out[263], _19365_);
  not g_27154_(out[262], _19376_);
  not g_27155_(out[261], _19387_);
  not g_27156_(out[260], _19398_);
  not g_27157_(out[257], _19409_);
  not g_27158_(out[256], _19420_);
  not g_27159_(out[258], _19431_);
  not g_27160_(out[259], _19442_);
  not g_27161_(out[264], _19453_);
  not g_27162_(out[265], _19464_);
  not g_27163_(out[266], _19475_);
  not g_27164_(out[283], _19486_);
  not g_27165_(out[279], _19497_);
  not g_27166_(out[278], _19508_);
  not g_27167_(out[277], _19519_);
  not g_27168_(out[276], _19530_);
  not g_27169_(out[273], _19541_);
  not g_27170_(out[272], _19552_);
  not g_27171_(out[274], _19563_);
  not g_27172_(out[275], _19574_);
  not g_27173_(out[280], _19585_);
  not g_27174_(out[281], _19596_);
  not g_27175_(out[282], _19607_);
  not g_27176_(out[299], _19618_);
  not g_27177_(out[295], _19629_);
  not g_27178_(out[294], _19640_);
  not g_27179_(out[293], _19651_);
  not g_27180_(out[292], _19662_);
  not g_27181_(out[289], _19673_);
  not g_27182_(out[290], _19684_);
  not g_27183_(out[291], _19695_);
  not g_27184_(out[296], _19706_);
  not g_27185_(out[297], _19717_);
  not g_27186_(out[298], _19728_);
  not g_27187_(out[315], _19739_);
  not g_27188_(out[311], _19750_);
  not g_27189_(out[310], _19761_);
  not g_27190_(out[308], _19772_);
  not g_27191_(out[309], _19783_);
  not g_27192_(out[305], _19794_);
  not g_27193_(out[306], _19805_);
  not g_27194_(out[307], _19816_);
  not g_27195_(out[312], _19827_);
  not g_27196_(out[313], _19838_);
  not g_27197_(out[314], _19849_);
  not g_27198_(out[112], _19860_);
  not g_27199_(out[11], _19871_);
  not g_27200_(out[6], _19882_);
  not g_27201_(out[7], _19893_);
  not g_27202_(out[5], _19904_);
  not g_27203_(out[4], _19915_);
  not g_27204_(out[1], _19926_);
  not g_27205_(out[0], _19937_);
  not g_27206_(out[2], _19948_);
  not g_27207_(out[3], _19959_);
  not g_27208_(out[8], _19970_);
  not g_27209_(out[9], _19981_);
  not g_27210_(out[10], _19992_);
  not g_27211_(out[27], _20003_);
  not g_27212_(out[23], _20014_);
  not g_27213_(out[22], _20025_);
  not g_27214_(out[21], _20036_);
  not g_27215_(out[20], _20047_);
  not g_27216_(out[17], _20058_);
  not g_27217_(out[16], _20069_);
  not g_27218_(out[18], _20080_);
  not g_27219_(out[19], _20091_);
  not g_27220_(out[24], _20102_);
  not g_27221_(out[25], _20113_);
  not g_27222_(out[26], _20124_);
  not g_27223_(out[43], _20135_);
  not g_27224_(out[39], _20146_);
  not g_27225_(out[38], _20157_);
  not g_27226_(out[37], _20168_);
  not g_27227_(out[36], _20179_);
  not g_27228_(out[33], _20190_);
  not g_27229_(out[32], _20201_);
  not g_27230_(out[34], _20212_);
  not g_27231_(out[35], _20223_);
  not g_27232_(out[40], _20234_);
  not g_27233_(out[41], _20245_);
  not g_27234_(out[42], _20256_);
  not g_27235_(out[59], _20267_);
  not g_27236_(out[55], _20278_);
  not g_27237_(out[54], _20289_);
  not g_27238_(out[53], _20300_);
  not g_27239_(out[52], _20311_);
  not g_27240_(out[49], _20322_);
  not g_27241_(out[48], _20333_);
  not g_27242_(out[50], _20344_);
  not g_27243_(out[51], _20355_);
  not g_27244_(out[56], _20366_);
  not g_27245_(out[57], _20377_);
  not g_27246_(out[58], _20388_);
  not g_27247_(out[75], _20399_);
  not g_27248_(out[71], _20410_);
  not g_27249_(out[70], _20421_);
  not g_27250_(out[69], _20432_);
  not g_27251_(out[68], _20443_);
  not g_27252_(out[65], _20454_);
  not g_27253_(out[64], _20465_);
  not g_27254_(out[66], _20476_);
  not g_27255_(out[67], _20487_);
  not g_27256_(out[72], _20498_);
  not g_27257_(out[73], _20509_);
  not g_27258_(out[74], _20520_);
  not g_27259_(out[91], _20531_);
  not g_27260_(out[87], _20542_);
  not g_27261_(out[86], _20553_);
  not g_27262_(out[85], _20564_);
  not g_27263_(out[84], _20575_);
  not g_27264_(out[81], _20586_);
  not g_27265_(out[80], _20597_);
  not g_27266_(out[82], _20608_);
  not g_27267_(out[83], _20619_);
  not g_27268_(out[88], _20630_);
  not g_27269_(out[89], _20641_);
  not g_27270_(out[90], _20652_);
  not g_27271_(out[107], _20663_);
  not g_27272_(out[103], _20674_);
  not g_27273_(out[102], _20685_);
  not g_27274_(out[101], _20696_);
  not g_27275_(out[100], _20707_);
  not g_27276_(out[97], _20718_);
  not g_27277_(out[96], _20729_);
  not g_27278_(out[98], _20740_);
  not g_27279_(out[99], _20751_);
  not g_27280_(out[104], _20762_);
  not g_27281_(out[105], _20773_);
  not g_27282_(out[106], _20784_);
  not g_27283_(out[123], _20795_);
  not g_27284_(out[119], _20806_);
  not g_27285_(out[118], _20817_);
  not g_27286_(out[117], _20828_);
  not g_27287_(out[116], _20839_);
  not g_27288_(out[113], _20850_);
  not g_27289_(out[114], _20861_);
  not g_27290_(out[115], _20872_);
  not g_27291_(out[120], _20883_);
  not g_27292_(out[121], _20894_);
  not g_27293_(out[122], _20905_);
  not g_27294_(out[139], _20916_);
  not g_27295_(out[135], _20927_);
  not g_27296_(out[134], _20938_);
  not g_27297_(out[133], _20949_);
  not g_27298_(out[132], _20960_);
  not g_27299_(out[129], _20971_);
  not g_27300_(out[128], _20982_);
  not g_27301_(out[130], _20993_);
  not g_27302_(out[131], _21004_);
  not g_27303_(out[136], _21015_);
  not g_27304_(out[137], _21026_);
  not g_27305_(out[138], _21037_);
  not g_27306_(out[155], _21048_);
  not g_27307_(out[151], _21059_);
  not g_27308_(out[150], _21070_);
  not g_27309_(out[148], _21081_);
  not g_27310_(out[149], _21092_);
  not g_27311_(out[145], _21103_);
  not g_27312_(out[144], _21114_);
  not g_27313_(out[146], _21125_);
  not g_27314_(out[147], _21136_);
  not g_27315_(out[152], _21147_);
  not g_27316_(out[153], _21158_);
  not g_27317_(out[154], _21169_);
  and g_27318_(out[145], out[146], _21180_);
  or g_27319_(out[148], out[147], _21191_);
  or g_27320_(out[147], _21180_, _21202_);
  or g_27321_(_21180_, _21191_, _21213_);
  or g_27322_(out[149], _21213_, _21224_);
  and g_27323_(out[150], _21224_, _21235_);
  and g_27324_(out[151], _21235_, _21246_);
  or g_27325_(out[152], _21246_, _21257_);
  or g_27326_(out[153], _21257_, _21268_);
  xor g_27327_(out[153], _21257_, _21279_);
  not g_27328_(_21279_, _21290_);
  or g_27329_(out[154], _21268_, _21301_);
  xor g_27330_(out[154], _21268_, _21312_);
  xor g_27331_(_21169_, _21268_, _21323_);
  and g_27332_(out[129], out[130], _21334_);
  or g_27333_(out[132], out[131], _21345_);
  or g_27334_(out[131], _21334_, _21356_);
  or g_27335_(_21334_, _21345_, _21367_);
  or g_27336_(out[133], _21367_, _21378_);
  and g_27337_(out[134], _21378_, _21389_);
  and g_27338_(out[135], _21389_, _21400_);
  or g_27339_(out[136], _21400_, _21411_);
  or g_27340_(out[137], _21411_, _21422_);
  or g_27341_(out[138], _21422_, _21433_);
  xor g_27342_(out[138], _21422_, _21444_);
  and g_27343_(out[81], out[82], _21455_);
  or g_27344_(out[84], out[83], _21466_);
  or g_27345_(out[83], _21455_, _21477_);
  or g_27346_(_21455_, _21466_, _21488_);
  or g_27347_(out[85], _21488_, _21499_);
  and g_27348_(out[86], _21499_, _21510_);
  and g_27349_(out[87], _21510_, _21521_);
  or g_27350_(out[88], _21521_, _21532_);
  or g_27351_(out[89], _21532_, _21543_);
  or g_27352_(out[90], _21543_, _21554_);
  xor g_27353_(out[90], _21543_, _21565_);
  xor g_27354_(_20652_, _21543_, _21576_);
  and g_27355_(out[65], out[66], _21587_);
  or g_27356_(out[68], out[67], _21598_);
  or g_27357_(out[67], _21587_, _21609_);
  or g_27358_(_21587_, _21598_, _21620_);
  or g_27359_(out[69], _21620_, _21631_);
  and g_27360_(out[70], _21631_, _21642_);
  and g_27361_(out[71], _21642_, _21653_);
  or g_27362_(out[72], _21653_, _21664_);
  or g_27363_(out[73], _21664_, _21675_);
  or g_27364_(out[74], _21675_, _21686_);
  xor g_27365_(out[75], _21686_, _21697_);
  not g_27366_(_21697_, _21708_);
  and g_27367_(out[49], out[50], _21719_);
  or g_27368_(out[52], out[51], _21730_);
  or g_27369_(out[51], _21719_, _21741_);
  or g_27370_(_21719_, _21730_, _21752_);
  or g_27371_(out[53], _21752_, _21763_);
  and g_27372_(out[54], _21763_, _21774_);
  and g_27373_(out[55], _21774_, _21785_);
  or g_27374_(out[56], _21785_, _21796_);
  or g_27375_(out[57], _21796_, _21807_);
  or g_27376_(out[58], _21807_, _21818_);
  xor g_27377_(_20267_, _21818_, _21829_);
  xor g_27378_(out[59], _21818_, _21840_);
  and g_27379_(out[1], out[2], _21851_);
  or g_27380_(out[4], out[3], _21862_);
  or g_27381_(out[3], _21851_, _21873_);
  or g_27382_(_21851_, _21862_, _21884_);
  or g_27383_(out[5], _21884_, _21895_);
  and g_27384_(out[6], _21895_, _21906_);
  and g_27385_(out[7], _21906_, _21917_);
  or g_27386_(out[8], _21917_, _21928_);
  or g_27387_(out[9], _21928_, _21939_);
  or g_27388_(out[10], _21939_, _21950_);
  xor g_27389_(out[10], _21939_, _21961_);
  xor g_27390_(_19992_, _21939_, _21972_);
  xor g_27391_(out[7], _21906_, _21983_);
  not g_27392_(_21983_, _21994_);
  and g_27393_(out[17], out[18], _22005_);
  or g_27394_(out[20], out[19], _22016_);
  or g_27395_(out[19], _22005_, _22027_);
  or g_27396_(_22005_, _22016_, _22038_);
  or g_27397_(out[21], _22038_, _22049_);
  and g_27398_(out[22], _22049_, _22060_);
  and g_27399_(out[23], _22060_, _22071_);
  xor g_27400_(out[23], _22060_, _22082_);
  not g_27401_(_22082_, _22093_);
  and g_27402_(_21994_, _22082_, _22104_);
  or g_27403_(_21983_, _22093_, _22115_);
  xor g_27404_(out[6], _21895_, _22126_);
  not g_27405_(_22126_, _22137_);
  xor g_27406_(out[22], _22049_, _22148_);
  not g_27407_(_22148_, _22159_);
  and g_27408_(_22126_, _22159_, _22170_);
  or g_27409_(_22137_, _22148_, _22181_);
  xor g_27410_(out[4], _21873_, _22192_);
  xor g_27411_(_19915_, _21873_, _22203_);
  xor g_27412_(out[20], _22027_, _22214_);
  xor g_27413_(_20047_, _22027_, _22225_);
  and g_27414_(_22203_, _22214_, _22236_);
  or g_27415_(_22192_, _22225_, _22247_);
  xor g_27416_(out[5], _21884_, _22258_);
  xor g_27417_(_19904_, _21884_, _22269_);
  xor g_27418_(out[21], _22038_, _22280_);
  xor g_27419_(_20036_, _22038_, _22291_);
  and g_27420_(_22269_, _22280_, _22302_);
  or g_27421_(_22258_, _22291_, _22313_);
  and g_27422_(_22247_, _22313_, _22324_);
  or g_27423_(_22236_, _22302_, _22335_);
  xor g_27424_(out[3], _21851_, _22346_);
  xor g_27425_(_19959_, _21851_, _22357_);
  xor g_27426_(out[19], _22005_, _22368_);
  or g_27427_(_22357_, _22368_, _22379_);
  or g_27428_(out[17], out[18], _22390_);
  xor g_27429_(out[17], out[18], _22401_);
  xor g_27430_(_20058_, out[18], _22412_);
  or g_27431_(out[1], out[2], _22423_);
  xor g_27432_(out[1], out[2], _22434_);
  xor g_27433_(_19926_, out[2], _22445_);
  and g_27434_(_22412_, _22434_, _22456_);
  and g_27435_(_22401_, _22445_, _22467_);
  or g_27436_(_22412_, _22434_, _22478_);
  xor g_27437_(_22412_, _22434_, _22489_);
  or g_27438_(_22456_, _22467_, _22500_);
  and g_27439_(_22357_, _22368_, _22511_);
  xor g_27440_(_22357_, _22368_, _22522_);
  xor g_27441_(_22346_, _22368_, _22533_);
  and g_27442_(_22489_, _22522_, _22544_);
  or g_27443_(_22500_, _22533_, _22555_);
  and g_27444_(_19926_, out[17], _22566_);
  or g_27445_(out[1], _20058_, _22577_);
  and g_27446_(out[1], _20058_, _22588_);
  or g_27447_(_19926_, out[17], _22599_);
  and g_27448_(_19937_, out[16], _22610_);
  or g_27449_(out[0], _20069_, _22621_);
  and g_27450_(_22599_, _22621_, _22632_);
  or g_27451_(_22588_, _22610_, _22643_);
  and g_27452_(_22577_, _22643_, _22654_);
  or g_27453_(_22566_, _22632_, _22665_);
  and g_27454_(_22544_, _22665_, _22676_);
  or g_27455_(_22555_, _22654_, _22687_);
  and g_27456_(_22379_, _22456_, _22698_);
  or g_27457_(_22511_, _22698_, _22709_);
  not g_27458_(_22709_, _22720_);
  and g_27459_(_22687_, _22720_, _22731_);
  or g_27460_(_22676_, _22709_, _22742_);
  and g_27461_(out[0], _20069_, _22753_);
  or g_27462_(_19937_, out[16], _22764_);
  and g_27463_(_22577_, _22632_, _22775_);
  or g_27464_(_22566_, _22643_, _22786_);
  and g_27465_(_22764_, _22775_, _22797_);
  or g_27466_(_22753_, _22786_, _22808_);
  and g_27467_(_22544_, _22797_, _22819_);
  or g_27468_(_22555_, _22808_, _22830_);
  and g_27469_(_22192_, _22225_, _22841_);
  or g_27470_(_22203_, _22214_, _22852_);
  and g_27471_(_22830_, _22852_, _22863_);
  or g_27472_(_22819_, _22841_, _22874_);
  and g_27473_(_22742_, _22863_, _22885_);
  or g_27474_(_22731_, _22874_, _22896_);
  and g_27475_(_22324_, _22896_, _22907_);
  or g_27476_(_22335_, _22885_, _22918_);
  and g_27477_(_22137_, _22148_, _22929_);
  or g_27478_(_22126_, _22159_, _22940_);
  and g_27479_(_22258_, _22291_, _22951_);
  or g_27480_(_22269_, _22280_, _22962_);
  and g_27481_(_22940_, _22962_, _22973_);
  or g_27482_(_22929_, _22951_, _22984_);
  and g_27483_(_22918_, _22973_, _22995_);
  or g_27484_(_22907_, _22984_, _23006_);
  or g_27485_(out[1], out[0], _23017_);
  not g_27486_(_23017_, _23028_);
  or g_27487_(out[2], _23017_, _23039_);
  and g_27488_(out[4], out[3], _23050_);
  and g_27489_(out[3], _23039_, _23061_);
  and g_27490_(_23039_, _23050_, _23072_);
  xor g_27491_(out[4], _23061_, _23083_);
  xor g_27492_(_19915_, _23061_, _23094_);
  or g_27493_(out[17], out[16], _23105_);
  not g_27494_(_23105_, _23116_);
  or g_27495_(out[16], _22390_, _23127_);
  and g_27496_(out[20], out[19], _23138_);
  and g_27497_(out[19], _23127_, _23149_);
  and g_27498_(_23127_, _23138_, _23160_);
  xor g_27499_(out[20], _23149_, _23171_);
  xor g_27500_(_20047_, _23149_, _23182_);
  and g_27501_(_23094_, _23171_, _23193_);
  or g_27502_(_23083_, _23182_, _23204_);
  and g_27503_(out[5], _23072_, _23215_);
  xor g_27504_(out[5], _23072_, _23226_);
  xor g_27505_(_19904_, _23072_, _23237_);
  and g_27506_(out[21], _23160_, _23248_);
  xor g_27507_(out[21], _23160_, _23259_);
  xor g_27508_(_20036_, _23160_, _23270_);
  and g_27509_(_23237_, _23259_, _23281_);
  or g_27510_(_23226_, _23270_, _23292_);
  and g_27511_(_23226_, _23270_, _23303_);
  or g_27512_(_23237_, _23259_, _23314_);
  and g_27513_(_23083_, _23182_, _23325_);
  or g_27514_(_23094_, _23171_, _23336_);
  and g_27515_(_23314_, _23336_, _23347_);
  or g_27516_(_23303_, _23325_, _23358_);
  and g_27517_(_22181_, _23006_, _23369_);
  or g_27518_(_22170_, _22995_, _23380_);
  and g_27519_(_22115_, _23380_, _23391_);
  or g_27520_(_22104_, _23369_, _23402_);
  xor g_27521_(out[8], _21917_, _23413_);
  xor g_27522_(_19970_, _21917_, _23424_);
  or g_27523_(out[24], _22071_, _23435_);
  xor g_27524_(out[24], _22071_, _23446_);
  xor g_27525_(_20102_, _22071_, _23457_);
  and g_27526_(_23424_, _23446_, _23468_);
  or g_27527_(_23413_, _23457_, _23479_);
  and g_27528_(_21983_, _22093_, _23490_);
  or g_27529_(_21994_, _22082_, _23501_);
  and g_27530_(_23479_, _23501_, _23512_);
  or g_27531_(_23468_, _23490_, _23523_);
  and g_27532_(_23402_, _23512_, _23534_);
  or g_27533_(_23391_, _23523_, _23545_);
  xor g_27534_(out[9], _21928_, _23556_);
  xor g_27535_(_19981_, _21928_, _23567_);
  or g_27536_(out[25], _23435_, _23578_);
  xor g_27537_(out[25], _23435_, _23589_);
  xor g_27538_(_20113_, _23435_, _23600_);
  and g_27539_(_23556_, _23600_, _23611_);
  or g_27540_(_23567_, _23589_, _23622_);
  and g_27541_(_23413_, _23457_, _23633_);
  or g_27542_(_23424_, _23446_, _23644_);
  and g_27543_(_23622_, _23644_, _23655_);
  or g_27544_(_23611_, _23633_, _23666_);
  and g_27545_(_23545_, _23655_, _23677_);
  or g_27546_(_23534_, _23666_, _23688_);
  or g_27547_(out[26], _23578_, _23699_);
  xor g_27548_(out[26], _23578_, _23710_);
  xor g_27549_(_20124_, _23578_, _23721_);
  and g_27550_(_21972_, _23710_, _23732_);
  or g_27551_(_21961_, _23721_, _23743_);
  and g_27552_(_23567_, _23589_, _23754_);
  or g_27553_(_23556_, _23600_, _23765_);
  and g_27554_(_23743_, _23765_, _23776_);
  or g_27555_(_23732_, _23754_, _23787_);
  and g_27556_(_23688_, _23776_, _23798_);
  or g_27557_(_23677_, _23787_, _23809_);
  and g_27558_(_21961_, _23721_, _23820_);
  or g_27559_(_21972_, _23710_, _23831_);
  xor g_27560_(_20003_, _23699_, _23842_);
  xor g_27561_(out[27], _23699_, _23853_);
  xor g_27562_(_19871_, _21950_, _23864_);
  xor g_27563_(out[11], _21950_, _23875_);
  and g_27564_(_23842_, _23875_, _23886_);
  or g_27565_(_23853_, _23864_, _23897_);
  and g_27566_(_23831_, _23897_, _23908_);
  or g_27567_(_23820_, _23886_, _23919_);
  and g_27568_(_23809_, _23908_, _23930_);
  or g_27569_(_23798_, _23919_, _23941_);
  and g_27570_(_23853_, _23864_, _23952_);
  or g_27571_(_23842_, _23875_, _23963_);
  and g_27572_(_23941_, _23963_, _23974_);
  or g_27573_(_23930_, _23952_, _23985_);
  and g_27574_(_21961_, _23974_, _23996_);
  or g_27575_(_21972_, _23985_, _24007_);
  and g_27576_(_23710_, _23985_, _24018_);
  or g_27577_(_23721_, _23974_, _24029_);
  and g_27578_(_24007_, _24029_, _24040_);
  or g_27579_(_23996_, _24018_, _24051_);
  and g_27580_(out[33], out[34], _24062_);
  or g_27581_(out[35], _24062_, _24073_);
  xor g_27582_(out[35], _24062_, _24084_);
  xor g_27583_(_20223_, _24062_, _24095_);
  and g_27584_(_22346_, _23974_, _24106_);
  and g_27585_(_22368_, _23985_, _24117_);
  or g_27586_(_24106_, _24117_, _24128_);
  not g_27587_(_24128_, _24139_);
  and g_27588_(_24084_, _24139_, _24150_);
  or g_27589_(_24095_, _24128_, _24161_);
  or g_27590_(out[33], out[34], _24172_);
  xor g_27591_(out[33], out[34], _24183_);
  xor g_27592_(_20190_, out[34], _24194_);
  or g_27593_(_22401_, _23974_, _24205_);
  or g_27594_(_22434_, _23985_, _24216_);
  and g_27595_(_24205_, _24216_, _24227_);
  not g_27596_(_24227_, _24238_);
  and g_27597_(_24194_, _24227_, _24249_);
  or g_27598_(_24183_, _24238_, _24260_);
  and g_27599_(_24161_, _24260_, _24271_);
  or g_27600_(_24150_, _24249_, _24282_);
  and g_27601_(_24095_, _24128_, _24293_);
  or g_27602_(_24084_, _24139_, _24304_);
  and g_27603_(_24183_, _24238_, _24315_);
  or g_27604_(_24194_, _24227_, _24326_);
  and g_27605_(_24304_, _24326_, _24337_);
  or g_27606_(_24293_, _24315_, _24348_);
  and g_27607_(_24271_, _24337_, _24359_);
  or g_27608_(_24282_, _24348_, _24370_);
  and g_27609_(out[17], _23985_, _24381_);
  or g_27610_(_20058_, _23974_, _24392_);
  and g_27611_(out[1], _23974_, _24403_);
  or g_27612_(_19926_, _23985_, _24414_);
  and g_27613_(_24392_, _24414_, _24425_);
  or g_27614_(_24381_, _24403_, _24436_);
  and g_27615_(out[33], _24425_, _24447_);
  or g_27616_(_20190_, _24436_, _24458_);
  and g_27617_(_19937_, _23974_, _24469_);
  or g_27618_(out[0], _23985_, _24480_);
  and g_27619_(_20069_, _23985_, _24491_);
  or g_27620_(out[16], _23974_, _24502_);
  and g_27621_(_24480_, _24502_, _24513_);
  or g_27622_(_24469_, _24491_, _24524_);
  and g_27623_(out[32], _24524_, _24535_);
  or g_27624_(_20201_, _24513_, _24546_);
  xor g_27625_(out[33], _24425_, _24557_);
  xor g_27626_(_20190_, _24425_, _24568_);
  and g_27627_(_24546_, _24557_, _24579_);
  or g_27628_(_24535_, _24568_, _24590_);
  and g_27629_(_24458_, _24590_, _24601_);
  or g_27630_(_24447_, _24579_, _24612_);
  and g_27631_(_24359_, _24612_, _24623_);
  or g_27632_(_24370_, _24601_, _24634_);
  and g_27633_(_24282_, _24304_, _24645_);
  or g_27634_(_24271_, _24293_, _24656_);
  and g_27635_(_24634_, _24656_, _24667_);
  or g_27636_(_24623_, _24645_, _24678_);
  and g_27637_(_23842_, _23864_, _24689_);
  or g_27638_(_23853_, _23875_, _24700_);
  or g_27639_(out[36], out[35], _24711_);
  or g_27640_(_24062_, _24711_, _24722_);
  or g_27641_(out[37], _24722_, _24733_);
  and g_27642_(out[38], _24733_, _24744_);
  and g_27643_(out[39], _24744_, _24755_);
  or g_27644_(out[40], _24755_, _24766_);
  or g_27645_(out[41], _24766_, _24777_);
  or g_27646_(out[42], _24777_, _24788_);
  xor g_27647_(_20135_, _24788_, _24799_);
  xor g_27648_(out[43], _24788_, _24810_);
  and g_27649_(_24689_, _24810_, _24821_);
  or g_27650_(_24700_, _24799_, _24832_);
  xor g_27651_(out[42], _24777_, _24843_);
  xor g_27652_(_20256_, _24777_, _24854_);
  and g_27653_(_24040_, _24843_, _24865_);
  or g_27654_(_24051_, _24854_, _24876_);
  and g_27655_(_24832_, _24876_, _24887_);
  or g_27656_(_24821_, _24865_, _24898_);
  and g_27657_(_24051_, _24854_, _24909_);
  or g_27658_(_24040_, _24843_, _24920_);
  and g_27659_(_24700_, _24799_, _24931_);
  or g_27660_(_24689_, _24810_, _24942_);
  xor g_27661_(out[41], _24766_, _24953_);
  xor g_27662_(_20245_, _24766_, _24964_);
  and g_27663_(_23556_, _23974_, _24975_);
  or g_27664_(_23567_, _23985_, _24986_);
  and g_27665_(_23589_, _23985_, _24997_);
  or g_27666_(_23600_, _23974_, _25008_);
  and g_27667_(_24986_, _25008_, _25019_);
  or g_27668_(_24975_, _24997_, _25030_);
  and g_27669_(_24964_, _25030_, _25041_);
  or g_27670_(_24953_, _25019_, _25052_);
  and g_27671_(_24920_, _24942_, _25063_);
  or g_27672_(_24909_, _24931_, _25074_);
  and g_27673_(_24887_, _25063_, _25085_);
  or g_27674_(_24898_, _25074_, _25096_);
  and g_27675_(_25052_, _25085_, _25107_);
  or g_27676_(_25041_, _25096_, _25118_);
  and g_27677_(_24953_, _25019_, _25129_);
  or g_27678_(_24964_, _25030_, _25140_);
  xor g_27679_(out[40], _24755_, _25151_);
  xor g_27680_(_20234_, _24755_, _25162_);
  and g_27681_(_23446_, _23985_, _25173_);
  or g_27682_(_23457_, _23974_, _25184_);
  and g_27683_(_23413_, _23974_, _25195_);
  or g_27684_(_23424_, _23985_, _25206_);
  and g_27685_(_25184_, _25206_, _25217_);
  or g_27686_(_25173_, _25195_, _25228_);
  and g_27687_(_25151_, _25217_, _25239_);
  or g_27688_(_25162_, _25228_, _25250_);
  and g_27689_(_25140_, _25250_, _25261_);
  or g_27690_(_25129_, _25239_, _25272_);
  and g_27691_(_25162_, _25228_, _25283_);
  or g_27692_(_25151_, _25217_, _25294_);
  and g_27693_(_25261_, _25294_, _25305_);
  or g_27694_(_25272_, _25283_, _25316_);
  and g_27695_(_25107_, _25305_, _25327_);
  or g_27696_(_25118_, _25316_, _25338_);
  xor g_27697_(out[39], _24744_, _25349_);
  xor g_27698_(_20146_, _24744_, _25360_);
  or g_27699_(_21983_, _23985_, _25371_);
  or g_27700_(_22082_, _23974_, _25382_);
  and g_27701_(_25371_, _25382_, _25393_);
  not g_27702_(_25393_, _25404_);
  and g_27703_(_25360_, _25393_, _25415_);
  xor g_27704_(out[38], _24733_, _25426_);
  xor g_27705_(_20157_, _24733_, _25437_);
  or g_27706_(_22126_, _23985_, _25448_);
  or g_27707_(_22148_, _23974_, _25459_);
  and g_27708_(_25448_, _25459_, _25470_);
  not g_27709_(_25470_, _25481_);
  and g_27710_(_25437_, _25470_, _25492_);
  or g_27711_(_25360_, _25393_, _25503_);
  xor g_27712_(_25437_, _25470_, _25514_);
  xor g_27713_(_25426_, _25470_, _25525_);
  xor g_27714_(_25360_, _25393_, _25536_);
  xor g_27715_(_25349_, _25393_, _25547_);
  and g_27716_(_25514_, _25536_, _25558_);
  or g_27717_(_25525_, _25547_, _25569_);
  xor g_27718_(out[37], _24722_, _25580_);
  xor g_27719_(_20168_, _24722_, _25591_);
  and g_27720_(_22258_, _23974_, _25602_);
  or g_27721_(_22269_, _23985_, _25613_);
  and g_27722_(_22280_, _23985_, _25624_);
  or g_27723_(_22291_, _23974_, _25635_);
  and g_27724_(_25613_, _25635_, _25646_);
  or g_27725_(_25602_, _25624_, _25657_);
  and g_27726_(_25580_, _25646_, _25668_);
  or g_27727_(_25591_, _25657_, _25679_);
  xor g_27728_(out[36], _24073_, _25690_);
  xor g_27729_(_20179_, _24073_, _25701_);
  and g_27730_(_22192_, _23974_, _25712_);
  or g_27731_(_22203_, _23985_, _25723_);
  and g_27732_(_22214_, _23985_, _25734_);
  or g_27733_(_22225_, _23974_, _25745_);
  and g_27734_(_25723_, _25745_, _25756_);
  or g_27735_(_25712_, _25734_, _25767_);
  and g_27736_(_25690_, _25756_, _25778_);
  or g_27737_(_25701_, _25767_, _25789_);
  and g_27738_(_25679_, _25789_, _25800_);
  or g_27739_(_25668_, _25778_, _25811_);
  and g_27740_(_25591_, _25657_, _25822_);
  or g_27741_(_25580_, _25646_, _25833_);
  and g_27742_(_25701_, _25767_, _25844_);
  or g_27743_(_25690_, _25756_, _25855_);
  and g_27744_(_25833_, _25855_, _25866_);
  or g_27745_(_25822_, _25844_, _25877_);
  and g_27746_(_25800_, _25866_, _25888_);
  or g_27747_(_25811_, _25877_, _25899_);
  and g_27748_(_25558_, _25888_, _25910_);
  or g_27749_(_25569_, _25899_, _25921_);
  and g_27750_(_25327_, _25910_, _25932_);
  or g_27751_(_25338_, _25921_, _25943_);
  and g_27752_(_24678_, _25932_, _25954_);
  or g_27753_(_24667_, _25943_, _25965_);
  and g_27754_(_24898_, _24942_, _25976_);
  or g_27755_(_24887_, _24931_, _25987_);
  and g_27756_(_25107_, _25272_, _25998_);
  or g_27757_(_25118_, _25261_, _26009_);
  and g_27758_(_25987_, _26009_, _26020_);
  or g_27759_(_25976_, _25998_, _26031_);
  and g_27760_(_25558_, _25811_, _26042_);
  or g_27761_(_25569_, _25800_, _26053_);
  and g_27762_(_25833_, _26042_, _26064_);
  or g_27763_(_25822_, _26053_, _26075_);
  and g_27764_(_25492_, _25503_, _26086_);
  or g_27765_(_25415_, _26086_, _26097_);
  not g_27766_(_26097_, _26108_);
  and g_27767_(_26075_, _26108_, _26119_);
  or g_27768_(_26064_, _26097_, _26130_);
  and g_27769_(_25327_, _26130_, _26141_);
  or g_27770_(_25338_, _26119_, _26152_);
  and g_27771_(_26020_, _26152_, _26163_);
  or g_27772_(_26031_, _26141_, _26174_);
  and g_27773_(_25965_, _26163_, _26185_);
  or g_27774_(_25954_, _26174_, _26196_);
  and g_27775_(_20201_, _24513_, _26207_);
  or g_27776_(_24370_, _26207_, _26218_);
  not g_27777_(_26218_, _26229_);
  and g_27778_(_24579_, _26229_, _26240_);
  or g_27779_(_24590_, _26218_, _26251_);
  and g_27780_(_25932_, _26240_, _26262_);
  or g_27781_(_25943_, _26251_, _26273_);
  and g_27782_(_26196_, _26273_, _26284_);
  or g_27783_(_26185_, _26262_, _26295_);
  and g_27784_(_24051_, _26295_, _26306_);
  or g_27785_(_24040_, _26284_, _26317_);
  and g_27786_(_24843_, _26284_, _26328_);
  or g_27787_(_24854_, _26295_, _26339_);
  and g_27788_(_26317_, _26339_, _26350_);
  or g_27789_(_26306_, _26328_, _26361_);
  xor g_27790_(out[58], _21807_, _26372_);
  xor g_27791_(_20388_, _21807_, _26383_);
  and g_27792_(_26350_, _26372_, _26394_);
  or g_27793_(_26361_, _26383_, _26405_);
  and g_27794_(_24810_, _26284_, _26416_);
  or g_27795_(_24799_, _26295_, _26427_);
  and g_27796_(_24700_, _26295_, _26438_);
  or g_27797_(_24689_, _26284_, _26449_);
  and g_27798_(_26427_, _26449_, _26460_);
  or g_27799_(_26416_, _26438_, _26471_);
  and g_27800_(_21840_, _26460_, _26482_);
  or g_27801_(_21829_, _26471_, _26493_);
  and g_27802_(_26405_, _26493_, _26504_);
  or g_27803_(_26394_, _26482_, _26515_);
  xor g_27804_(out[57], _21796_, _26526_);
  xor g_27805_(_20377_, _21796_, _26537_);
  and g_27806_(_24953_, _26284_, _26548_);
  not g_27807_(_26548_, _26559_);
  or g_27808_(_25019_, _26284_, _26570_);
  not g_27809_(_26570_, _26581_);
  and g_27810_(_26559_, _26570_, _26592_);
  or g_27811_(_26548_, _26581_, _26603_);
  and g_27812_(_26537_, _26603_, _26614_);
  or g_27813_(_26526_, _26592_, _26625_);
  and g_27814_(_21829_, _26471_, _26636_);
  or g_27815_(_21840_, _26460_, _26647_);
  and g_27816_(_26361_, _26383_, _26658_);
  or g_27817_(_26350_, _26372_, _26669_);
  and g_27818_(_26647_, _26669_, _26680_);
  or g_27819_(_26636_, _26658_, _26691_);
  and g_27820_(_26625_, _26680_, _26702_);
  or g_27821_(_26614_, _26691_, _26713_);
  and g_27822_(_26504_, _26702_, _26724_);
  or g_27823_(_26515_, _26713_, _26735_);
  xor g_27824_(out[56], _21785_, _26746_);
  xor g_27825_(_20366_, _21785_, _26757_);
  and g_27826_(_25151_, _26284_, _26768_);
  not g_27827_(_26768_, _26779_);
  or g_27828_(_25217_, _26284_, _26790_);
  not g_27829_(_26790_, _26801_);
  and g_27830_(_26779_, _26790_, _26812_);
  or g_27831_(_26768_, _26801_, _26823_);
  and g_27832_(_26757_, _26823_, _26834_);
  or g_27833_(_26746_, _26812_, _09284_);
  and g_27834_(_26526_, _26592_, _09295_);
  or g_27835_(_26537_, _26603_, _09306_);
  and g_27836_(_26746_, _26812_, _09317_);
  or g_27837_(_26757_, _26823_, _09328_);
  and g_27838_(_09306_, _09328_, _09339_);
  or g_27839_(_09295_, _09317_, _09350_);
  and g_27840_(_09284_, _09339_, _09361_);
  or g_27841_(_26834_, _09350_, _09372_);
  and g_27842_(_26724_, _09361_, _09383_);
  or g_27843_(_26735_, _09372_, _09394_);
  xor g_27844_(out[54], _21763_, _09405_);
  xor g_27845_(_20289_, _21763_, _09416_);
  and g_27846_(_25437_, _26284_, _09427_);
  or g_27847_(_25426_, _26295_, _09438_);
  and g_27848_(_25481_, _26295_, _09449_);
  or g_27849_(_25470_, _26284_, _09460_);
  and g_27850_(_09438_, _09460_, _09471_);
  or g_27851_(_09427_, _09449_, _09482_);
  and g_27852_(_09416_, _09471_, _09493_);
  or g_27853_(_09405_, _09482_, _09504_);
  xor g_27854_(out[55], _21774_, _09515_);
  xor g_27855_(_20278_, _21774_, _09526_);
  and g_27856_(_25349_, _26284_, _09537_);
  or g_27857_(_25360_, _26295_, _09548_);
  and g_27858_(_25393_, _26295_, _09559_);
  or g_27859_(_25404_, _26284_, _09570_);
  and g_27860_(_09548_, _09570_, _09581_);
  or g_27861_(_09537_, _09559_, _09592_);
  and g_27862_(_09526_, _09592_, _09603_);
  or g_27863_(_09515_, _09581_, _09614_);
  and g_27864_(_09504_, _09614_, _09625_);
  or g_27865_(_09493_, _09603_, _09636_);
  and g_27866_(_09515_, _09581_, _09647_);
  or g_27867_(_09526_, _09592_, _09658_);
  and g_27868_(_09405_, _09482_, _09669_);
  or g_27869_(_09416_, _09471_, _09680_);
  and g_27870_(_09658_, _09680_, _09691_);
  or g_27871_(_09647_, _09669_, _09702_);
  and g_27872_(_09625_, _09691_, _09713_);
  or g_27873_(_09636_, _09702_, _09724_);
  xor g_27874_(out[52], _21741_, _09735_);
  xor g_27875_(_20311_, _21741_, _09746_);
  and g_27876_(_25690_, _26284_, _09757_);
  or g_27877_(_25701_, _26295_, _09768_);
  and g_27878_(_25767_, _26295_, _09779_);
  or g_27879_(_25756_, _26284_, _09790_);
  and g_27880_(_09768_, _09790_, _09801_);
  or g_27881_(_09757_, _09779_, _09812_);
  and g_27882_(_09735_, _09801_, _09823_);
  or g_27883_(_09746_, _09812_, _09834_);
  xor g_27884_(out[53], _21752_, _09845_);
  xor g_27885_(_20300_, _21752_, _09856_);
  and g_27886_(_25591_, _26284_, _09867_);
  or g_27887_(_25580_, _26295_, _09878_);
  and g_27888_(_25646_, _26295_, _09889_);
  or g_27889_(_25657_, _26284_, _09900_);
  and g_27890_(_09878_, _09900_, _09911_);
  or g_27891_(_09867_, _09889_, _09922_);
  and g_27892_(_09845_, _09922_, _09933_);
  or g_27893_(_09856_, _09911_, _09944_);
  and g_27894_(_09834_, _09944_, _09955_);
  or g_27895_(_09823_, _09933_, _09966_);
  and g_27896_(_09856_, _09911_, _09977_);
  or g_27897_(_09845_, _09922_, _09988_);
  and g_27898_(_09746_, _09812_, _09999_);
  or g_27899_(_09735_, _09801_, _10010_);
  and g_27900_(_09988_, _10010_, _10021_);
  or g_27901_(_09977_, _09999_, _10032_);
  and g_27902_(_09955_, _10021_, _10043_);
  or g_27903_(_09966_, _10032_, _10054_);
  and g_27904_(_09713_, _10043_, _10065_);
  or g_27905_(_09724_, _10054_, _10076_);
  and g_27906_(_09383_, _10065_, _10087_);
  or g_27907_(_09394_, _10076_, _10098_);
  xor g_27908_(out[51], _21719_, _10109_);
  xor g_27909_(_20355_, _21719_, _10120_);
  and g_27910_(_24139_, _26295_, _10131_);
  or g_27911_(_24128_, _26284_, _10142_);
  and g_27912_(_24095_, _26284_, _10153_);
  or g_27913_(_24084_, _26295_, _10164_);
  and g_27914_(_10142_, _10164_, _10175_);
  or g_27915_(_10131_, _10153_, _10186_);
  and g_27916_(_10109_, _10186_, _10197_);
  or g_27917_(_10120_, _10175_, _10208_);
  or g_27918_(out[49], out[50], _10219_);
  xor g_27919_(out[49], out[50], _10230_);
  xor g_27920_(_20322_, out[50], _10241_);
  or g_27921_(_24227_, _26284_, _10252_);
  or g_27922_(_24183_, _26295_, _10263_);
  and g_27923_(_10252_, _10263_, _10274_);
  not g_27924_(_10274_, _10285_);
  and g_27925_(_10230_, _10285_, _10296_);
  or g_27926_(_10197_, _10296_, _10307_);
  and g_27927_(_10120_, _10175_, _10318_);
  or g_27928_(_10109_, _10186_, _10329_);
  and g_27929_(_10241_, _10274_, _10340_);
  or g_27930_(_10230_, _10285_, _10351_);
  or g_27931_(_10318_, _10340_, _10362_);
  xor g_27932_(_10241_, _10274_, _10373_);
  and g_27933_(_10208_, _10329_, _10384_);
  and g_27934_(_10373_, _10384_, _10395_);
  or g_27935_(_10307_, _10362_, _10406_);
  and g_27936_(out[33], _26284_, _10417_);
  not g_27937_(_10417_, _10428_);
  and g_27938_(_24436_, _26295_, _10439_);
  or g_27939_(_24425_, _26284_, _10450_);
  and g_27940_(_10428_, _10450_, _10461_);
  or g_27941_(_10417_, _10439_, _10472_);
  and g_27942_(out[49], _10461_, _10483_);
  or g_27943_(_20322_, _10472_, _10494_);
  xor g_27944_(_20322_, _10472_, _10505_);
  xor g_27945_(out[49], _10472_, _10516_);
  or g_27946_(_24513_, _26284_, _10527_);
  not g_27947_(_10527_, _10538_);
  and g_27948_(_20201_, _26284_, _10549_);
  or g_27949_(out[32], _26295_, _10560_);
  and g_27950_(_10527_, _10560_, _10571_);
  or g_27951_(_10538_, _10549_, _10582_);
  and g_27952_(out[48], _10582_, _10593_);
  or g_27953_(_20333_, _10571_, _10604_);
  and g_27954_(_10505_, _10604_, _10615_);
  or g_27955_(_10516_, _10593_, _10626_);
  and g_27956_(_10395_, _10615_, _10637_);
  or g_27957_(_10406_, _10626_, _10648_);
  and g_27958_(_10329_, _10340_, _10659_);
  or g_27959_(_10318_, _10351_, _10670_);
  and g_27960_(_10208_, _10670_, _10681_);
  or g_27961_(_10197_, _10659_, _10692_);
  and g_27962_(_10395_, _10483_, _10703_);
  or g_27963_(_10406_, _10494_, _10714_);
  and g_27964_(_10681_, _10714_, _10725_);
  or g_27965_(_10692_, _10703_, _10736_);
  and g_27966_(_10648_, _10725_, _10747_);
  or g_27967_(_10637_, _10736_, _10758_);
  and g_27968_(_10087_, _10758_, _10769_);
  or g_27969_(_10098_, _10747_, _10780_);
  and g_27970_(_09636_, _09658_, _10791_);
  or g_27971_(_09625_, _09647_, _10802_);
  and g_27972_(_09966_, _09988_, _10813_);
  or g_27973_(_09955_, _09977_, _10824_);
  and g_27974_(_09713_, _10813_, _10835_);
  or g_27975_(_09724_, _10824_, _10846_);
  and g_27976_(_10802_, _10846_, _10857_);
  or g_27977_(_10791_, _10835_, _10868_);
  and g_27978_(_09383_, _10868_, _10879_);
  or g_27979_(_09394_, _10857_, _10890_);
  and g_27980_(_26515_, _26647_, _10901_);
  or g_27981_(_26504_, _26636_, _10912_);
  and g_27982_(_26724_, _09350_, _10923_);
  or g_27983_(_26735_, _09339_, _10934_);
  and g_27984_(_10912_, _10934_, _10945_);
  or g_27985_(_10901_, _10923_, _10956_);
  and g_27986_(_10890_, _10945_, _10967_);
  or g_27987_(_10879_, _10956_, _10978_);
  and g_27988_(_10780_, _10967_, _10989_);
  or g_27989_(_10769_, _10978_, _11000_);
  and g_27990_(_20333_, _10571_, _11011_);
  or g_27991_(out[48], _10582_, _11022_);
  and g_27992_(_10637_, _11022_, _11033_);
  or g_27993_(_10648_, _11011_, _11044_);
  and g_27994_(_10087_, _11033_, _11055_);
  or g_27995_(_10098_, _11044_, _11066_);
  and g_27996_(_11000_, _11066_, _11077_);
  or g_27997_(_10989_, _11055_, _11088_);
  and g_27998_(_21840_, _11077_, _11099_);
  not g_27999_(_11099_, _11110_);
  or g_28000_(_26460_, _11077_, _11121_);
  not g_28001_(_11121_, _11132_);
  and g_28002_(_11110_, _11121_, _11143_);
  or g_28003_(_11099_, _11132_, _11154_);
  and g_28004_(_21708_, _11143_, _11165_);
  or g_28005_(_21697_, _11154_, _11176_);
  xor g_28006_(_20531_, _21554_, _11187_);
  xor g_28007_(out[91], _21554_, _11198_);
  and g_28008_(_11165_, _11198_, _11209_);
  or g_28009_(_11176_, _11187_, _11220_);
  or g_28010_(_26350_, _11077_, _11231_);
  not g_28011_(_11231_, _11242_);
  and g_28012_(_26372_, _11077_, _11253_);
  not g_28013_(_11253_, _11264_);
  and g_28014_(_11231_, _11264_, _11275_);
  or g_28015_(_11242_, _11253_, _11286_);
  xor g_28016_(out[74], _21675_, _11297_);
  and g_28017_(_11275_, _11297_, _11308_);
  and g_28018_(_21697_, _11143_, _11319_);
  or g_28019_(_11308_, _11319_, _11330_);
  or g_28020_(_21697_, _11143_, _11341_);
  xor g_28021_(_11275_, _11297_, _11352_);
  xor g_28022_(_11286_, _11297_, _11363_);
  xor g_28023_(_21697_, _11143_, _11374_);
  xor g_28024_(_21708_, _11143_, _11385_);
  and g_28025_(_11352_, _11374_, _11396_);
  or g_28026_(_11363_, _11385_, _11407_);
  xor g_28027_(out[72], _21653_, _11418_);
  xor g_28028_(_20498_, _21653_, _11429_);
  and g_28029_(_26746_, _11077_, _11440_);
  or g_28030_(_26757_, _11088_, _11451_);
  and g_28031_(_26823_, _11088_, _11462_);
  or g_28032_(_26812_, _11077_, _11473_);
  and g_28033_(_11451_, _11473_, _11484_);
  or g_28034_(_11440_, _11462_, _11495_);
  and g_28035_(_11429_, _11495_, _11506_);
  or g_28036_(_11418_, _11484_, _11517_);
  xor g_28037_(out[73], _21664_, _11528_);
  xor g_28038_(_20509_, _21664_, _11539_);
  and g_28039_(_26537_, _11077_, _11550_);
  or g_28040_(_26526_, _11088_, _11561_);
  and g_28041_(_26592_, _11088_, _11572_);
  or g_28042_(_26603_, _11077_, _11583_);
  and g_28043_(_11561_, _11583_, _11594_);
  or g_28044_(_11550_, _11572_, _11605_);
  and g_28045_(_11539_, _11594_, _11616_);
  or g_28046_(_11528_, _11605_, _11627_);
  and g_28047_(_11517_, _11627_, _11638_);
  or g_28048_(_11506_, _11616_, _11649_);
  and g_28049_(_11528_, _11605_, _11660_);
  or g_28050_(_11539_, _11594_, _11671_);
  and g_28051_(_11418_, _11484_, _11682_);
  or g_28052_(_11429_, _11495_, _11693_);
  and g_28053_(_11671_, _11693_, _11704_);
  or g_28054_(_11660_, _11682_, _11715_);
  and g_28055_(_11638_, _11704_, _11726_);
  or g_28056_(_11649_, _11715_, _11737_);
  and g_28057_(_11396_, _11726_, _11748_);
  or g_28058_(_11407_, _11737_, _11759_);
  xor g_28059_(out[70], _21631_, _11770_);
  not g_28060_(_11770_, _11781_);
  and g_28061_(_09416_, _11077_, _11792_);
  not g_28062_(_11792_, _11803_);
  or g_28063_(_09471_, _11077_, _11814_);
  not g_28064_(_11814_, _11825_);
  and g_28065_(_11803_, _11814_, _11836_);
  or g_28066_(_11792_, _11825_, _11847_);
  or g_28067_(_11770_, _11847_, _11858_);
  xor g_28068_(out[71], _21642_, _11869_);
  and g_28069_(_09515_, _11077_, _11880_);
  not g_28070_(_11880_, _11891_);
  or g_28071_(_09581_, _11077_, _11902_);
  not g_28072_(_11902_, _11913_);
  and g_28073_(_11891_, _11902_, _11924_);
  or g_28074_(_11880_, _11913_, _11935_);
  or g_28075_(_11869_, _11924_, _11946_);
  and g_28076_(_11858_, _11946_, _11957_);
  and g_28077_(_11869_, _11924_, _11968_);
  xor g_28078_(_11781_, _11836_, _11979_);
  xor g_28079_(_11770_, _11836_, _11990_);
  xor g_28080_(_11869_, _11924_, _12001_);
  xor g_28081_(_11869_, _11935_, _12012_);
  and g_28082_(_11979_, _12001_, _12023_);
  or g_28083_(_11990_, _12012_, _12034_);
  xor g_28084_(out[69], _21620_, _12045_);
  xor g_28085_(_20432_, _21620_, _12056_);
  and g_28086_(_09856_, _11077_, _12067_);
  not g_28087_(_12067_, _12078_);
  or g_28088_(_09911_, _11077_, _12089_);
  not g_28089_(_12089_, _12100_);
  and g_28090_(_12078_, _12089_, _12111_);
  or g_28091_(_12067_, _12100_, _12122_);
  and g_28092_(_12045_, _12122_, _12133_);
  or g_28093_(_12056_, _12111_, _12144_);
  xor g_28094_(out[68], _21609_, _12155_);
  xor g_28095_(_20443_, _21609_, _12166_);
  and g_28096_(_09735_, _11077_, _12177_);
  not g_28097_(_12177_, _12188_);
  or g_28098_(_09801_, _11077_, _12199_);
  not g_28099_(_12199_, _12210_);
  and g_28100_(_12188_, _12199_, _12221_);
  or g_28101_(_12177_, _12210_, _12232_);
  and g_28102_(_12155_, _12221_, _12243_);
  or g_28103_(_12166_, _12232_, _12254_);
  and g_28104_(_12144_, _12254_, _12265_);
  or g_28105_(_12133_, _12243_, _12276_);
  and g_28106_(_12166_, _12232_, _12287_);
  or g_28107_(_12155_, _12221_, _12298_);
  and g_28108_(_12056_, _12111_, _12309_);
  or g_28109_(_12045_, _12122_, _12320_);
  and g_28110_(_12298_, _12320_, _12331_);
  or g_28111_(_12287_, _12309_, _12342_);
  and g_28112_(_12265_, _12331_, _12353_);
  or g_28113_(_12276_, _12342_, _12364_);
  and g_28114_(_12023_, _12353_, _12375_);
  or g_28115_(_12034_, _12364_, _12386_);
  and g_28116_(_11748_, _12375_, _12397_);
  or g_28117_(_11759_, _12386_, _12408_);
  xor g_28118_(out[67], _21587_, _12419_);
  xor g_28119_(_20487_, _21587_, _12430_);
  or g_28120_(_10175_, _11077_, _12441_);
  not g_28121_(_12441_, _12452_);
  and g_28122_(_10120_, _11077_, _12463_);
  not g_28123_(_12463_, _12474_);
  and g_28124_(_12441_, _12474_, _12485_);
  or g_28125_(_12452_, _12463_, _12496_);
  or g_28126_(_12419_, _12496_, _12507_);
  or g_28127_(out[65], out[66], _12518_);
  xor g_28128_(out[65], out[66], _12529_);
  xor g_28129_(_20454_, out[66], _12540_);
  or g_28130_(_10230_, _11088_, _12551_);
  or g_28131_(_10274_, _11077_, _12562_);
  and g_28132_(_12551_, _12562_, _12573_);
  not g_28133_(_12573_, _12584_);
  and g_28134_(_12540_, _12573_, _12595_);
  and g_28135_(_12419_, _12496_, _12606_);
  xor g_28136_(_12430_, _12485_, _12617_);
  xor g_28137_(_12419_, _12485_, _12628_);
  xor g_28138_(_12540_, _12573_, _12639_);
  xor g_28139_(_12529_, _12573_, _12650_);
  and g_28140_(_12617_, _12639_, _12661_);
  or g_28141_(_12628_, _12650_, _12672_);
  or g_28142_(_20322_, _11088_, _12683_);
  or g_28143_(_10461_, _11077_, _12694_);
  and g_28144_(_12683_, _12694_, _12705_);
  and g_28145_(out[65], _12705_, _12716_);
  or g_28146_(_10571_, _11077_, _12727_);
  not g_28147_(_12727_, _12738_);
  and g_28148_(_20333_, _11077_, _12749_);
  or g_28149_(out[48], _11088_, _12760_);
  and g_28150_(_12727_, _12760_, _12771_);
  or g_28151_(_12738_, _12749_, _12782_);
  and g_28152_(out[64], _12782_, _12793_);
  or g_28153_(_20465_, _12771_, _12804_);
  xor g_28154_(out[65], _12705_, _12815_);
  xor g_28155_(_20454_, _12705_, _12826_);
  and g_28156_(_12804_, _12815_, _12837_);
  or g_28157_(_12793_, _12826_, _12848_);
  or g_28158_(_12716_, _12837_, _12859_);
  and g_28159_(_12661_, _12859_, _12870_);
  or g_28160_(_12595_, _12606_, _12881_);
  and g_28161_(_12507_, _12881_, _12892_);
  or g_28162_(_12870_, _12892_, _12903_);
  and g_28163_(_12397_, _12903_, _12914_);
  and g_28164_(_12023_, _12276_, _12925_);
  or g_28165_(_12034_, _12265_, _12936_);
  and g_28166_(_12320_, _12925_, _12947_);
  or g_28167_(_12309_, _12936_, _12958_);
  or g_28168_(_11957_, _11968_, _12969_);
  not g_28169_(_12969_, _12980_);
  and g_28170_(_12958_, _12969_, _12991_);
  or g_28171_(_12947_, _12980_, _13002_);
  and g_28172_(_11748_, _13002_, _13013_);
  or g_28173_(_11759_, _12991_, _13024_);
  and g_28174_(_11330_, _11341_, _13035_);
  and g_28175_(_11396_, _11715_, _13046_);
  or g_28176_(_11407_, _11704_, _13057_);
  and g_28177_(_11627_, _13046_, _13068_);
  or g_28178_(_11616_, _13057_, _13079_);
  or g_28179_(_12914_, _13035_, _13090_);
  not g_28180_(_13090_, _13101_);
  and g_28181_(_13024_, _13079_, _13112_);
  or g_28182_(_13013_, _13068_, _13123_);
  and g_28183_(_13101_, _13112_, _13134_);
  or g_28184_(_13090_, _13123_, _13145_);
  and g_28185_(_20465_, _12771_, _13156_);
  or g_28186_(out[64], _12782_, _13167_);
  and g_28187_(_12661_, _12837_, _13178_);
  or g_28188_(_12672_, _12848_, _13189_);
  and g_28189_(_13167_, _13178_, _13200_);
  or g_28190_(_13156_, _13189_, _13211_);
  and g_28191_(_12397_, _13200_, _13222_);
  or g_28192_(_12408_, _13211_, _13233_);
  and g_28193_(_13145_, _13233_, _13244_);
  or g_28194_(_13134_, _13222_, _13255_);
  or g_28195_(_11275_, _13244_, _13266_);
  not g_28196_(_13266_, _13277_);
  and g_28197_(_11297_, _13244_, _13288_);
  not g_28198_(_13288_, _13299_);
  and g_28199_(_13266_, _13299_, _13310_);
  or g_28200_(_13277_, _13288_, _13321_);
  and g_28201_(_21565_, _13310_, _13332_);
  or g_28202_(_21576_, _13321_, _13343_);
  and g_28203_(_11220_, _13343_, _13354_);
  or g_28204_(_11209_, _13332_, _13365_);
  and g_28205_(_11176_, _11187_, _13376_);
  or g_28206_(_11165_, _11198_, _13387_);
  and g_28207_(_21576_, _13321_, _13398_);
  or g_28208_(_21565_, _13310_, _13409_);
  and g_28209_(_13387_, _13409_, _13420_);
  or g_28210_(_13376_, _13398_, _13431_);
  xor g_28211_(out[89], _21532_, _13442_);
  xor g_28212_(_20641_, _21532_, _13453_);
  and g_28213_(_11539_, _13244_, _13464_);
  not g_28214_(_13464_, _13475_);
  or g_28215_(_11594_, _13244_, _13486_);
  not g_28216_(_13486_, _13497_);
  and g_28217_(_13475_, _13486_, _13508_);
  or g_28218_(_13464_, _13497_, _13519_);
  and g_28219_(_13453_, _13508_, _13530_);
  or g_28220_(_13442_, _13519_, _13541_);
  and g_28221_(_13354_, _13420_, _13552_);
  or g_28222_(_13365_, _13431_, _13563_);
  and g_28223_(_13541_, _13552_, _13574_);
  or g_28224_(_13530_, _13563_, _13585_);
  xor g_28225_(out[88], _21521_, _13596_);
  xor g_28226_(_20630_, _21521_, _13607_);
  and g_28227_(_11418_, _13244_, _13618_);
  not g_28228_(_13618_, _13629_);
  or g_28229_(_11484_, _13244_, _13640_);
  not g_28230_(_13640_, _13651_);
  and g_28231_(_13629_, _13640_, _13662_);
  or g_28232_(_13618_, _13651_, _13673_);
  and g_28233_(_13607_, _13673_, _13684_);
  or g_28234_(_13596_, _13662_, _13695_);
  and g_28235_(_13442_, _13519_, _13706_);
  or g_28236_(_13453_, _13508_, _13717_);
  and g_28237_(_13596_, _13662_, _13728_);
  or g_28238_(_13607_, _13673_, _13739_);
  and g_28239_(_13717_, _13739_, _13750_);
  or g_28240_(_13706_, _13728_, _13761_);
  and g_28241_(_13695_, _13750_, _13772_);
  or g_28242_(_13684_, _13761_, _13783_);
  and g_28243_(_13574_, _13772_, _13794_);
  or g_28244_(_13585_, _13783_, _13805_);
  xor g_28245_(out[87], _21510_, _13816_);
  xor g_28246_(_20542_, _21510_, _13827_);
  and g_28247_(_11869_, _13244_, _13838_);
  not g_28248_(_13838_, _13849_);
  or g_28249_(_11924_, _13244_, _13860_);
  not g_28250_(_13860_, _13871_);
  and g_28251_(_13849_, _13860_, _13882_);
  or g_28252_(_13838_, _13871_, _13893_);
  and g_28253_(_13816_, _13882_, _13904_);
  or g_28254_(_13827_, _13893_, _13915_);
  and g_28255_(_13827_, _13893_, _13926_);
  or g_28256_(_13816_, _13882_, _13937_);
  xor g_28257_(out[86], _21499_, _13948_);
  xor g_28258_(_20553_, _21499_, _13959_);
  and g_28259_(_11781_, _13244_, _13970_);
  not g_28260_(_13970_, _13981_);
  or g_28261_(_11836_, _13244_, _13992_);
  not g_28262_(_13992_, _14003_);
  and g_28263_(_13981_, _13992_, _14014_);
  or g_28264_(_13970_, _14003_, _14025_);
  and g_28265_(_13959_, _14014_, _14036_);
  or g_28266_(_13948_, _14025_, _14047_);
  and g_28267_(_13937_, _14047_, _14058_);
  or g_28268_(_13926_, _14036_, _14069_);
  and g_28269_(_13915_, _14069_, _14080_);
  or g_28270_(_13904_, _14058_, _14091_);
  and g_28271_(_13948_, _14025_, _14102_);
  or g_28272_(_13959_, _14014_, _14113_);
  and g_28273_(_13915_, _14113_, _14124_);
  or g_28274_(_13904_, _14102_, _14135_);
  and g_28275_(_14058_, _14124_, _14146_);
  or g_28276_(_14069_, _14135_, _14157_);
  xor g_28277_(out[85], _21488_, _14168_);
  xor g_28278_(_20564_, _21488_, _14179_);
  and g_28279_(_12056_, _13244_, _14190_);
  not g_28280_(_14190_, _14201_);
  or g_28281_(_12111_, _13244_, _14212_);
  not g_28282_(_14212_, _14223_);
  and g_28283_(_14201_, _14212_, _14234_);
  or g_28284_(_14190_, _14223_, _14245_);
  and g_28285_(_14179_, _14234_, _14256_);
  or g_28286_(_14168_, _14245_, _14267_);
  and g_28287_(_14146_, _14267_, _14278_);
  or g_28288_(_14157_, _14256_, _14289_);
  and g_28289_(_14168_, _14245_, _14300_);
  or g_28290_(_14179_, _14234_, _14311_);
  xor g_28291_(out[84], _21477_, _14322_);
  xor g_28292_(_20575_, _21477_, _14333_);
  and g_28293_(_12155_, _13244_, _14344_);
  not g_28294_(_14344_, _14355_);
  or g_28295_(_12221_, _13244_, _14366_);
  not g_28296_(_14366_, _14377_);
  and g_28297_(_14355_, _14366_, _14388_);
  or g_28298_(_14344_, _14377_, _14399_);
  and g_28299_(_14322_, _14388_, _14410_);
  or g_28300_(_14333_, _14399_, _14421_);
  and g_28301_(_14311_, _14421_, _14432_);
  or g_28302_(_14300_, _14410_, _14443_);
  xor g_28303_(out[83], _21455_, _14454_);
  xor g_28304_(_20619_, _21455_, _14465_);
  and g_28305_(_12496_, _13255_, _14476_);
  or g_28306_(_12485_, _13244_, _14487_);
  and g_28307_(_12430_, _13244_, _14498_);
  or g_28308_(_12419_, _13255_, _14509_);
  and g_28309_(_14487_, _14509_, _14520_);
  or g_28310_(_14476_, _14498_, _14531_);
  and g_28311_(_14454_, _14531_, _14542_);
  or g_28312_(_14465_, _14520_, _14553_);
  or g_28313_(out[81], out[82], _14564_);
  xor g_28314_(out[81], out[82], _14575_);
  xor g_28315_(_20586_, out[82], _14586_);
  and g_28316_(_12540_, _13244_, _14597_);
  or g_28317_(_12529_, _13255_, _14608_);
  and g_28318_(_12584_, _13255_, _14619_);
  or g_28319_(_12573_, _13244_, _14630_);
  and g_28320_(_14608_, _14630_, _14641_);
  or g_28321_(_14597_, _14619_, _14652_);
  and g_28322_(_14586_, _14641_, _14663_);
  or g_28323_(_14575_, _14652_, _14674_);
  and g_28324_(_14465_, _14520_, _14685_);
  or g_28325_(_14454_, _14531_, _14696_);
  and g_28326_(_14553_, _14674_, _14707_);
  or g_28327_(_14542_, _14663_, _14718_);
  or g_28328_(_14685_, _14707_, _14729_);
  and g_28329_(_14696_, _14718_, _14740_);
  and g_28330_(_14575_, _14652_, _14751_);
  or g_28331_(_14586_, _14641_, _14762_);
  and g_28332_(_14696_, _14762_, _14773_);
  or g_28333_(_14685_, _14751_, _14784_);
  and g_28334_(_14707_, _14773_, _14795_);
  or g_28335_(_14718_, _14784_, _14806_);
  and g_28336_(out[65], _13244_, _14817_);
  not g_28337_(_14817_, _14828_);
  or g_28338_(_12705_, _13244_, _14839_);
  not g_28339_(_14839_, _14850_);
  and g_28340_(_14828_, _14839_, _14861_);
  or g_28341_(_14817_, _14850_, _14872_);
  and g_28342_(out[81], _14861_, _14883_);
  or g_28343_(_20586_, _14872_, _14894_);
  and g_28344_(_20586_, _14872_, _14905_);
  or g_28345_(out[81], _14861_, _14916_);
  and g_28346_(out[64], _13244_, _14927_);
  not g_28347_(_14927_, _14938_);
  and g_28348_(_12771_, _13255_, _14949_);
  or g_28349_(_12782_, _13244_, _14960_);
  or g_28350_(_14927_, _14949_, _14971_);
  and g_28351_(_14938_, _14960_, _14982_);
  and g_28352_(out[80], _14982_, _14993_);
  or g_28353_(_20597_, _14971_, _15004_);
  and g_28354_(_14916_, _15004_, _15015_);
  or g_28355_(_14905_, _14993_, _15026_);
  and g_28356_(_14894_, _15026_, _15037_);
  or g_28357_(_14883_, _15015_, _15048_);
  and g_28358_(_14795_, _15048_, _15059_);
  or g_28359_(_14806_, _15037_, _15070_);
  and g_28360_(_14795_, _14894_, _15081_);
  or g_28361_(_14806_, _14883_, _15092_);
  and g_28362_(_15015_, _15081_, _15103_);
  or g_28363_(_15026_, _15092_, _15114_);
  and g_28364_(_14729_, _15070_, _15125_);
  or g_28365_(_14740_, _15059_, _15136_);
  and g_28366_(_14333_, _14399_, _15147_);
  or g_28367_(_14322_, _14388_, _15158_);
  and g_28368_(_14267_, _15158_, _15169_);
  or g_28369_(_14256_, _15147_, _15180_);
  and g_28370_(_14146_, _15169_, _15191_);
  or g_28371_(_14157_, _15180_, _15202_);
  and g_28372_(_14432_, _15191_, _15213_);
  or g_28373_(_14443_, _15202_, _15224_);
  and g_28374_(_15136_, _15213_, _15235_);
  or g_28375_(_15125_, _15224_, _15246_);
  and g_28376_(_14278_, _14443_, _15257_);
  or g_28377_(_14289_, _14432_, _15268_);
  and g_28378_(_14091_, _15268_, _15279_);
  or g_28379_(_14080_, _15257_, _15290_);
  and g_28380_(_15246_, _15279_, _15301_);
  or g_28381_(_15235_, _15290_, _15312_);
  and g_28382_(_13794_, _15312_, _15323_);
  or g_28383_(_13805_, _15301_, _15334_);
  and g_28384_(_13365_, _13387_, _15345_);
  or g_28385_(_13354_, _13376_, _15356_);
  and g_28386_(_13574_, _13761_, _15367_);
  or g_28387_(_13585_, _13750_, _15378_);
  and g_28388_(_15356_, _15378_, _15389_);
  or g_28389_(_15345_, _15367_, _15400_);
  and g_28390_(_15334_, _15389_, _15411_);
  or g_28391_(_15323_, _15400_, _15422_);
  or g_28392_(out[80], _14982_, _15433_);
  not g_28393_(_15433_, _15444_);
  and g_28394_(_15103_, _15433_, _15455_);
  or g_28395_(_15114_, _15444_, _15466_);
  and g_28396_(_13794_, _15455_, _15477_);
  or g_28397_(_13805_, _15466_, _15488_);
  and g_28398_(_15213_, _15477_, _15499_);
  or g_28399_(_15224_, _15488_, _15510_);
  and g_28400_(_15422_, _15510_, _15521_);
  or g_28401_(_15411_, _15499_, _15532_);
  and g_28402_(_21565_, _15521_, _15543_);
  or g_28403_(_21576_, _15532_, _15554_);
  and g_28404_(_13321_, _15532_, _15565_);
  or g_28405_(_13310_, _15521_, _15576_);
  and g_28406_(_15554_, _15576_, _15587_);
  or g_28407_(_15543_, _15565_, _15598_);
  and g_28408_(out[97], out[98], _15609_);
  or g_28409_(out[100], out[99], _15620_);
  or g_28410_(out[99], _15609_, _15631_);
  or g_28411_(_15609_, _15620_, _15642_);
  or g_28412_(out[101], _15642_, _15653_);
  and g_28413_(out[102], _15653_, _15664_);
  and g_28414_(out[103], _15664_, _15675_);
  or g_28415_(out[104], _15675_, _15686_);
  or g_28416_(out[105], _15686_, _15697_);
  or g_28417_(out[106], _15697_, _15708_);
  xor g_28418_(out[106], _15697_, _15719_);
  xor g_28419_(_20784_, _15697_, _15730_);
  and g_28420_(_15587_, _15719_, _15741_);
  or g_28421_(_15598_, _15730_, _15752_);
  and g_28422_(_11165_, _11187_, _15763_);
  or g_28423_(_11176_, _11198_, _15774_);
  xor g_28424_(_20663_, _15708_, _15785_);
  xor g_28425_(out[107], _15708_, _15796_);
  and g_28426_(_15763_, _15796_, _15807_);
  or g_28427_(_15774_, _15785_, _15818_);
  and g_28428_(_15752_, _15818_, _15829_);
  or g_28429_(_15741_, _15807_, _15840_);
  and g_28430_(_15774_, _15785_, _15851_);
  or g_28431_(_15763_, _15796_, _15862_);
  and g_28432_(_15598_, _15730_, _15873_);
  or g_28433_(_15587_, _15719_, _15884_);
  and g_28434_(_15862_, _15884_, _15895_);
  or g_28435_(_15851_, _15873_, _15906_);
  and g_28436_(_15829_, _15895_, _15917_);
  or g_28437_(_15840_, _15906_, _15928_);
  xor g_28438_(out[105], _15686_, _15939_);
  xor g_28439_(_20773_, _15686_, _15950_);
  or g_28440_(_13508_, _15521_, _15961_);
  or g_28441_(_13442_, _15532_, _15972_);
  and g_28442_(_15961_, _15972_, _15983_);
  not g_28443_(_15983_, _15994_);
  or g_28444_(_15950_, _15983_, _16005_);
  not g_28445_(_16005_, _16016_);
  xor g_28446_(out[104], _15675_, _16027_);
  or g_28447_(_13662_, _15521_, _16038_);
  or g_28448_(_13607_, _15532_, _16049_);
  and g_28449_(_16038_, _16049_, _16060_);
  and g_28450_(_16027_, _16060_, _16071_);
  not g_28451_(_16071_, _16082_);
  and g_28452_(_16005_, _16082_, _16093_);
  or g_28453_(_16016_, _16071_, _16104_);
  and g_28454_(_15950_, _15983_, _16115_);
  or g_28455_(_15939_, _15994_, _16126_);
  or g_28456_(_16027_, _16060_, _16137_);
  not g_28457_(_16137_, _16148_);
  and g_28458_(_16126_, _16137_, _16159_);
  or g_28459_(_16115_, _16148_, _16170_);
  and g_28460_(_16093_, _16159_, _16181_);
  or g_28461_(_16104_, _16170_, _16192_);
  and g_28462_(_15917_, _16181_, _16203_);
  or g_28463_(_15928_, _16192_, _16214_);
  xor g_28464_(out[103], _15664_, _16225_);
  not g_28465_(_16225_, _16236_);
  or g_28466_(_13882_, _15521_, _16247_);
  or g_28467_(_13827_, _15532_, _16258_);
  and g_28468_(_16247_, _16258_, _16269_);
  not g_28469_(_16269_, _16280_);
  and g_28470_(_16236_, _16280_, _16291_);
  or g_28471_(_16225_, _16269_, _16302_);
  xor g_28472_(out[102], _15653_, _16313_);
  xor g_28473_(_20685_, _15653_, _16324_);
  or g_28474_(_14014_, _15521_, _16335_);
  or g_28475_(_13948_, _15532_, _16346_);
  and g_28476_(_16335_, _16346_, _16357_);
  not g_28477_(_16357_, _16368_);
  and g_28478_(_16324_, _16357_, _16379_);
  or g_28479_(_16313_, _16368_, _16390_);
  and g_28480_(_16302_, _16390_, _16401_);
  or g_28481_(_16291_, _16379_, _16412_);
  and g_28482_(_16225_, _16269_, _16423_);
  or g_28483_(_16236_, _16280_, _16434_);
  or g_28484_(_16324_, _16357_, _16445_);
  or g_28485_(_16379_, _16423_, _16456_);
  not g_28486_(_16456_, _16467_);
  and g_28487_(_16302_, _16445_, _16478_);
  not g_28488_(_16478_, _16489_);
  and g_28489_(_16467_, _16478_, _16500_);
  or g_28490_(_16456_, _16489_, _16511_);
  xor g_28491_(out[100], _15631_, _16522_);
  or g_28492_(_14333_, _15532_, _16533_);
  or g_28493_(_14388_, _15521_, _16544_);
  and g_28494_(_16533_, _16544_, _16555_);
  and g_28495_(_16522_, _16555_, _16566_);
  not g_28496_(_16566_, _16577_);
  or g_28497_(_16522_, _16555_, _16588_);
  xor g_28498_(out[101], _15642_, _16599_);
  xor g_28499_(_20696_, _15642_, _16610_);
  or g_28500_(_14234_, _15521_, _16621_);
  or g_28501_(_14168_, _15532_, _16632_);
  and g_28502_(_16621_, _16632_, _16643_);
  not g_28503_(_16643_, _16654_);
  and g_28504_(_16610_, _16643_, _16665_);
  or g_28505_(_16599_, _16654_, _16676_);
  or g_28506_(_16610_, _16643_, _16687_);
  not g_28507_(_16687_, _16698_);
  and g_28508_(_16577_, _16687_, _16709_);
  or g_28509_(_16566_, _16698_, _16720_);
  and g_28510_(_16588_, _16676_, _16731_);
  and g_28511_(_16709_, _16731_, _16742_);
  not g_28512_(_16742_, _16753_);
  and g_28513_(_16500_, _16742_, _16764_);
  or g_28514_(_16511_, _16753_, _16775_);
  and g_28515_(_16203_, _16764_, _16786_);
  or g_28516_(_16214_, _16775_, _16797_);
  or g_28517_(_20586_, _15532_, _16808_);
  or g_28518_(_14861_, _15521_, _16819_);
  and g_28519_(_16808_, _16819_, _16830_);
  and g_28520_(out[97], _16830_, _16841_);
  xor g_28521_(out[99], _15609_, _16852_);
  xor g_28522_(_20751_, _15609_, _16863_);
  or g_28523_(_14520_, _15521_, _16874_);
  or g_28524_(_14454_, _15532_, _16885_);
  and g_28525_(_16874_, _16885_, _16896_);
  or g_28526_(_16863_, _16896_, _16907_);
  and g_28527_(_16863_, _16896_, _16918_);
  xor g_28528_(_16863_, _16896_, _16929_);
  xor g_28529_(_16852_, _16896_, _16940_);
  or g_28530_(_14575_, _15532_, _16951_);
  or g_28531_(_14641_, _15521_, _16962_);
  and g_28532_(_16951_, _16962_, _16973_);
  or g_28533_(out[97], out[98], _16984_);
  xor g_28534_(out[97], out[98], _16995_);
  xor g_28535_(_20718_, out[98], _17006_);
  and g_28536_(_16973_, _17006_, _17017_);
  not g_28537_(_17017_, _17028_);
  xor g_28538_(_16973_, _17006_, _17039_);
  xor g_28539_(_16973_, _16995_, _17050_);
  and g_28540_(_16929_, _17039_, _17061_);
  or g_28541_(_16940_, _17050_, _17072_);
  and g_28542_(_16841_, _17061_, _17083_);
  not g_28543_(_17083_, _17094_);
  and g_28544_(_14982_, _15532_, _17105_);
  not g_28545_(_17105_, _17116_);
  or g_28546_(out[80], _15532_, _17127_);
  not g_28547_(_17127_, _17138_);
  and g_28548_(_17116_, _17127_, _17149_);
  or g_28549_(_17105_, _17138_, _17160_);
  and g_28550_(out[96], _17160_, _17171_);
  or g_28551_(_20729_, _17149_, _17182_);
  xor g_28552_(out[97], _16830_, _17193_);
  xor g_28553_(_20718_, _16830_, _17204_);
  and g_28554_(_17061_, _17182_, _17215_);
  or g_28555_(_17072_, _17171_, _17226_);
  and g_28556_(_17193_, _17215_, _17237_);
  or g_28557_(_17204_, _17226_, _17248_);
  and g_28558_(_16907_, _17028_, _17259_);
  or g_28559_(_16918_, _17259_, _17270_);
  not g_28560_(_17270_, _17281_);
  and g_28561_(_17248_, _17270_, _17292_);
  or g_28562_(_17237_, _17281_, _17303_);
  and g_28563_(_17094_, _17292_, _17314_);
  or g_28564_(_17083_, _17303_, _17325_);
  and g_28565_(_16786_, _17325_, _17336_);
  or g_28566_(_16797_, _17314_, _17347_);
  and g_28567_(_16676_, _16720_, _17358_);
  or g_28568_(_16665_, _16709_, _17369_);
  and g_28569_(_16500_, _17358_, _17380_);
  or g_28570_(_16511_, _17369_, _17391_);
  and g_28571_(_16412_, _16434_, _17402_);
  or g_28572_(_16401_, _16423_, _17413_);
  and g_28573_(_17391_, _17413_, _17424_);
  or g_28574_(_17380_, _17402_, _17435_);
  and g_28575_(_16203_, _17435_, _17446_);
  or g_28576_(_16214_, _17424_, _17457_);
  and g_28577_(_15840_, _15862_, _17468_);
  or g_28578_(_15829_, _15851_, _17479_);
  and g_28579_(_15917_, _16104_, _17490_);
  or g_28580_(_15928_, _16093_, _17501_);
  and g_28581_(_16126_, _17490_, _17512_);
  or g_28582_(_16115_, _17501_, _17523_);
  and g_28583_(_17479_, _17523_, _17534_);
  or g_28584_(_17468_, _17512_, _17545_);
  and g_28585_(_17457_, _17534_, _17556_);
  or g_28586_(_17446_, _17545_, _17567_);
  and g_28587_(_17347_, _17556_, _17578_);
  or g_28588_(_17336_, _17567_, _17589_);
  or g_28589_(out[96], _17160_, _17600_);
  and g_28590_(_17237_, _17600_, _17611_);
  and g_28591_(_16786_, _17611_, _17622_);
  not g_28592_(_17622_, _17633_);
  and g_28593_(_17589_, _17633_, _17644_);
  or g_28594_(_17578_, _17622_, _17655_);
  and g_28595_(_15598_, _17655_, _17666_);
  or g_28596_(_15587_, _17644_, _17677_);
  and g_28597_(_15719_, _17644_, _17688_);
  or g_28598_(_15730_, _17655_, _17699_);
  and g_28599_(_17677_, _17699_, _17710_);
  or g_28600_(_17666_, _17688_, _17721_);
  and g_28601_(out[113], out[114], _17732_);
  or g_28602_(out[116], out[115], _17743_);
  or g_28603_(out[115], _17732_, _17754_);
  or g_28604_(_17732_, _17743_, _17765_);
  or g_28605_(out[117], _17765_, _17776_);
  and g_28606_(out[118], _17776_, _17787_);
  and g_28607_(out[119], _17787_, _17798_);
  or g_28608_(out[120], _17798_, _17809_);
  or g_28609_(out[121], _17809_, _17820_);
  or g_28610_(out[122], _17820_, _17831_);
  xor g_28611_(out[122], _17820_, _17842_);
  xor g_28612_(_20905_, _17820_, _17853_);
  and g_28613_(_17710_, _17842_, _17862_);
  or g_28614_(_17721_, _17853_, _17863_);
  and g_28615_(_15763_, _15785_, _17864_);
  or g_28616_(_15774_, _15796_, _17865_);
  xor g_28617_(_20795_, _17831_, _17866_);
  xor g_28618_(out[123], _17831_, _17867_);
  and g_28619_(_17864_, _17867_, _17868_);
  or g_28620_(_17865_, _17866_, _17869_);
  and g_28621_(_17863_, _17869_, _17870_);
  or g_28622_(_17862_, _17868_, _17871_);
  and g_28623_(_17721_, _17853_, _17872_);
  or g_28624_(_17710_, _17842_, _17873_);
  and g_28625_(_17865_, _17866_, _17874_);
  or g_28626_(_17864_, _17867_, _17875_);
  and g_28627_(_17873_, _17875_, _17876_);
  or g_28628_(_17872_, _17874_, _17877_);
  and g_28629_(_17870_, _17876_, _17878_);
  or g_28630_(_17871_, _17877_, _17879_);
  xor g_28631_(out[121], _17809_, _17880_);
  xor g_28632_(_20894_, _17809_, _17881_);
  and g_28633_(_15950_, _17644_, _17882_);
  not g_28634_(_17882_, _17883_);
  or g_28635_(_15983_, _17644_, _17884_);
  not g_28636_(_17884_, _17885_);
  and g_28637_(_17883_, _17884_, _17886_);
  or g_28638_(_17882_, _17885_, _17887_);
  and g_28639_(_17880_, _17887_, _17888_);
  or g_28640_(_17881_, _17886_, _17889_);
  xor g_28641_(out[120], _17798_, _17890_);
  xor g_28642_(_20883_, _17798_, _17891_);
  and g_28643_(_16027_, _17644_, _17892_);
  not g_28644_(_17892_, _17893_);
  or g_28645_(_16060_, _17644_, _17894_);
  not g_28646_(_17894_, _17895_);
  and g_28647_(_17893_, _17894_, _17896_);
  or g_28648_(_17892_, _17895_, _17897_);
  and g_28649_(_17890_, _17896_, _17898_);
  or g_28650_(_17891_, _17897_, _17899_);
  and g_28651_(_17889_, _17899_, _17900_);
  or g_28652_(_17888_, _17898_, _17901_);
  and g_28653_(_17881_, _17886_, _17902_);
  or g_28654_(_17880_, _17887_, _17903_);
  and g_28655_(_17891_, _17897_, _17904_);
  or g_28656_(_17890_, _17896_, _17905_);
  and g_28657_(_17903_, _17905_, _17906_);
  or g_28658_(_17902_, _17904_, _17907_);
  and g_28659_(_17878_, _17906_, _17908_);
  or g_28660_(_17879_, _17907_, _17909_);
  and g_28661_(_17900_, _17908_, _17910_);
  or g_28662_(_17901_, _17909_, _17911_);
  xor g_28663_(out[116], _17754_, _17912_);
  not g_28664_(_17912_, _17913_);
  and g_28665_(_16522_, _17644_, _17914_);
  not g_28666_(_17914_, _17915_);
  or g_28667_(_16555_, _17644_, _17916_);
  not g_28668_(_17916_, _17917_);
  and g_28669_(_17915_, _17916_, _17918_);
  or g_28670_(_17914_, _17917_, _17919_);
  or g_28671_(_17913_, _17919_, _17920_);
  not g_28672_(_17920_, _17921_);
  xor g_28673_(out[117], _17765_, _17922_);
  xor g_28674_(_20828_, _17765_, _17923_);
  and g_28675_(_16610_, _17644_, _17924_);
  not g_28676_(_17924_, _17925_);
  or g_28677_(_16643_, _17644_, _17926_);
  not g_28678_(_17926_, _17927_);
  and g_28679_(_17925_, _17926_, _17928_);
  or g_28680_(_17924_, _17927_, _17929_);
  and g_28681_(_17922_, _17929_, _17930_);
  or g_28682_(_17923_, _17928_, _17931_);
  and g_28683_(_17920_, _17931_, _17932_);
  or g_28684_(_17921_, _17930_, _17933_);
  xor g_28685_(out[119], _17787_, _17934_);
  xor g_28686_(_20806_, _17787_, _17935_);
  and g_28687_(_16225_, _17644_, _17936_);
  not g_28688_(_17936_, _17937_);
  or g_28689_(_16269_, _17644_, _17938_);
  not g_28690_(_17938_, _17939_);
  and g_28691_(_17937_, _17938_, _17940_);
  or g_28692_(_17936_, _17939_, _17941_);
  and g_28693_(_17934_, _17940_, _17942_);
  or g_28694_(_17935_, _17941_, _17943_);
  or g_28695_(_17912_, _17918_, _17944_);
  and g_28696_(_17943_, _17944_, _17945_);
  and g_28697_(_17932_, _17945_, _17946_);
  xor g_28698_(out[118], _17776_, _17947_);
  xor g_28699_(_20817_, _17776_, _17948_);
  and g_28700_(_16324_, _17644_, _17949_);
  not g_28701_(_17949_, _17950_);
  or g_28702_(_16357_, _17644_, _17951_);
  not g_28703_(_17951_, _17952_);
  and g_28704_(_17950_, _17951_, _17953_);
  or g_28705_(_17949_, _17952_, _17954_);
  and g_28706_(_17948_, _17953_, _17955_);
  or g_28707_(_17947_, _17954_, _17956_);
  and g_28708_(_17935_, _17941_, _17957_);
  or g_28709_(_17934_, _17940_, _17958_);
  and g_28710_(_17956_, _17958_, _17959_);
  or g_28711_(_17955_, _17957_, _17960_);
  and g_28712_(_17947_, _17954_, _17961_);
  or g_28713_(_17948_, _17953_, _17962_);
  and g_28714_(_17923_, _17928_, _17963_);
  or g_28715_(_17922_, _17929_, _17964_);
  and g_28716_(_17962_, _17964_, _17965_);
  or g_28717_(_17961_, _17963_, _17966_);
  and g_28718_(_17959_, _17965_, _17967_);
  and g_28719_(_17946_, _17967_, _17968_);
  and g_28720_(_17910_, _17968_, _17969_);
  not g_28721_(_17969_, _17970_);
  xor g_28722_(out[115], _17732_, _17971_);
  xor g_28723_(_20872_, _17732_, _17972_);
  or g_28724_(_16896_, _17644_, _17973_);
  not g_28725_(_17973_, _17974_);
  and g_28726_(_16863_, _17644_, _17975_);
  not g_28727_(_17975_, _17976_);
  and g_28728_(_17973_, _17976_, _17977_);
  or g_28729_(_17974_, _17975_, _17978_);
  and g_28730_(_17971_, _17978_, _17979_);
  or g_28731_(_17972_, _17977_, _17980_);
  or g_28732_(_16973_, _17644_, _17981_);
  not g_28733_(_17981_, _17982_);
  and g_28734_(_17006_, _17644_, _17983_);
  not g_28735_(_17983_, _17984_);
  and g_28736_(_17981_, _17984_, _17985_);
  or g_28737_(_17982_, _17983_, _17986_);
  or g_28738_(out[113], out[114], _17987_);
  xor g_28739_(out[113], out[114], _17988_);
  xor g_28740_(_20850_, out[114], _17989_);
  and g_28741_(_17985_, _17989_, _17990_);
  or g_28742_(_17986_, _17988_, _17991_);
  and g_28743_(_17972_, _17977_, _17992_);
  or g_28744_(_17971_, _17978_, _17993_);
  xor g_28745_(_17986_, _17988_, _17994_);
  xor g_28746_(_17985_, _17988_, _17995_);
  and g_28747_(_17980_, _17993_, _17996_);
  or g_28748_(_17979_, _17992_, _17997_);
  and g_28749_(_17994_, _17996_, _17998_);
  or g_28750_(_17995_, _17997_, _17999_);
  and g_28751_(out[97], _17644_, _18000_);
  not g_28752_(_18000_, _18001_);
  or g_28753_(_16830_, _17644_, _18002_);
  not g_28754_(_18002_, _18003_);
  and g_28755_(_18001_, _18002_, _18004_);
  or g_28756_(_18000_, _18003_, _18005_);
  and g_28757_(out[113], _18004_, _18006_);
  or g_28758_(_20850_, _18005_, _18007_);
  and g_28759_(out[96], _17644_, _18008_);
  not g_28760_(_18008_, _18009_);
  and g_28761_(_17149_, _17655_, _18010_);
  or g_28762_(_17160_, _17644_, _18011_);
  or g_28763_(_18008_, _18010_, _18012_);
  and g_28764_(_18009_, _18011_, _18013_);
  and g_28765_(out[112], _18013_, _18014_);
  or g_28766_(_19860_, _18012_, _18015_);
  xor g_28767_(out[113], _18004_, _18016_);
  xor g_28768_(_20850_, _18004_, _18017_);
  and g_28769_(_18015_, _18016_, _18018_);
  or g_28770_(_18014_, _18017_, _18019_);
  and g_28771_(_18007_, _18019_, _18020_);
  or g_28772_(_18006_, _18018_, _18021_);
  and g_28773_(_17998_, _18021_, _18022_);
  or g_28774_(_17999_, _18020_, _18023_);
  and g_28775_(_17990_, _17993_, _18024_);
  or g_28776_(_17991_, _17992_, _18025_);
  and g_28777_(_17980_, _18025_, _18026_);
  or g_28778_(_17979_, _18024_, _18027_);
  and g_28779_(_18023_, _18026_, _18028_);
  or g_28780_(_18022_, _18027_, _18029_);
  and g_28781_(_17969_, _18029_, _18030_);
  or g_28782_(_17970_, _18028_, _18031_);
  and g_28783_(_17933_, _17965_, _18032_);
  or g_28784_(_17932_, _17966_, _18033_);
  and g_28785_(_17959_, _18033_, _18034_);
  or g_28786_(_17960_, _18032_, _18035_);
  and g_28787_(_17910_, _17943_, _18036_);
  or g_28788_(_17911_, _17942_, _18037_);
  and g_28789_(_18035_, _18036_, _18038_);
  or g_28790_(_18034_, _18037_, _18039_);
  and g_28791_(_17878_, _17901_, _18040_);
  or g_28792_(_17879_, _17900_, _18041_);
  and g_28793_(_17903_, _18040_, _18042_);
  or g_28794_(_17902_, _18041_, _18043_);
  and g_28795_(_17871_, _17875_, _18044_);
  or g_28796_(_17870_, _17874_, _18045_);
  and g_28797_(_18043_, _18045_, _18046_);
  or g_28798_(_18042_, _18044_, _18047_);
  and g_28799_(_18039_, _18046_, _18048_);
  or g_28800_(_18038_, _18047_, _18049_);
  and g_28801_(_18031_, _18048_, _18050_);
  or g_28802_(_18030_, _18049_, _18051_);
  or g_28803_(out[112], _18013_, _18052_);
  or g_28804_(_17999_, _18019_, _18053_);
  not g_28805_(_18053_, _18054_);
  and g_28806_(_17969_, _18052_, _18055_);
  not g_28807_(_18055_, _18056_);
  and g_28808_(_18054_, _18055_, _18057_);
  or g_28809_(_18053_, _18056_, _18058_);
  and g_28810_(_18051_, _18058_, _18059_);
  or g_28811_(_18050_, _18057_, _18060_);
  or g_28812_(_17710_, _18059_, _18061_);
  not g_28813_(_18061_, _18062_);
  and g_28814_(_17842_, _18059_, _18063_);
  not g_28815_(_18063_, _18064_);
  and g_28816_(_18061_, _18064_, _18065_);
  or g_28817_(_18062_, _18063_, _18066_);
  and g_28818_(_21444_, _18065_, _18067_);
  and g_28819_(_17864_, _17866_, _18068_);
  or g_28820_(_17865_, _17867_, _18069_);
  xor g_28821_(_20916_, _21433_, _18070_);
  xor g_28822_(out[139], _21433_, _18071_);
  and g_28823_(_18068_, _18071_, _18072_);
  or g_28824_(_18067_, _18072_, _18073_);
  not g_28825_(_18073_, _18074_);
  or g_28826_(_18068_, _18071_, _18075_);
  or g_28827_(_21444_, _18065_, _18076_);
  and g_28828_(_18075_, _18076_, _18077_);
  not g_28829_(_18077_, _18078_);
  and g_28830_(_18074_, _18077_, _18079_);
  or g_28831_(_18073_, _18078_, _18080_);
  xor g_28832_(out[135], _21389_, _18081_);
  not g_28833_(_18081_, _18082_);
  and g_28834_(_17934_, _18059_, _18083_);
  not g_28835_(_18083_, _18084_);
  or g_28836_(_17940_, _18059_, _18085_);
  not g_28837_(_18085_, _18086_);
  and g_28838_(_18084_, _18085_, _18087_);
  or g_28839_(_18083_, _18086_, _18088_);
  or g_28840_(_18082_, _18088_, _18089_);
  xor g_28841_(out[134], _21378_, _18090_);
  not g_28842_(_18090_, _18091_);
  and g_28843_(_17948_, _18059_, _18092_);
  or g_28844_(_17947_, _18060_, _18093_);
  or g_28845_(_17953_, _18059_, _18094_);
  not g_28846_(_18094_, _18095_);
  and g_28847_(_18093_, _18094_, _18096_);
  or g_28848_(_18092_, _18095_, _18097_);
  and g_28849_(_18091_, _18096_, _18098_);
  and g_28850_(_18082_, _18088_, _18099_);
  or g_28851_(_18098_, _18099_, _18100_);
  and g_28852_(_18089_, _18100_, _18101_);
  xor g_28853_(out[133], _21367_, _18102_);
  and g_28854_(_17923_, _18059_, _18103_);
  and g_28855_(_17929_, _18060_, _18104_);
  or g_28856_(_18103_, _18104_, _18105_);
  or g_28857_(_18102_, _18105_, _18106_);
  and g_28858_(_18090_, _18097_, _18107_);
  and g_28859_(_18089_, _18106_, _18108_);
  not g_28860_(_18108_, _18109_);
  or g_28861_(_18100_, _18107_, _18110_);
  not g_28862_(_18110_, _18111_);
  and g_28863_(_18108_, _18111_, _18112_);
  or g_28864_(_18109_, _18110_, _18113_);
  xor g_28865_(out[132], _21356_, _18114_);
  not g_28866_(_18114_, _18115_);
  and g_28867_(_17912_, _18059_, _18116_);
  and g_28868_(_17919_, _18060_, _18117_);
  or g_28869_(_18116_, _18117_, _18118_);
  not g_28870_(_18118_, _18119_);
  and g_28871_(_18114_, _18119_, _18120_);
  and g_28872_(_18102_, _18105_, _18121_);
  or g_28873_(_18120_, _18121_, _18122_);
  or g_28874_(_17985_, _18059_, _18123_);
  or g_28875_(_17988_, _18060_, _18124_);
  and g_28876_(_18123_, _18124_, _18125_);
  or g_28877_(out[129], out[130], _18126_);
  xor g_28878_(out[129], out[130], _18127_);
  xor g_28879_(_20971_, out[130], _18128_);
  and g_28880_(_18125_, _18128_, _18129_);
  xor g_28881_(out[131], _21334_, _18130_);
  and g_28882_(_17978_, _18060_, _18131_);
  and g_28883_(_17972_, _18059_, _18132_);
  or g_28884_(_18131_, _18132_, _18133_);
  and g_28885_(_18130_, _18133_, _18134_);
  or g_28886_(_18129_, _18134_, _18135_);
  or g_28887_(_18130_, _18133_, _18136_);
  xor g_28888_(_18125_, _18128_, _18137_);
  xor g_28889_(_18130_, _18133_, _18138_);
  and g_28890_(_18137_, _18138_, _18139_);
  not g_28891_(_18139_, _18140_);
  and g_28892_(out[113], _18059_, _18141_);
  not g_28893_(_18141_, _18142_);
  or g_28894_(_18004_, _18059_, _18143_);
  not g_28895_(_18143_, _18144_);
  and g_28896_(_18142_, _18143_, _18145_);
  or g_28897_(_18141_, _18144_, _18146_);
  and g_28898_(_20971_, _18146_, _18147_);
  and g_28899_(out[129], _18145_, _18148_);
  or g_28900_(_18012_, _18059_, _18149_);
  or g_28901_(out[112], _18060_, _18150_);
  and g_28902_(_18149_, _18150_, _18151_);
  not g_28903_(_18151_, _18152_);
  and g_28904_(out[128], _18152_, _18153_);
  or g_28905_(_20982_, _18151_, _18154_);
  or g_28906_(_18148_, _18153_, _18155_);
  or g_28907_(_18147_, _18155_, _18156_);
  xor g_28908_(out[129], _18145_, _18157_);
  and g_28909_(_18139_, _18154_, _18158_);
  and g_28910_(_18157_, _18158_, _18159_);
  or g_28911_(_18140_, _18156_, _18160_);
  and g_28912_(_18139_, _18148_, _18161_);
  and g_28913_(_18135_, _18136_, _18162_);
  or g_28914_(_18161_, _18162_, _18163_);
  or g_28915_(_18159_, _18163_, _18164_);
  and g_28916_(_18115_, _18118_, _18165_);
  or g_28917_(_18114_, _18119_, _18166_);
  and g_28918_(_18164_, _18166_, _18167_);
  or g_28919_(_18122_, _18167_, _18168_);
  and g_28920_(_18112_, _18168_, _18169_);
  or g_28921_(_18101_, _18169_, _18170_);
  xor g_28922_(out[137], _21411_, _18171_);
  or g_28923_(_17880_, _18060_, _18172_);
  or g_28924_(_17886_, _18059_, _18173_);
  and g_28925_(_18172_, _18173_, _18174_);
  not g_28926_(_18174_, _18175_);
  or g_28927_(_18171_, _18175_, _18176_);
  not g_28928_(_18176_, _18177_);
  xor g_28929_(out[136], _21400_, _18178_);
  not g_28930_(_18178_, _18179_);
  and g_28931_(_17890_, _18059_, _18180_);
  not g_28932_(_18180_, _18181_);
  or g_28933_(_17896_, _18059_, _18182_);
  not g_28934_(_18182_, _18183_);
  and g_28935_(_18181_, _18182_, _18184_);
  or g_28936_(_18180_, _18183_, _18185_);
  and g_28937_(_18178_, _18184_, _18186_);
  not g_28938_(_18186_, _18187_);
  and g_28939_(_18176_, _18187_, _18188_);
  or g_28940_(_18177_, _18186_, _18189_);
  and g_28941_(_18171_, _18175_, _18190_);
  not g_28942_(_18190_, _18191_);
  and g_28943_(_18179_, _18185_, _18192_);
  or g_28944_(_18178_, _18184_, _18193_);
  and g_28945_(_18191_, _18193_, _18194_);
  or g_28946_(_18190_, _18192_, _18195_);
  and g_28947_(_18188_, _18194_, _18196_);
  or g_28948_(_18189_, _18195_, _18197_);
  and g_28949_(_18170_, _18196_, _18198_);
  or g_28950_(_18186_, _18190_, _18199_);
  and g_28951_(_18176_, _18199_, _18200_);
  or g_28952_(_18198_, _18200_, _18201_);
  and g_28953_(_18079_, _18201_, _18202_);
  and g_28954_(_18073_, _18075_, _18203_);
  or g_28955_(_18202_, _18203_, _18204_);
  and g_28956_(_20982_, _18151_, _18205_);
  or g_28957_(_18165_, _18205_, _18206_);
  or g_28958_(_18122_, _18206_, _18207_);
  or g_28959_(_18080_, _18207_, _18208_);
  or g_28960_(_18197_, _18208_, _18209_);
  or g_28961_(_18113_, _18160_, _18210_);
  or g_28962_(_18209_, _18210_, _18211_);
  and g_28963_(_18204_, _18211_, _18212_);
  not g_28964_(_18212_, _18213_);
  and g_28965_(_21444_, _18212_, _18214_);
  not g_28966_(_18214_, _18215_);
  and g_28967_(_18066_, _18213_, _18216_);
  or g_28968_(_18065_, _18212_, _18217_);
  and g_28969_(_18215_, _18217_, _18218_);
  or g_28970_(_18214_, _18216_, _18219_);
  and g_28971_(_21312_, _18218_, _18220_);
  or g_28972_(_21323_, _18219_, _18221_);
  and g_28973_(_18068_, _18070_, _18222_);
  or g_28974_(_18069_, _18071_, _18223_);
  xor g_28975_(_21048_, _21301_, _18224_);
  xor g_28976_(out[155], _21301_, _18225_);
  and g_28977_(_18222_, _18225_, _18226_);
  or g_28978_(_18223_, _18224_, _18227_);
  and g_28979_(_18221_, _18227_, _18228_);
  or g_28980_(_18220_, _18226_, _18229_);
  and g_28981_(_18223_, _18224_, _18230_);
  or g_28982_(_18222_, _18225_, _18231_);
  and g_28983_(_21323_, _18219_, _18232_);
  or g_28984_(_21312_, _18218_, _18233_);
  and g_28985_(_18231_, _18233_, _18234_);
  or g_28986_(_18230_, _18232_, _18235_);
  or g_28987_(_18174_, _18212_, _18236_);
  or g_28988_(_18171_, _18213_, _18237_);
  and g_28989_(_18236_, _18237_, _18238_);
  not g_28990_(_18238_, _18239_);
  and g_28991_(_21290_, _18238_, _18240_);
  or g_28992_(_21279_, _18239_, _18241_);
  and g_28993_(_18228_, _18234_, _18242_);
  or g_28994_(_18229_, _18235_, _18243_);
  and g_28995_(_18241_, _18242_, _18244_);
  or g_28996_(_18240_, _18243_, _18245_);
  xor g_28997_(out[152], _21246_, _18246_);
  xor g_28998_(_21147_, _21246_, _18247_);
  and g_28999_(_18185_, _18213_, _18248_);
  or g_29000_(_18184_, _18212_, _18249_);
  and g_29001_(_18178_, _18212_, _18250_);
  not g_29002_(_18250_, _18251_);
  and g_29003_(_18249_, _18251_, _18252_);
  or g_29004_(_18248_, _18250_, _18253_);
  and g_29005_(_18247_, _18253_, _18254_);
  or g_29006_(_18246_, _18252_, _18255_);
  and g_29007_(_21279_, _18239_, _18256_);
  or g_29008_(_21290_, _18238_, _18257_);
  and g_29009_(_18246_, _18252_, _18258_);
  or g_29010_(_18247_, _18253_, _18259_);
  and g_29011_(_18257_, _18259_, _18260_);
  or g_29012_(_18256_, _18258_, _18261_);
  and g_29013_(_18255_, _18260_, _18262_);
  or g_29014_(_18254_, _18261_, _18263_);
  and g_29015_(_18244_, _18262_, _18264_);
  or g_29016_(_18245_, _18263_, _18265_);
  xor g_29017_(out[150], _21224_, _18266_);
  and g_29018_(_18096_, _18213_, _18267_);
  or g_29019_(_18097_, _18212_, _18268_);
  and g_29020_(_18090_, _18212_, _18269_);
  not g_29021_(_18269_, _18270_);
  or g_29022_(_18267_, _18269_, _18271_);
  and g_29023_(_18268_, _18270_, _18272_);
  or g_29024_(_18266_, _18272_, _18273_);
  xor g_29025_(out[151], _21235_, _18274_);
  not g_29026_(_18274_, _18275_);
  and g_29027_(_18088_, _18213_, _18276_);
  or g_29028_(_18087_, _18212_, _18277_);
  and g_29029_(_18081_, _18212_, _18278_);
  not g_29030_(_18278_, _18279_);
  and g_29031_(_18277_, _18279_, _18280_);
  or g_29032_(_18276_, _18278_, _18281_);
  or g_29033_(_18274_, _18280_, _18282_);
  and g_29034_(_18273_, _18282_, _18283_);
  and g_29035_(_18274_, _18280_, _18284_);
  xor g_29036_(_18266_, _18272_, _18285_);
  xor g_29037_(_18266_, _18271_, _18286_);
  xor g_29038_(_18274_, _18280_, _18287_);
  xor g_29039_(_18275_, _18280_, _18288_);
  and g_29040_(_18285_, _18287_, _18289_);
  or g_29041_(_18286_, _18288_, _18290_);
  xor g_29042_(out[148], _21202_, _18291_);
  not g_29043_(_18291_, _18292_);
  and g_29044_(_18118_, _18213_, _18293_);
  and g_29045_(_18114_, _18212_, _18294_);
  or g_29046_(_18293_, _18294_, _18295_);
  not g_29047_(_18295_, _18296_);
  and g_29048_(_18291_, _18296_, _18297_);
  or g_29049_(_18292_, _18295_, _18298_);
  xor g_29050_(out[149], _21213_, _18299_);
  xor g_29051_(_21092_, _21213_, _18300_);
  or g_29052_(_18105_, _18212_, _18301_);
  not g_29053_(_18301_, _18302_);
  and g_29054_(_18102_, _18212_, _18303_);
  not g_29055_(_18303_, _18304_);
  or g_29056_(_18302_, _18303_, _18305_);
  and g_29057_(_18301_, _18304_, _18306_);
  and g_29058_(_18299_, _18306_, _18307_);
  or g_29059_(_18300_, _18305_, _18308_);
  and g_29060_(_18298_, _18308_, _18309_);
  or g_29061_(_18297_, _18307_, _18310_);
  and g_29062_(_18292_, _18295_, _18311_);
  or g_29063_(_18291_, _18296_, _18312_);
  and g_29064_(_18300_, _18305_, _18313_);
  or g_29065_(_18299_, _18306_, _18314_);
  and g_29066_(_18312_, _18314_, _18315_);
  or g_29067_(_18311_, _18313_, _18316_);
  and g_29068_(_18309_, _18315_, _18317_);
  or g_29069_(_18310_, _18316_, _18318_);
  and g_29070_(_18289_, _18317_, _18319_);
  or g_29071_(_18290_, _18318_, _18320_);
  xor g_29072_(out[147], _21180_, _18321_);
  xor g_29073_(_21136_, _21180_, _18322_);
  and g_29074_(_18130_, _18212_, _18323_);
  not g_29075_(_18323_, _18324_);
  or g_29076_(_18133_, _18212_, _18325_);
  not g_29077_(_18325_, _18326_);
  or g_29078_(_18323_, _18326_, _18327_);
  and g_29079_(_18324_, _18325_, _18328_);
  and g_29080_(_18321_, _18328_, _18329_);
  or g_29081_(_18125_, _18212_, _18330_);
  not g_29082_(_18330_, _18331_);
  and g_29083_(_18128_, _18212_, _18332_);
  or g_29084_(_18127_, _18213_, _18333_);
  and g_29085_(_18330_, _18333_, _18334_);
  or g_29086_(_18331_, _18332_, _18335_);
  or g_29087_(out[145], out[146], _18336_);
  xor g_29088_(out[145], out[146], _18337_);
  xor g_29089_(_21103_, out[146], _18338_);
  and g_29090_(_18334_, _18338_, _18339_);
  or g_29091_(_18329_, _18339_, _18340_);
  and g_29092_(_18322_, _18327_, _18341_);
  or g_29093_(_18321_, _18328_, _18342_);
  and g_29094_(_18335_, _18337_, _18343_);
  or g_29095_(_18341_, _18343_, _18344_);
  xor g_29096_(_18322_, _18327_, _18345_);
  xor g_29097_(_18335_, _18337_, _18346_);
  and g_29098_(_18345_, _18346_, _18347_);
  or g_29099_(_18340_, _18344_, _18348_);
  and g_29100_(out[129], _18212_, _18349_);
  and g_29101_(_18146_, _18213_, _18350_);
  or g_29102_(_18349_, _18350_, _18351_);
  not g_29103_(_18351_, _18352_);
  and g_29104_(out[145], _18352_, _18353_);
  or g_29105_(_21103_, _18351_, _18354_);
  or g_29106_(_18151_, _18212_, _18355_);
  or g_29107_(out[128], _18213_, _18356_);
  and g_29108_(_18355_, _18356_, _18357_);
  not g_29109_(_18357_, _18358_);
  and g_29110_(out[144], _18358_, _18359_);
  or g_29111_(_21114_, _18357_, _18360_);
  xor g_29112_(_21103_, _18351_, _18361_);
  xor g_29113_(out[145], _18351_, _18362_);
  and g_29114_(_18360_, _18361_, _18363_);
  or g_29115_(_18359_, _18362_, _18364_);
  and g_29116_(_18354_, _18364_, _18365_);
  or g_29117_(_18353_, _18363_, _18366_);
  and g_29118_(_18347_, _18366_, _18367_);
  or g_29119_(_18348_, _18365_, _18368_);
  and g_29120_(_18340_, _18342_, _18369_);
  not g_29121_(_18369_, _18370_);
  and g_29122_(_18368_, _18370_, _18371_);
  or g_29123_(_18367_, _18369_, _18372_);
  and g_29124_(_18319_, _18372_, _18373_);
  or g_29125_(_18320_, _18371_, _18374_);
  or g_29126_(_18283_, _18284_, _18375_);
  not g_29127_(_18375_, _18376_);
  and g_29128_(_18289_, _18310_, _18377_);
  or g_29129_(_18290_, _18309_, _18378_);
  and g_29130_(_18314_, _18377_, _18379_);
  or g_29131_(_18313_, _18378_, _18380_);
  and g_29132_(_18375_, _18380_, _18381_);
  or g_29133_(_18376_, _18379_, _18382_);
  and g_29134_(_18374_, _18381_, _18383_);
  or g_29135_(_18373_, _18382_, _18384_);
  and g_29136_(_18264_, _18384_, _18385_);
  or g_29137_(_18265_, _18383_, _18386_);
  and g_29138_(_18244_, _18261_, _18387_);
  or g_29139_(_18245_, _18260_, _18388_);
  and g_29140_(_18229_, _18231_, _18389_);
  or g_29141_(_18228_, _18230_, _18390_);
  and g_29142_(_18388_, _18390_, _18391_);
  or g_29143_(_18387_, _18389_, _18392_);
  and g_29144_(_18386_, _18391_, _18393_);
  or g_29145_(_18385_, _18392_, _18394_);
  and g_29146_(_21114_, _18357_, _18395_);
  or g_29147_(_18348_, _18364_, _18396_);
  or g_29148_(_18395_, _18396_, _18397_);
  or g_29149_(_18320_, _18397_, _18398_);
  not g_29150_(_18398_, _18399_);
  and g_29151_(_18264_, _18399_, _18400_);
  or g_29152_(_18265_, _18398_, _18401_);
  and g_29153_(_18394_, _18401_, _18402_);
  or g_29154_(_18393_, _18400_, _18403_);
  or g_29155_(_21279_, _18403_, _18404_);
  or g_29156_(_18238_, _18402_, _18405_);
  and g_29157_(_18404_, _18405_, _18406_);
  and g_29158_(out[305], out[306], _18407_);
  or g_29159_(out[308], out[307], _18408_);
  or g_29160_(out[307], _18407_, _18409_);
  or g_29161_(_18407_, _18408_, _18410_);
  or g_29162_(out[309], _18410_, _18411_);
  and g_29163_(out[310], _18411_, _18412_);
  and g_29164_(out[311], _18412_, _18413_);
  or g_29165_(out[312], _18413_, _18414_);
  or g_29166_(out[313], _18414_, _18415_);
  xor g_29167_(out[313], _18414_, _18416_);
  not g_29168_(_18416_, _18417_);
  or g_29169_(out[314], _18415_, _18418_);
  xor g_29170_(out[314], _18415_, _18419_);
  not g_29171_(_18419_, _18420_);
  and g_29172_(out[177], out[178], _18421_);
  or g_29173_(out[180], out[179], _18422_);
  or g_29174_(out[179], _18421_, _18423_);
  or g_29175_(_18421_, _18422_, _18424_);
  or g_29176_(out[181], _18424_, _18425_);
  and g_29177_(out[182], _18425_, _18426_);
  and g_29178_(out[183], _18426_, _18427_);
  or g_29179_(out[184], _18427_, _18428_);
  or g_29180_(out[185], _18428_, _18429_);
  or g_29181_(out[186], _18429_, _18430_);
  xor g_29182_(out[186], _18429_, _18431_);
  xor g_29183_(_18837_, _18429_, _18432_);
  and g_29184_(out[161], out[162], _18433_);
  or g_29185_(out[164], out[163], _18434_);
  or g_29186_(out[163], _18433_, _18435_);
  or g_29187_(_18433_, _18434_, _18436_);
  or g_29188_(out[165], _18436_, _18437_);
  and g_29189_(out[166], _18437_, _18438_);
  and g_29190_(out[167], _18438_, _18439_);
  or g_29191_(out[168], _18439_, _18440_);
  or g_29192_(out[169], _18440_, _18441_);
  or g_29193_(out[170], _18441_, _18442_);
  xor g_29194_(_18595_, _18442_, _18443_);
  xor g_29195_(out[171], _18442_, _18444_);
  xor g_29196_(_18716_, _18430_, _18445_);
  xor g_29197_(out[187], _18430_, _18446_);
  and g_29198_(_18443_, _18446_, _18447_);
  or g_29199_(_18444_, _18445_, _18448_);
  xor g_29200_(out[166], _18437_, _18449_);
  xor g_29201_(_18617_, _18437_, _18450_);
  xor g_29202_(out[182], _18425_, _18451_);
  xor g_29203_(_18738_, _18425_, _18452_);
  and g_29204_(_18449_, _18452_, _18453_);
  or g_29205_(_18450_, _18451_, _18454_);
  xor g_29206_(out[163], _18433_, _18455_);
  xor g_29207_(_18672_, _18433_, _18456_);
  xor g_29208_(out[179], _18421_, _18457_);
  xor g_29209_(_18804_, _18421_, _18458_);
  and g_29210_(_18455_, _18458_, _18459_);
  or g_29211_(_18456_, _18457_, _18460_);
  and g_29212_(_18456_, _18457_, _18461_);
  or g_29213_(_18455_, _18458_, _18462_);
  or g_29214_(out[177], out[178], _18463_);
  not g_29215_(_18463_, _18464_);
  xor g_29216_(out[177], out[178], _18465_);
  or g_29217_(_18421_, _18464_, _18466_);
  or g_29218_(out[161], out[162], _18467_);
  xor g_29219_(out[161], out[162], _18468_);
  xor g_29220_(_18650_, out[162], _18469_);
  and g_29221_(_18466_, _18468_, _18470_);
  or g_29222_(_18465_, _18469_, _18471_);
  and g_29223_(_18465_, _18469_, _18472_);
  not g_29224_(_18472_, _18473_);
  and g_29225_(_18460_, _18471_, _18474_);
  or g_29226_(_18459_, _18470_, _18475_);
  and g_29227_(_18462_, _18473_, _18476_);
  or g_29228_(_18461_, _18472_, _18477_);
  and g_29229_(_18474_, _18476_, _18478_);
  or g_29230_(_18475_, _18477_, _18479_);
  and g_29231_(_18650_, out[177], _18480_);
  or g_29232_(out[161], _18771_, _18481_);
  and g_29233_(_18584_, out[176], _18482_);
  or g_29234_(out[160], _18782_, _18483_);
  and g_29235_(out[161], _18771_, _18484_);
  or g_29236_(_18650_, out[177], _18485_);
  xor g_29237_(_18650_, out[177], _18486_);
  xor g_29238_(out[161], out[177], _18487_);
  and g_29239_(_18483_, _18486_, _18488_);
  or g_29240_(_18482_, _18487_, _18489_);
  and g_29241_(_18481_, _18489_, _18490_);
  or g_29242_(_18480_, _18488_, _18491_);
  and g_29243_(_18478_, _18491_, _18492_);
  or g_29244_(_18479_, _18490_, _18493_);
  and g_29245_(_18460_, _18470_, _18494_);
  or g_29246_(_18459_, _18471_, _18495_);
  and g_29247_(_18462_, _18495_, _18496_);
  or g_29248_(_18461_, _18494_, _18497_);
  and g_29249_(_18493_, _18496_, _18498_);
  or g_29250_(_18492_, _18497_, _18499_);
  xor g_29251_(out[164], _18435_, _18500_);
  xor g_29252_(_18639_, _18435_, _18501_);
  xor g_29253_(out[180], _18423_, _18502_);
  xor g_29254_(_18760_, _18423_, _18503_);
  and g_29255_(_18500_, _18503_, _18504_);
  or g_29256_(_18501_, _18502_, _18505_);
  and g_29257_(out[160], _18782_, _18506_);
  or g_29258_(_18584_, out[176], _18507_);
  and g_29259_(_18488_, _18507_, _18508_);
  or g_29260_(_18489_, _18506_, _18509_);
  and g_29261_(_18478_, _18508_, _18510_);
  or g_29262_(_18479_, _18509_, _18511_);
  and g_29263_(_18505_, _18511_, _18512_);
  or g_29264_(_18504_, _18510_, _18513_);
  and g_29265_(_18499_, _18512_, _18514_);
  or g_29266_(_18498_, _18513_, _18515_);
  xor g_29267_(out[165], _18436_, _18516_);
  xor g_29268_(_18628_, _18436_, _18517_);
  xor g_29269_(out[181], _18424_, _18518_);
  xor g_29270_(_18749_, _18424_, _18519_);
  and g_29271_(_18517_, _18518_, _18520_);
  or g_29272_(_18516_, _18519_, _18521_);
  and g_29273_(_18501_, _18502_, _18522_);
  or g_29274_(_18500_, _18503_, _18523_);
  and g_29275_(_18521_, _18523_, _18524_);
  or g_29276_(_18520_, _18522_, _18525_);
  and g_29277_(_18515_, _18524_, _18526_);
  or g_29278_(_18514_, _18525_, _18527_);
  and g_29279_(_18516_, _18519_, _18528_);
  or g_29280_(_18517_, _18518_, _18529_);
  xor g_29281_(out[167], _18438_, _18530_);
  xor g_29282_(_18606_, _18438_, _18531_);
  xor g_29283_(out[183], _18426_, _18532_);
  xor g_29284_(_18727_, _18426_, _18533_);
  and g_29285_(_18531_, _18532_, _18534_);
  or g_29286_(_18530_, _18533_, _18535_);
  and g_29287_(_18450_, _18451_, _18536_);
  or g_29288_(_18449_, _18452_, _18537_);
  and g_29289_(_18529_, _18537_, _18538_);
  or g_29290_(_18528_, _18536_, _18539_);
  and g_29291_(_18527_, _18538_, _18540_);
  or g_29292_(_18526_, _18539_, _18541_);
  and g_29293_(_18454_, _18541_, _18542_);
  or g_29294_(_18453_, _18540_, _18543_);
  and g_29295_(_18535_, _18543_, _18544_);
  or g_29296_(_18534_, _18542_, _18545_);
  and g_29297_(_18530_, _18533_, _18546_);
  or g_29298_(_18531_, _18532_, _18547_);
  xor g_29299_(out[184], _18427_, _18548_);
  xor g_29300_(_18815_, _18427_, _18549_);
  xor g_29301_(out[168], _18439_, _18550_);
  xor g_29302_(_18683_, _18439_, _18551_);
  and g_29303_(_18548_, _18551_, _18552_);
  or g_29304_(_18549_, _18550_, _18553_);
  and g_29305_(_18547_, _18553_, _18554_);
  or g_29306_(_18546_, _18552_, _18555_);
  and g_29307_(_18545_, _18554_, _18556_);
  or g_29308_(_18544_, _18555_, _18557_);
  xor g_29309_(out[185], _18428_, _18558_);
  xor g_29310_(_18826_, _18428_, _18559_);
  xor g_29311_(out[169], _18440_, _18560_);
  xor g_29312_(_18694_, _18440_, _18561_);
  and g_29313_(_18559_, _18560_, _18563_);
  or g_29314_(_18558_, _18561_, _18564_);
  and g_29315_(_18549_, _18550_, _18565_);
  or g_29316_(_18548_, _18551_, _18566_);
  and g_29317_(_18564_, _18566_, _18567_);
  or g_29318_(_18563_, _18565_, _18568_);
  and g_29319_(_18557_, _18567_, _18569_);
  or g_29320_(_18556_, _18568_, _18570_);
  xor g_29321_(out[170], _18441_, _18571_);
  xor g_29322_(_18705_, _18441_, _18572_);
  and g_29323_(_18431_, _18572_, _18574_);
  or g_29324_(_18432_, _18571_, _18575_);
  and g_29325_(_18558_, _18561_, _18576_);
  or g_29326_(_18559_, _18560_, _18577_);
  and g_29327_(_18575_, _18577_, _18578_);
  or g_29328_(_18574_, _18576_, _18579_);
  and g_29329_(_18570_, _18578_, _18580_);
  or g_29330_(_18569_, _18579_, _18581_);
  and g_29331_(_18444_, _18445_, _18582_);
  or g_29332_(_18443_, _18446_, _18583_);
  and g_29333_(_18432_, _18571_, _18585_);
  or g_29334_(_18431_, _18572_, _18586_);
  and g_29335_(_18583_, _18586_, _18587_);
  or g_29336_(_18582_, _18585_, _18588_);
  and g_29337_(_18581_, _18587_, _18589_);
  or g_29338_(_18580_, _18588_, _18590_);
  and g_29339_(_18448_, _18590_, _18591_);
  or g_29340_(_18447_, _18589_, _18592_);
  and g_29341_(_18431_, _18592_, _18593_);
  or g_29342_(_18432_, _18591_, _18594_);
  and g_29343_(_18571_, _18591_, _18596_);
  or g_29344_(_18572_, _18592_, _18597_);
  and g_29345_(_18594_, _18597_, _18598_);
  or g_29346_(_18593_, _18596_, _18599_);
  and g_29347_(out[193], out[194], _18600_);
  or g_29348_(out[196], out[195], _18601_);
  or g_29349_(out[195], _18600_, _18602_);
  or g_29350_(_18600_, _18601_, _18603_);
  or g_29351_(out[197], _18603_, _18604_);
  and g_29352_(out[198], _18604_, _18605_);
  and g_29353_(out[199], _18605_, _18607_);
  or g_29354_(out[200], _18607_, _18608_);
  or g_29355_(out[201], _18608_, _18609_);
  not g_29356_(_18609_, _18610_);
  or g_29357_(out[202], _18609_, _18611_);
  xor g_29358_(out[202], _18609_, _18612_);
  xor g_29359_(out[202], _18610_, _18613_);
  and g_29360_(_18598_, _18612_, _18614_);
  or g_29361_(_18599_, _18613_, _18615_);
  and g_29362_(_18443_, _18445_, _18616_);
  or g_29363_(_18444_, _18446_, _18618_);
  xor g_29364_(_18848_, _18611_, _18619_);
  xor g_29365_(out[203], _18611_, _18620_);
  and g_29366_(_18616_, _18620_, _18621_);
  or g_29367_(_18618_, _18619_, _18622_);
  and g_29368_(_18615_, _18622_, _18623_);
  or g_29369_(_18614_, _18621_, _18624_);
  and g_29370_(_18618_, _18619_, _18625_);
  or g_29371_(_18616_, _18620_, _18626_);
  and g_29372_(_18599_, _18613_, _18627_);
  or g_29373_(_18598_, _18612_, _18629_);
  and g_29374_(_18626_, _18629_, _18630_);
  or g_29375_(_18625_, _18627_, _18631_);
  and g_29376_(out[201], _18608_, _18632_);
  xor g_29377_(out[201], _18608_, _18633_);
  or g_29378_(_18610_, _18632_, _18634_);
  and g_29379_(_18558_, _18592_, _18635_);
  or g_29380_(_18559_, _18591_, _18636_);
  and g_29381_(_18560_, _18591_, _18637_);
  or g_29382_(_18561_, _18592_, _18638_);
  and g_29383_(_18636_, _18638_, _18640_);
  or g_29384_(_18635_, _18637_, _18641_);
  and g_29385_(_18634_, _18641_, _18642_);
  or g_29386_(_18633_, _18640_, _18643_);
  and g_29387_(_18633_, _18640_, _18644_);
  or g_29388_(_18634_, _18641_, _18645_);
  xor g_29389_(out[200], _18607_, _18646_);
  xor g_29390_(_18947_, _18607_, _18647_);
  and g_29391_(_18550_, _18591_, _18648_);
  or g_29392_(_18551_, _18592_, _18649_);
  and g_29393_(_18548_, _18592_, _18651_);
  or g_29394_(_18549_, _18591_, _18652_);
  and g_29395_(_18649_, _18652_, _18653_);
  or g_29396_(_18648_, _18651_, _18654_);
  and g_29397_(_18646_, _18653_, _18655_);
  or g_29398_(_18647_, _18654_, _18656_);
  and g_29399_(_18645_, _18656_, _18657_);
  or g_29400_(_18644_, _18655_, _18658_);
  and g_29401_(_18647_, _18654_, _18659_);
  or g_29402_(_18646_, _18653_, _18660_);
  and g_29403_(_18623_, _18630_, _18662_);
  or g_29404_(_18624_, _18631_, _18663_);
  and g_29405_(_18643_, _18660_, _18664_);
  or g_29406_(_18642_, _18659_, _18665_);
  and g_29407_(_18657_, _18664_, _18666_);
  or g_29408_(_18658_, _18665_, _18667_);
  and g_29409_(_18662_, _18666_, _18668_);
  or g_29410_(_18663_, _18667_, _18669_);
  xor g_29411_(out[198], _18604_, _18670_);
  xor g_29412_(_18870_, _18604_, _18671_);
  and g_29413_(_18452_, _18592_, _18673_);
  or g_29414_(_18451_, _18591_, _18674_);
  and g_29415_(_18450_, _18591_, _18675_);
  or g_29416_(_18449_, _18592_, _18676_);
  and g_29417_(_18674_, _18676_, _18677_);
  or g_29418_(_18673_, _18675_, _18678_);
  and g_29419_(_18671_, _18677_, _18679_);
  or g_29420_(_18670_, _18678_, _18680_);
  xor g_29421_(out[199], _18605_, _18681_);
  xor g_29422_(_18859_, _18605_, _18682_);
  and g_29423_(_18533_, _18592_, _18684_);
  or g_29424_(_18532_, _18591_, _18685_);
  and g_29425_(_18531_, _18591_, _18686_);
  or g_29426_(_18530_, _18592_, _18687_);
  and g_29427_(_18685_, _18687_, _18688_);
  or g_29428_(_18684_, _18686_, _18689_);
  and g_29429_(_18682_, _18688_, _18690_);
  or g_29430_(_18681_, _18689_, _18691_);
  and g_29431_(_18680_, _18691_, _18692_);
  or g_29432_(_18679_, _18690_, _18693_);
  and g_29433_(_18681_, _18689_, _18695_);
  or g_29434_(_18682_, _18688_, _18696_);
  and g_29435_(_18670_, _18678_, _18697_);
  or g_29436_(_18671_, _18677_, _18698_);
  and g_29437_(_18696_, _18698_, _18699_);
  or g_29438_(_18695_, _18697_, _18700_);
  and g_29439_(_18692_, _18699_, _18701_);
  or g_29440_(_18693_, _18700_, _18702_);
  xor g_29441_(out[197], _18603_, _18703_);
  xor g_29442_(_18881_, _18603_, _18704_);
  and g_29443_(_18518_, _18592_, _18706_);
  or g_29444_(_18519_, _18591_, _18707_);
  and g_29445_(_18516_, _18591_, _18708_);
  or g_29446_(_18517_, _18592_, _18709_);
  and g_29447_(_18707_, _18709_, _18710_);
  or g_29448_(_18706_, _18708_, _18711_);
  and g_29449_(_18703_, _18710_, _18712_);
  or g_29450_(_18704_, _18711_, _18713_);
  xor g_29451_(out[196], _18602_, _18714_);
  xor g_29452_(_18892_, _18602_, _18715_);
  and g_29453_(_18502_, _18592_, _18717_);
  or g_29454_(_18503_, _18591_, _18718_);
  and g_29455_(_18500_, _18591_, _18719_);
  or g_29456_(_18501_, _18592_, _18720_);
  and g_29457_(_18718_, _18720_, _18721_);
  or g_29458_(_18717_, _18719_, _18722_);
  and g_29459_(_18714_, _18721_, _18723_);
  or g_29460_(_18715_, _18722_, _18724_);
  and g_29461_(_18713_, _18724_, _18725_);
  or g_29462_(_18712_, _18723_, _18726_);
  and g_29463_(_18704_, _18711_, _18728_);
  or g_29464_(_18703_, _18710_, _18729_);
  and g_29465_(_18715_, _18722_, _18730_);
  or g_29466_(_18714_, _18721_, _18731_);
  and g_29467_(_18729_, _18731_, _18732_);
  or g_29468_(_18728_, _18730_, _18733_);
  and g_29469_(_18725_, _18732_, _18734_);
  or g_29470_(_18726_, _18733_, _18735_);
  and g_29471_(_18701_, _18734_, _18736_);
  or g_29472_(_18702_, _18735_, _18737_);
  and g_29473_(_18668_, _18736_, _18739_);
  or g_29474_(_18669_, _18737_, _18740_);
  or g_29475_(out[193], out[194], _18741_);
  xor g_29476_(out[193], out[194], _18742_);
  xor g_29477_(_18903_, out[194], _18743_);
  or g_29478_(_18465_, _18591_, _18744_);
  or g_29479_(_18468_, _18592_, _18745_);
  and g_29480_(_18744_, _18745_, _18746_);
  not g_29481_(_18746_, _18747_);
  and g_29482_(_18743_, _18746_, _18748_);
  or g_29483_(_18742_, _18747_, _18750_);
  xor g_29484_(out[195], _18600_, _18751_);
  xor g_29485_(_18936_, _18600_, _18752_);
  and g_29486_(_18457_, _18592_, _18753_);
  or g_29487_(_18458_, _18591_, _18754_);
  and g_29488_(_18455_, _18591_, _18755_);
  or g_29489_(_18456_, _18592_, _18756_);
  and g_29490_(_18754_, _18756_, _18757_);
  or g_29491_(_18753_, _18755_, _18758_);
  and g_29492_(_18751_, _18757_, _18759_);
  or g_29493_(_18752_, _18758_, _18761_);
  or g_29494_(_18748_, _18759_, _18762_);
  and g_29495_(_18752_, _18758_, _18763_);
  or g_29496_(_18751_, _18757_, _18764_);
  and g_29497_(_18742_, _18747_, _18765_);
  or g_29498_(_18763_, _18765_, _18766_);
  and g_29499_(_18761_, _18764_, _18767_);
  xor g_29500_(_18743_, _18746_, _18768_);
  and g_29501_(_18767_, _18768_, _18769_);
  or g_29502_(_18762_, _18766_, _18770_);
  and g_29503_(out[161], _18591_, _18772_);
  or g_29504_(_18650_, _18592_, _18773_);
  and g_29505_(out[177], _18592_, _18774_);
  or g_29506_(_18771_, _18591_, _18775_);
  and g_29507_(_18773_, _18775_, _18776_);
  or g_29508_(_18772_, _18774_, _18777_);
  and g_29509_(out[193], _18776_, _18778_);
  or g_29510_(_18903_, _18777_, _18779_);
  and g_29511_(_18782_, _18592_, _18780_);
  or g_29512_(out[176], _18591_, _18781_);
  and g_29513_(_18584_, _18591_, _18783_);
  or g_29514_(out[160], _18592_, _18784_);
  and g_29515_(_18781_, _18784_, _18785_);
  or g_29516_(_18780_, _18783_, _18786_);
  and g_29517_(out[192], _18786_, _18787_);
  or g_29518_(_18914_, _18785_, _18788_);
  xor g_29519_(out[193], _18776_, _18789_);
  xor g_29520_(_18903_, _18776_, _18790_);
  and g_29521_(_18788_, _18789_, _18791_);
  or g_29522_(_18787_, _18790_, _18792_);
  and g_29523_(_18779_, _18792_, _18794_);
  or g_29524_(_18778_, _18791_, _18795_);
  and g_29525_(_18769_, _18795_, _18796_);
  or g_29526_(_18770_, _18794_, _18797_);
  or g_29527_(_18750_, _18763_, _18798_);
  and g_29528_(_18761_, _18798_, _18799_);
  and g_29529_(_18762_, _18764_, _18800_);
  and g_29530_(_18797_, _18799_, _18801_);
  or g_29531_(_18796_, _18800_, _18802_);
  and g_29532_(_18739_, _18802_, _18803_);
  or g_29533_(_18740_, _18801_, _18805_);
  and g_29534_(_18693_, _18696_, _18806_);
  or g_29535_(_18692_, _18695_, _18807_);
  and g_29536_(_18726_, _18729_, _18808_);
  or g_29537_(_18725_, _18728_, _18809_);
  and g_29538_(_18701_, _18808_, _18810_);
  or g_29539_(_18702_, _18809_, _18811_);
  and g_29540_(_18807_, _18811_, _18812_);
  or g_29541_(_18806_, _18810_, _18813_);
  and g_29542_(_18668_, _18813_, _18814_);
  or g_29543_(_18669_, _18812_, _18816_);
  and g_29544_(_18624_, _18626_, _18817_);
  or g_29545_(_18623_, _18625_, _18818_);
  and g_29546_(_18658_, _18662_, _18819_);
  or g_29547_(_18657_, _18663_, _18820_);
  and g_29548_(_18643_, _18819_, _18821_);
  or g_29549_(_18642_, _18820_, _18822_);
  and g_29550_(_18818_, _18822_, _18823_);
  or g_29551_(_18817_, _18821_, _18824_);
  and g_29552_(_18816_, _18823_, _18825_);
  or g_29553_(_18814_, _18824_, _18827_);
  and g_29554_(_18805_, _18825_, _18828_);
  or g_29555_(_18803_, _18827_, _18829_);
  and g_29556_(_18914_, _18785_, _18830_);
  or g_29557_(out[192], _18786_, _18831_);
  and g_29558_(_18769_, _18831_, _18832_);
  or g_29559_(_18770_, _18830_, _18833_);
  and g_29560_(_18791_, _18832_, _18834_);
  or g_29561_(_18792_, _18833_, _18835_);
  and g_29562_(_18739_, _18834_, _18836_);
  or g_29563_(_18740_, _18835_, _18838_);
  and g_29564_(_18829_, _18838_, _18839_);
  or g_29565_(_18828_, _18836_, _18840_);
  and g_29566_(_18599_, _18840_, _18841_);
  or g_29567_(_18598_, _18839_, _18842_);
  and g_29568_(_18612_, _18839_, _18843_);
  not g_29569_(_18843_, _18844_);
  and g_29570_(_18842_, _18844_, _18845_);
  or g_29571_(_18841_, _18843_, _18846_);
  and g_29572_(out[209], out[210], _18847_);
  or g_29573_(out[209], out[210], _18849_);
  xor g_29574_(out[209], out[210], _18850_);
  xor g_29575_(_19013_, out[210], _18851_);
  or g_29576_(_18746_, _18839_, _18852_);
  or g_29577_(_18742_, _18840_, _18853_);
  and g_29578_(_18852_, _18853_, _18854_);
  and g_29579_(_18851_, _18854_, _18855_);
  or g_29580_(out[211], _18847_, _18856_);
  xor g_29581_(out[211], _18847_, _18857_);
  xor g_29582_(_19046_, _18847_, _18858_);
  or g_29583_(_18758_, _18839_, _18860_);
  not g_29584_(_18860_, _18861_);
  and g_29585_(_18752_, _18839_, _18862_);
  or g_29586_(_18751_, _18840_, _18863_);
  and g_29587_(_18860_, _18863_, _18864_);
  or g_29588_(_18861_, _18862_, _18865_);
  and g_29589_(_18857_, _18865_, _18866_);
  or g_29590_(_18858_, _18864_, _18867_);
  or g_29591_(_18855_, _18866_, _18868_);
  and g_29592_(out[193], _18839_, _18869_);
  not g_29593_(_18869_, _18871_);
  and g_29594_(_18777_, _18840_, _18872_);
  or g_29595_(_18776_, _18839_, _18873_);
  and g_29596_(_18871_, _18873_, _18874_);
  or g_29597_(_18869_, _18872_, _18875_);
  and g_29598_(out[209], _18874_, _18876_);
  or g_29599_(_18785_, _18839_, _18877_);
  not g_29600_(_18877_, _18878_);
  and g_29601_(_18914_, _18839_, _18879_);
  or g_29602_(out[192], _18840_, _18880_);
  and g_29603_(_18877_, _18880_, _18882_);
  or g_29604_(_18878_, _18879_, _18883_);
  and g_29605_(out[208], _18883_, _18884_);
  or g_29606_(_19024_, _18882_, _18885_);
  xor g_29607_(_19013_, _18875_, _18886_);
  xor g_29608_(out[209], _18875_, _18887_);
  and g_29609_(_18885_, _18886_, _18888_);
  or g_29610_(_18884_, _18887_, _18889_);
  or g_29611_(_18876_, _18888_, _18890_);
  xor g_29612_(_18851_, _18854_, _18891_);
  xor g_29613_(_18850_, _18854_, _18893_);
  and g_29614_(_18890_, _18891_, _18894_);
  or g_29615_(_18868_, _18894_, _18895_);
  not g_29616_(_18895_, _18896_);
  or g_29617_(out[212], out[211], _18897_);
  or g_29618_(_18847_, _18897_, _18898_);
  or g_29619_(out[213], _18898_, _18899_);
  and g_29620_(out[214], _18899_, _18900_);
  and g_29621_(out[215], _18900_, _18901_);
  or g_29622_(out[216], _18901_, _18902_);
  or g_29623_(out[217], _18902_, _18904_);
  or g_29624_(out[218], _18904_, _18905_);
  xor g_29625_(out[218], _18904_, _18906_);
  not g_29626_(_18906_, _18907_);
  and g_29627_(_18845_, _18906_, _18908_);
  and g_29628_(_18620_, _18839_, _18909_);
  not g_29629_(_18909_, _18910_);
  and g_29630_(_18618_, _18840_, _18911_);
  or g_29631_(_18616_, _18839_, _18912_);
  and g_29632_(_18910_, _18912_, _18913_);
  or g_29633_(_18909_, _18911_, _18915_);
  xor g_29634_(out[219], _18905_, _18916_);
  not g_29635_(_18916_, _18917_);
  and g_29636_(_18913_, _18916_, _18918_);
  or g_29637_(_18908_, _18918_, _18919_);
  and g_29638_(_18846_, _18907_, _18920_);
  and g_29639_(_18915_, _18917_, _18921_);
  or g_29640_(_18913_, _18916_, _18922_);
  xor g_29641_(out[217], _18902_, _18923_);
  xor g_29642_(_19068_, _18902_, _18924_);
  and g_29643_(_18641_, _18840_, _18926_);
  or g_29644_(_18640_, _18839_, _18927_);
  and g_29645_(_18633_, _18839_, _18928_);
  not g_29646_(_18928_, _18929_);
  and g_29647_(_18927_, _18929_, _18930_);
  or g_29648_(_18926_, _18928_, _18931_);
  and g_29649_(_18924_, _18931_, _18932_);
  or g_29650_(_18923_, _18930_, _18933_);
  or g_29651_(_18921_, _18932_, _18934_);
  or g_29652_(_18920_, _18934_, _18935_);
  xor g_29653_(_18846_, _18907_, _18937_);
  xor g_29654_(_18915_, _18917_, _18938_);
  and g_29655_(_18937_, _18938_, _18939_);
  and g_29656_(_18933_, _18939_, _18940_);
  or g_29657_(_18919_, _18935_, _18941_);
  xor g_29658_(out[216], _18901_, _18942_);
  xor g_29659_(_19057_, _18901_, _18943_);
  and g_29660_(_18646_, _18839_, _18944_);
  not g_29661_(_18944_, _18945_);
  and g_29662_(_18654_, _18840_, _18946_);
  or g_29663_(_18653_, _18839_, _18948_);
  and g_29664_(_18945_, _18948_, _18949_);
  or g_29665_(_18944_, _18946_, _18950_);
  and g_29666_(_18943_, _18950_, _18951_);
  or g_29667_(_18942_, _18949_, _18952_);
  and g_29668_(_18923_, _18930_, _18953_);
  or g_29669_(_18924_, _18931_, _18954_);
  and g_29670_(_18942_, _18949_, _18955_);
  or g_29671_(_18943_, _18950_, _18956_);
  and g_29672_(_18954_, _18956_, _18957_);
  or g_29673_(_18953_, _18955_, _18959_);
  and g_29674_(_18952_, _18957_, _18960_);
  or g_29675_(_18951_, _18959_, _18961_);
  and g_29676_(_18940_, _18960_, _18962_);
  or g_29677_(_18941_, _18961_, _18963_);
  xor g_29678_(out[214], _18899_, _18964_);
  xor g_29679_(_18980_, _18899_, _18965_);
  and g_29680_(_18678_, _18840_, _18966_);
  or g_29681_(_18677_, _18839_, _18967_);
  and g_29682_(_18671_, _18839_, _18968_);
  or g_29683_(_18670_, _18840_, _18970_);
  and g_29684_(_18967_, _18970_, _18971_);
  or g_29685_(_18966_, _18968_, _18972_);
  and g_29686_(_18965_, _18971_, _18973_);
  or g_29687_(_18964_, _18972_, _18974_);
  xor g_29688_(out[215], _18900_, _18975_);
  xor g_29689_(_18969_, _18900_, _18976_);
  and g_29690_(_18688_, _18840_, _18977_);
  or g_29691_(_18689_, _18839_, _18978_);
  and g_29692_(_18681_, _18839_, _18979_);
  or g_29693_(_18682_, _18840_, _18981_);
  and g_29694_(_18978_, _18981_, _18982_);
  or g_29695_(_18977_, _18979_, _18983_);
  and g_29696_(_18976_, _18983_, _18984_);
  or g_29697_(_18975_, _18982_, _18985_);
  and g_29698_(_18974_, _18985_, _18986_);
  or g_29699_(_18973_, _18984_, _18987_);
  and g_29700_(_18975_, _18982_, _18988_);
  or g_29701_(_18976_, _18983_, _18989_);
  and g_29702_(_18964_, _18972_, _18990_);
  or g_29703_(_18965_, _18971_, _18992_);
  and g_29704_(_18989_, _18992_, _18993_);
  or g_29705_(_18988_, _18990_, _18994_);
  and g_29706_(_18986_, _18993_, _18995_);
  or g_29707_(_18987_, _18994_, _18996_);
  xor g_29708_(out[212], _18856_, _18997_);
  xor g_29709_(_19002_, _18856_, _18998_);
  and g_29710_(_18722_, _18840_, _18999_);
  or g_29711_(_18721_, _18839_, _19000_);
  and g_29712_(_18714_, _18839_, _19001_);
  or g_29713_(_18715_, _18840_, _19003_);
  and g_29714_(_19000_, _19003_, _19004_);
  or g_29715_(_18999_, _19001_, _19005_);
  and g_29716_(_18997_, _19004_, _19006_);
  or g_29717_(_18998_, _19005_, _19007_);
  xor g_29718_(out[213], _18898_, _19008_);
  xor g_29719_(_18991_, _18898_, _19009_);
  and g_29720_(_18710_, _18840_, _19010_);
  or g_29721_(_18711_, _18839_, _19011_);
  and g_29722_(_18704_, _18839_, _19012_);
  or g_29723_(_18703_, _18840_, _19014_);
  and g_29724_(_19011_, _19014_, _19015_);
  or g_29725_(_19010_, _19012_, _19016_);
  and g_29726_(_19008_, _19016_, _19017_);
  or g_29727_(_19009_, _19015_, _19018_);
  and g_29728_(_19007_, _19018_, _19019_);
  or g_29729_(_19006_, _19017_, _19020_);
  and g_29730_(_18998_, _19005_, _19021_);
  or g_29731_(_18997_, _19004_, _19022_);
  and g_29732_(_19009_, _19015_, _19023_);
  or g_29733_(_19008_, _19016_, _19025_);
  and g_29734_(_18858_, _18864_, _19026_);
  or g_29735_(_18857_, _18865_, _19027_);
  and g_29736_(_19025_, _19027_, _19028_);
  or g_29737_(_19023_, _19026_, _19029_);
  and g_29738_(_19022_, _19028_, _19030_);
  or g_29739_(_19021_, _19029_, _19031_);
  and g_29740_(_19019_, _19030_, _19032_);
  or g_29741_(_19020_, _19031_, _19033_);
  and g_29742_(_18995_, _19032_, _19034_);
  or g_29743_(_18996_, _19033_, _19036_);
  and g_29744_(_18962_, _19034_, _19037_);
  or g_29745_(_18963_, _19036_, _19038_);
  and g_29746_(_18895_, _19037_, _19039_);
  or g_29747_(_18896_, _19038_, _19040_);
  and g_29748_(_18987_, _18989_, _19041_);
  or g_29749_(_18986_, _18988_, _19042_);
  and g_29750_(_19020_, _19025_, _19043_);
  or g_29751_(_19019_, _19023_, _19044_);
  and g_29752_(_18995_, _19043_, _19045_);
  or g_29753_(_18996_, _19044_, _19047_);
  and g_29754_(_19042_, _19047_, _19048_);
  or g_29755_(_19041_, _19045_, _19049_);
  and g_29756_(_18962_, _19049_, _19050_);
  or g_29757_(_18963_, _19048_, _19051_);
  and g_29758_(_18940_, _18959_, _19052_);
  and g_29759_(_18919_, _18922_, _19053_);
  or g_29760_(_19052_, _19053_, _19054_);
  not g_29761_(_19054_, _19055_);
  and g_29762_(_19051_, _19055_, _19056_);
  or g_29763_(_19050_, _19054_, _19058_);
  and g_29764_(_19040_, _19056_, _19059_);
  or g_29765_(_19039_, _19058_, _19060_);
  and g_29766_(_19024_, _18882_, _19061_);
  or g_29767_(out[208], _18883_, _19062_);
  and g_29768_(_18867_, _19062_, _19063_);
  or g_29769_(_18866_, _19061_, _19064_);
  and g_29770_(_18891_, _19063_, _19065_);
  or g_29771_(_18893_, _19064_, _19066_);
  and g_29772_(_18888_, _19065_, _19067_);
  or g_29773_(_18889_, _19066_, _19069_);
  and g_29774_(_19037_, _19067_, _19070_);
  or g_29775_(_19038_, _19069_, _19071_);
  and g_29776_(_19060_, _19071_, _19072_);
  or g_29777_(_19059_, _19070_, _19073_);
  and g_29778_(_18846_, _19073_, _19074_);
  or g_29779_(_18845_, _19072_, _19075_);
  and g_29780_(_18906_, _19072_, _19076_);
  or g_29781_(_18907_, _19073_, _19077_);
  and g_29782_(_19075_, _19077_, _19078_);
  or g_29783_(_19074_, _19076_, _19080_);
  and g_29784_(out[225], out[226], _19081_);
  or g_29785_(out[228], out[227], _19082_);
  or g_29786_(out[227], _19081_, _19083_);
  or g_29787_(_19081_, _19082_, _19084_);
  or g_29788_(out[229], _19084_, _19085_);
  and g_29789_(out[230], _19085_, _19086_);
  and g_29790_(out[231], _19086_, _19087_);
  or g_29791_(out[232], _19087_, _19088_);
  or g_29792_(out[233], _19088_, _19089_);
  or g_29793_(out[234], _19089_, _19091_);
  xor g_29794_(out[234], _19089_, _19092_);
  xor g_29795_(_19211_, _19089_, _19093_);
  and g_29796_(_19078_, _19092_, _19094_);
  or g_29797_(_19080_, _19093_, _19095_);
  xor g_29798_(_19090_, _19091_, _19096_);
  xor g_29799_(out[235], _19091_, _19097_);
  and g_29800_(_18916_, _19072_, _19098_);
  or g_29801_(_18917_, _19073_, _19099_);
  and g_29802_(_18915_, _19073_, _19100_);
  or g_29803_(_18913_, _19072_, _19102_);
  and g_29804_(_19099_, _19102_, _19103_);
  or g_29805_(_19098_, _19100_, _19104_);
  and g_29806_(_19097_, _19103_, _19105_);
  or g_29807_(_19096_, _19104_, _19106_);
  and g_29808_(_19095_, _19106_, _19107_);
  or g_29809_(_19094_, _19105_, _19108_);
  and g_29810_(_19096_, _19104_, _19109_);
  or g_29811_(_19097_, _19103_, _19110_);
  and g_29812_(_19080_, _19093_, _19111_);
  or g_29813_(_19078_, _19092_, _19113_);
  and g_29814_(_19110_, _19113_, _19114_);
  or g_29815_(_19109_, _19111_, _19115_);
  xor g_29816_(out[233], _19088_, _19116_);
  xor g_29817_(_19200_, _19088_, _19117_);
  and g_29818_(_18924_, _19072_, _19118_);
  or g_29819_(_18923_, _19073_, _19119_);
  or g_29820_(_18931_, _19072_, _19120_);
  not g_29821_(_19120_, _19121_);
  and g_29822_(_19119_, _19120_, _19122_);
  or g_29823_(_19118_, _19121_, _19124_);
  and g_29824_(_19117_, _19122_, _19125_);
  or g_29825_(_19116_, _19124_, _19126_);
  and g_29826_(_19114_, _19126_, _19127_);
  or g_29827_(_19115_, _19125_, _19128_);
  and g_29828_(_19107_, _19127_, _19129_);
  or g_29829_(_19108_, _19128_, _19130_);
  xor g_29830_(out[232], _19087_, _19131_);
  xor g_29831_(_19189_, _19087_, _19132_);
  and g_29832_(_18942_, _19072_, _19133_);
  not g_29833_(_19133_, _19135_);
  and g_29834_(_18950_, _19073_, _19136_);
  or g_29835_(_18949_, _19072_, _19137_);
  and g_29836_(_19135_, _19137_, _19138_);
  or g_29837_(_19133_, _19136_, _19139_);
  and g_29838_(_19132_, _19139_, _19140_);
  or g_29839_(_19131_, _19138_, _19141_);
  and g_29840_(_19116_, _19124_, _19142_);
  or g_29841_(_19117_, _19122_, _19143_);
  and g_29842_(_19131_, _19138_, _19144_);
  or g_29843_(_19132_, _19139_, _19146_);
  and g_29844_(_19143_, _19146_, _19147_);
  or g_29845_(_19142_, _19144_, _19148_);
  and g_29846_(_19141_, _19147_, _19149_);
  or g_29847_(_19140_, _19148_, _19150_);
  and g_29848_(_19129_, _19149_, _19151_);
  or g_29849_(_19130_, _19150_, _19152_);
  and g_29850_(_18965_, _19072_, _19153_);
  or g_29851_(_18964_, _19073_, _19154_);
  or g_29852_(_18971_, _19072_, _19155_);
  not g_29853_(_19155_, _19157_);
  and g_29854_(_19154_, _19155_, _19158_);
  or g_29855_(_19153_, _19157_, _19159_);
  xor g_29856_(out[230], _19085_, _19160_);
  not g_29857_(_19160_, _19161_);
  or g_29858_(_19159_, _19160_, _19162_);
  xor g_29859_(out[231], _19086_, _19163_);
  and g_29860_(_18975_, _19072_, _19164_);
  not g_29861_(_19164_, _19165_);
  and g_29862_(_18983_, _19073_, _19166_);
  or g_29863_(_18982_, _19072_, _19168_);
  and g_29864_(_19165_, _19168_, _19169_);
  or g_29865_(_19164_, _19166_, _19170_);
  or g_29866_(_19163_, _19169_, _19171_);
  and g_29867_(_19162_, _19171_, _19172_);
  and g_29868_(_19163_, _19169_, _19173_);
  xor g_29869_(_19158_, _19161_, _19174_);
  xor g_29870_(_19158_, _19160_, _19175_);
  xor g_29871_(_19163_, _19169_, _19176_);
  xor g_29872_(_19163_, _19170_, _19177_);
  and g_29873_(_19174_, _19176_, _19179_);
  or g_29874_(_19175_, _19177_, _19180_);
  xor g_29875_(out[229], _19084_, _19181_);
  xor g_29876_(_19123_, _19084_, _19182_);
  and g_29877_(_19009_, _19072_, _19183_);
  or g_29878_(_19008_, _19073_, _19184_);
  or g_29879_(_19015_, _19072_, _19185_);
  not g_29880_(_19185_, _19186_);
  and g_29881_(_19184_, _19185_, _19187_);
  or g_29882_(_19183_, _19186_, _19188_);
  and g_29883_(_19181_, _19188_, _19190_);
  or g_29884_(_19182_, _19187_, _19191_);
  xor g_29885_(out[228], _19083_, _19192_);
  xor g_29886_(_19134_, _19083_, _19193_);
  and g_29887_(_18997_, _19072_, _19194_);
  not g_29888_(_19194_, _19195_);
  and g_29889_(_19005_, _19073_, _19196_);
  or g_29890_(_19004_, _19072_, _19197_);
  and g_29891_(_19195_, _19197_, _19198_);
  or g_29892_(_19194_, _19196_, _19199_);
  and g_29893_(_19192_, _19198_, _19201_);
  or g_29894_(_19193_, _19199_, _19202_);
  and g_29895_(_19191_, _19202_, _19203_);
  or g_29896_(_19190_, _19201_, _19204_);
  and g_29897_(_19193_, _19199_, _19205_);
  or g_29898_(_19192_, _19198_, _19206_);
  and g_29899_(_19182_, _19187_, _19207_);
  or g_29900_(_19181_, _19188_, _19208_);
  and g_29901_(_19206_, _19208_, _19209_);
  or g_29902_(_19205_, _19207_, _19210_);
  and g_29903_(_19203_, _19209_, _19212_);
  or g_29904_(_19204_, _19210_, _19213_);
  and g_29905_(_19179_, _19212_, _19214_);
  or g_29906_(_19180_, _19213_, _19215_);
  and g_29907_(_19151_, _19214_, _19216_);
  or g_29908_(_19152_, _19215_, _19217_);
  xor g_29909_(out[227], _19081_, _19218_);
  xor g_29910_(_19178_, _19081_, _19219_);
  or g_29911_(_18864_, _19072_, _19220_);
  not g_29912_(_19220_, _19221_);
  and g_29913_(_18858_, _19072_, _19223_);
  or g_29914_(_18857_, _19073_, _19224_);
  and g_29915_(_19220_, _19224_, _19225_);
  or g_29916_(_19221_, _19223_, _19226_);
  and g_29917_(_19219_, _19225_, _19227_);
  or g_29918_(_19218_, _19226_, _19228_);
  or g_29919_(out[225], out[226], _19229_);
  xor g_29920_(out[225], out[226], _19230_);
  xor g_29921_(_19145_, out[226], _19231_);
  or g_29922_(_18850_, _19073_, _19232_);
  or g_29923_(_18854_, _19072_, _19234_);
  and g_29924_(_19232_, _19234_, _19235_);
  and g_29925_(_19231_, _19235_, _19236_);
  and g_29926_(_19218_, _19226_, _19237_);
  or g_29927_(_19236_, _19237_, _19238_);
  not g_29928_(_19238_, _19239_);
  and g_29929_(out[209], _19072_, _19240_);
  not g_29930_(_19240_, _19241_);
  and g_29931_(_18875_, _19073_, _19242_);
  or g_29932_(_18874_, _19072_, _19243_);
  and g_29933_(_19241_, _19243_, _19245_);
  or g_29934_(_19240_, _19242_, _19246_);
  and g_29935_(out[225], _19245_, _19247_);
  or g_29936_(_19145_, _19246_, _19248_);
  or g_29937_(_18882_, _19072_, _19249_);
  or g_29938_(out[208], _19073_, _19250_);
  and g_29939_(_19249_, _19250_, _19251_);
  not g_29940_(_19251_, _19252_);
  and g_29941_(out[224], _19252_, _19253_);
  or g_29942_(_19156_, _19251_, _19254_);
  xor g_29943_(_19145_, _19246_, _19256_);
  xor g_29944_(out[225], _19246_, _19257_);
  and g_29945_(_19254_, _19256_, _19258_);
  or g_29946_(_19253_, _19257_, _19259_);
  and g_29947_(_19248_, _19259_, _19260_);
  or g_29948_(_19247_, _19258_, _19261_);
  xor g_29949_(_19231_, _19235_, _19262_);
  xor g_29950_(_19230_, _19235_, _19263_);
  and g_29951_(_19261_, _19262_, _19264_);
  or g_29952_(_19260_, _19263_, _19265_);
  and g_29953_(_19239_, _19265_, _19267_);
  or g_29954_(_19238_, _19264_, _19268_);
  or g_29955_(_19227_, _19263_, _19269_);
  xor g_29956_(_19219_, _19225_, _19270_);
  and g_29957_(_19228_, _19268_, _19271_);
  or g_29958_(_19227_, _19267_, _19272_);
  and g_29959_(_19216_, _19271_, _19273_);
  or g_29960_(_19217_, _19272_, _19274_);
  or g_29961_(_19172_, _19173_, _19275_);
  not g_29962_(_19275_, _19276_);
  and g_29963_(_19179_, _19204_, _19278_);
  or g_29964_(_19180_, _19203_, _19279_);
  and g_29965_(_19208_, _19278_, _19280_);
  or g_29966_(_19207_, _19279_, _19281_);
  and g_29967_(_19275_, _19281_, _19282_);
  or g_29968_(_19276_, _19280_, _19283_);
  and g_29969_(_19151_, _19283_, _19284_);
  or g_29970_(_19152_, _19282_, _19285_);
  and g_29971_(_19108_, _19110_, _19286_);
  or g_29972_(_19107_, _19109_, _19287_);
  and g_29973_(_19129_, _19148_, _19289_);
  or g_29974_(_19130_, _19147_, _19290_);
  and g_29975_(_19287_, _19290_, _19291_);
  or g_29976_(_19286_, _19289_, _19292_);
  and g_29977_(_19285_, _19291_, _19293_);
  or g_29978_(_19284_, _19292_, _19294_);
  and g_29979_(_19274_, _19293_, _19295_);
  or g_29980_(_19273_, _19294_, _19296_);
  and g_29981_(_19156_, _19251_, _19297_);
  or g_29982_(out[224], _19252_, _19298_);
  and g_29983_(_19270_, _19298_, _19300_);
  or g_29984_(_19237_, _19297_, _19301_);
  and g_29985_(_19262_, _19300_, _19302_);
  or g_29986_(_19269_, _19301_, _19303_);
  and g_29987_(_19258_, _19302_, _19304_);
  or g_29988_(_19259_, _19303_, _19305_);
  and g_29989_(_19216_, _19304_, _19306_);
  or g_29990_(_19217_, _19305_, _19307_);
  and g_29991_(_19296_, _19307_, _19308_);
  or g_29992_(_19295_, _19306_, _19309_);
  or g_29993_(_19078_, _19308_, _19311_);
  not g_29994_(_19311_, _19312_);
  and g_29995_(_19092_, _19308_, _19313_);
  not g_29996_(_19313_, _19314_);
  and g_29997_(_19311_, _19314_, _19315_);
  or g_29998_(_19312_, _19313_, _19316_);
  and g_29999_(out[241], out[242], _19317_);
  or g_30000_(out[244], out[243], _19318_);
  or g_30001_(out[243], _19317_, _19319_);
  or g_30002_(_19317_, _19318_, _19320_);
  or g_30003_(out[245], _19320_, _19322_);
  and g_30004_(out[246], _19322_, _19323_);
  and g_30005_(out[247], _19323_, _19324_);
  or g_30006_(out[248], _19324_, _19325_);
  or g_30007_(out[249], _19325_, _19326_);
  or g_30008_(out[250], _19326_, _19327_);
  xor g_30009_(out[250], _19326_, _19328_);
  xor g_30010_(_19343_, _19326_, _19329_);
  and g_30011_(_19315_, _19328_, _19330_);
  or g_30012_(_19316_, _19329_, _19331_);
  and g_30013_(_19096_, _19103_, _19333_);
  or g_30014_(_19097_, _19104_, _19334_);
  xor g_30015_(_19222_, _19327_, _19335_);
  xor g_30016_(out[251], _19327_, _19336_);
  and g_30017_(_19333_, _19336_, _19337_);
  or g_30018_(_19334_, _19335_, _19338_);
  and g_30019_(_19331_, _19338_, _19339_);
  or g_30020_(_19330_, _19337_, _19340_);
  and g_30021_(_19334_, _19335_, _19341_);
  or g_30022_(_19333_, _19336_, _19342_);
  and g_30023_(_19316_, _19329_, _19344_);
  or g_30024_(_19315_, _19328_, _19345_);
  and g_30025_(_19342_, _19345_, _19346_);
  or g_30026_(_19341_, _19344_, _19347_);
  xor g_30027_(out[249], _19325_, _19348_);
  not g_30028_(_19348_, _19349_);
  and g_30029_(_19117_, _19308_, _19350_);
  not g_30030_(_19350_, _19351_);
  or g_30031_(_19122_, _19308_, _19352_);
  not g_30032_(_19352_, _19353_);
  and g_30033_(_19351_, _19352_, _19355_);
  or g_30034_(_19350_, _19353_, _19356_);
  and g_30035_(_19349_, _19355_, _19357_);
  or g_30036_(_19348_, _19356_, _19358_);
  and g_30037_(_19339_, _19346_, _19359_);
  or g_30038_(_19340_, _19347_, _19360_);
  and g_30039_(_19358_, _19359_, _19361_);
  or g_30040_(_19357_, _19360_, _19362_);
  xor g_30041_(out[248], _19324_, _19363_);
  xor g_30042_(_19321_, _19324_, _19364_);
  and g_30043_(_19131_, _19308_, _19366_);
  not g_30044_(_19366_, _19367_);
  or g_30045_(_19138_, _19308_, _19368_);
  not g_30046_(_19368_, _19369_);
  and g_30047_(_19367_, _19368_, _19370_);
  or g_30048_(_19366_, _19369_, _19371_);
  and g_30049_(_19364_, _19371_, _19372_);
  or g_30050_(_19363_, _19370_, _19373_);
  and g_30051_(_19348_, _19356_, _19374_);
  or g_30052_(_19349_, _19355_, _19375_);
  and g_30053_(_19363_, _19370_, _19377_);
  or g_30054_(_19364_, _19371_, _19378_);
  and g_30055_(_19375_, _19378_, _19379_);
  or g_30056_(_19374_, _19377_, _19380_);
  and g_30057_(_19373_, _19379_, _19381_);
  or g_30058_(_19372_, _19380_, _19382_);
  and g_30059_(_19361_, _19381_, _19383_);
  or g_30060_(_19362_, _19382_, _19384_);
  xor g_30061_(out[247], _19323_, _19385_);
  xor g_30062_(_19233_, _19323_, _19386_);
  and g_30063_(_19163_, _19308_, _19388_);
  not g_30064_(_19388_, _19389_);
  or g_30065_(_19169_, _19308_, _19390_);
  not g_30066_(_19390_, _19391_);
  and g_30067_(_19389_, _19390_, _19392_);
  or g_30068_(_19388_, _19391_, _19393_);
  and g_30069_(_19385_, _19392_, _19394_);
  or g_30070_(_19385_, _19392_, _19395_);
  xor g_30071_(_19385_, _19392_, _19396_);
  xor g_30072_(_19386_, _19392_, _19397_);
  and g_30073_(_19161_, _19308_, _19399_);
  not g_30074_(_19399_, _19400_);
  or g_30075_(_19158_, _19308_, _19401_);
  not g_30076_(_19401_, _19402_);
  and g_30077_(_19400_, _19401_, _19403_);
  or g_30078_(_19399_, _19402_, _19404_);
  xor g_30079_(out[246], _19322_, _19405_);
  or g_30080_(_19404_, _19405_, _19406_);
  xor g_30081_(_19404_, _19405_, _19407_);
  xor g_30082_(_19403_, _19405_, _19408_);
  and g_30083_(_19396_, _19407_, _19410_);
  or g_30084_(_19397_, _19408_, _19411_);
  xor g_30085_(out[244], _19319_, _19412_);
  not g_30086_(_19412_, _19413_);
  and g_30087_(_19192_, _19308_, _19414_);
  not g_30088_(_19414_, _19415_);
  or g_30089_(_19198_, _19308_, _19416_);
  not g_30090_(_19416_, _19417_);
  and g_30091_(_19415_, _19416_, _19418_);
  or g_30092_(_19414_, _19417_, _19419_);
  or g_30093_(_19412_, _19418_, _19421_);
  xor g_30094_(out[245], _19320_, _19422_);
  not g_30095_(_19422_, _19423_);
  or g_30096_(_19181_, _19309_, _19424_);
  or g_30097_(_19187_, _19308_, _19425_);
  and g_30098_(_19424_, _19425_, _19426_);
  not g_30099_(_19426_, _19427_);
  or g_30100_(_19422_, _19427_, _19428_);
  not g_30101_(_19428_, _19429_);
  and g_30102_(_19421_, _19428_, _19430_);
  or g_30103_(_19413_, _19419_, _19432_);
  or g_30104_(_19423_, _19426_, _19433_);
  and g_30105_(_19432_, _19433_, _19434_);
  and g_30106_(_19430_, _19434_, _19435_);
  xor g_30107_(_19413_, _19418_, _19436_);
  xor g_30108_(_19422_, _19426_, _19437_);
  or g_30109_(_19411_, _19437_, _19438_);
  and g_30110_(_19410_, _19435_, _19439_);
  or g_30111_(_19436_, _19438_, _19440_);
  or g_30112_(out[241], out[242], _19441_);
  xor g_30113_(out[241], out[242], _19443_);
  xor g_30114_(_19277_, out[242], _19444_);
  or g_30115_(_19235_, _19308_, _19445_);
  not g_30116_(_19445_, _19446_);
  and g_30117_(_19231_, _19308_, _19447_);
  not g_30118_(_19447_, _19448_);
  and g_30119_(_19445_, _19448_, _19449_);
  or g_30120_(_19446_, _19447_, _19450_);
  xor g_30121_(out[243], _19317_, _19451_);
  xor g_30122_(_19310_, _19317_, _19452_);
  and g_30123_(_19226_, _19309_, _19454_);
  or g_30124_(_19225_, _19308_, _19455_);
  and g_30125_(_19219_, _19308_, _19456_);
  or g_30126_(_19218_, _19309_, _19457_);
  and g_30127_(_19455_, _19457_, _19458_);
  or g_30128_(_19454_, _19456_, _19459_);
  and g_30129_(_19452_, _19458_, _19460_);
  or g_30130_(_19443_, _19450_, _19461_);
  or g_30131_(_19452_, _19458_, _19462_);
  xor g_30132_(_19444_, _19449_, _19463_);
  xor g_30133_(_19443_, _19449_, _19465_);
  xor g_30134_(_19452_, _19458_, _19466_);
  xor g_30135_(_19451_, _19458_, _19467_);
  and g_30136_(_19463_, _19466_, _19468_);
  or g_30137_(_19465_, _19467_, _19469_);
  and g_30138_(out[225], _19308_, _19470_);
  not g_30139_(_19470_, _19471_);
  or g_30140_(_19245_, _19308_, _19472_);
  not g_30141_(_19472_, _19473_);
  and g_30142_(_19471_, _19472_, _19474_);
  or g_30143_(_19470_, _19473_, _19476_);
  or g_30144_(_19277_, _19476_, _19477_);
  or g_30145_(out[241], _19474_, _19478_);
  or g_30146_(_19251_, _19308_, _19479_);
  not g_30147_(_19479_, _19480_);
  and g_30148_(_19156_, _19308_, _19481_);
  not g_30149_(_19481_, _19482_);
  and g_30150_(_19479_, _19482_, _19483_);
  or g_30151_(_19480_, _19481_, _19484_);
  and g_30152_(out[240], _19484_, _19485_);
  or g_30153_(_19288_, _19483_, _19487_);
  and g_30154_(_19478_, _19487_, _19488_);
  and g_30155_(_19477_, _19488_, _19489_);
  xor g_30156_(_19277_, _19474_, _19490_);
  or g_30157_(_19469_, _19485_, _19491_);
  and g_30158_(_19468_, _19489_, _19492_);
  or g_30159_(_19490_, _19491_, _19493_);
  and g_30160_(_19439_, _19492_, _19494_);
  or g_30161_(out[240], _19484_, _19495_);
  and g_30162_(_19383_, _19495_, _19496_);
  and g_30163_(_19494_, _19496_, _19498_);
  or g_30164_(_19469_, _19477_, _19499_);
  or g_30165_(_19460_, _19461_, _19500_);
  and g_30166_(_19462_, _19500_, _19501_);
  and g_30167_(_19499_, _19501_, _19502_);
  or g_30168_(_19411_, _19434_, _19503_);
  or g_30169_(_19429_, _19503_, _19504_);
  or g_30170_(_19394_, _19406_, _19505_);
  and g_30171_(_19395_, _19505_, _19506_);
  and g_30172_(_19504_, _19506_, _19507_);
  and g_30173_(_19493_, _19502_, _19509_);
  or g_30174_(_19440_, _19509_, _19510_);
  and g_30175_(_19507_, _19510_, _19511_);
  or g_30176_(_19384_, _19511_, _19512_);
  and g_30177_(_19361_, _19380_, _19513_);
  and g_30178_(_19340_, _19342_, _19514_);
  or g_30179_(_19513_, _19514_, _19515_);
  not g_30180_(_19515_, _19516_);
  and g_30181_(_19512_, _19516_, _19517_);
  or g_30182_(_19498_, _19517_, _19518_);
  not g_30183_(_19518_, _19520_);
  and g_30184_(_19316_, _19518_, _19521_);
  or g_30185_(_19315_, _19520_, _19522_);
  and g_30186_(_19328_, _19520_, _19523_);
  or g_30187_(_19329_, _19518_, _19524_);
  and g_30188_(_19522_, _19524_, _19525_);
  or g_30189_(_19521_, _19523_, _19526_);
  and g_30190_(out[257], out[258], _19527_);
  or g_30191_(out[260], out[259], _19528_);
  or g_30192_(out[259], _19527_, _19529_);
  or g_30193_(_19527_, _19528_, _19531_);
  or g_30194_(out[261], _19531_, _19532_);
  and g_30195_(out[262], _19532_, _19533_);
  and g_30196_(out[263], _19533_, _19534_);
  or g_30197_(out[264], _19534_, _19535_);
  or g_30198_(out[265], _19535_, _19536_);
  or g_30199_(out[266], _19536_, _19537_);
  xor g_30200_(out[266], _19536_, _19538_);
  not g_30201_(_19538_, _19539_);
  and g_30202_(_19525_, _19538_, _19540_);
  or g_30203_(_19526_, _19539_, _19542_);
  and g_30204_(_19333_, _19335_, _19543_);
  or g_30205_(_19334_, _19336_, _19544_);
  xor g_30206_(_19354_, _19537_, _19545_);
  xor g_30207_(out[267], _19537_, _19546_);
  and g_30208_(_19543_, _19546_, _19547_);
  or g_30209_(_19540_, _19547_, _19548_);
  xor g_30210_(out[265], _19535_, _19549_);
  xor g_30211_(_19464_, _19535_, _19550_);
  or g_30212_(_19348_, _19518_, _19551_);
  not g_30213_(_19551_, _19553_);
  and g_30214_(_19356_, _19518_, _19554_);
  or g_30215_(_19355_, _19520_, _19555_);
  and g_30216_(_19551_, _19555_, _19556_);
  or g_30217_(_19553_, _19554_, _19557_);
  and g_30218_(_19550_, _19556_, _19558_);
  or g_30219_(_19549_, _19557_, _19559_);
  and g_30220_(_19526_, _19539_, _19560_);
  or g_30221_(_19525_, _19538_, _19561_);
  and g_30222_(_19544_, _19545_, _19562_);
  or g_30223_(_19543_, _19546_, _19564_);
  or g_30224_(_19560_, _19562_, _19565_);
  or g_30225_(_19558_, _19565_, _19566_);
  and g_30226_(_19559_, _19561_, _19567_);
  xor g_30227_(_19544_, _19545_, _19568_);
  and g_30228_(_19542_, _19568_, _19569_);
  and g_30229_(_19567_, _19569_, _19570_);
  or g_30230_(_19548_, _19566_, _19571_);
  xor g_30231_(out[264], _19534_, _19572_);
  not g_30232_(_19572_, _19573_);
  and g_30233_(_19363_, _19520_, _19575_);
  or g_30234_(_19364_, _19518_, _19576_);
  and g_30235_(_19371_, _19518_, _19577_);
  or g_30236_(_19370_, _19520_, _19578_);
  and g_30237_(_19576_, _19578_, _19579_);
  or g_30238_(_19575_, _19577_, _19580_);
  and g_30239_(_19573_, _19580_, _19581_);
  or g_30240_(_19572_, _19579_, _19582_);
  and g_30241_(_19572_, _19579_, _19583_);
  or g_30242_(_19573_, _19580_, _19584_);
  and g_30243_(_19549_, _19557_, _19586_);
  or g_30244_(_19550_, _19556_, _19587_);
  and g_30245_(_19584_, _19587_, _19588_);
  or g_30246_(_19583_, _19586_, _19589_);
  and g_30247_(_19582_, _19588_, _19590_);
  or g_30248_(_19581_, _19589_, _19591_);
  and g_30249_(_19570_, _19590_, _19592_);
  or g_30250_(_19571_, _19591_, _19593_);
  xor g_30251_(out[262], _19532_, _19594_);
  xor g_30252_(_19376_, _19532_, _19595_);
  or g_30253_(_19405_, _19518_, _19597_);
  or g_30254_(_19403_, _19520_, _19598_);
  and g_30255_(_19597_, _19598_, _19599_);
  not g_30256_(_19599_, _19600_);
  and g_30257_(_19595_, _19599_, _19601_);
  or g_30258_(_19594_, _19600_, _19602_);
  xor g_30259_(out[263], _19533_, _19603_);
  not g_30260_(_19603_, _19604_);
  and g_30261_(_19385_, _19520_, _19605_);
  or g_30262_(_19386_, _19518_, _19606_);
  and g_30263_(_19393_, _19518_, _19608_);
  or g_30264_(_19392_, _19520_, _19609_);
  and g_30265_(_19606_, _19609_, _19610_);
  or g_30266_(_19605_, _19608_, _19611_);
  and g_30267_(_19604_, _19611_, _19612_);
  or g_30268_(_19603_, _19610_, _19613_);
  and g_30269_(_19602_, _19613_, _19614_);
  or g_30270_(_19601_, _19612_, _19615_);
  and g_30271_(_19594_, _19600_, _19616_);
  or g_30272_(_19595_, _19599_, _19617_);
  and g_30273_(_19603_, _19610_, _19619_);
  or g_30274_(_19604_, _19611_, _19620_);
  xor g_30275_(out[261], _19531_, _19621_);
  xor g_30276_(_19387_, _19531_, _19622_);
  or g_30277_(_19422_, _19518_, _19623_);
  not g_30278_(_19623_, _19624_);
  and g_30279_(_19427_, _19518_, _19625_);
  or g_30280_(_19426_, _19520_, _19626_);
  and g_30281_(_19623_, _19626_, _19627_);
  or g_30282_(_19624_, _19625_, _19628_);
  and g_30283_(_19622_, _19627_, _19630_);
  or g_30284_(_19621_, _19628_, _19631_);
  and g_30285_(_19620_, _19631_, _19632_);
  or g_30286_(_19619_, _19630_, _19633_);
  and g_30287_(_19617_, _19632_, _19634_);
  or g_30288_(_19616_, _19633_, _19635_);
  and g_30289_(_19614_, _19634_, _19636_);
  or g_30290_(_19615_, _19635_, _19637_);
  xor g_30291_(out[260], _19529_, _19638_);
  not g_30292_(_19638_, _19639_);
  and g_30293_(_19412_, _19520_, _19641_);
  or g_30294_(_19413_, _19518_, _19642_);
  and g_30295_(_19419_, _19518_, _19643_);
  or g_30296_(_19418_, _19520_, _19644_);
  and g_30297_(_19642_, _19644_, _19645_);
  or g_30298_(_19641_, _19643_, _19646_);
  and g_30299_(_19639_, _19646_, _19647_);
  or g_30300_(_19638_, _19645_, _19648_);
  and g_30301_(_19621_, _19628_, _19649_);
  or g_30302_(_19622_, _19627_, _19650_);
  and g_30303_(_19638_, _19645_, _19652_);
  or g_30304_(_19639_, _19646_, _19653_);
  and g_30305_(_19650_, _19653_, _19654_);
  or g_30306_(_19649_, _19652_, _19655_);
  and g_30307_(_19648_, _19654_, _19656_);
  or g_30308_(_19647_, _19655_, _19657_);
  and g_30309_(_19636_, _19656_, _19658_);
  or g_30310_(_19637_, _19657_, _19659_);
  and g_30311_(_19592_, _19658_, _19660_);
  or g_30312_(_19593_, _19659_, _19661_);
  xor g_30313_(out[259], _19527_, _19663_);
  xor g_30314_(_19442_, _19527_, _19664_);
  and g_30315_(_19459_, _19518_, _19665_);
  or g_30316_(_19458_, _19520_, _19666_);
  or g_30317_(_19451_, _19518_, _19667_);
  not g_30318_(_19667_, _19668_);
  and g_30319_(_19666_, _19667_, _19669_);
  or g_30320_(_19665_, _19668_, _19670_);
  and g_30321_(_19663_, _19670_, _19671_);
  or g_30322_(out[257], out[258], _19672_);
  xor g_30323_(out[257], out[258], _19674_);
  xor g_30324_(_19409_, out[258], _19675_);
  or g_30325_(_19443_, _19518_, _19676_);
  or g_30326_(_19449_, _19520_, _19677_);
  and g_30327_(_19676_, _19677_, _19678_);
  and g_30328_(_19675_, _19678_, _19679_);
  or g_30329_(_19671_, _19679_, _19680_);
  or g_30330_(_19663_, _19670_, _19681_);
  xor g_30331_(_19664_, _19669_, _19682_);
  xor g_30332_(_19663_, _19669_, _19683_);
  xor g_30333_(_19675_, _19678_, _19685_);
  xor g_30334_(_19674_, _19678_, _19686_);
  and g_30335_(_19682_, _19685_, _19687_);
  or g_30336_(_19683_, _19686_, _19688_);
  or g_30337_(_19277_, _19518_, _19689_);
  or g_30338_(_19474_, _19520_, _19690_);
  and g_30339_(_19689_, _19690_, _19691_);
  and g_30340_(out[257], _19691_, _19692_);
  or g_30341_(_19483_, _19520_, _19693_);
  or g_30342_(out[240], _19518_, _19694_);
  and g_30343_(_19693_, _19694_, _19696_);
  not g_30344_(_19696_, _19697_);
  and g_30345_(out[256], _19697_, _19698_);
  or g_30346_(_19420_, _19696_, _19699_);
  xor g_30347_(out[257], _19691_, _19700_);
  xor g_30348_(_19409_, _19691_, _19701_);
  and g_30349_(_19699_, _19700_, _19702_);
  or g_30350_(_19698_, _19701_, _19703_);
  or g_30351_(_19692_, _19702_, _19704_);
  and g_30352_(_19687_, _19704_, _19705_);
  and g_30353_(_19680_, _19681_, _19707_);
  or g_30354_(_19705_, _19707_, _19708_);
  not g_30355_(_19708_, _19709_);
  and g_30356_(_19660_, _19708_, _19710_);
  or g_30357_(_19661_, _19709_, _19711_);
  and g_30358_(_19615_, _19620_, _19712_);
  or g_30359_(_19614_, _19619_, _19713_);
  and g_30360_(_19636_, _19655_, _19714_);
  or g_30361_(_19637_, _19654_, _19715_);
  and g_30362_(_19713_, _19715_, _19716_);
  or g_30363_(_19712_, _19714_, _19718_);
  and g_30364_(_19592_, _19718_, _19719_);
  or g_30365_(_19593_, _19716_, _19720_);
  and g_30366_(_19570_, _19589_, _19721_);
  and g_30367_(_19548_, _19564_, _19722_);
  or g_30368_(_19721_, _19722_, _19723_);
  not g_30369_(_19723_, _19724_);
  and g_30370_(_19720_, _19724_, _19725_);
  or g_30371_(_19719_, _19723_, _19726_);
  and g_30372_(_19711_, _19725_, _19727_);
  or g_30373_(_19710_, _19726_, _19729_);
  and g_30374_(_19420_, _19696_, _19730_);
  or g_30375_(out[256], _19697_, _19731_);
  and g_30376_(_19687_, _19731_, _19732_);
  or g_30377_(_19688_, _19730_, _19733_);
  and g_30378_(_19702_, _19732_, _19734_);
  or g_30379_(_19703_, _19733_, _19735_);
  and g_30380_(_19660_, _19734_, _19736_);
  or g_30381_(_19661_, _19735_, _19737_);
  and g_30382_(_19729_, _19737_, _19738_);
  or g_30383_(_19727_, _19736_, _19740_);
  or g_30384_(_19525_, _19738_, _19741_);
  not g_30385_(_19741_, _19742_);
  and g_30386_(_19538_, _19738_, _19743_);
  not g_30387_(_19743_, _19744_);
  and g_30388_(_19741_, _19744_, _19745_);
  or g_30389_(_19742_, _19743_, _19746_);
  and g_30390_(out[273], out[274], _19747_);
  or g_30391_(out[276], out[275], _19748_);
  or g_30392_(out[275], _19747_, _19749_);
  or g_30393_(_19747_, _19748_, _19751_);
  or g_30394_(out[277], _19751_, _19752_);
  and g_30395_(out[278], _19752_, _19753_);
  and g_30396_(out[279], _19753_, _19754_);
  or g_30397_(out[280], _19754_, _19755_);
  or g_30398_(out[281], _19755_, _19756_);
  or g_30399_(out[282], _19756_, _19757_);
  xor g_30400_(out[282], _19756_, _19758_);
  not g_30401_(_19758_, _19759_);
  and g_30402_(_19745_, _19758_, _19760_);
  or g_30403_(_19746_, _19759_, _19762_);
  and g_30404_(_19543_, _19545_, _19763_);
  or g_30405_(_19544_, _19546_, _19764_);
  xor g_30406_(_19486_, _19757_, _19765_);
  xor g_30407_(out[283], _19757_, _19766_);
  and g_30408_(_19763_, _19766_, _19767_);
  or g_30409_(_19764_, _19765_, _19768_);
  and g_30410_(_19762_, _19768_, _19769_);
  or g_30411_(_19760_, _19767_, _19770_);
  and g_30412_(_19764_, _19765_, _19771_);
  or g_30413_(_19763_, _19766_, _19773_);
  or g_30414_(_19745_, _19758_, _19774_);
  and g_30415_(_19773_, _19774_, _19775_);
  xor g_30416_(out[281], _19755_, _19776_);
  not g_30417_(_19776_, _19777_);
  and g_30418_(_19550_, _19738_, _19778_);
  not g_30419_(_19778_, _19779_);
  or g_30420_(_19556_, _19738_, _19780_);
  not g_30421_(_19780_, _19781_);
  and g_30422_(_19779_, _19780_, _19782_);
  or g_30423_(_19778_, _19781_, _19784_);
  or g_30424_(_19776_, _19784_, _19785_);
  and g_30425_(_19775_, _19785_, _19786_);
  not g_30426_(_19786_, _19787_);
  and g_30427_(_19769_, _19786_, _19788_);
  or g_30428_(_19770_, _19787_, _19789_);
  xor g_30429_(out[280], _19754_, _19790_);
  not g_30430_(_19790_, _19791_);
  and g_30431_(_19572_, _19738_, _19792_);
  not g_30432_(_19792_, _19793_);
  or g_30433_(_19579_, _19738_, _19795_);
  not g_30434_(_19795_, _19796_);
  and g_30435_(_19793_, _19795_, _19797_);
  or g_30436_(_19792_, _19796_, _19798_);
  and g_30437_(_19790_, _19797_, _19799_);
  or g_30438_(_19791_, _19798_, _19800_);
  and g_30439_(_19776_, _19784_, _19801_);
  or g_30440_(_19777_, _19782_, _19802_);
  and g_30441_(_19800_, _19802_, _19803_);
  or g_30442_(_19799_, _19801_, _19804_);
  xor g_30443_(out[278], _19752_, _19806_);
  and g_30444_(_19595_, _19738_, _19807_);
  not g_30445_(_19807_, _19808_);
  or g_30446_(_19599_, _19738_, _19809_);
  not g_30447_(_19809_, _19810_);
  and g_30448_(_19808_, _19809_, _19811_);
  or g_30449_(_19807_, _19810_, _19812_);
  or g_30450_(_19806_, _19812_, _19813_);
  xor g_30451_(out[279], _19753_, _19814_);
  and g_30452_(_19603_, _19738_, _19815_);
  not g_30453_(_19815_, _19817_);
  or g_30454_(_19610_, _19738_, _19818_);
  not g_30455_(_19818_, _19819_);
  and g_30456_(_19817_, _19818_, _19820_);
  or g_30457_(_19815_, _19819_, _19821_);
  or g_30458_(_19814_, _19820_, _19822_);
  and g_30459_(_19813_, _19822_, _19823_);
  and g_30460_(_19814_, _19820_, _19824_);
  xor g_30461_(_19806_, _19812_, _19825_);
  xor g_30462_(_19806_, _19811_, _19826_);
  xor g_30463_(_19814_, _19820_, _19828_);
  xor g_30464_(_19814_, _19821_, _19829_);
  and g_30465_(_19825_, _19828_, _19830_);
  or g_30466_(_19826_, _19829_, _19831_);
  xor g_30467_(out[276], _19749_, _19832_);
  not g_30468_(_19832_, _19833_);
  and g_30469_(_19638_, _19738_, _19834_);
  not g_30470_(_19834_, _19835_);
  or g_30471_(_19645_, _19738_, _19836_);
  not g_30472_(_19836_, _19837_);
  and g_30473_(_19835_, _19836_, _19839_);
  or g_30474_(_19834_, _19837_, _19840_);
  and g_30475_(_19832_, _19839_, _19841_);
  or g_30476_(_19833_, _19840_, _19842_);
  xor g_30477_(out[277], _19751_, _19843_);
  not g_30478_(_19843_, _19844_);
  and g_30479_(_19622_, _19738_, _19845_);
  not g_30480_(_19845_, _19846_);
  or g_30481_(_19627_, _19738_, _19847_);
  not g_30482_(_19847_, _19848_);
  and g_30483_(_19846_, _19847_, _19850_);
  or g_30484_(_19845_, _19848_, _19851_);
  and g_30485_(_19843_, _19851_, _19852_);
  or g_30486_(_19844_, _19850_, _19853_);
  and g_30487_(_19842_, _19853_, _19854_);
  or g_30488_(_19841_, _19852_, _19855_);
  and g_30489_(_19844_, _19850_, _19856_);
  or g_30490_(_19843_, _19851_, _19857_);
  and g_30491_(_19833_, _19840_, _19858_);
  or g_30492_(_19832_, _19839_, _19859_);
  and g_30493_(_19857_, _19859_, _19861_);
  or g_30494_(_19856_, _19858_, _19862_);
  and g_30495_(_19854_, _19861_, _19863_);
  or g_30496_(_19855_, _19862_, _19864_);
  and g_30497_(_19830_, _19863_, _19865_);
  or g_30498_(_19831_, _19864_, _19866_);
  xor g_30499_(out[275], _19747_, _19867_);
  not g_30500_(_19867_, _19868_);
  and g_30501_(_19670_, _19740_, _19869_);
  or g_30502_(_19669_, _19738_, _19870_);
  and g_30503_(_19664_, _19738_, _19872_);
  or g_30504_(_19663_, _19740_, _19873_);
  and g_30505_(_19870_, _19873_, _19874_);
  or g_30506_(_19869_, _19872_, _19875_);
  and g_30507_(_19868_, _19874_, _19876_);
  or g_30508_(_19867_, _19875_, _19877_);
  and g_30509_(_19675_, _19738_, _19878_);
  not g_30510_(_19878_, _19879_);
  or g_30511_(_19678_, _19738_, _19880_);
  not g_30512_(_19880_, _19881_);
  and g_30513_(_19879_, _19880_, _19883_);
  or g_30514_(_19878_, _19881_, _19884_);
  or g_30515_(out[273], out[274], _19885_);
  xor g_30516_(out[273], out[274], _19886_);
  xor g_30517_(_19541_, out[274], _19887_);
  and g_30518_(_19883_, _19887_, _19888_);
  or g_30519_(_19884_, _19886_, _19889_);
  or g_30520_(_19876_, _19888_, _19890_);
  and g_30521_(_19867_, _19875_, _19891_);
  or g_30522_(_19868_, _19874_, _19892_);
  and g_30523_(_19884_, _19886_, _19894_);
  or g_30524_(_19891_, _19894_, _19895_);
  and g_30525_(_19877_, _19892_, _19896_);
  xor g_30526_(_19884_, _19886_, _19897_);
  and g_30527_(_19896_, _19897_, _19898_);
  or g_30528_(_19890_, _19895_, _19899_);
  and g_30529_(out[257], _19738_, _19900_);
  not g_30530_(_19900_, _19901_);
  or g_30531_(_19691_, _19738_, _19902_);
  not g_30532_(_19902_, _19903_);
  and g_30533_(_19901_, _19902_, _19905_);
  or g_30534_(_19900_, _19903_, _19906_);
  and g_30535_(out[273], _19905_, _19907_);
  or g_30536_(_19541_, _19906_, _19908_);
  and g_30537_(_19898_, _19907_, _19909_);
  or g_30538_(_19899_, _19908_, _19910_);
  and g_30539_(_19889_, _19892_, _19911_);
  or g_30540_(_19888_, _19891_, _19912_);
  and g_30541_(_19877_, _19912_, _19913_);
  or g_30542_(_19876_, _19911_, _19914_);
  and g_30543_(_19910_, _19914_, _19916_);
  or g_30544_(_19909_, _19913_, _19917_);
  and g_30545_(_19865_, _19917_, _19918_);
  or g_30546_(_19866_, _19916_, _19919_);
  or g_30547_(_19823_, _19824_, _19920_);
  not g_30548_(_19920_, _19921_);
  and g_30549_(_19830_, _19855_, _19922_);
  or g_30550_(_19831_, _19854_, _19923_);
  and g_30551_(_19857_, _19922_, _19924_);
  or g_30552_(_19856_, _19923_, _19925_);
  and g_30553_(_19920_, _19925_, _19927_);
  or g_30554_(_19921_, _19924_, _19928_);
  xor g_30555_(out[273], _19905_, _19929_);
  xor g_30556_(_19541_, _19905_, _19930_);
  or g_30557_(_19696_, _19738_, _19931_);
  or g_30558_(out[256], _19740_, _19932_);
  and g_30559_(_19931_, _19932_, _19933_);
  not g_30560_(_19933_, _19934_);
  and g_30561_(out[272], _19934_, _19935_);
  or g_30562_(_19552_, _19933_, _19936_);
  and g_30563_(_19929_, _19936_, _19938_);
  or g_30564_(_19930_, _19935_, _19939_);
  and g_30565_(_19898_, _19938_, _19940_);
  or g_30566_(_19899_, _19939_, _19941_);
  and g_30567_(_19865_, _19940_, _19942_);
  or g_30568_(_19866_, _19941_, _19943_);
  and g_30569_(_19927_, _19943_, _19944_);
  or g_30570_(_19918_, _19928_, _19945_);
  and g_30571_(_19919_, _19944_, _19946_);
  or g_30572_(_19942_, _19945_, _19947_);
  and g_30573_(_19791_, _19798_, _19949_);
  or g_30574_(_19790_, _19797_, _19950_);
  and g_30575_(_19947_, _19950_, _19951_);
  or g_30576_(_19946_, _19949_, _19952_);
  and g_30577_(_19803_, _19952_, _19953_);
  or g_30578_(_19804_, _19951_, _19954_);
  and g_30579_(_19788_, _19954_, _19955_);
  or g_30580_(_19789_, _19953_, _19956_);
  and g_30581_(_19770_, _19773_, _19957_);
  or g_30582_(_19769_, _19771_, _19958_);
  and g_30583_(_19956_, _19958_, _19960_);
  or g_30584_(_19955_, _19957_, _19961_);
  and g_30585_(_19552_, _19933_, _19962_);
  or g_30586_(out[272], _19934_, _19963_);
  and g_30587_(_19950_, _19963_, _19964_);
  or g_30588_(_19949_, _19962_, _19965_);
  and g_30589_(_19803_, _19964_, _19966_);
  or g_30590_(_19804_, _19965_, _19967_);
  and g_30591_(_19788_, _19966_, _19968_);
  or g_30592_(_19789_, _19967_, _19969_);
  and g_30593_(_19942_, _19968_, _19971_);
  or g_30594_(_19943_, _19969_, _19972_);
  and g_30595_(_19961_, _19972_, _19973_);
  or g_30596_(_19960_, _19971_, _19974_);
  and g_30597_(_19746_, _19974_, _19975_);
  or g_30598_(_19745_, _19973_, _19976_);
  and g_30599_(_19758_, _19973_, _19977_);
  not g_30600_(_19977_, _19978_);
  and g_30601_(_19976_, _19978_, _19979_);
  or g_30602_(_19975_, _19977_, _19980_);
  and g_30603_(out[289], out[290], _19982_);
  or g_30604_(out[292], out[291], _19983_);
  or g_30605_(out[291], _19982_, _19984_);
  or g_30606_(_19982_, _19983_, _19985_);
  or g_30607_(out[293], _19985_, _19986_);
  and g_30608_(out[294], _19986_, _19987_);
  and g_30609_(out[295], _19987_, _19988_);
  or g_30610_(out[296], _19988_, _19989_);
  or g_30611_(out[297], _19989_, _19990_);
  or g_30612_(out[298], _19990_, _19991_);
  xor g_30613_(out[298], _19990_, _19993_);
  not g_30614_(_19993_, _19994_);
  and g_30615_(_19979_, _19993_, _19995_);
  or g_30616_(_19980_, _19994_, _19996_);
  or g_30617_(_19764_, _19766_, _19997_);
  not g_30618_(_19997_, _19998_);
  xor g_30619_(out[299], _19991_, _19999_);
  not g_30620_(_19999_, _20000_);
  and g_30621_(_19998_, _19999_, _20001_);
  or g_30622_(_19997_, _20000_, _20002_);
  and g_30623_(_19996_, _20002_, _20004_);
  or g_30624_(_19995_, _20001_, _20005_);
  or g_30625_(_19998_, _19999_, _20006_);
  or g_30626_(_19979_, _19993_, _20007_);
  and g_30627_(_20006_, _20007_, _20008_);
  and g_30628_(_20004_, _20008_, _20009_);
  not g_30629_(_20009_, _20010_);
  xor g_30630_(out[297], _19989_, _20011_);
  not g_30631_(_20011_, _20012_);
  or g_30632_(_19776_, _19974_, _20013_);
  or g_30633_(_19782_, _19973_, _20015_);
  and g_30634_(_20013_, _20015_, _20016_);
  not g_30635_(_20016_, _20017_);
  and g_30636_(_20011_, _20017_, _20018_);
  or g_30637_(_20012_, _20016_, _20019_);
  xor g_30638_(out[296], _19988_, _20020_);
  not g_30639_(_20020_, _20021_);
  and g_30640_(_19790_, _19973_, _20022_);
  not g_30641_(_20022_, _20023_);
  or g_30642_(_19797_, _19973_, _20024_);
  not g_30643_(_20024_, _20026_);
  and g_30644_(_20023_, _20024_, _20027_);
  or g_30645_(_20022_, _20026_, _20028_);
  and g_30646_(_20020_, _20027_, _20029_);
  or g_30647_(_20021_, _20028_, _20030_);
  and g_30648_(_20019_, _20030_, _20031_);
  or g_30649_(_20018_, _20029_, _20032_);
  or g_30650_(_20020_, _20027_, _20033_);
  or g_30651_(_20011_, _20017_, _20034_);
  and g_30652_(_20033_, _20034_, _20035_);
  not g_30653_(_20035_, _20037_);
  and g_30654_(_20031_, _20035_, _20038_);
  or g_30655_(_20032_, _20037_, _20039_);
  and g_30656_(_20009_, _20038_, _20040_);
  or g_30657_(_20010_, _20039_, _20041_);
  xor g_30658_(out[293], _19985_, _20042_);
  not g_30659_(_20042_, _20043_);
  and g_30660_(_19843_, _19973_, _20044_);
  not g_30661_(_20044_, _20045_);
  and g_30662_(_19850_, _19974_, _20046_);
  or g_30663_(_19851_, _19973_, _20048_);
  or g_30664_(_20044_, _20046_, _20049_);
  and g_30665_(_20045_, _20048_, _20050_);
  or g_30666_(_20042_, _20050_, _20051_);
  xor g_30667_(out[294], _19986_, _20052_);
  not g_30668_(_20052_, _20053_);
  or g_30669_(_19806_, _19974_, _20054_);
  or g_30670_(_19811_, _19973_, _20055_);
  and g_30671_(_20054_, _20055_, _20056_);
  not g_30672_(_20056_, _20057_);
  or g_30673_(_20053_, _20056_, _20059_);
  and g_30674_(_20051_, _20059_, _20060_);
  xor g_30675_(out[295], _19987_, _20061_);
  not g_30676_(_20061_, _20062_);
  and g_30677_(_19814_, _19973_, _20063_);
  not g_30678_(_20063_, _20064_);
  or g_30679_(_19820_, _19973_, _20065_);
  not g_30680_(_20065_, _20066_);
  and g_30681_(_20064_, _20065_, _20067_);
  or g_30682_(_20063_, _20066_, _20068_);
  and g_30683_(_20061_, _20067_, _20070_);
  or g_30684_(_20062_, _20068_, _20071_);
  xor g_30685_(out[292], _19984_, _20072_);
  not g_30686_(_20072_, _20073_);
  and g_30687_(_19832_, _19973_, _20074_);
  not g_30688_(_20074_, _20075_);
  or g_30689_(_19839_, _19973_, _20076_);
  not g_30690_(_20076_, _20077_);
  and g_30691_(_20075_, _20076_, _20078_);
  or g_30692_(_20074_, _20077_, _20079_);
  or g_30693_(_20072_, _20078_, _20081_);
  and g_30694_(_20071_, _20081_, _20082_);
  and g_30695_(_20060_, _20082_, _20083_);
  or g_30696_(_20052_, _20057_, _20084_);
  or g_30697_(_20061_, _20067_, _20085_);
  and g_30698_(_20084_, _20085_, _20086_);
  and g_30699_(_20072_, _20078_, _20087_);
  or g_30700_(_20073_, _20079_, _20088_);
  and g_30701_(_20042_, _20050_, _20089_);
  or g_30702_(_20043_, _20049_, _20090_);
  and g_30703_(_20088_, _20090_, _20092_);
  or g_30704_(_20087_, _20089_, _20093_);
  and g_30705_(_20086_, _20092_, _20094_);
  and g_30706_(_20083_, _20094_, _20095_);
  and g_30707_(_20040_, _20095_, _20096_);
  xor g_30708_(out[291], _19982_, _20097_);
  and g_30709_(_19868_, _19973_, _20098_);
  and g_30710_(_19875_, _19974_, _20099_);
  or g_30711_(_20098_, _20099_, _20100_);
  and g_30712_(_20097_, _20100_, _20101_);
  or g_30713_(_19883_, _19973_, _20103_);
  or g_30714_(_19886_, _19974_, _20104_);
  and g_30715_(_20103_, _20104_, _20105_);
  or g_30716_(out[289], out[290], _20106_);
  xor g_30717_(out[289], out[290], _20107_);
  xor g_30718_(_19673_, out[290], _20108_);
  and g_30719_(_20105_, _20108_, _20109_);
  or g_30720_(_20101_, _20109_, _20110_);
  or g_30721_(_20097_, _20100_, _20111_);
  xor g_30722_(_20097_, _20100_, _20112_);
  xor g_30723_(_20105_, _20108_, _20114_);
  and g_30724_(_20112_, _20114_, _20115_);
  or g_30725_(_19905_, _19973_, _20116_);
  not g_30726_(_20116_, _20117_);
  and g_30727_(out[273], _19973_, _20118_);
  not g_30728_(_20118_, _20119_);
  and g_30729_(_20116_, _20119_, _20120_);
  or g_30730_(_20117_, _20118_, _20121_);
  and g_30731_(out[289], _20120_, _20122_);
  or g_30732_(_19933_, _19973_, _20123_);
  or g_30733_(out[272], _19974_, _20125_);
  and g_30734_(_20123_, _20125_, _20126_);
  or g_30735_(_18573_, _20126_, _20127_);
  xor g_30736_(out[289], _20120_, _20128_);
  and g_30737_(_20127_, _20128_, _20129_);
  or g_30738_(_20122_, _20129_, _20130_);
  and g_30739_(_20115_, _20130_, _20131_);
  and g_30740_(_20110_, _20111_, _20132_);
  or g_30741_(_20131_, _20132_, _20133_);
  and g_30742_(_20096_, _20133_, _20134_);
  and g_30743_(_20060_, _20093_, _20136_);
  not g_30744_(_20136_, _20137_);
  and g_30745_(_20086_, _20137_, _20138_);
  or g_30746_(_20070_, _20138_, _20139_);
  or g_30747_(_20041_, _20139_, _20140_);
  not g_30748_(_20140_, _20141_);
  and g_30749_(_20005_, _20006_, _20142_);
  and g_30750_(_20032_, _20034_, _20143_);
  and g_30751_(_20009_, _20143_, _20144_);
  or g_30752_(_20142_, _20144_, _20145_);
  or g_30753_(_20134_, _20145_, _20147_);
  or g_30754_(_20141_, _20147_, _20148_);
  and g_30755_(_18573_, _20126_, _20149_);
  and g_30756_(_20115_, _20129_, _20150_);
  and g_30757_(_20096_, _20150_, _20151_);
  not g_30758_(_20151_, _20152_);
  or g_30759_(_20149_, _20152_, _20153_);
  and g_30760_(_20148_, _20153_, _20154_);
  not g_30761_(_20154_, _20155_);
  or g_30762_(_19979_, _20154_, _20156_);
  not g_30763_(_20156_, _20158_);
  and g_30764_(_19993_, _20154_, _20159_);
  not g_30765_(_20159_, _20160_);
  and g_30766_(_20156_, _20160_, _20161_);
  or g_30767_(_20158_, _20159_, _20162_);
  and g_30768_(_18419_, _20161_, _20163_);
  or g_30769_(_18420_, _20162_, _20164_);
  or g_30770_(_19997_, _19999_, _20165_);
  not g_30771_(_20165_, _20166_);
  xor g_30772_(out[315], _18418_, _20167_);
  not g_30773_(_20167_, _20169_);
  and g_30774_(_20166_, _20167_, _20170_);
  or g_30775_(_20165_, _20169_, _20171_);
  and g_30776_(_20164_, _20171_, _20172_);
  or g_30777_(_20163_, _20170_, _20173_);
  and g_30778_(_20165_, _20169_, _20174_);
  or g_30779_(_20166_, _20167_, _20175_);
  and g_30780_(_18420_, _20162_, _20176_);
  or g_30781_(_18419_, _20161_, _20177_);
  and g_30782_(_20175_, _20177_, _20178_);
  or g_30783_(_20174_, _20176_, _20180_);
  and g_30784_(_20172_, _20178_, _20181_);
  or g_30785_(_20173_, _20180_, _20182_);
  or g_30786_(_20011_, _20155_, _20183_);
  or g_30787_(_20016_, _20154_, _20184_);
  and g_30788_(_20183_, _20184_, _20185_);
  not g_30789_(_20185_, _20186_);
  and g_30790_(_18416_, _20186_, _20187_);
  or g_30791_(_18417_, _20185_, _20188_);
  and g_30792_(_20020_, _20154_, _20189_);
  not g_30793_(_20189_, _20191_);
  and g_30794_(_20028_, _20155_, _20192_);
  or g_30795_(_20027_, _20154_, _20193_);
  and g_30796_(_20191_, _20193_, _20194_);
  or g_30797_(_20189_, _20192_, _20195_);
  xor g_30798_(out[312], _18413_, _20196_);
  xor g_30799_(_19827_, _18413_, _20197_);
  and g_30800_(_20194_, _20196_, _20198_);
  or g_30801_(_20195_, _20197_, _20199_);
  and g_30802_(_20188_, _20199_, _20200_);
  or g_30803_(_20187_, _20198_, _20202_);
  and g_30804_(_20195_, _20197_, _20203_);
  or g_30805_(_20194_, _20196_, _20204_);
  and g_30806_(_18417_, _20185_, _20205_);
  or g_30807_(_18416_, _20186_, _20206_);
  and g_30808_(_20204_, _20206_, _20207_);
  or g_30809_(_20203_, _20205_, _20208_);
  and g_30810_(_20200_, _20207_, _20209_);
  or g_30811_(_20202_, _20208_, _20210_);
  and g_30812_(_20181_, _20209_, _20211_);
  or g_30813_(_20182_, _20210_, _20213_);
  xor g_30814_(out[310], _18411_, _20214_);
  not g_30815_(_20214_, _20215_);
  or g_30816_(_20052_, _20155_, _20216_);
  or g_30817_(_20056_, _20154_, _20217_);
  and g_30818_(_20216_, _20217_, _20218_);
  and g_30819_(_20215_, _20218_, _20219_);
  xor g_30820_(out[311], _18412_, _20220_);
  xor g_30821_(_19750_, _18412_, _20221_);
  and g_30822_(_20061_, _20154_, _20222_);
  and g_30823_(_20068_, _20155_, _20224_);
  or g_30824_(_20222_, _20224_, _20225_);
  not g_30825_(_20225_, _20226_);
  and g_30826_(_20221_, _20225_, _20227_);
  or g_30827_(_20219_, _20227_, _20228_);
  or g_30828_(_20221_, _20225_, _20229_);
  xor g_30829_(_20215_, _20218_, _20230_);
  xor g_30830_(_20214_, _20218_, _20231_);
  xor g_30831_(_20221_, _20225_, _20232_);
  xor g_30832_(_20220_, _20225_, _20233_);
  and g_30833_(_20230_, _20232_, _20235_);
  or g_30834_(_20231_, _20233_, _20236_);
  xor g_30835_(out[309], _18410_, _20237_);
  xor g_30836_(_19783_, _18410_, _20238_);
  or g_30837_(_20050_, _20154_, _20239_);
  not g_30838_(_20239_, _20240_);
  and g_30839_(_20042_, _20154_, _20241_);
  not g_30840_(_20241_, _20242_);
  or g_30841_(_20240_, _20241_, _20243_);
  and g_30842_(_20239_, _20242_, _20244_);
  and g_30843_(_20237_, _20244_, _20246_);
  or g_30844_(_20238_, _20243_, _20247_);
  and g_30845_(_20072_, _20154_, _20248_);
  not g_30846_(_20248_, _20249_);
  and g_30847_(_20079_, _20155_, _20250_);
  or g_30848_(_20078_, _20154_, _20251_);
  and g_30849_(_20249_, _20251_, _20252_);
  or g_30850_(_20248_, _20250_, _20253_);
  xor g_30851_(out[308], _18409_, _20254_);
  xor g_30852_(_19772_, _18409_, _20255_);
  and g_30853_(_20252_, _20254_, _20257_);
  or g_30854_(_20253_, _20255_, _20258_);
  and g_30855_(_20247_, _20258_, _20259_);
  or g_30856_(_20246_, _20257_, _20260_);
  and g_30857_(_20238_, _20243_, _20261_);
  or g_30858_(_20237_, _20244_, _20262_);
  and g_30859_(_20253_, _20255_, _20263_);
  or g_30860_(_20252_, _20254_, _20264_);
  and g_30861_(_20262_, _20264_, _20265_);
  or g_30862_(_20261_, _20263_, _20266_);
  and g_30863_(_20259_, _20265_, _20268_);
  or g_30864_(_20260_, _20266_, _20269_);
  and g_30865_(_20235_, _20268_, _20270_);
  or g_30866_(_20236_, _20269_, _20271_);
  xor g_30867_(out[307], _18407_, _20272_);
  xor g_30868_(_19816_, _18407_, _20273_);
  and g_30869_(_20097_, _20154_, _20274_);
  not g_30870_(_20274_, _20275_);
  or g_30871_(_20100_, _20154_, _20276_);
  not g_30872_(_20276_, _20277_);
  or g_30873_(_20274_, _20277_, _20279_);
  and g_30874_(_20275_, _20276_, _20280_);
  and g_30875_(_20273_, _20279_, _20281_);
  or g_30876_(_20272_, _20280_, _20282_);
  and g_30877_(_20272_, _20280_, _20283_);
  or g_30878_(_20273_, _20279_, _20284_);
  or g_30879_(_20105_, _20154_, _20285_);
  not g_30880_(_20285_, _20286_);
  and g_30881_(_20108_, _20154_, _20287_);
  not g_30882_(_20287_, _20288_);
  and g_30883_(_20285_, _20288_, _20290_);
  or g_30884_(_20286_, _20287_, _20291_);
  or g_30885_(out[305], out[306], _20292_);
  xor g_30886_(out[305], out[306], _20293_);
  xor g_30887_(_19794_, out[306], _20294_);
  and g_30888_(_20290_, _20294_, _20295_);
  or g_30889_(_20291_, _20293_, _20296_);
  and g_30890_(_20284_, _20296_, _20297_);
  or g_30891_(_20283_, _20295_, _20298_);
  and g_30892_(_20282_, _20298_, _20299_);
  or g_30893_(_20281_, _20297_, _20301_);
  and g_30894_(_20282_, _20284_, _20302_);
  or g_30895_(_20281_, _20283_, _20303_);
  xor g_30896_(_20291_, _20293_, _20304_);
  xor g_30897_(_20290_, _20293_, _20305_);
  and g_30898_(_20302_, _20304_, _20306_);
  or g_30899_(_20303_, _20305_, _20307_);
  and g_30900_(out[289], _20154_, _20308_);
  and g_30901_(_20121_, _20155_, _20309_);
  or g_30902_(_20308_, _20309_, _20310_);
  not g_30903_(_20310_, _20312_);
  and g_30904_(out[305], _20312_, _20313_);
  or g_30905_(_19794_, _20310_, _20314_);
  or g_30906_(_20126_, _20154_, _20315_);
  or g_30907_(out[288], _20155_, _20316_);
  and g_30908_(_20315_, _20316_, _20317_);
  not g_30909_(_20317_, _20318_);
  and g_30910_(out[304], _20318_, _20319_);
  or g_30911_(_18562_, _20317_, _20320_);
  xor g_30912_(_19794_, _20310_, _20321_);
  xor g_30913_(out[305], _20310_, _20323_);
  and g_30914_(_20320_, _20321_, _20324_);
  or g_30915_(_20319_, _20323_, _20325_);
  and g_30916_(_20306_, _20324_, _20326_);
  or g_30917_(_20307_, _20325_, _20327_);
  and g_30918_(_20306_, _20313_, _20328_);
  or g_30919_(_20307_, _20314_, _20329_);
  and g_30920_(_20301_, _20329_, _20330_);
  or g_30921_(_20299_, _20328_, _20331_);
  and g_30922_(_20327_, _20330_, _20332_);
  or g_30923_(_20326_, _20331_, _20334_);
  and g_30924_(_20270_, _20334_, _20335_);
  or g_30925_(_20271_, _20332_, _20336_);
  and g_30926_(_20228_, _20229_, _20337_);
  not g_30927_(_20337_, _20338_);
  and g_30928_(_20235_, _20260_, _20339_);
  or g_30929_(_20236_, _20259_, _20340_);
  and g_30930_(_20262_, _20339_, _20341_);
  or g_30931_(_20261_, _20340_, _20342_);
  and g_30932_(_20338_, _20342_, _20343_);
  or g_30933_(_20337_, _20341_, _20345_);
  and g_30934_(_20336_, _20343_, _20346_);
  or g_30935_(_20335_, _20345_, _20347_);
  and g_30936_(_20211_, _20347_, _20348_);
  or g_30937_(_20213_, _20346_, _20349_);
  or g_30938_(_20200_, _20205_, _20350_);
  and g_30939_(_20181_, _20202_, _20351_);
  and g_30940_(_20206_, _20351_, _20352_);
  or g_30941_(_20182_, _20350_, _20353_);
  and g_30942_(_20173_, _20175_, _20354_);
  or g_30943_(_20172_, _20174_, _20356_);
  and g_30944_(_20353_, _20356_, _20357_);
  or g_30945_(_20352_, _20354_, _20358_);
  and g_30946_(_20349_, _20357_, _20359_);
  or g_30947_(_20348_, _20358_, _20360_);
  and g_30948_(_18562_, _20317_, _20361_);
  or g_30949_(out[304], _20318_, _20362_);
  and g_30950_(_20211_, _20362_, _20363_);
  or g_30951_(_20213_, _20361_, _20364_);
  and g_30952_(_20270_, _20363_, _20365_);
  or g_30953_(_20271_, _20364_, _20367_);
  and g_30954_(_20326_, _20365_, _20368_);
  or g_30955_(_20327_, _20367_, _20369_);
  and g_30956_(_20360_, _20369_, _20370_);
  or g_30957_(_20359_, _20368_, _20371_);
  or g_30958_(_18417_, _20371_, _20372_);
  or g_30959_(_20186_, _20370_, _20373_);
  and g_30960_(_20372_, _20373_, _20374_);
  and g_30961_(_18246_, _18402_, _20375_);
  or g_30962_(_18247_, _18403_, _20376_);
  and g_30963_(_18253_, _18403_, _20378_);
  or g_30964_(_18252_, _18402_, _20379_);
  and g_30965_(_20376_, _20379_, _20380_);
  or g_30966_(_20375_, _20378_, _20381_);
  and g_30967_(_20195_, _20371_, _20382_);
  or g_30968_(_20194_, _20370_, _20383_);
  and g_30969_(_20196_, _20370_, _20384_);
  or g_30970_(_20197_, _20371_, _20385_);
  and g_30971_(_20383_, _20385_, _20386_);
  or g_30972_(_20382_, _20384_, _20387_);
  or g_30973_(_20381_, _20386_, _20389_);
  and g_30974_(_18219_, _18403_, _20390_);
  or g_30975_(_18218_, _18402_, _20391_);
  and g_30976_(_21312_, _18402_, _20392_);
  or g_30977_(_21323_, _18403_, _20393_);
  and g_30978_(_20391_, _20393_, _20394_);
  or g_30979_(_20390_, _20392_, _20395_);
  and g_30980_(_18419_, _20370_, _20396_);
  not g_30981_(_20396_, _20397_);
  and g_30982_(_20162_, _20371_, _20398_);
  or g_30983_(_20161_, _20370_, _20400_);
  and g_30984_(_20397_, _20400_, _20401_);
  or g_30985_(_20396_, _20398_, _20402_);
  or g_30986_(_20394_, _20402_, _20403_);
  or g_30987_(_18292_, _18403_, _20404_);
  or g_30988_(_18296_, _18402_, _20405_);
  and g_30989_(_20404_, _20405_, _20406_);
  or g_30990_(_20253_, _20370_, _20407_);
  or g_30991_(_20254_, _20371_, _20408_);
  and g_30992_(_20407_, _20408_, _20409_);
  xor g_30993_(_20406_, _20409_, _20411_);
  and g_30994_(_18222_, _18224_, _20412_);
  or g_30995_(_20165_, _20167_, _20413_);
  xor g_30996_(_20412_, _20413_, _20414_);
  and g_30997_(_18335_, _18403_, _20415_);
  or g_30998_(_18334_, _18402_, _20416_);
  and g_30999_(_18338_, _18402_, _20417_);
  or g_31000_(_18337_, _18403_, _20418_);
  and g_31001_(_20416_, _20418_, _20419_);
  or g_31002_(_20415_, _20417_, _20420_);
  and g_31003_(_20291_, _20371_, _20422_);
  or g_31004_(_20290_, _20370_, _20423_);
  and g_31005_(_20294_, _20370_, _20424_);
  or g_31006_(_20293_, _20371_, _20425_);
  and g_31007_(_20423_, _20425_, _20426_);
  or g_31008_(_20422_, _20424_, _20427_);
  or g_31009_(_20420_, _20426_, _20428_);
  and g_31010_(_18274_, _18402_, _20429_);
  or g_31011_(_18275_, _18403_, _20430_);
  and g_31012_(_18281_, _18403_, _20431_);
  or g_31013_(_18280_, _18402_, _20433_);
  and g_31014_(_20430_, _20433_, _20434_);
  or g_31015_(_20429_, _20431_, _20435_);
  and g_31016_(_20225_, _20371_, _20436_);
  or g_31017_(_20226_, _20370_, _20437_);
  and g_31018_(_20220_, _20370_, _20438_);
  or g_31019_(_20221_, _20371_, _20439_);
  and g_31020_(_20437_, _20439_, _20440_);
  or g_31021_(_20436_, _20438_, _20441_);
  or g_31022_(_20434_, _20441_, _20442_);
  and g_31023_(_18358_, _18403_, _20444_);
  and g_31024_(_21114_, _18402_, _20445_);
  or g_31025_(_20444_, _20445_, _20446_);
  or g_31026_(_20317_, _20370_, _20447_);
  or g_31027_(out[304], _20371_, _20448_);
  and g_31028_(_20447_, _20448_, _20449_);
  or g_31029_(_20395_, _20401_, _20450_);
  and g_31030_(_18300_, _18402_, _20451_);
  or g_31031_(_18299_, _18403_, _20452_);
  and g_31032_(_18306_, _18403_, _20453_);
  or g_31033_(_18305_, _18402_, _20455_);
  and g_31034_(_20452_, _20455_, _20456_);
  or g_31035_(_20451_, _20453_, _20457_);
  and g_31036_(_20244_, _20371_, _20458_);
  or g_31037_(_20243_, _20370_, _20459_);
  and g_31038_(_20238_, _20370_, _20460_);
  or g_31039_(_20237_, _20371_, _20461_);
  and g_31040_(_20459_, _20461_, _20462_);
  or g_31041_(_20458_, _20460_, _20463_);
  or g_31042_(_20456_, _20463_, _20464_);
  and g_31043_(_18328_, _18403_, _20466_);
  or g_31044_(_18327_, _18402_, _20467_);
  and g_31045_(_18322_, _18402_, _20468_);
  or g_31046_(_18321_, _18403_, _20469_);
  and g_31047_(_20467_, _20469_, _20470_);
  or g_31048_(_20466_, _20468_, _20471_);
  and g_31049_(_20280_, _20371_, _20472_);
  or g_31050_(_20279_, _20370_, _20473_);
  and g_31051_(_20273_, _20370_, _20474_);
  or g_31052_(_20272_, _20371_, _20475_);
  and g_31053_(_20473_, _20475_, _20477_);
  or g_31054_(_20472_, _20474_, _20478_);
  or g_31055_(_20470_, _20478_, _20479_);
  or g_31056_(_20419_, _20427_, _20480_);
  or g_31057_(_20380_, _20387_, _20481_);
  or g_31058_(_18266_, _18403_, _20482_);
  or g_31059_(_18271_, _18402_, _20483_);
  and g_31060_(_20482_, _20483_, _20484_);
  not g_31061_(_20484_, _20485_);
  and g_31062_(_20214_, _20370_, _20486_);
  and g_31063_(_20218_, _20371_, _20488_);
  or g_31064_(_20486_, _20488_, _20489_);
  or g_31065_(_20457_, _20462_, _20490_);
  and g_31066_(out[145], _18402_, _20491_);
  and g_31067_(_18351_, _18403_, _20492_);
  or g_31068_(_20491_, _20492_, _20493_);
  or g_31069_(_19794_, _20371_, _20494_);
  or g_31070_(_20312_, _20370_, _20495_);
  and g_31071_(_20494_, _20495_, _20496_);
  or g_31072_(_20471_, _20477_, _20497_);
  or g_31073_(_20435_, _20440_, _20499_);
  and g_31074_(_20389_, _20479_, _20500_);
  and g_31075_(_20428_, _20500_, _20501_);
  and g_31076_(_20442_, _20464_, _20502_);
  and g_31077_(_20411_, _20502_, _20503_);
  and g_31078_(_20501_, _20503_, _20504_);
  xor g_31079_(_18406_, _20374_, _20505_);
  xor g_31080_(_20446_, _20449_, _20506_);
  and g_31081_(_20505_, _20506_, _20507_);
  xor g_31082_(_20493_, _20496_, _20508_);
  and g_31083_(_20414_, _20490_, _20510_);
  and g_31084_(_20508_, _20510_, _20511_);
  and g_31085_(_20507_, _20511_, _20512_);
  xor g_31086_(_20485_, _20489_, _20513_);
  and g_31087_(_20403_, _20481_, _20514_);
  and g_31088_(_20513_, _20514_, _20515_);
  and g_31089_(_20480_, _20497_, _20516_);
  and g_31090_(_20450_, _20499_, _20517_);
  and g_31091_(_20516_, _20517_, _20518_);
  and g_31092_(_20515_, _20518_, _20519_);
  and g_31093_(_20512_, _20519_, _20521_);
  and g_31094_(_20504_, _20521_, _20522_);
  or g_31095_(out[147], _18336_, _20523_);
  not g_31096_(_20523_, _20524_);
  xor g_31097_(out[147], _18336_, _20525_);
  xor g_31098_(_21136_, _18336_, _20526_);
  or g_31099_(out[131], _18126_, _20527_);
  not g_31100_(_20527_, _20528_);
  xor g_31101_(out[131], _18126_, _20529_);
  xor g_31102_(_21004_, _18126_, _20530_);
  and g_31103_(out[132], _20527_, _20532_);
  or g_31104_(_20960_, _20528_, _20533_);
  or g_31105_(_21345_, _18126_, _20534_);
  not g_31106_(_20534_, _20535_);
  and g_31107_(_20533_, _20534_, _20536_);
  or g_31108_(_20532_, _20535_, _20537_);
  or g_31109_(out[3], _22423_, _20538_);
  and g_31110_(out[4], _20538_, _20539_);
  not g_31111_(_20539_, _20540_);
  or g_31112_(_21862_, _22423_, _20541_);
  not g_31113_(_20541_, _20543_);
  and g_31114_(_20540_, _20541_, _20544_);
  or g_31115_(_20539_, _20543_, _20545_);
  and g_31116_(out[5], _20539_, _20546_);
  and g_31117_(out[6], _20546_, _20547_);
  or g_31118_(out[7], _20547_, _20548_);
  and g_31119_(out[8], _20548_, _20549_);
  or g_31120_(out[9], _20549_, _20550_);
  or g_31121_(out[10], _20550_, _20551_);
  xor g_31122_(out[10], _20550_, _20552_);
  xor g_31123_(_19992_, _20550_, _20554_);
  or g_31124_(out[19], _22390_, _20555_);
  and g_31125_(out[20], _20555_, _20556_);
  not g_31126_(_20556_, _20557_);
  and g_31127_(out[21], _20556_, _20558_);
  and g_31128_(out[22], _20558_, _20559_);
  or g_31129_(out[23], _20559_, _20560_);
  and g_31130_(out[24], _20560_, _20561_);
  or g_31131_(out[25], _20561_, _20562_);
  or g_31132_(out[26], _20562_, _20563_);
  xor g_31133_(out[26], _20562_, _20565_);
  xor g_31134_(_20124_, _20562_, _20566_);
  and g_31135_(_20554_, _20565_, _20567_);
  or g_31136_(_20552_, _20566_, _20568_);
  xor g_31137_(out[11], _20551_, _20569_);
  xor g_31138_(_19871_, _20551_, _20570_);
  xor g_31139_(out[27], _20563_, _20571_);
  xor g_31140_(_20003_, _20563_, _20572_);
  and g_31141_(_20569_, _20572_, _20573_);
  or g_31142_(_20570_, _20571_, _20574_);
  and g_31143_(_20568_, _20574_, _20576_);
  or g_31144_(_20567_, _20573_, _20577_);
  and g_31145_(_20570_, _20571_, _20578_);
  or g_31146_(_20569_, _20572_, _20579_);
  and g_31147_(out[9], _20549_, _20580_);
  xor g_31148_(out[9], _20549_, _20581_);
  xor g_31149_(_19981_, _20549_, _20582_);
  and g_31150_(out[25], _20561_, _20583_);
  xor g_31151_(out[25], _20561_, _20584_);
  xor g_31152_(_20113_, _20561_, _20585_);
  and g_31153_(_20582_, _20584_, _20587_);
  or g_31154_(_20581_, _20585_, _20588_);
  and g_31155_(_20581_, _20585_, _20589_);
  or g_31156_(_20582_, _20584_, _20590_);
  xor g_31157_(_20582_, _20584_, _20591_);
  xor g_31158_(_20581_, _20584_, _20592_);
  xor g_31159_(out[8], _20548_, _20593_);
  xor g_31160_(_19970_, _20548_, _20594_);
  xor g_31161_(out[24], _20560_, _20595_);
  xor g_31162_(_20102_, _20560_, _20596_);
  and g_31163_(_20593_, _20596_, _20598_);
  or g_31164_(_20594_, _20595_, _20599_);
  xor g_31165_(_20594_, _20595_, _20600_);
  xor g_31166_(_20593_, _20595_, _20601_);
  and g_31167_(_20591_, _20600_, _20602_);
  or g_31168_(_20592_, _20601_, _20603_);
  and g_31169_(_20552_, _20566_, _20604_);
  or g_31170_(_20554_, _20565_, _20605_);
  and g_31171_(_20602_, _20605_, _20606_);
  or g_31172_(_20603_, _20604_, _20607_);
  and g_31173_(_20579_, _20606_, _20609_);
  or g_31174_(_20578_, _20607_, _20610_);
  and g_31175_(_20576_, _20609_, _20611_);
  or g_31176_(_20577_, _20610_, _20612_);
  xor g_31177_(out[6], _20546_, _20613_);
  xor g_31178_(_19882_, _20546_, _20614_);
  xor g_31179_(out[22], _20558_, _20615_);
  not g_31180_(_20615_, _20616_);
  and g_31181_(_20613_, _20616_, _20617_);
  or g_31182_(_20614_, _20615_, _20618_);
  xor g_31183_(out[7], _20547_, _20620_);
  xor g_31184_(_19893_, _20547_, _20621_);
  xor g_31185_(out[23], _20559_, _20622_);
  xor g_31186_(_20014_, _20559_, _20623_);
  and g_31187_(_20621_, _20622_, _20624_);
  or g_31188_(_20620_, _20623_, _20625_);
  and g_31189_(_20618_, _20625_, _20626_);
  or g_31190_(_20617_, _20624_, _20627_);
  and g_31191_(_20614_, _20615_, _20628_);
  or g_31192_(_20613_, _20616_, _20629_);
  and g_31193_(_20620_, _20623_, _20631_);
  or g_31194_(_20621_, _20622_, _20632_);
  and g_31195_(_20629_, _20632_, _20633_);
  or g_31196_(_20628_, _20631_, _20634_);
  and g_31197_(_20626_, _20633_, _20635_);
  or g_31198_(_20627_, _20634_, _20636_);
  or g_31199_(_22016_, _22390_, _20637_);
  not g_31200_(_20637_, _20638_);
  and g_31201_(_20557_, _20637_, _20639_);
  or g_31202_(_20556_, _20638_, _20640_);
  and g_31203_(_20544_, _20640_, _20642_);
  or g_31204_(_20545_, _20639_, _20643_);
  xor g_31205_(out[5], _20539_, _20644_);
  xor g_31206_(_19904_, _20539_, _20645_);
  xor g_31207_(out[21], _20556_, _20646_);
  xor g_31208_(_20036_, _20556_, _20647_);
  and g_31209_(_20644_, _20647_, _20648_);
  or g_31210_(_20645_, _20646_, _20649_);
  and g_31211_(_20643_, _20649_, _20650_);
  or g_31212_(_20642_, _20648_, _20651_);
  and g_31213_(_20645_, _20646_, _20653_);
  or g_31214_(_20644_, _20647_, _20654_);
  and g_31215_(_20545_, _20639_, _20655_);
  or g_31216_(_20544_, _20640_, _20656_);
  and g_31217_(_20654_, _20656_, _20657_);
  or g_31218_(_20653_, _20655_, _20658_);
  and g_31219_(_20650_, _20657_, _20659_);
  or g_31220_(_20651_, _20658_, _20660_);
  and g_31221_(_20635_, _20659_, _20661_);
  or g_31222_(_20636_, _20660_, _20662_);
  or g_31223_(out[6], _23215_, _20664_);
  and g_31224_(out[7], _20664_, _20665_);
  xor g_31225_(out[7], _20664_, _20666_);
  xor g_31226_(_19893_, _20664_, _20667_);
  or g_31227_(out[22], _23248_, _20668_);
  and g_31228_(out[23], _20668_, _20669_);
  xor g_31229_(out[23], _20668_, _20670_);
  xor g_31230_(_20014_, _20668_, _20671_);
  and g_31231_(_20666_, _20671_, _20672_);
  or g_31232_(_20667_, _20670_, _20673_);
  and g_31233_(_20667_, _20670_, _20675_);
  or g_31234_(_20666_, _20671_, _20676_);
  xor g_31235_(out[6], _23215_, _20677_);
  xor g_31236_(_19882_, _23215_, _20678_);
  xor g_31237_(out[22], _23248_, _20679_);
  xor g_31238_(_20025_, _23248_, _20680_);
  and g_31239_(_20678_, _20679_, _20681_);
  or g_31240_(_20677_, _20680_, _20682_);
  and g_31241_(_20677_, _20680_, _20683_);
  or g_31242_(_20678_, _20679_, _20684_);
  and g_31243_(_22819_, _20661_, _20686_);
  or g_31244_(_22830_, _20662_, _20687_);
  and g_31245_(_20611_, _20686_, _20688_);
  or g_31246_(_20612_, _20687_, _20689_);
  xor g_31247_(out[3], _22423_, _20690_);
  xor g_31248_(_19959_, _22423_, _20691_);
  xor g_31249_(out[19], _22390_, _20692_);
  xor g_31250_(_20091_, _22390_, _20693_);
  and g_31251_(_20690_, _20693_, _20694_);
  or g_31252_(_20691_, _20692_, _20695_);
  and g_31253_(_20691_, _20692_, _20697_);
  or g_31254_(_20690_, _20693_, _20698_);
  and g_31255_(_22478_, _20698_, _20699_);
  or g_31256_(_22467_, _20697_, _20700_);
  and g_31257_(_20695_, _20700_, _20701_);
  or g_31258_(_20694_, _20699_, _20702_);
  and g_31259_(_22687_, _20702_, _20703_);
  or g_31260_(_22676_, _20701_, _20704_);
  and g_31261_(_20661_, _20704_, _20705_);
  or g_31262_(_20662_, _20703_, _20706_);
  and g_31263_(_20627_, _20632_, _20708_);
  or g_31264_(_20626_, _20631_, _20709_);
  and g_31265_(_20651_, _20654_, _20710_);
  or g_31266_(_20650_, _20653_, _20711_);
  and g_31267_(_20635_, _20710_, _20712_);
  or g_31268_(_20636_, _20711_, _20713_);
  and g_31269_(_20709_, _20713_, _20714_);
  or g_31270_(_20708_, _20712_, _20715_);
  and g_31271_(_20706_, _20714_, _20716_);
  or g_31272_(_20705_, _20715_, _20717_);
  and g_31273_(_20611_, _20717_, _20719_);
  or g_31274_(_20612_, _20716_, _20720_);
  and g_31275_(_20591_, _20598_, _20721_);
  or g_31276_(_20592_, _20599_, _20722_);
  and g_31277_(_20588_, _20722_, _20723_);
  or g_31278_(_20587_, _20721_, _20724_);
  and g_31279_(_20605_, _20724_, _20725_);
  or g_31280_(_20604_, _20723_, _20726_);
  and g_31281_(_20576_, _20726_, _20727_);
  or g_31282_(_20577_, _20725_, _20728_);
  and g_31283_(_20579_, _20728_, _20730_);
  or g_31284_(_20578_, _20727_, _20731_);
  and g_31285_(_20720_, _20731_, _20732_);
  or g_31286_(_20719_, _20730_, _20733_);
  and g_31287_(_20689_, _20733_, _20734_);
  or g_31288_(_20688_, _20732_, _20735_);
  and g_31289_(_20545_, _20735_, _20736_);
  or g_31290_(_20544_, _20734_, _20737_);
  and g_31291_(_20640_, _20734_, _20738_);
  or g_31292_(_20639_, _20735_, _20739_);
  and g_31293_(_20737_, _20739_, _20741_);
  or g_31294_(_20736_, _20738_, _20742_);
  or g_31295_(out[35], _24172_, _20743_);
  not g_31296_(_20743_, _20744_);
  and g_31297_(out[36], _20743_, _20745_);
  or g_31298_(_20179_, _20744_, _20746_);
  and g_31299_(out[37], _20745_, _20747_);
  and g_31300_(out[38], _20747_, _20748_);
  or g_31301_(out[39], _20748_, _20749_);
  and g_31302_(out[40], _20749_, _20750_);
  or g_31303_(out[41], _20750_, _20752_);
  or g_31304_(out[42], _20752_, _20753_);
  xor g_31305_(out[42], _20752_, _20754_);
  not g_31306_(_20754_, _20755_);
  and g_31307_(_20552_, _20735_, _20756_);
  or g_31308_(_20554_, _20734_, _20757_);
  and g_31309_(_20565_, _20734_, _20758_);
  or g_31310_(_20566_, _20735_, _20759_);
  and g_31311_(_20757_, _20759_, _20760_);
  or g_31312_(_20756_, _20758_, _20761_);
  or g_31313_(_20755_, _20761_, _20763_);
  and g_31314_(_20569_, _20571_, _20764_);
  or g_31315_(_20570_, _20572_, _20765_);
  xor g_31316_(out[43], _20753_, _20766_);
  not g_31317_(_20766_, _20767_);
  or g_31318_(_20765_, _20766_, _20768_);
  and g_31319_(_20763_, _20768_, _20769_);
  or g_31320_(_20754_, _20760_, _20770_);
  and g_31321_(_20765_, _20766_, _20771_);
  or g_31322_(_20764_, _20767_, _20772_);
  and g_31323_(_20770_, _20772_, _20774_);
  xor g_31324_(_20755_, _20760_, _20775_);
  xor g_31325_(_20764_, _20766_, _20776_);
  and g_31326_(_20769_, _20774_, _20777_);
  or g_31327_(_20775_, _20776_, _20778_);
  and g_31328_(_20581_, _20735_, _20779_);
  or g_31329_(_20582_, _20734_, _20780_);
  and g_31330_(_20584_, _20734_, _20781_);
  or g_31331_(_20585_, _20735_, _20782_);
  and g_31332_(_20780_, _20782_, _20783_);
  or g_31333_(_20779_, _20781_, _20785_);
  and g_31334_(out[41], _20750_, _20786_);
  xor g_31335_(out[41], _20750_, _20787_);
  xor g_31336_(_20245_, _20750_, _20788_);
  and g_31337_(_20783_, _20787_, _20789_);
  or g_31338_(_20785_, _20788_, _20790_);
  xor g_31339_(out[40], _20749_, _20791_);
  xor g_31340_(_20234_, _20749_, _20792_);
  and g_31341_(_20594_, _20735_, _20793_);
  or g_31342_(_20593_, _20734_, _20794_);
  and g_31343_(_20596_, _20734_, _20796_);
  or g_31344_(_20595_, _20735_, _20797_);
  and g_31345_(_20794_, _20797_, _20798_);
  or g_31346_(_20793_, _20796_, _20799_);
  and g_31347_(_20792_, _20798_, _20800_);
  or g_31348_(_20791_, _20799_, _20801_);
  and g_31349_(_20790_, _20801_, _20802_);
  or g_31350_(_20789_, _20800_, _20803_);
  and g_31351_(_20785_, _20788_, _20804_);
  or g_31352_(_20783_, _20787_, _20805_);
  and g_31353_(_20791_, _20799_, _20807_);
  or g_31354_(_20792_, _20798_, _20808_);
  and g_31355_(_20805_, _20808_, _20809_);
  or g_31356_(_20804_, _20807_, _20810_);
  and g_31357_(_20802_, _20809_, _20811_);
  or g_31358_(_20803_, _20810_, _20812_);
  and g_31359_(_20777_, _20811_, _20813_);
  or g_31360_(_20778_, _20812_, _20814_);
  xor g_31361_(out[38], _20747_, _20815_);
  not g_31362_(_20815_, _20816_);
  or g_31363_(_20613_, _20734_, _20818_);
  or g_31364_(_20615_, _20735_, _20819_);
  and g_31365_(_20818_, _20819_, _20820_);
  and g_31366_(_20816_, _20820_, _20821_);
  xor g_31367_(_20816_, _20820_, _20822_);
  xor g_31368_(_20815_, _20820_, _20823_);
  xor g_31369_(out[39], _20748_, _20824_);
  xor g_31370_(_20146_, _20748_, _20825_);
  or g_31371_(_20623_, _20735_, _20826_);
  or g_31372_(_20621_, _20734_, _20827_);
  and g_31373_(_20826_, _20827_, _20829_);
  or g_31374_(_20824_, _20829_, _20830_);
  and g_31375_(_20824_, _20829_, _20831_);
  xor g_31376_(_20824_, _20829_, _20832_);
  xor g_31377_(_20825_, _20829_, _20833_);
  and g_31378_(_20822_, _20832_, _20834_);
  or g_31379_(_20823_, _20833_, _20835_);
  or g_31380_(_24172_, _24711_, _20836_);
  not g_31381_(_20836_, _20837_);
  and g_31382_(_20746_, _20836_, _20838_);
  or g_31383_(_20745_, _20837_, _20840_);
  and g_31384_(_20741_, _20840_, _20841_);
  or g_31385_(_20742_, _20838_, _20842_);
  xor g_31386_(out[37], _20745_, _20843_);
  xor g_31387_(_20168_, _20745_, _20844_);
  and g_31388_(_20645_, _20735_, _20845_);
  or g_31389_(_20644_, _20734_, _20846_);
  and g_31390_(_20647_, _20734_, _20847_);
  or g_31391_(_20646_, _20735_, _20848_);
  and g_31392_(_20846_, _20848_, _20849_);
  or g_31393_(_20845_, _20847_, _20851_);
  and g_31394_(_20844_, _20849_, _20852_);
  or g_31395_(_20843_, _20851_, _20853_);
  and g_31396_(_20842_, _20853_, _20854_);
  or g_31397_(_20841_, _20852_, _20855_);
  and g_31398_(_20742_, _20838_, _20856_);
  or g_31399_(_20741_, _20840_, _20857_);
  and g_31400_(_20843_, _20851_, _20858_);
  or g_31401_(_20844_, _20849_, _20859_);
  and g_31402_(_20857_, _20859_, _20860_);
  or g_31403_(_20856_, _20858_, _20862_);
  and g_31404_(_20854_, _20860_, _20863_);
  or g_31405_(_20855_, _20862_, _20864_);
  and g_31406_(_20834_, _20863_, _20865_);
  or g_31407_(_20835_, _20864_, _20866_);
  and g_31408_(_20813_, _20865_, _20867_);
  or g_31409_(_20814_, _20866_, _20868_);
  and g_31410_(_22434_, _20735_, _20869_);
  and g_31411_(_22401_, _20734_, _20870_);
  or g_31412_(_20869_, _20870_, _20871_);
  not g_31413_(_20871_, _20873_);
  and g_31414_(_24183_, _20873_, _20874_);
  or g_31415_(_24194_, _20871_, _20875_);
  xor g_31416_(out[35], _24172_, _20876_);
  xor g_31417_(_20223_, _24172_, _20877_);
  and g_31418_(_20690_, _20735_, _20878_);
  or g_31419_(_20691_, _20734_, _20879_);
  and g_31420_(_20692_, _20734_, _20880_);
  or g_31421_(_20693_, _20735_, _20881_);
  and g_31422_(_20879_, _20881_, _20882_);
  or g_31423_(_20878_, _20880_, _20884_);
  and g_31424_(_20876_, _20882_, _20885_);
  or g_31425_(_20877_, _20884_, _20886_);
  and g_31426_(_20875_, _20886_, _20887_);
  or g_31427_(_20874_, _20885_, _20888_);
  and g_31428_(_24194_, _20871_, _20889_);
  or g_31429_(_24183_, _20873_, _20890_);
  and g_31430_(_20877_, _20884_, _20891_);
  or g_31431_(_20876_, _20882_, _20892_);
  and g_31432_(_20890_, _20892_, _20893_);
  or g_31433_(_20889_, _20891_, _20895_);
  and g_31434_(_20887_, _20893_, _20896_);
  or g_31435_(_20888_, _20895_, _20897_);
  or g_31436_(_20058_, _20735_, _20898_);
  or g_31437_(_19926_, _20734_, _20899_);
  and g_31438_(_20898_, _20899_, _20900_);
  or g_31439_(out[0], _20734_, _20901_);
  not g_31440_(_20901_, _20902_);
  and g_31441_(_20069_, _20734_, _20903_);
  or g_31442_(out[16], _20735_, _20904_);
  and g_31443_(_20901_, _20904_, _20906_);
  or g_31444_(_20902_, _20903_, _20907_);
  and g_31445_(out[32], _20907_, _20908_);
  or g_31446_(_20201_, _20906_, _20909_);
  and g_31447_(out[33], _20900_, _20910_);
  not g_31448_(_20910_, _20911_);
  xor g_31449_(out[33], _20900_, _20912_);
  xor g_31450_(_20190_, _20900_, _20913_);
  and g_31451_(_20909_, _20912_, _20914_);
  or g_31452_(_20908_, _20913_, _20915_);
  and g_31453_(_20201_, _20906_, _20917_);
  or g_31454_(out[32], _20907_, _20918_);
  and g_31455_(_20914_, _20918_, _20919_);
  or g_31456_(_20915_, _20917_, _20920_);
  and g_31457_(_20896_, _20919_, _20921_);
  or g_31458_(_20897_, _20920_, _20922_);
  and g_31459_(_20867_, _20921_, _20923_);
  or g_31460_(_20868_, _20922_, _20924_);
  and g_31461_(_20911_, _20915_, _20925_);
  or g_31462_(_20910_, _20914_, _20926_);
  and g_31463_(_20896_, _20926_, _20928_);
  or g_31464_(_20897_, _20925_, _20929_);
  and g_31465_(_20888_, _20892_, _20930_);
  or g_31466_(_20887_, _20891_, _20931_);
  and g_31467_(_20929_, _20931_, _20932_);
  or g_31468_(_20928_, _20930_, _20933_);
  and g_31469_(_20867_, _20933_, _20934_);
  or g_31470_(_20868_, _20932_, _20935_);
  and g_31471_(_20834_, _20855_, _20936_);
  or g_31472_(_20835_, _20854_, _20937_);
  and g_31473_(_20859_, _20936_, _20939_);
  or g_31474_(_20858_, _20937_, _20940_);
  and g_31475_(_20821_, _20830_, _20941_);
  or g_31476_(_20831_, _20941_, _20942_);
  not g_31477_(_20942_, _20943_);
  and g_31478_(_20940_, _20943_, _20944_);
  or g_31479_(_20939_, _20942_, _20945_);
  and g_31480_(_20813_, _20945_, _20946_);
  or g_31481_(_20814_, _20944_, _20947_);
  or g_31482_(_20769_, _20771_, _20948_);
  or g_31483_(_20778_, _20802_, _20950_);
  or g_31484_(_20804_, _20950_, _20951_);
  and g_31485_(_20948_, _20951_, _20952_);
  not g_31486_(_20952_, _20953_);
  and g_31487_(_20947_, _20952_, _20954_);
  or g_31488_(_20946_, _20953_, _20955_);
  and g_31489_(_20935_, _20954_, _20956_);
  or g_31490_(_20934_, _20955_, _20957_);
  and g_31491_(_20924_, _20957_, _20958_);
  or g_31492_(_20923_, _20956_, _20959_);
  or g_31493_(_20741_, _20958_, _20961_);
  or g_31494_(_20838_, _20959_, _20962_);
  and g_31495_(_20961_, _20962_, _20963_);
  not g_31496_(_20963_, _20964_);
  or g_31497_(out[51], _10219_, _20965_);
  not g_31498_(_20965_, _20966_);
  and g_31499_(out[52], _20965_, _20967_);
  or g_31500_(_20311_, _20966_, _20968_);
  and g_31501_(out[53], _20967_, _20969_);
  and g_31502_(out[54], _20969_, _20970_);
  or g_31503_(out[55], _20970_, _20972_);
  and g_31504_(out[56], _20972_, _20973_);
  or g_31505_(out[57], _20973_, _20974_);
  or g_31506_(out[58], _20974_, _20975_);
  xor g_31507_(out[58], _20974_, _20976_);
  or g_31508_(_20760_, _20958_, _20977_);
  or g_31509_(_20755_, _20959_, _20978_);
  and g_31510_(_20977_, _20978_, _20979_);
  and g_31511_(_20976_, _20979_, _20980_);
  not g_31512_(_20980_, _20981_);
  and g_31513_(_20764_, _20766_, _20983_);
  or g_31514_(_20765_, _20767_, _20984_);
  xor g_31515_(out[59], _20975_, _20985_);
  xor g_31516_(_20267_, _20975_, _20986_);
  and g_31517_(_20983_, _20986_, _20987_);
  or g_31518_(_20984_, _20985_, _20988_);
  and g_31519_(_20981_, _20988_, _20989_);
  or g_31520_(_20980_, _20987_, _20990_);
  or g_31521_(_20976_, _20979_, _20991_);
  and g_31522_(_20984_, _20985_, _20992_);
  or g_31523_(_20983_, _20986_, _20994_);
  and g_31524_(_20991_, _20994_, _20995_);
  not g_31525_(_20995_, _20996_);
  and g_31526_(_20989_, _20995_, _20997_);
  or g_31527_(_20990_, _20996_, _20998_);
  or g_31528_(_20787_, _20959_, _20999_);
  or g_31529_(_20785_, _20958_, _21000_);
  and g_31530_(_20999_, _21000_, _21001_);
  not g_31531_(_21001_, _21002_);
  and g_31532_(out[57], _20973_, _21003_);
  xor g_31533_(out[57], _20973_, _21005_);
  xor g_31534_(_20377_, _20973_, _21006_);
  or g_31535_(_21001_, _21006_, _21007_);
  not g_31536_(_21007_, _21008_);
  xor g_31537_(out[56], _20972_, _21009_);
  xor g_31538_(_20366_, _20972_, _21010_);
  or g_31539_(_20791_, _20959_, _21011_);
  or g_31540_(_20798_, _20958_, _21012_);
  and g_31541_(_21011_, _21012_, _21013_);
  not g_31542_(_21013_, _21014_);
  and g_31543_(_21010_, _21013_, _21016_);
  not g_31544_(_21016_, _21017_);
  and g_31545_(_21007_, _21017_, _21018_);
  or g_31546_(_21008_, _21016_, _21019_);
  and g_31547_(_21001_, _21006_, _21020_);
  or g_31548_(_21002_, _21005_, _21021_);
  and g_31549_(_21009_, _21014_, _21022_);
  or g_31550_(_21010_, _21013_, _21023_);
  and g_31551_(_21021_, _21023_, _21024_);
  or g_31552_(_21020_, _21022_, _21025_);
  and g_31553_(_21018_, _21024_, _21027_);
  or g_31554_(_21019_, _21025_, _21028_);
  and g_31555_(_20997_, _21027_, _21029_);
  or g_31556_(_20998_, _21028_, _21030_);
  xor g_31557_(out[54], _20969_, _21031_);
  xor g_31558_(_20289_, _20969_, _21032_);
  or g_31559_(_20815_, _20959_, _21033_);
  or g_31560_(_20820_, _20958_, _21034_);
  and g_31561_(_21033_, _21034_, _21035_);
  xor g_31562_(out[55], _20970_, _21036_);
  xor g_31563_(_20278_, _20970_, _21038_);
  or g_31564_(_20829_, _20958_, _21039_);
  or g_31565_(_20825_, _20959_, _21040_);
  and g_31566_(_21039_, _21040_, _21041_);
  not g_31567_(_21041_, _21042_);
  and g_31568_(_21036_, _21041_, _21043_);
  or g_31569_(_21036_, _21041_, _21044_);
  and g_31570_(_21032_, _21035_, _21045_);
  xor g_31571_(out[53], _20967_, _21046_);
  xor g_31572_(_20300_, _20967_, _21047_);
  or g_31573_(_20849_, _20958_, _21049_);
  or g_31574_(_20843_, _20959_, _21050_);
  and g_31575_(_21049_, _21050_, _21051_);
  or g_31576_(_21047_, _21051_, _21052_);
  not g_31577_(_21052_, _21053_);
  xor g_31578_(_21032_, _21035_, _21054_);
  xor g_31579_(_21031_, _21035_, _21055_);
  xor g_31580_(_21036_, _21041_, _21056_);
  xor g_31581_(_21038_, _21041_, _21057_);
  and g_31582_(_21054_, _21056_, _21058_);
  or g_31583_(_21055_, _21057_, _21060_);
  and g_31584_(_21052_, _21058_, _21061_);
  or g_31585_(_21053_, _21060_, _21062_);
  or g_31586_(_21730_, _10219_, _21063_);
  not g_31587_(_21063_, _21064_);
  and g_31588_(_20968_, _21063_, _21065_);
  or g_31589_(_20967_, _21064_, _21066_);
  and g_31590_(_20963_, _21066_, _21067_);
  or g_31591_(_20964_, _21065_, _21068_);
  and g_31592_(_21047_, _21051_, _21069_);
  not g_31593_(_21069_, _21071_);
  and g_31594_(_21068_, _21071_, _21072_);
  or g_31595_(_21067_, _21069_, _21073_);
  and g_31596_(_20964_, _21065_, _21074_);
  or g_31597_(_20963_, _21066_, _21075_);
  and g_31598_(_21072_, _21075_, _21076_);
  or g_31599_(_21073_, _21074_, _21077_);
  and g_31600_(_21061_, _21076_, _21078_);
  or g_31601_(_21062_, _21077_, _21079_);
  xor g_31602_(out[51], _10219_, _21080_);
  xor g_31603_(_20355_, _10219_, _21082_);
  and g_31604_(_20884_, _20959_, _21083_);
  or g_31605_(_20882_, _20958_, _21084_);
  and g_31606_(_20876_, _20958_, _21085_);
  or g_31607_(_20877_, _20959_, _21086_);
  and g_31608_(_21084_, _21086_, _21087_);
  or g_31609_(_21083_, _21085_, _21088_);
  and g_31610_(_21080_, _21087_, _21089_);
  or g_31611_(_21082_, _21088_, _21090_);
  and g_31612_(_20871_, _20959_, _21091_);
  or g_31613_(_20873_, _20958_, _21093_);
  and g_31614_(_24183_, _20958_, _21094_);
  or g_31615_(_24194_, _20959_, _21095_);
  and g_31616_(_21093_, _21095_, _21096_);
  or g_31617_(_21091_, _21094_, _21097_);
  and g_31618_(_10230_, _21096_, _21098_);
  or g_31619_(_10241_, _21097_, _21099_);
  and g_31620_(_21090_, _21099_, _21100_);
  or g_31621_(_21089_, _21098_, _21101_);
  or g_31622_(_21080_, _21087_, _21102_);
  not g_31623_(_21102_, _21104_);
  and g_31624_(_10241_, _21097_, _21105_);
  or g_31625_(_10230_, _21096_, _21106_);
  and g_31626_(_21102_, _21106_, _21107_);
  or g_31627_(_21104_, _21105_, _21108_);
  and g_31628_(_21100_, _21107_, _21109_);
  or g_31629_(_21101_, _21108_, _21110_);
  or g_31630_(_20190_, _20959_, _21111_);
  or g_31631_(_20900_, _20958_, _21112_);
  and g_31632_(_21111_, _21112_, _21113_);
  and g_31633_(out[49], _21113_, _21115_);
  and g_31634_(_21109_, _21115_, _21116_);
  not g_31635_(_21116_, _21117_);
  and g_31636_(_21101_, _21102_, _21118_);
  or g_31637_(_21100_, _21104_, _21119_);
  and g_31638_(out[32], _20958_, _21120_);
  or g_31639_(_20201_, _20959_, _21121_);
  and g_31640_(_20906_, _20959_, _21122_);
  or g_31641_(_20907_, _20958_, _21123_);
  and g_31642_(_21121_, _21123_, _21124_);
  or g_31643_(_21120_, _21122_, _21126_);
  and g_31644_(out[48], _21124_, _21127_);
  or g_31645_(_20333_, _21126_, _21128_);
  xor g_31646_(out[49], _21113_, _21129_);
  xor g_31647_(_20322_, _21113_, _21130_);
  and g_31648_(_21128_, _21129_, _21131_);
  or g_31649_(_21127_, _21130_, _21132_);
  and g_31650_(_21109_, _21131_, _21133_);
  or g_31651_(_21110_, _21132_, _21134_);
  and g_31652_(_21119_, _21134_, _21135_);
  or g_31653_(_21118_, _21133_, _21137_);
  and g_31654_(_21117_, _21135_, _21138_);
  or g_31655_(_21116_, _21137_, _21139_);
  and g_31656_(_21078_, _21139_, _21140_);
  or g_31657_(_21079_, _21138_, _21141_);
  and g_31658_(_21061_, _21073_, _21142_);
  not g_31659_(_21142_, _21143_);
  and g_31660_(_21044_, _21045_, _21144_);
  or g_31661_(_21043_, _21144_, _21145_);
  not g_31662_(_21145_, _21146_);
  and g_31663_(_21143_, _21146_, _21148_);
  or g_31664_(_21142_, _21145_, _21149_);
  and g_31665_(_21141_, _21148_, _21150_);
  or g_31666_(_21140_, _21149_, _21151_);
  and g_31667_(_21029_, _21151_, _21152_);
  or g_31668_(_21030_, _21150_, _21153_);
  and g_31669_(_21019_, _21021_, _21154_);
  or g_31670_(_21018_, _21020_, _21155_);
  and g_31671_(_20997_, _21154_, _21156_);
  or g_31672_(_20998_, _21155_, _21157_);
  and g_31673_(_20990_, _20994_, _21159_);
  or g_31674_(_20989_, _20992_, _21160_);
  and g_31675_(_21157_, _21160_, _21161_);
  or g_31676_(_21156_, _21159_, _21162_);
  and g_31677_(_21153_, _21161_, _21163_);
  or g_31678_(_21152_, _21162_, _21164_);
  or g_31679_(out[48], _21124_, _21165_);
  and g_31680_(_21029_, _21165_, _21166_);
  and g_31681_(_21078_, _21133_, _21167_);
  and g_31682_(_21166_, _21167_, _21168_);
  not g_31683_(_21168_, _21170_);
  and g_31684_(_21164_, _21170_, _21171_);
  or g_31685_(_21163_, _21168_, _21172_);
  or g_31686_(_20963_, _21171_, _21173_);
  not g_31687_(_21173_, _21174_);
  and g_31688_(_21066_, _21171_, _21175_);
  not g_31689_(_21175_, _21176_);
  and g_31690_(_21173_, _21176_, _21177_);
  or g_31691_(_21174_, _21175_, _21178_);
  or g_31692_(out[67], _12518_, _21179_);
  not g_31693_(_21179_, _21181_);
  and g_31694_(out[68], _21179_, _21182_);
  or g_31695_(_20443_, _21181_, _21183_);
  and g_31696_(out[69], _21182_, _21184_);
  and g_31697_(out[70], _21184_, _21185_);
  or g_31698_(out[71], _21185_, _21186_);
  and g_31699_(out[72], _21186_, _21187_);
  or g_31700_(out[73], _21187_, _21188_);
  not g_31701_(_21188_, _21189_);
  or g_31702_(out[74], _21188_, _21190_);
  xor g_31703_(out[74], _21188_, _21192_);
  xor g_31704_(_20520_, _21188_, _21193_);
  or g_31705_(_20979_, _21171_, _21194_);
  not g_31706_(_21194_, _21195_);
  and g_31707_(_20976_, _21171_, _21196_);
  not g_31708_(_21196_, _21197_);
  and g_31709_(_21194_, _21197_, _21198_);
  or g_31710_(_21195_, _21196_, _21199_);
  and g_31711_(_21192_, _21198_, _21200_);
  or g_31712_(_21193_, _21199_, _21201_);
  and g_31713_(_20983_, _20985_, _21203_);
  or g_31714_(_20984_, _20986_, _21204_);
  xor g_31715_(out[75], _21190_, _21205_);
  xor g_31716_(_20399_, _21190_, _21206_);
  and g_31717_(_21203_, _21206_, _21207_);
  or g_31718_(_21204_, _21205_, _21208_);
  and g_31719_(_21201_, _21208_, _21209_);
  or g_31720_(_21200_, _21207_, _21210_);
  and g_31721_(_21193_, _21199_, _21211_);
  or g_31722_(_21192_, _21198_, _21212_);
  and g_31723_(_21204_, _21205_, _21214_);
  or g_31724_(_21203_, _21206_, _21215_);
  and g_31725_(out[73], _21187_, _21216_);
  xor g_31726_(out[73], _21187_, _21217_);
  or g_31727_(_21189_, _21216_, _21218_);
  or g_31728_(_21001_, _21171_, _21219_);
  not g_31729_(_21219_, _21220_);
  and g_31730_(_21006_, _21171_, _21221_);
  not g_31731_(_21221_, _21222_);
  and g_31732_(_21219_, _21222_, _21223_);
  or g_31733_(_21220_, _21221_, _21225_);
  and g_31734_(_21217_, _21225_, _21226_);
  or g_31735_(_21218_, _21223_, _21227_);
  xor g_31736_(out[72], _21186_, _21228_);
  xor g_31737_(_20498_, _21186_, _21229_);
  and g_31738_(_21010_, _21171_, _21230_);
  not g_31739_(_21230_, _21231_);
  or g_31740_(_21013_, _21171_, _21232_);
  not g_31741_(_21232_, _21233_);
  and g_31742_(_21231_, _21232_, _21234_);
  or g_31743_(_21230_, _21233_, _21236_);
  and g_31744_(_21229_, _21234_, _21237_);
  or g_31745_(_21228_, _21236_, _21238_);
  and g_31746_(_21218_, _21223_, _21239_);
  or g_31747_(_21217_, _21225_, _21240_);
  and g_31748_(_21238_, _21240_, _21241_);
  or g_31749_(_21237_, _21239_, _21242_);
  and g_31750_(_21228_, _21236_, _21243_);
  or g_31751_(_21229_, _21234_, _21244_);
  and g_31752_(_21212_, _21215_, _21245_);
  or g_31753_(_21211_, _21214_, _21247_);
  and g_31754_(_21209_, _21245_, _21248_);
  or g_31755_(_21210_, _21247_, _21249_);
  and g_31756_(_21227_, _21244_, _21250_);
  or g_31757_(_21226_, _21243_, _21251_);
  and g_31758_(_21241_, _21250_, _21252_);
  or g_31759_(_21242_, _21251_, _21253_);
  and g_31760_(_21248_, _21252_, _21254_);
  or g_31761_(_21249_, _21253_, _21255_);
  xor g_31762_(out[70], _21184_, _21256_);
  xor g_31763_(_20421_, _21184_, _21258_);
  or g_31764_(_21031_, _21172_, _21259_);
  or g_31765_(_21035_, _21171_, _21260_);
  and g_31766_(_21259_, _21260_, _21261_);
  not g_31767_(_21261_, _21262_);
  and g_31768_(_21258_, _21261_, _21263_);
  or g_31769_(_21256_, _21262_, _21264_);
  xor g_31770_(_21258_, _21261_, _21265_);
  xor g_31771_(_21256_, _21261_, _21266_);
  xor g_31772_(out[71], _21185_, _21267_);
  xor g_31773_(_20410_, _21185_, _21269_);
  and g_31774_(_21036_, _21171_, _21270_);
  or g_31775_(_21038_, _21172_, _21271_);
  and g_31776_(_21042_, _21172_, _21272_);
  or g_31777_(_21041_, _21171_, _21273_);
  and g_31778_(_21271_, _21273_, _21274_);
  or g_31779_(_21270_, _21272_, _21275_);
  and g_31780_(_21267_, _21274_, _21276_);
  or g_31781_(_21269_, _21275_, _21277_);
  and g_31782_(_21269_, _21275_, _21278_);
  or g_31783_(_21267_, _21274_, _21280_);
  and g_31784_(_21265_, _21277_, _21281_);
  or g_31785_(_21266_, _21276_, _21282_);
  and g_31786_(_21280_, _21281_, _21283_);
  or g_31787_(_21278_, _21282_, _21284_);
  or g_31788_(_21598_, _12518_, _21285_);
  not g_31789_(_21285_, _21286_);
  and g_31790_(_21183_, _21285_, _21287_);
  or g_31791_(_21182_, _21286_, _21288_);
  and g_31792_(_21177_, _21288_, _21289_);
  or g_31793_(_21178_, _21287_, _21291_);
  xor g_31794_(out[69], _21182_, _21292_);
  xor g_31795_(_20432_, _21182_, _21293_);
  and g_31796_(_21047_, _21171_, _21294_);
  not g_31797_(_21294_, _21295_);
  or g_31798_(_21051_, _21171_, _21296_);
  not g_31799_(_21296_, _21297_);
  and g_31800_(_21295_, _21296_, _21298_);
  or g_31801_(_21294_, _21297_, _21299_);
  and g_31802_(_21293_, _21298_, _21300_);
  or g_31803_(_21292_, _21299_, _21302_);
  and g_31804_(_21291_, _21302_, _21303_);
  or g_31805_(_21289_, _21300_, _21304_);
  and g_31806_(_21292_, _21299_, _21305_);
  or g_31807_(_21293_, _21298_, _21306_);
  and g_31808_(_21178_, _21287_, _21307_);
  or g_31809_(_21177_, _21288_, _21308_);
  and g_31810_(_21306_, _21308_, _21309_);
  or g_31811_(_21305_, _21307_, _21310_);
  and g_31812_(_21303_, _21309_, _21311_);
  or g_31813_(_21304_, _21310_, _21313_);
  and g_31814_(_21283_, _21311_, _21314_);
  or g_31815_(_21284_, _21313_, _21315_);
  and g_31816_(_21254_, _21314_, _21316_);
  or g_31817_(_21255_, _21315_, _21317_);
  xor g_31818_(out[67], _12518_, _21318_);
  xor g_31819_(_20487_, _12518_, _21319_);
  and g_31820_(_21080_, _21171_, _21320_);
  not g_31821_(_21320_, _21321_);
  or g_31822_(_21087_, _21171_, _21322_);
  not g_31823_(_21322_, _21324_);
  and g_31824_(_21321_, _21322_, _21325_);
  or g_31825_(_21320_, _21324_, _21326_);
  and g_31826_(_21318_, _21325_, _21327_);
  or g_31827_(_21319_, _21326_, _21328_);
  and g_31828_(_21319_, _21326_, _21329_);
  or g_31829_(_21318_, _21325_, _21330_);
  and g_31830_(_21328_, _21330_, _21331_);
  or g_31831_(_21327_, _21329_, _21332_);
  or g_31832_(_21096_, _21171_, _21333_);
  or g_31833_(_10241_, _21172_, _21335_);
  and g_31834_(_21333_, _21335_, _21336_);
  not g_31835_(_21336_, _21337_);
  and g_31836_(_12529_, _21336_, _21338_);
  or g_31837_(_12540_, _21337_, _21339_);
  xor g_31838_(_12529_, _21336_, _21340_);
  xor g_31839_(_12540_, _21336_, _21341_);
  and g_31840_(_21331_, _21340_, _21342_);
  or g_31841_(_21332_, _21341_, _21343_);
  and g_31842_(out[49], _21171_, _21344_);
  not g_31843_(_21344_, _21346_);
  or g_31844_(_21113_, _21171_, _21347_);
  not g_31845_(_21347_, _21348_);
  and g_31846_(_21346_, _21347_, _21349_);
  or g_31847_(_21344_, _21348_, _21350_);
  and g_31848_(out[65], _21349_, _21351_);
  or g_31849_(_20454_, _21350_, _21352_);
  and g_31850_(_21328_, _21339_, _21353_);
  or g_31851_(_21327_, _21338_, _21354_);
  and g_31852_(_21330_, _21354_, _21355_);
  or g_31853_(_21329_, _21353_, _21357_);
  and g_31854_(out[48], _21171_, _21358_);
  not g_31855_(_21358_, _21359_);
  or g_31856_(_21124_, _21171_, _21360_);
  not g_31857_(_21360_, _21361_);
  and g_31858_(_21359_, _21360_, _21362_);
  or g_31859_(_21358_, _21361_, _21363_);
  and g_31860_(out[64], _21362_, _21364_);
  or g_31861_(_20465_, _21363_, _21365_);
  xor g_31862_(out[65], _21349_, _21366_);
  xor g_31863_(_20454_, _21349_, _21368_);
  and g_31864_(_21365_, _21366_, _21369_);
  or g_31865_(_21364_, _21368_, _21370_);
  and g_31866_(_21342_, _21369_, _21371_);
  or g_31867_(_21343_, _21370_, _21372_);
  and g_31868_(_21352_, _21370_, _21373_);
  or g_31869_(_21351_, _21369_, _21374_);
  and g_31870_(_21342_, _21374_, _21375_);
  or g_31871_(_21343_, _21373_, _21376_);
  and g_31872_(_21357_, _21376_, _21377_);
  or g_31873_(_21355_, _21375_, _21379_);
  and g_31874_(_21316_, _21379_, _21380_);
  or g_31875_(_21317_, _21377_, _21381_);
  and g_31876_(_21304_, _21306_, _21382_);
  or g_31877_(_21303_, _21305_, _21383_);
  and g_31878_(_21283_, _21382_, _21384_);
  or g_31879_(_21284_, _21383_, _21385_);
  and g_31880_(_21263_, _21280_, _21386_);
  or g_31881_(_21264_, _21278_, _21387_);
  and g_31882_(_21277_, _21387_, _21388_);
  or g_31883_(_21276_, _21386_, _21390_);
  and g_31884_(_21385_, _21388_, _21391_);
  or g_31885_(_21384_, _21390_, _21392_);
  and g_31886_(_21254_, _21392_, _21393_);
  or g_31887_(_21255_, _21391_, _21394_);
  and g_31888_(_21227_, _21238_, _21395_);
  or g_31889_(_21226_, _21237_, _21396_);
  and g_31890_(_21240_, _21396_, _21397_);
  or g_31891_(_21239_, _21395_, _21398_);
  and g_31892_(_21248_, _21397_, _21399_);
  or g_31893_(_21249_, _21398_, _21401_);
  and g_31894_(_21394_, _21401_, _21402_);
  or g_31895_(_21393_, _21399_, _21403_);
  and g_31896_(_21210_, _21215_, _21404_);
  or g_31897_(_21209_, _21214_, _21405_);
  and g_31898_(_21381_, _21405_, _21406_);
  or g_31899_(_21380_, _21404_, _21407_);
  and g_31900_(_21402_, _21406_, _21408_);
  or g_31901_(_21403_, _21407_, _21409_);
  and g_31902_(_20465_, _21363_, _21410_);
  or g_31903_(out[64], _21362_, _21412_);
  and g_31904_(_21371_, _21412_, _21413_);
  or g_31905_(_21372_, _21410_, _21414_);
  and g_31906_(_21316_, _21413_, _21415_);
  or g_31907_(_21317_, _21414_, _21416_);
  and g_31908_(_21409_, _21416_, _21417_);
  or g_31909_(_21408_, _21415_, _21418_);
  or g_31910_(_21177_, _21417_, _21419_);
  not g_31911_(_21419_, _21420_);
  and g_31912_(_21288_, _21417_, _21421_);
  not g_31913_(_21421_, _21423_);
  and g_31914_(_21419_, _21423_, _21424_);
  or g_31915_(_21420_, _21421_, _21425_);
  and g_31916_(_21203_, _21205_, _21426_);
  or g_31917_(_21204_, _21206_, _21427_);
  or g_31918_(out[83], _14564_, _21428_);
  not g_31919_(_21428_, _21429_);
  and g_31920_(out[84], _21428_, _21430_);
  or g_31921_(_20575_, _21429_, _21431_);
  and g_31922_(out[85], _21430_, _21432_);
  and g_31923_(out[86], _21432_, _21434_);
  or g_31924_(out[87], _21434_, _21435_);
  and g_31925_(out[88], _21435_, _21436_);
  or g_31926_(out[89], _21436_, _21437_);
  not g_31927_(_21437_, _21438_);
  or g_31928_(out[90], _21437_, _21439_);
  xor g_31929_(out[91], _21439_, _21440_);
  xor g_31930_(_20531_, _21439_, _21441_);
  and g_31931_(_21427_, _21440_, _21442_);
  or g_31932_(_21426_, _21441_, _21443_);
  xor g_31933_(out[90], _21437_, _21445_);
  xor g_31934_(_20652_, _21437_, _21446_);
  or g_31935_(_21198_, _21417_, _21447_);
  not g_31936_(_21447_, _21448_);
  and g_31937_(_21192_, _21417_, _21449_);
  not g_31938_(_21449_, _21450_);
  and g_31939_(_21447_, _21450_, _21451_);
  or g_31940_(_21448_, _21449_, _21452_);
  and g_31941_(_21445_, _21451_, _21453_);
  or g_31942_(_21446_, _21452_, _21454_);
  and g_31943_(_21426_, _21441_, _21456_);
  or g_31944_(_21427_, _21440_, _21457_);
  and g_31945_(_21454_, _21457_, _21458_);
  or g_31946_(_21453_, _21456_, _21459_);
  and g_31947_(_21225_, _21418_, _21460_);
  or g_31948_(_21223_, _21417_, _21461_);
  and g_31949_(_21218_, _21417_, _21462_);
  or g_31950_(_21217_, _21418_, _21463_);
  and g_31951_(_21461_, _21463_, _21464_);
  or g_31952_(_21460_, _21462_, _21465_);
  and g_31953_(out[89], _21436_, _21467_);
  xor g_31954_(out[89], _21436_, _21468_);
  or g_31955_(_21438_, _21467_, _21469_);
  and g_31956_(_21464_, _21469_, _21470_);
  or g_31957_(_21465_, _21468_, _21471_);
  and g_31958_(_21465_, _21468_, _21472_);
  or g_31959_(_21464_, _21469_, _21473_);
  xor g_31960_(out[88], _21435_, _21474_);
  xor g_31961_(_20630_, _21435_, _21475_);
  and g_31962_(_21229_, _21417_, _21476_);
  not g_31963_(_21476_, _21478_);
  or g_31964_(_21234_, _21417_, _21479_);
  not g_31965_(_21479_, _21480_);
  and g_31966_(_21478_, _21479_, _21481_);
  or g_31967_(_21476_, _21480_, _21482_);
  and g_31968_(_21475_, _21481_, _21483_);
  or g_31969_(_21474_, _21482_, _21484_);
  and g_31970_(_21473_, _21484_, _21485_);
  or g_31971_(_21472_, _21483_, _21486_);
  and g_31972_(_21471_, _21486_, _21487_);
  or g_31973_(_21470_, _21485_, _21489_);
  and g_31974_(_21446_, _21452_, _21490_);
  or g_31975_(_21445_, _21451_, _21491_);
  and g_31976_(_21458_, _21491_, _21492_);
  or g_31977_(_21459_, _21490_, _21493_);
  and g_31978_(_21487_, _21492_, _21494_);
  or g_31979_(_21489_, _21493_, _21495_);
  and g_31980_(_21458_, _21495_, _21496_);
  or g_31981_(_21459_, _21494_, _21497_);
  and g_31982_(_21443_, _21497_, _21498_);
  or g_31983_(_21442_, _21496_, _21500_);
  and g_31984_(_21474_, _21482_, _21501_);
  or g_31985_(_21475_, _21481_, _21502_);
  and g_31986_(_21443_, _21471_, _21503_);
  or g_31987_(_21442_, _21470_, _21504_);
  and g_31988_(_21502_, _21503_, _21505_);
  or g_31989_(_21501_, _21504_, _21506_);
  and g_31990_(_21485_, _21505_, _21507_);
  or g_31991_(_21486_, _21506_, _21508_);
  and g_31992_(_21492_, _21507_, _21509_);
  or g_31993_(_21493_, _21508_, _21511_);
  xor g_31994_(out[87], _21434_, _21512_);
  xor g_31995_(_20542_, _21434_, _21513_);
  and g_31996_(_21267_, _21417_, _21514_);
  or g_31997_(_21269_, _21418_, _21515_);
  and g_31998_(_21275_, _21418_, _21516_);
  or g_31999_(_21274_, _21417_, _21517_);
  and g_32000_(_21515_, _21517_, _21518_);
  or g_32001_(_21514_, _21516_, _21519_);
  and g_32002_(_21513_, _21519_, _21520_);
  or g_32003_(_21512_, _21518_, _21522_);
  and g_32004_(_21512_, _21518_, _21523_);
  or g_32005_(_21513_, _21519_, _21524_);
  xor g_32006_(out[86], _21432_, _21525_);
  xor g_32007_(_20553_, _21432_, _21526_);
  and g_32008_(_21262_, _21418_, _21527_);
  or g_32009_(_21261_, _21417_, _21528_);
  and g_32010_(_21258_, _21417_, _21529_);
  or g_32011_(_21256_, _21418_, _21530_);
  and g_32012_(_21528_, _21530_, _21531_);
  or g_32013_(_21527_, _21529_, _21533_);
  and g_32014_(_21526_, _21531_, _21534_);
  or g_32015_(_21525_, _21533_, _21535_);
  and g_32016_(_21524_, _21535_, _21536_);
  or g_32017_(_21523_, _21534_, _21537_);
  and g_32018_(_21522_, _21537_, _21538_);
  or g_32019_(_21520_, _21536_, _21539_);
  xor g_32020_(_21526_, _21531_, _21540_);
  xor g_32021_(_21525_, _21531_, _21541_);
  and g_32022_(_21524_, _21540_, _21542_);
  or g_32023_(_21523_, _21541_, _21544_);
  and g_32024_(_21522_, _21542_, _21545_);
  or g_32025_(_21520_, _21544_, _21546_);
  xor g_32026_(out[85], _21430_, _21547_);
  xor g_32027_(_20564_, _21430_, _21548_);
  and g_32028_(_21293_, _21417_, _21549_);
  not g_32029_(_21549_, _21550_);
  or g_32030_(_21298_, _21417_, _21551_);
  not g_32031_(_21551_, _21552_);
  and g_32032_(_21550_, _21551_, _21553_);
  or g_32033_(_21549_, _21552_, _21555_);
  and g_32034_(_21547_, _21555_, _21556_);
  or g_32035_(_21548_, _21553_, _21557_);
  or g_32036_(_21466_, _14564_, _21558_);
  not g_32037_(_21558_, _21559_);
  and g_32038_(_21431_, _21558_, _21560_);
  or g_32039_(_21430_, _21559_, _21561_);
  and g_32040_(_21424_, _21561_, _21562_);
  or g_32041_(_21425_, _21560_, _21563_);
  and g_32042_(_21548_, _21553_, _21564_);
  or g_32043_(_21547_, _21555_, _21566_);
  and g_32044_(_21563_, _21566_, _21567_);
  or g_32045_(_21562_, _21564_, _21568_);
  and g_32046_(_21557_, _21568_, _21569_);
  or g_32047_(_21556_, _21567_, _21570_);
  xor g_32048_(out[83], _14564_, _21571_);
  xor g_32049_(_20619_, _14564_, _21572_);
  and g_32050_(_21318_, _21417_, _21573_);
  not g_32051_(_21573_, _21574_);
  or g_32052_(_21325_, _21417_, _21575_);
  not g_32053_(_21575_, _21577_);
  and g_32054_(_21574_, _21575_, _21578_);
  or g_32055_(_21573_, _21577_, _21579_);
  and g_32056_(_21571_, _21578_, _21580_);
  or g_32057_(_21572_, _21579_, _21581_);
  or g_32058_(_21336_, _21417_, _21582_);
  or g_32059_(_12540_, _21418_, _21583_);
  and g_32060_(_21582_, _21583_, _21584_);
  not g_32061_(_21584_, _21585_);
  and g_32062_(_14575_, _21584_, _21586_);
  or g_32063_(_14586_, _21585_, _21588_);
  and g_32064_(_21581_, _21588_, _21589_);
  or g_32065_(_21580_, _21586_, _21590_);
  and g_32066_(_21572_, _21579_, _21591_);
  or g_32067_(_21571_, _21578_, _21592_);
  and g_32068_(_14586_, _21585_, _21593_);
  or g_32069_(_14575_, _21584_, _21594_);
  and g_32070_(_21592_, _21594_, _21595_);
  or g_32071_(_21591_, _21593_, _21596_);
  and g_32072_(_21589_, _21595_, _21597_);
  or g_32073_(_21590_, _21596_, _21599_);
  and g_32074_(out[65], _21417_, _21600_);
  not g_32075_(_21600_, _21601_);
  or g_32076_(_21349_, _21417_, _21602_);
  not g_32077_(_21602_, _21603_);
  and g_32078_(_21601_, _21602_, _21604_);
  or g_32079_(_21600_, _21603_, _21605_);
  and g_32080_(out[81], _21604_, _21606_);
  or g_32081_(_20586_, _21605_, _21607_);
  and g_32082_(out[64], _21417_, _21608_);
  not g_32083_(_21608_, _21610_);
  or g_32084_(_21362_, _21417_, _21611_);
  not g_32085_(_21611_, _21612_);
  and g_32086_(_21610_, _21611_, _21613_);
  or g_32087_(_21608_, _21612_, _21614_);
  and g_32088_(out[80], _21613_, _21615_);
  or g_32089_(_20597_, _21614_, _21616_);
  xor g_32090_(out[81], _21604_, _21617_);
  xor g_32091_(_20586_, _21604_, _21618_);
  and g_32092_(_21616_, _21617_, _21619_);
  or g_32093_(_21615_, _21618_, _21621_);
  and g_32094_(_21607_, _21621_, _21622_);
  or g_32095_(_21606_, _21619_, _21623_);
  and g_32096_(_21597_, _21623_, _21624_);
  or g_32097_(_21599_, _21622_, _21625_);
  and g_32098_(_21586_, _21592_, _21626_);
  or g_32099_(_21588_, _21591_, _21627_);
  and g_32100_(_21581_, _21627_, _21628_);
  or g_32101_(_21580_, _21626_, _21629_);
  and g_32102_(_21625_, _21628_, _21630_);
  or g_32103_(_21624_, _21629_, _21632_);
  and g_32104_(_21425_, _21560_, _21633_);
  or g_32105_(_21424_, _21561_, _21634_);
  and g_32106_(_21557_, _21634_, _21635_);
  or g_32107_(_21556_, _21633_, _21636_);
  and g_32108_(_21567_, _21635_, _21637_);
  or g_32109_(_21568_, _21636_, _21638_);
  and g_32110_(_21632_, _21637_, _21639_);
  or g_32111_(_21630_, _21638_, _21640_);
  and g_32112_(_21570_, _21640_, _21641_);
  or g_32113_(_21569_, _21639_, _21643_);
  and g_32114_(_21545_, _21643_, _21644_);
  or g_32115_(_21546_, _21641_, _21645_);
  and g_32116_(_21539_, _21645_, _21646_);
  or g_32117_(_21538_, _21644_, _21647_);
  and g_32118_(_21509_, _21647_, _21648_);
  or g_32119_(_21511_, _21646_, _21649_);
  and g_32120_(_21500_, _21649_, _21650_);
  or g_32121_(_21498_, _21648_, _21651_);
  and g_32122_(_20597_, _21614_, _21652_);
  or g_32123_(out[80], _21613_, _21654_);
  and g_32124_(_21545_, _21654_, _21655_);
  or g_32125_(_21546_, _21652_, _21656_);
  and g_32126_(_21597_, _21637_, _21657_);
  or g_32127_(_21599_, _21638_, _21658_);
  and g_32128_(_21619_, _21657_, _21659_);
  or g_32129_(_21621_, _21658_, _21660_);
  and g_32130_(_21655_, _21659_, _21661_);
  or g_32131_(_21656_, _21660_, _21662_);
  and g_32132_(_21509_, _21661_, _21663_);
  or g_32133_(_21511_, _21662_, _21665_);
  and g_32134_(_21651_, _21665_, _21666_);
  or g_32135_(_21650_, _21663_, _21667_);
  or g_32136_(_21424_, _21666_, _21668_);
  or g_32137_(_21560_, _21667_, _21669_);
  and g_32138_(_21668_, _21669_, _21670_);
  not g_32139_(_21670_, _21671_);
  or g_32140_(out[99], _16984_, _21672_);
  not g_32141_(_21672_, _21673_);
  and g_32142_(out[100], _21672_, _21674_);
  or g_32143_(_20707_, _21673_, _21676_);
  and g_32144_(out[101], _21674_, _21677_);
  and g_32145_(out[102], _21677_, _21678_);
  or g_32146_(out[103], _21678_, _21679_);
  and g_32147_(out[104], _21679_, _21680_);
  or g_32148_(out[105], _21680_, _21681_);
  or g_32149_(out[106], _21681_, _21682_);
  xor g_32150_(out[106], _21681_, _21683_);
  not g_32151_(_21683_, _21684_);
  and g_32152_(_21452_, _21667_, _21685_);
  or g_32153_(_21451_, _21666_, _21687_);
  and g_32154_(_21445_, _21666_, _21688_);
  or g_32155_(_21446_, _21667_, _21689_);
  and g_32156_(_21687_, _21689_, _21690_);
  or g_32157_(_21685_, _21688_, _21691_);
  and g_32158_(_21683_, _21690_, _21692_);
  or g_32159_(_21684_, _21691_, _21693_);
  and g_32160_(_21426_, _21440_, _21694_);
  or g_32161_(_21427_, _21441_, _21695_);
  xor g_32162_(out[107], _21682_, _21696_);
  xor g_32163_(_20663_, _21682_, _21698_);
  and g_32164_(_21694_, _21698_, _21699_);
  or g_32165_(_21695_, _21696_, _21700_);
  and g_32166_(_21693_, _21700_, _21701_);
  or g_32167_(_21692_, _21699_, _21702_);
  and g_32168_(_21695_, _21696_, _21703_);
  or g_32169_(_21694_, _21698_, _21704_);
  and g_32170_(_21684_, _21691_, _21705_);
  or g_32171_(_21683_, _21690_, _21706_);
  and g_32172_(_21704_, _21706_, _21707_);
  or g_32173_(_21703_, _21705_, _21709_);
  and g_32174_(out[105], _21680_, _21710_);
  xor g_32175_(out[105], _21680_, _21711_);
  xor g_32176_(_20773_, _21680_, _21712_);
  or g_32177_(_21464_, _21666_, _21713_);
  or g_32178_(_21468_, _21667_, _21714_);
  and g_32179_(_21713_, _21714_, _21715_);
  not g_32180_(_21715_, _21716_);
  or g_32181_(_21711_, _21716_, _21717_);
  xor g_32182_(out[104], _21679_, _21718_);
  xor g_32183_(_20762_, _21679_, _21720_);
  or g_32184_(_21474_, _21667_, _21721_);
  or g_32185_(_21481_, _21666_, _21722_);
  and g_32186_(_21721_, _21722_, _21723_);
  and g_32187_(_21711_, _21716_, _21724_);
  and g_32188_(_21720_, _21723_, _21725_);
  or g_32189_(_21724_, _21725_, _21726_);
  xor g_32190_(_21720_, _21723_, _21727_);
  xor g_32191_(_21718_, _21723_, _21728_);
  and g_32192_(_21701_, _21707_, _21729_);
  or g_32193_(_21702_, _21709_, _21731_);
  xor g_32194_(_21712_, _21715_, _21732_);
  xor g_32195_(_21711_, _21715_, _21733_);
  and g_32196_(_21729_, _21732_, _21734_);
  or g_32197_(_21731_, _21733_, _21735_);
  and g_32198_(_21727_, _21734_, _21736_);
  or g_32199_(_21728_, _21735_, _21737_);
  xor g_32200_(out[101], _21674_, _21738_);
  xor g_32201_(_20696_, _21674_, _21739_);
  or g_32202_(_21547_, _21667_, _21740_);
  or g_32203_(_21553_, _21666_, _21742_);
  and g_32204_(_21740_, _21742_, _21743_);
  not g_32205_(_21743_, _21744_);
  and g_32206_(_21738_, _21744_, _21745_);
  or g_32207_(_21739_, _21743_, _21746_);
  xor g_32208_(out[102], _21677_, _21747_);
  xor g_32209_(_20685_, _21677_, _21748_);
  or g_32210_(_21525_, _21667_, _21749_);
  or g_32211_(_21531_, _21666_, _21750_);
  and g_32212_(_21749_, _21750_, _21751_);
  and g_32213_(_21748_, _21751_, _21753_);
  xor g_32214_(out[103], _21678_, _21754_);
  xor g_32215_(_20674_, _21678_, _21755_);
  or g_32216_(_21518_, _21666_, _21756_);
  or g_32217_(_21513_, _21667_, _21757_);
  and g_32218_(_21756_, _21757_, _21758_);
  not g_32219_(_21758_, _21759_);
  or g_32220_(_21754_, _21758_, _21760_);
  and g_32221_(_21754_, _21758_, _21761_);
  xor g_32222_(_21748_, _21751_, _21762_);
  xor g_32223_(_21754_, _21758_, _21764_);
  and g_32224_(_21762_, _21764_, _21765_);
  not g_32225_(_21765_, _21766_);
  and g_32226_(_21736_, _21746_, _21767_);
  or g_32227_(_21737_, _21745_, _21768_);
  and g_32228_(_21765_, _21767_, _21769_);
  or g_32229_(_21766_, _21768_, _21770_);
  or g_32230_(_15620_, _16984_, _21771_);
  not g_32231_(_21771_, _21772_);
  and g_32232_(_21676_, _21771_, _21773_);
  or g_32233_(_21674_, _21772_, _21775_);
  and g_32234_(_21670_, _21775_, _21776_);
  or g_32235_(_21671_, _21773_, _21777_);
  and g_32236_(_21739_, _21743_, _21778_);
  or g_32237_(_21738_, _21744_, _21779_);
  and g_32238_(_21777_, _21779_, _21780_);
  or g_32239_(_21776_, _21778_, _21781_);
  and g_32240_(_21671_, _21773_, _21782_);
  or g_32241_(_21670_, _21775_, _21783_);
  or g_32242_(_21584_, _21666_, _21784_);
  or g_32243_(_14586_, _21667_, _21786_);
  and g_32244_(_21784_, _21786_, _21787_);
  and g_32245_(_16995_, _21787_, _21788_);
  xor g_32246_(out[99], _16984_, _21789_);
  xor g_32247_(_20751_, _16984_, _21790_);
  and g_32248_(_21579_, _21667_, _21791_);
  or g_32249_(_21578_, _21666_, _21792_);
  and g_32250_(_21571_, _21666_, _21793_);
  or g_32251_(_21572_, _21667_, _21794_);
  and g_32252_(_21792_, _21794_, _21795_);
  or g_32253_(_21791_, _21793_, _21797_);
  and g_32254_(_21789_, _21795_, _21798_);
  or g_32255_(_21788_, _21798_, _21799_);
  or g_32256_(_21789_, _21795_, _21800_);
  xor g_32257_(_16995_, _21787_, _21801_);
  xor g_32258_(_17006_, _21787_, _21802_);
  xor g_32259_(_21789_, _21795_, _21803_);
  xor g_32260_(_21790_, _21795_, _21804_);
  and g_32261_(_21801_, _21803_, _21805_);
  or g_32262_(_21802_, _21804_, _21806_);
  or g_32263_(_20586_, _21667_, _21808_);
  or g_32264_(_21604_, _21666_, _21809_);
  and g_32265_(_21808_, _21809_, _21810_);
  and g_32266_(out[97], _21810_, _21811_);
  not g_32267_(_21811_, _21812_);
  and g_32268_(out[80], _21666_, _21813_);
  or g_32269_(_20597_, _21667_, _21814_);
  and g_32270_(_21614_, _21667_, _21815_);
  or g_32271_(_21613_, _21666_, _21816_);
  and g_32272_(_21814_, _21816_, _21817_);
  or g_32273_(_21813_, _21815_, _21819_);
  and g_32274_(out[96], _21817_, _21820_);
  or g_32275_(_20729_, _21819_, _21821_);
  xor g_32276_(out[97], _21810_, _21822_);
  xor g_32277_(_20718_, _21810_, _21823_);
  and g_32278_(_21821_, _21822_, _21824_);
  or g_32279_(_21820_, _21823_, _21825_);
  and g_32280_(_21812_, _21825_, _21826_);
  or g_32281_(_21811_, _21824_, _21827_);
  and g_32282_(_21805_, _21827_, _21828_);
  or g_32283_(_21806_, _21826_, _21830_);
  and g_32284_(_21799_, _21800_, _21831_);
  not g_32285_(_21831_, _21832_);
  and g_32286_(_21830_, _21832_, _21833_);
  or g_32287_(_21828_, _21831_, _21834_);
  and g_32288_(_21783_, _21834_, _21835_);
  or g_32289_(_21782_, _21833_, _21836_);
  and g_32290_(_21780_, _21836_, _21837_);
  or g_32291_(_21781_, _21835_, _21838_);
  and g_32292_(_21769_, _21838_, _21839_);
  or g_32293_(_21770_, _21837_, _21841_);
  and g_32294_(_21753_, _21760_, _21842_);
  or g_32295_(_21761_, _21842_, _21843_);
  and g_32296_(_21736_, _21843_, _21844_);
  and g_32297_(_21702_, _21704_, _21845_);
  and g_32298_(_21726_, _21729_, _21846_);
  and g_32299_(_21717_, _21846_, _21847_);
  or g_32300_(_21845_, _21847_, _21848_);
  or g_32301_(_21844_, _21848_, _21849_);
  not g_32302_(_21849_, _21850_);
  and g_32303_(_21841_, _21850_, _21852_);
  or g_32304_(_21839_, _21849_, _21853_);
  or g_32305_(out[96], _21817_, _21854_);
  and g_32306_(_21783_, _21854_, _21855_);
  not g_32307_(_21855_, _21856_);
  or g_32308_(_21781_, _21856_, _21857_);
  or g_32309_(_21806_, _21857_, _21858_);
  or g_32310_(_21825_, _21858_, _21859_);
  not g_32311_(_21859_, _21860_);
  and g_32312_(_21769_, _21860_, _21861_);
  or g_32313_(_21770_, _21859_, _21863_);
  and g_32314_(_21853_, _21863_, _21864_);
  or g_32315_(_21852_, _21861_, _21865_);
  and g_32316_(_21671_, _21865_, _21866_);
  and g_32317_(_21775_, _21864_, _21867_);
  or g_32318_(_21866_, _21867_, _21868_);
  and g_32319_(_21694_, _21696_, _21869_);
  or g_32320_(_21695_, _21698_, _21870_);
  or g_32321_(out[115], _17987_, _21871_);
  not g_32322_(_21871_, _21872_);
  and g_32323_(out[116], _21871_, _21874_);
  or g_32324_(_20839_, _21872_, _21875_);
  and g_32325_(out[117], _21874_, _21876_);
  and g_32326_(out[118], _21876_, _21877_);
  or g_32327_(out[119], _21877_, _21878_);
  and g_32328_(out[120], _21878_, _21879_);
  or g_32329_(out[121], _21879_, _21880_);
  or g_32330_(out[122], _21880_, _21881_);
  xor g_32331_(out[123], _21881_, _21882_);
  xor g_32332_(_20795_, _21881_, _21883_);
  or g_32333_(_21870_, _21882_, _21885_);
  xor g_32334_(out[122], _21880_, _21886_);
  not g_32335_(_21886_, _21887_);
  and g_32336_(_21683_, _21864_, _21888_);
  and g_32337_(_21691_, _21865_, _21889_);
  or g_32338_(_21888_, _21889_, _21890_);
  or g_32339_(_21887_, _21890_, _21891_);
  and g_32340_(_21885_, _21891_, _21892_);
  not g_32341_(_21892_, _21893_);
  and g_32342_(_21870_, _21882_, _21894_);
  and g_32343_(_21887_, _21890_, _21896_);
  or g_32344_(_21894_, _21896_, _21897_);
  or g_32345_(_21893_, _21897_, _21898_);
  not g_32346_(_21898_, _21899_);
  and g_32347_(out[121], _21879_, _21900_);
  xor g_32348_(out[121], _21879_, _21901_);
  xor g_32349_(_20894_, _21879_, _21902_);
  or g_32350_(_21715_, _21864_, _21903_);
  not g_32351_(_21903_, _21904_);
  and g_32352_(_21712_, _21864_, _21905_);
  not g_32353_(_21905_, _21907_);
  and g_32354_(_21903_, _21907_, _21908_);
  or g_32355_(_21904_, _21905_, _21909_);
  and g_32356_(_21902_, _21908_, _21910_);
  xor g_32357_(out[120], _21878_, _21911_);
  not g_32358_(_21911_, _21912_);
  and g_32359_(_21720_, _21864_, _21913_);
  or g_32360_(_21723_, _21864_, _21914_);
  not g_32361_(_21914_, _21915_);
  or g_32362_(_21913_, _21915_, _21916_);
  or g_32363_(_21911_, _21916_, _21918_);
  or g_32364_(_21902_, _21908_, _21919_);
  xor g_32365_(_21902_, _21908_, _21920_);
  xor g_32366_(_21901_, _21908_, _21921_);
  xor g_32367_(_21911_, _21916_, _21922_);
  xor g_32368_(_21912_, _21916_, _21923_);
  and g_32369_(_21899_, _21922_, _21924_);
  or g_32370_(_21898_, _21923_, _21925_);
  and g_32371_(_21920_, _21924_, _21926_);
  or g_32372_(_21921_, _21925_, _21927_);
  xor g_32373_(out[118], _21876_, _21929_);
  not g_32374_(_21929_, _21930_);
  or g_32375_(_21751_, _21864_, _21931_);
  not g_32376_(_21931_, _21932_);
  and g_32377_(_21748_, _21864_, _21933_);
  not g_32378_(_21933_, _21934_);
  and g_32379_(_21931_, _21934_, _21935_);
  or g_32380_(_21932_, _21933_, _21936_);
  or g_32381_(_21929_, _21936_, _21937_);
  xor g_32382_(out[119], _21877_, _21938_);
  xor g_32383_(_20806_, _21877_, _21940_);
  and g_32384_(_21754_, _21864_, _21941_);
  and g_32385_(_21759_, _21865_, _21942_);
  or g_32386_(_21941_, _21942_, _21943_);
  or g_32387_(_21940_, _21943_, _21944_);
  and g_32388_(_21937_, _21944_, _21945_);
  xor g_32389_(out[117], _21874_, _21946_);
  xor g_32390_(_20828_, _21874_, _21947_);
  and g_32391_(_21744_, _21865_, _21948_);
  and g_32392_(_21739_, _21864_, _21949_);
  or g_32393_(_21948_, _21949_, _21951_);
  and g_32394_(_21946_, _21951_, _21952_);
  and g_32395_(_21940_, _21943_, _21953_);
  xor g_32396_(_21938_, _21943_, _21954_);
  xor g_32397_(_21929_, _21935_, _21955_);
  or g_32398_(_21952_, _21955_, _21956_);
  or g_32399_(_21954_, _21956_, _21957_);
  or g_32400_(_17743_, _17987_, _21958_);
  not g_32401_(_21958_, _21959_);
  and g_32402_(_21875_, _21958_, _21960_);
  or g_32403_(_21874_, _21959_, _21962_);
  and g_32404_(_21868_, _21960_, _21963_);
  or g_32405_(_21957_, _21963_, _21964_);
  not g_32406_(_21964_, _21965_);
  xor g_32407_(out[115], _17987_, _21966_);
  xor g_32408_(_20872_, _17987_, _21967_);
  and g_32409_(_21789_, _21864_, _21968_);
  or g_32410_(_21790_, _21865_, _21969_);
  and g_32411_(_21797_, _21865_, _21970_);
  or g_32412_(_21795_, _21864_, _21971_);
  and g_32413_(_21969_, _21971_, _21973_);
  or g_32414_(_21968_, _21970_, _21974_);
  or g_32415_(_21967_, _21974_, _21975_);
  or g_32416_(_21787_, _21864_, _21976_);
  not g_32417_(_21976_, _21977_);
  and g_32418_(_16995_, _21864_, _21978_);
  or g_32419_(_21977_, _21978_, _21979_);
  and g_32420_(_21967_, _21974_, _21980_);
  or g_32421_(_17989_, _21979_, _21981_);
  xor g_32422_(_21967_, _21973_, _21982_);
  xor g_32423_(_17988_, _21979_, _21984_);
  or g_32424_(_21982_, _21984_, _21985_);
  and g_32425_(out[97], _21864_, _21986_);
  or g_32426_(_21810_, _21864_, _21987_);
  not g_32427_(_21987_, _21988_);
  or g_32428_(_21986_, _21988_, _21989_);
  or g_32429_(_20850_, _21989_, _21990_);
  xor g_32430_(out[113], _21989_, _21991_);
  or g_32431_(_20729_, _21865_, _21992_);
  or g_32432_(_21817_, _21864_, _21993_);
  and g_32433_(_21992_, _21993_, _21995_);
  and g_32434_(out[112], _21995_, _21996_);
  or g_32435_(_21991_, _21996_, _21997_);
  or g_32436_(_21985_, _21997_, _21998_);
  not g_32437_(_21998_, _21999_);
  or g_32438_(_21985_, _21990_, _22000_);
  or g_32439_(_21980_, _21981_, _22001_);
  and g_32440_(_21975_, _22001_, _22002_);
  and g_32441_(_22000_, _22002_, _22003_);
  and g_32442_(_21998_, _22003_, _22004_);
  or g_32443_(_21964_, _22004_, _22006_);
  or g_32444_(_21945_, _21953_, _22007_);
  or g_32445_(_21868_, _21960_, _22008_);
  or g_32446_(_21946_, _21951_, _22009_);
  and g_32447_(_22008_, _22009_, _22010_);
  or g_32448_(_21957_, _22010_, _22011_);
  and g_32449_(_22007_, _22011_, _22012_);
  and g_32450_(_22006_, _22012_, _22013_);
  or g_32451_(_21927_, _22013_, _22014_);
  or g_32452_(_21892_, _21894_, _22015_);
  and g_32453_(_21918_, _21919_, _22017_);
  or g_32454_(_21897_, _21910_, _22018_);
  or g_32455_(_22017_, _22018_, _22019_);
  and g_32456_(_22015_, _22019_, _22020_);
  and g_32457_(_22014_, _22020_, _22021_);
  or g_32458_(out[112], _21995_, _22022_);
  and g_32459_(_22010_, _22022_, _22023_);
  and g_32460_(_21926_, _22023_, _22024_);
  and g_32461_(_21999_, _22024_, _22025_);
  and g_32462_(_21965_, _22025_, _22026_);
  or g_32463_(_22021_, _22026_, _22028_);
  not g_32464_(_22028_, _22029_);
  and g_32465_(_21868_, _22028_, _22030_);
  not g_32466_(_22030_, _22031_);
  or g_32467_(_21960_, _22028_, _22032_);
  not g_32468_(_22032_, _22033_);
  and g_32469_(_22031_, _22032_, _22034_);
  or g_32470_(_22030_, _22033_, _22035_);
  and g_32471_(_20537_, _22034_, _22036_);
  or g_32472_(_20536_, _22035_, _22037_);
  and g_32473_(out[133], _20532_, _22039_);
  xor g_32474_(out[133], _20532_, _22040_);
  xor g_32475_(_20949_, _20532_, _22041_);
  or g_32476_(_21946_, _22028_, _22042_);
  not g_32477_(_22042_, _22043_);
  and g_32478_(_21951_, _22028_, _22044_);
  not g_32479_(_22044_, _22045_);
  and g_32480_(_22042_, _22045_, _22046_);
  or g_32481_(_22043_, _22044_, _22047_);
  and g_32482_(_22041_, _22046_, _22048_);
  or g_32483_(_22040_, _22047_, _22050_);
  and g_32484_(_22037_, _22050_, _22051_);
  or g_32485_(_22036_, _22048_, _22052_);
  and g_32486_(_20536_, _22035_, _22053_);
  or g_32487_(_20537_, _22034_, _22054_);
  and g_32488_(_21979_, _22028_, _22055_);
  not g_32489_(_22055_, _22056_);
  and g_32490_(_17988_, _22029_, _22057_);
  or g_32491_(_17989_, _22028_, _22058_);
  and g_32492_(_22056_, _22058_, _22059_);
  or g_32493_(_22055_, _22057_, _22061_);
  and g_32494_(_21974_, _22028_, _22062_);
  or g_32495_(_21973_, _22029_, _22063_);
  and g_32496_(_21966_, _22029_, _22064_);
  or g_32497_(_21967_, _22028_, _22065_);
  and g_32498_(_22063_, _22065_, _22066_);
  or g_32499_(_22062_, _22064_, _22067_);
  and g_32500_(_20529_, _22066_, _22068_);
  or g_32501_(_20530_, _22067_, _22069_);
  and g_32502_(_18127_, _22059_, _22070_);
  or g_32503_(_18128_, _22061_, _22072_);
  and g_32504_(_20530_, _22067_, _22073_);
  or g_32505_(_20529_, _22066_, _22074_);
  xor g_32506_(_18127_, _22059_, _22075_);
  xor g_32507_(_18128_, _22059_, _22076_);
  and g_32508_(_22069_, _22075_, _22077_);
  or g_32509_(_22068_, _22076_, _22078_);
  and g_32510_(_22074_, _22077_, _22079_);
  or g_32511_(_22073_, _22078_, _22080_);
  and g_32512_(out[113], _22029_, _22081_);
  or g_32513_(_20850_, _22028_, _22083_);
  and g_32514_(_21989_, _22028_, _22084_);
  not g_32515_(_22084_, _22085_);
  and g_32516_(_22083_, _22085_, _22086_);
  or g_32517_(_22081_, _22084_, _22087_);
  and g_32518_(out[129], _22086_, _22088_);
  or g_32519_(_20971_, _22087_, _22089_);
  and g_32520_(_21995_, _22028_, _22090_);
  not g_32521_(_22090_, _22091_);
  or g_32522_(out[112], _22028_, _22092_);
  not g_32523_(_22092_, _22094_);
  or g_32524_(_22090_, _22094_, _22095_);
  and g_32525_(_22091_, _22092_, _22096_);
  and g_32526_(out[128], _22095_, _22097_);
  or g_32527_(_20982_, _22096_, _22098_);
  xor g_32528_(out[129], _22086_, _22099_);
  xor g_32529_(_20971_, _22086_, _22100_);
  and g_32530_(_22098_, _22099_, _22101_);
  or g_32531_(_22097_, _22100_, _22102_);
  and g_32532_(_22089_, _22102_, _22103_);
  or g_32533_(_22088_, _22101_, _22105_);
  and g_32534_(_22079_, _22105_, _22106_);
  or g_32535_(_22080_, _22103_, _22107_);
  and g_32536_(_22069_, _22072_, _22108_);
  or g_32537_(_22068_, _22070_, _22109_);
  and g_32538_(_22074_, _22109_, _22110_);
  or g_32539_(_22073_, _22108_, _22111_);
  and g_32540_(_22107_, _22111_, _22112_);
  or g_32541_(_22106_, _22110_, _22113_);
  and g_32542_(_22054_, _22113_, _22114_);
  or g_32543_(_22053_, _22112_, _22116_);
  and g_32544_(_22051_, _22116_, _22117_);
  or g_32545_(_22052_, _22114_, _22118_);
  and g_32546_(out[134], _22039_, _22119_);
  or g_32547_(out[135], _22119_, _22120_);
  and g_32548_(out[136], _22120_, _22121_);
  or g_32549_(out[137], _22121_, _22122_);
  or g_32550_(out[138], _22122_, _22123_);
  xor g_32551_(out[138], _22122_, _22124_);
  not g_32552_(_22124_, _22125_);
  and g_32553_(_21886_, _22029_, _22127_);
  and g_32554_(_21890_, _22028_, _22128_);
  or g_32555_(_22127_, _22128_, _22129_);
  or g_32556_(_22125_, _22129_, _22130_);
  and g_32557_(_21869_, _21882_, _22131_);
  or g_32558_(_21870_, _21883_, _22132_);
  xor g_32559_(out[139], _22123_, _22133_);
  or g_32560_(_22132_, _22133_, _22134_);
  and g_32561_(_22130_, _22134_, _22135_);
  and g_32562_(_22132_, _22133_, _22136_);
  xor g_32563_(_22124_, _22129_, _22138_);
  xor g_32564_(_22131_, _22133_, _22139_);
  or g_32565_(_22138_, _22139_, _22140_);
  and g_32566_(out[137], _22121_, _22141_);
  xor g_32567_(out[137], _22121_, _22142_);
  xor g_32568_(_21026_, _22121_, _22143_);
  and g_32569_(_21909_, _22028_, _22144_);
  or g_32570_(_21908_, _22029_, _22145_);
  or g_32571_(_21901_, _22028_, _22146_);
  not g_32572_(_22146_, _22147_);
  and g_32573_(_22145_, _22146_, _22149_);
  or g_32574_(_22144_, _22147_, _22150_);
  and g_32575_(_22143_, _22149_, _22151_);
  xor g_32576_(out[136], _22120_, _22152_);
  xor g_32577_(_21015_, _22120_, _22153_);
  or g_32578_(_21911_, _22028_, _22154_);
  not g_32579_(_22154_, _22155_);
  and g_32580_(_21916_, _22028_, _22156_);
  not g_32581_(_22156_, _22157_);
  and g_32582_(_22154_, _22157_, _22158_);
  or g_32583_(_22155_, _22156_, _22160_);
  and g_32584_(_22152_, _22160_, _22161_);
  or g_32585_(_22151_, _22161_, _22162_);
  and g_32586_(_22142_, _22150_, _22163_);
  or g_32587_(_22143_, _22149_, _22164_);
  and g_32588_(_22153_, _22158_, _22165_);
  or g_32589_(_22152_, _22160_, _22166_);
  and g_32590_(_22164_, _22166_, _22167_);
  or g_32591_(_22163_, _22165_, _22168_);
  or g_32592_(_22162_, _22168_, _22169_);
  or g_32593_(_22140_, _22169_, _22171_);
  xor g_32594_(out[135], _22119_, _22172_);
  xor g_32595_(_20927_, _22119_, _22173_);
  and g_32596_(_21938_, _22029_, _22174_);
  and g_32597_(_21943_, _22028_, _22175_);
  or g_32598_(_22174_, _22175_, _22176_);
  and g_32599_(_22173_, _22176_, _22177_);
  xor g_32600_(out[134], _22039_, _22178_);
  xor g_32601_(_20938_, _22039_, _22179_);
  or g_32602_(_21929_, _22028_, _22180_);
  or g_32603_(_21935_, _22029_, _22182_);
  and g_32604_(_22180_, _22182_, _22183_);
  not g_32605_(_22183_, _22184_);
  or g_32606_(_22178_, _22184_, _22185_);
  or g_32607_(_22173_, _22176_, _22186_);
  and g_32608_(_22040_, _22047_, _22187_);
  xor g_32609_(_22178_, _22183_, _22188_);
  xor g_32610_(_22173_, _22176_, _22189_);
  xor g_32611_(_22172_, _22176_, _22190_);
  or g_32612_(_22187_, _22188_, _22191_);
  or g_32613_(_22171_, _22191_, _22193_);
  not g_32614_(_22193_, _22194_);
  and g_32615_(_22189_, _22194_, _22195_);
  or g_32616_(_22190_, _22193_, _22196_);
  and g_32617_(_22118_, _22195_, _22197_);
  or g_32618_(_22117_, _22196_, _22198_);
  and g_32619_(_22185_, _22186_, _22199_);
  or g_32620_(_22177_, _22199_, _22200_);
  or g_32621_(_22171_, _22200_, _22201_);
  or g_32622_(_22135_, _22136_, _22202_);
  or g_32623_(_22140_, _22167_, _22204_);
  or g_32624_(_22151_, _22204_, _22205_);
  and g_32625_(_22202_, _22205_, _22206_);
  and g_32626_(_22201_, _22206_, _22207_);
  not g_32627_(_22207_, _22208_);
  and g_32628_(_22198_, _22207_, _22209_);
  or g_32629_(_22197_, _22208_, _22210_);
  and g_32630_(_20982_, _22096_, _22211_);
  or g_32631_(_22053_, _22211_, _22212_);
  not g_32632_(_22212_, _22213_);
  and g_32633_(_22051_, _22213_, _22215_);
  and g_32634_(_22079_, _22215_, _22216_);
  and g_32635_(_22101_, _22216_, _22217_);
  not g_32636_(_22217_, _22218_);
  and g_32637_(_22195_, _22217_, _22219_);
  or g_32638_(_22196_, _22218_, _22220_);
  and g_32639_(_22210_, _22220_, _22221_);
  or g_32640_(_22209_, _22219_, _22222_);
  or g_32641_(_20530_, _22222_, _22223_);
  not g_32642_(_22223_, _22224_);
  and g_32643_(_22067_, _22222_, _22226_);
  not g_32644_(_22226_, _22227_);
  and g_32645_(_22223_, _22227_, _22228_);
  or g_32646_(_22224_, _22226_, _22229_);
  or g_32647_(_20526_, _22229_, _22230_);
  and g_32648_(_22061_, _22222_, _22231_);
  and g_32649_(_18127_, _22221_, _22232_);
  or g_32650_(_22231_, _22232_, _22233_);
  and g_32651_(_20526_, _22229_, _22234_);
  or g_32652_(_18338_, _22233_, _22235_);
  xor g_32653_(_20525_, _22228_, _22237_);
  xor g_32654_(_20526_, _22228_, _22238_);
  xor g_32655_(_18338_, _22233_, _22239_);
  xor g_32656_(_18337_, _22233_, _22240_);
  and g_32657_(_22237_, _22239_, _22241_);
  or g_32658_(_22238_, _22240_, _22242_);
  or g_32659_(_20971_, _22222_, _22243_);
  or g_32660_(_22086_, _22221_, _22244_);
  and g_32661_(_22243_, _22244_, _22245_);
  and g_32662_(out[145], _22245_, _22246_);
  and g_32663_(out[128], _22221_, _22248_);
  and g_32664_(_22096_, _22222_, _22249_);
  or g_32665_(_22248_, _22249_, _22250_);
  not g_32666_(_22250_, _22251_);
  or g_32667_(_21114_, _22250_, _22252_);
  xor g_32668_(out[145], _22245_, _22253_);
  and g_32669_(_22252_, _22253_, _22254_);
  or g_32670_(_22246_, _22254_, _22255_);
  not g_32671_(_22255_, _22256_);
  or g_32672_(_22242_, _22256_, _22257_);
  or g_32673_(_22234_, _22235_, _22259_);
  and g_32674_(_22230_, _22259_, _22260_);
  and g_32675_(_22257_, _22260_, _22261_);
  and g_32676_(out[148], _20523_, _22262_);
  or g_32677_(_21081_, _20524_, _22263_);
  and g_32678_(out[149], _22262_, _22264_);
  and g_32679_(out[150], _22264_, _22265_);
  or g_32680_(out[151], _22265_, _22266_);
  xor g_32681_(out[151], _22265_, _22267_);
  xor g_32682_(_21059_, _22265_, _22268_);
  and g_32683_(_22172_, _22221_, _22270_);
  and g_32684_(_22176_, _22222_, _22271_);
  or g_32685_(_22270_, _22271_, _22272_);
  and g_32686_(_22268_, _22272_, _22273_);
  xor g_32687_(out[150], _22264_, _22274_);
  not g_32688_(_22274_, _22275_);
  and g_32689_(_22184_, _22222_, _22276_);
  and g_32690_(_22179_, _22221_, _22277_);
  or g_32691_(_22276_, _22277_, _22278_);
  or g_32692_(_22274_, _22278_, _22279_);
  or g_32693_(_22268_, _22272_, _22281_);
  xor g_32694_(out[149], _22262_, _22282_);
  xor g_32695_(_21092_, _22262_, _22283_);
  or g_32696_(_22040_, _22222_, _22284_);
  not g_32697_(_22284_, _22285_);
  and g_32698_(_22047_, _22222_, _22286_);
  not g_32699_(_22286_, _22287_);
  and g_32700_(_22284_, _22287_, _22288_);
  or g_32701_(_22285_, _22286_, _22289_);
  and g_32702_(_22282_, _22289_, _22290_);
  xor g_32703_(_22267_, _22272_, _22292_);
  xor g_32704_(_22275_, _22278_, _22293_);
  or g_32705_(_22292_, _22293_, _22294_);
  or g_32706_(_22290_, _22294_, _22295_);
  not g_32707_(_22295_, _22296_);
  and g_32708_(_22131_, _22133_, _22297_);
  not g_32709_(_22297_, _22298_);
  and g_32710_(out[152], _22266_, _22299_);
  or g_32711_(out[153], _22299_, _22300_);
  or g_32712_(out[154], _22300_, _22301_);
  xor g_32713_(out[155], _22301_, _22303_);
  not g_32714_(_22303_, _22304_);
  and g_32715_(_22297_, _22304_, _22305_);
  or g_32716_(_22298_, _22303_, _22306_);
  xor g_32717_(out[154], _22300_, _22307_);
  not g_32718_(_22307_, _22308_);
  and g_32719_(_22129_, _22222_, _22309_);
  and g_32720_(_22124_, _22221_, _22310_);
  or g_32721_(_22309_, _22310_, _22311_);
  not g_32722_(_22311_, _22312_);
  and g_32723_(_22307_, _22312_, _22314_);
  or g_32724_(_22308_, _22311_, _22315_);
  and g_32725_(_22306_, _22315_, _22316_);
  or g_32726_(_22305_, _22314_, _22317_);
  and g_32727_(_22298_, _22303_, _22318_);
  or g_32728_(_22297_, _22304_, _22319_);
  and g_32729_(_22308_, _22311_, _22320_);
  or g_32730_(_22307_, _22312_, _22321_);
  or g_32731_(_22318_, _22320_, _22322_);
  and g_32732_(_22316_, _22319_, _22323_);
  and g_32733_(_22321_, _22323_, _22325_);
  or g_32734_(_22317_, _22322_, _22326_);
  xor g_32735_(out[152], _22266_, _22327_);
  xor g_32736_(_21147_, _22266_, _22328_);
  or g_32737_(_22152_, _22222_, _22329_);
  not g_32738_(_22329_, _22330_);
  and g_32739_(_22160_, _22222_, _22331_);
  not g_32740_(_22331_, _22332_);
  and g_32741_(_22329_, _22332_, _22333_);
  or g_32742_(_22330_, _22331_, _22334_);
  or g_32743_(_22327_, _22334_, _22336_);
  xor g_32744_(_22328_, _22333_, _22337_);
  xor g_32745_(_22327_, _22333_, _22338_);
  and g_32746_(out[153], _22299_, _22339_);
  xor g_32747_(out[153], _22299_, _22340_);
  xor g_32748_(_21158_, _22299_, _22341_);
  and g_32749_(_22142_, _22221_, _22342_);
  and g_32750_(_22149_, _22222_, _22343_);
  or g_32751_(_22342_, _22343_, _22344_);
  and g_32752_(_22341_, _22344_, _22345_);
  or g_32753_(_22341_, _22344_, _22347_);
  xor g_32754_(_22341_, _22344_, _22348_);
  xor g_32755_(_22340_, _22344_, _22349_);
  and g_32756_(_22337_, _22348_, _22350_);
  or g_32757_(_22338_, _22349_, _22351_);
  and g_32758_(_22325_, _22350_, _22352_);
  or g_32759_(_22326_, _22351_, _22353_);
  or g_32760_(_21191_, _18336_, _22354_);
  not g_32761_(_22354_, _22355_);
  and g_32762_(_22263_, _22354_, _22356_);
  or g_32763_(_22262_, _22355_, _22358_);
  and g_32764_(_22035_, _22222_, _22359_);
  not g_32765_(_22359_, _22360_);
  or g_32766_(_20536_, _22222_, _22361_);
  not g_32767_(_22361_, _22362_);
  and g_32768_(_22360_, _22361_, _22363_);
  or g_32769_(_22359_, _22362_, _22364_);
  or g_32770_(_22356_, _22364_, _22365_);
  or g_32771_(_22282_, _22289_, _22366_);
  and g_32772_(_22365_, _22366_, _22367_);
  not g_32773_(_22367_, _22369_);
  and g_32774_(_22356_, _22364_, _22370_);
  or g_32775_(_22358_, _22363_, _22371_);
  and g_32776_(_22367_, _22371_, _22372_);
  or g_32777_(_22369_, _22370_, _22373_);
  and g_32778_(_22352_, _22372_, _22374_);
  or g_32779_(_22295_, _22373_, _22375_);
  and g_32780_(_22296_, _22374_, _22376_);
  or g_32781_(_22316_, _22318_, _22377_);
  and g_32782_(_22336_, _22347_, _22378_);
  or g_32783_(_22345_, _22378_, _22380_);
  or g_32784_(_22326_, _22380_, _22381_);
  and g_32785_(_22377_, _22381_, _22382_);
  or g_32786_(_22295_, _22367_, _22383_);
  or g_32787_(_22273_, _22279_, _22384_);
  and g_32788_(_22281_, _22384_, _22385_);
  and g_32789_(_22383_, _22385_, _22386_);
  or g_32790_(_22261_, _22375_, _22387_);
  and g_32791_(_22386_, _22387_, _22388_);
  or g_32792_(_22353_, _22388_, _22389_);
  and g_32793_(_22382_, _22389_, _22391_);
  or g_32794_(out[144], _22251_, _22392_);
  and g_32795_(_22241_, _22392_, _22393_);
  and g_32796_(_22254_, _22393_, _22394_);
  and g_32797_(_22376_, _22394_, _22395_);
  or g_32798_(_22391_, _22395_, _22396_);
  not g_32799_(_22396_, _22397_);
  and g_32800_(_22245_, _22396_, _22398_);
  not g_32801_(_22398_, _22399_);
  or g_32802_(out[145], _22396_, _22400_);
  not g_32803_(_22400_, _22402_);
  or g_32804_(_22398_, _22402_, _22403_);
  and g_32805_(_22399_, _22400_, _22404_);
  or g_32806_(out[307], _20292_, _22405_);
  not g_32807_(_22405_, _22406_);
  and g_32808_(out[308], _22405_, _22407_);
  or g_32809_(_19772_, _22406_, _22408_);
  and g_32810_(out[309], _22407_, _22409_);
  and g_32811_(out[310], _22409_, _22410_);
  xor g_32812_(out[310], _22409_, _22411_);
  not g_32813_(_22411_, _22413_);
  or g_32814_(out[291], _20106_, _22414_);
  not g_32815_(_22414_, _22415_);
  and g_32816_(out[292], _22414_, _22416_);
  or g_32817_(_19662_, _22415_, _22417_);
  and g_32818_(out[293], _22416_, _22418_);
  and g_32819_(out[294], _22418_, _22419_);
  xor g_32820_(out[294], _22418_, _22420_);
  not g_32821_(_22420_, _22421_);
  or g_32822_(out[295], _22419_, _22422_);
  and g_32823_(out[296], _22422_, _22424_);
  or g_32824_(out[297], _22424_, _22425_);
  not g_32825_(_22425_, _22426_);
  or g_32826_(out[298], _22425_, _22427_);
  xor g_32827_(out[298], _22425_, _22428_);
  xor g_32828_(_19728_, _22425_, _22429_);
  or g_32829_(out[195], _18741_, _22430_);
  not g_32830_(_22430_, _22431_);
  and g_32831_(out[196], _22430_, _22432_);
  or g_32832_(_18892_, _22431_, _22433_);
  and g_32833_(out[197], _22432_, _22435_);
  and g_32834_(out[198], _22435_, _22436_);
  or g_32835_(out[199], _22436_, _22437_);
  and g_32836_(out[200], _22437_, _22438_);
  or g_32837_(out[201], _22438_, _22439_);
  not g_32838_(_22439_, _22440_);
  or g_32839_(out[202], _22439_, _22441_);
  xor g_32840_(out[202], _22439_, _22442_);
  xor g_32841_(out[202], _22440_, _22443_);
  or g_32842_(out[163], _18467_, _22444_);
  and g_32843_(out[164], _22444_, _22446_);
  not g_32844_(_22446_, _22447_);
  and g_32845_(out[165], _22446_, _22448_);
  and g_32846_(out[166], _22448_, _22449_);
  or g_32847_(out[167], _22449_, _22450_);
  and g_32848_(out[168], _22450_, _22451_);
  or g_32849_(out[169], _22451_, _22452_);
  or g_32850_(out[170], _22452_, _22453_);
  xor g_32851_(out[171], _22453_, _22454_);
  xor g_32852_(_18595_, _22453_, _22455_);
  or g_32853_(out[179], _18463_, _22457_);
  and g_32854_(out[180], _22457_, _22458_);
  not g_32855_(_22458_, _22459_);
  and g_32856_(out[181], _22458_, _22460_);
  and g_32857_(out[182], _22460_, _22461_);
  or g_32858_(out[183], _22461_, _22462_);
  and g_32859_(out[184], _22462_, _22463_);
  or g_32860_(out[185], _22463_, _22464_);
  or g_32861_(out[186], _22464_, _22465_);
  xor g_32862_(out[187], _22465_, _22466_);
  xor g_32863_(_18716_, _22465_, _22468_);
  and g_32864_(_22454_, _22466_, _22469_);
  or g_32865_(_22455_, _22468_, _22470_);
  xor g_32866_(out[203], _22441_, _22471_);
  xor g_32867_(_18848_, _22441_, _22472_);
  and g_32868_(_22469_, _22472_, _22473_);
  or g_32869_(_22470_, _22471_, _22474_);
  xor g_32870_(out[170], _22452_, _22475_);
  xor g_32871_(_18705_, _22452_, _22476_);
  xor g_32872_(out[186], _22464_, _22477_);
  xor g_32873_(_18837_, _22464_, _22479_);
  and g_32874_(_22476_, _22477_, _22480_);
  or g_32875_(_22475_, _22479_, _22481_);
  and g_32876_(_22454_, _22468_, _22482_);
  or g_32877_(_22455_, _22466_, _22483_);
  and g_32878_(_22481_, _22483_, _22484_);
  or g_32879_(_22480_, _22482_, _22485_);
  and g_32880_(_22455_, _22466_, _22486_);
  or g_32881_(_22454_, _22468_, _22487_);
  and g_32882_(out[169], _22451_, _22488_);
  xor g_32883_(out[169], _22451_, _22490_);
  xor g_32884_(_18694_, _22451_, _22491_);
  and g_32885_(out[185], _22463_, _22492_);
  xor g_32886_(out[185], _22463_, _22493_);
  xor g_32887_(_18826_, _22463_, _22494_);
  and g_32888_(_22491_, _22493_, _22495_);
  or g_32889_(_22490_, _22494_, _22496_);
  and g_32890_(_22490_, _22494_, _22497_);
  or g_32891_(_22491_, _22493_, _22498_);
  and g_32892_(_22496_, _22498_, _22499_);
  or g_32893_(_22495_, _22497_, _22501_);
  xor g_32894_(out[168], _22450_, _22502_);
  xor g_32895_(_18683_, _22450_, _22503_);
  xor g_32896_(out[184], _22462_, _22504_);
  xor g_32897_(_18815_, _22462_, _22505_);
  and g_32898_(_22502_, _22505_, _22506_);
  or g_32899_(_22503_, _22504_, _22507_);
  xor g_32900_(_22503_, _22504_, _22508_);
  xor g_32901_(_22502_, _22504_, _22509_);
  and g_32902_(_22499_, _22508_, _22510_);
  or g_32903_(_22501_, _22509_, _22512_);
  and g_32904_(_22475_, _22479_, _22513_);
  or g_32905_(_22476_, _22477_, _22514_);
  and g_32906_(_22510_, _22514_, _22515_);
  or g_32907_(_22512_, _22513_, _22516_);
  and g_32908_(_22487_, _22515_, _22517_);
  or g_32909_(_22486_, _22516_, _22518_);
  and g_32910_(_22484_, _22517_, _22519_);
  or g_32911_(_22485_, _22518_, _22520_);
  xor g_32912_(out[166], _22448_, _22521_);
  not g_32913_(_22521_, _22523_);
  xor g_32914_(out[182], _22460_, _22524_);
  or g_32915_(_22523_, _22524_, _22525_);
  xor g_32916_(out[167], _22449_, _22526_);
  xor g_32917_(_18606_, _22449_, _22527_);
  xor g_32918_(_18727_, _22461_, _22528_);
  or g_32919_(_22526_, _22528_, _22529_);
  and g_32920_(_22525_, _22529_, _22530_);
  and g_32921_(_22526_, _22528_, _22531_);
  xor g_32922_(_22523_, _22524_, _22532_);
  xor g_32923_(_22521_, _22524_, _22534_);
  xor g_32924_(_22526_, _22528_, _22535_);
  xor g_32925_(_22527_, _22528_, _22536_);
  and g_32926_(_22532_, _22535_, _22537_);
  or g_32927_(_22534_, _22536_, _22538_);
  or g_32928_(_18434_, _18467_, _22539_);
  not g_32929_(_22539_, _22540_);
  and g_32930_(_22447_, _22539_, _22541_);
  or g_32931_(_22446_, _22540_, _22542_);
  or g_32932_(_18422_, _18463_, _22543_);
  not g_32933_(_22543_, _22545_);
  and g_32934_(_22459_, _22543_, _22546_);
  or g_32935_(_22458_, _22545_, _22547_);
  and g_32936_(_22541_, _22547_, _22548_);
  or g_32937_(_22542_, _22546_, _22549_);
  xor g_32938_(out[165], _22446_, _22550_);
  xor g_32939_(_18628_, _22446_, _22551_);
  xor g_32940_(out[181], _22458_, _22552_);
  xor g_32941_(_18749_, _22458_, _22553_);
  and g_32942_(_22550_, _22553_, _22554_);
  or g_32943_(_22551_, _22552_, _22556_);
  and g_32944_(_22549_, _22556_, _22557_);
  or g_32945_(_22548_, _22554_, _22558_);
  and g_32946_(_22551_, _22552_, _22559_);
  or g_32947_(_22550_, _22553_, _22560_);
  and g_32948_(_22542_, _22546_, _22561_);
  or g_32949_(_22541_, _22547_, _22562_);
  and g_32950_(_22560_, _22562_, _22563_);
  or g_32951_(_22559_, _22561_, _22564_);
  and g_32952_(_22557_, _22563_, _22565_);
  or g_32953_(_22558_, _22564_, _22567_);
  and g_32954_(_22537_, _22565_, _22568_);
  or g_32955_(_22538_, _22567_, _22569_);
  and g_32956_(_18510_, _22568_, _22570_);
  or g_32957_(_18511_, _22569_, _22571_);
  and g_32958_(_22519_, _22570_, _22572_);
  or g_32959_(_22520_, _22571_, _22573_);
  xor g_32960_(out[163], _18467_, _22574_);
  xor g_32961_(_18672_, _18467_, _22575_);
  xor g_32962_(out[179], _18463_, _22576_);
  xor g_32963_(_18804_, _18463_, _22578_);
  or g_32964_(_22574_, _22578_, _22579_);
  and g_32965_(_18473_, _22579_, _22580_);
  and g_32966_(_22574_, _22578_, _22581_);
  or g_32967_(_22580_, _22581_, _22582_);
  and g_32968_(_18493_, _22582_, _22583_);
  or g_32969_(_22569_, _22583_, _22584_);
  or g_32970_(_22530_, _22531_, _22585_);
  or g_32971_(_22557_, _22559_, _22586_);
  or g_32972_(_22538_, _22586_, _22587_);
  and g_32973_(_22585_, _22587_, _22589_);
  and g_32974_(_22584_, _22589_, _22590_);
  not g_32975_(_22590_, _22591_);
  and g_32976_(_22519_, _22591_, _22592_);
  or g_32977_(_22520_, _22590_, _22593_);
  and g_32978_(_22499_, _22506_, _22594_);
  or g_32979_(_22501_, _22507_, _22595_);
  and g_32980_(_22496_, _22595_, _22596_);
  or g_32981_(_22495_, _22594_, _22597_);
  and g_32982_(_22514_, _22597_, _22598_);
  or g_32983_(_22513_, _22596_, _22600_);
  and g_32984_(_22484_, _22600_, _22601_);
  or g_32985_(_22485_, _22598_, _22602_);
  and g_32986_(_22487_, _22602_, _22603_);
  or g_32987_(_22486_, _22601_, _22604_);
  and g_32988_(_22593_, _22604_, _22605_);
  or g_32989_(_22592_, _22603_, _22606_);
  and g_32990_(_22573_, _22606_, _22607_);
  or g_32991_(_22572_, _22605_, _22608_);
  and g_32992_(_22475_, _22608_, _22609_);
  or g_32993_(_22476_, _22607_, _22611_);
  and g_32994_(_22477_, _22607_, _22612_);
  or g_32995_(_22479_, _22608_, _22613_);
  and g_32996_(_22611_, _22613_, _22614_);
  or g_32997_(_22609_, _22612_, _22615_);
  and g_32998_(_22442_, _22614_, _22616_);
  or g_32999_(_22443_, _22615_, _22617_);
  and g_33000_(_22474_, _22617_, _22618_);
  or g_33001_(_22473_, _22616_, _22619_);
  and g_33002_(_22443_, _22615_, _22620_);
  or g_33003_(_22442_, _22614_, _22622_);
  and g_33004_(_22470_, _22471_, _22623_);
  or g_33005_(_22469_, _22472_, _22624_);
  and g_33006_(out[201], _22438_, _22625_);
  xor g_33007_(out[201], _22438_, _22626_);
  or g_33008_(_22440_, _22625_, _22627_);
  and g_33009_(_22490_, _22608_, _22628_);
  or g_33010_(_22491_, _22607_, _22629_);
  and g_33011_(_22493_, _22607_, _22630_);
  or g_33012_(_22494_, _22608_, _22631_);
  and g_33013_(_22629_, _22631_, _22633_);
  or g_33014_(_22628_, _22630_, _22634_);
  and g_33015_(_22627_, _22634_, _22635_);
  or g_33016_(_22626_, _22633_, _22636_);
  and g_33017_(_22624_, _22636_, _22637_);
  or g_33018_(_22623_, _22635_, _22638_);
  and g_33019_(_22622_, _22637_, _22639_);
  or g_33020_(_22620_, _22638_, _22640_);
  and g_33021_(_22618_, _22639_, _22641_);
  or g_33022_(_22619_, _22640_, _22642_);
  and g_33023_(_22626_, _22633_, _22644_);
  or g_33024_(_22627_, _22634_, _22645_);
  xor g_33025_(out[200], _22437_, _22646_);
  xor g_33026_(_18947_, _22437_, _22647_);
  and g_33027_(_22503_, _22608_, _22648_);
  or g_33028_(_22502_, _22607_, _22649_);
  or g_33029_(_22504_, _22608_, _22650_);
  not g_33030_(_22650_, _22651_);
  and g_33031_(_22649_, _22650_, _22652_);
  or g_33032_(_22648_, _22651_, _22653_);
  and g_33033_(_22647_, _22652_, _22655_);
  or g_33034_(_22646_, _22653_, _22656_);
  and g_33035_(_22645_, _22656_, _22657_);
  or g_33036_(_22644_, _22655_, _22658_);
  and g_33037_(_22646_, _22653_, _22659_);
  or g_33038_(_22647_, _22652_, _22660_);
  and g_33039_(_22657_, _22660_, _22661_);
  or g_33040_(_22658_, _22659_, _22662_);
  and g_33041_(_22641_, _22661_, _22663_);
  or g_33042_(_22642_, _22662_, _22664_);
  xor g_33043_(out[199], _22436_, _22666_);
  not g_33044_(_22666_, _22667_);
  or g_33045_(_22528_, _22608_, _22668_);
  or g_33046_(_22527_, _22607_, _22669_);
  and g_33047_(_22668_, _22669_, _22670_);
  and g_33048_(_22666_, _22670_, _22671_);
  or g_33049_(_22666_, _22670_, _22672_);
  xor g_33050_(_22666_, _22670_, _22673_);
  xor g_33051_(_22667_, _22670_, _22674_);
  xor g_33052_(out[198], _22435_, _22675_);
  xor g_33053_(_18870_, _22435_, _22677_);
  or g_33054_(_22521_, _22607_, _22678_);
  or g_33055_(_22524_, _22608_, _22679_);
  and g_33056_(_22678_, _22679_, _22680_);
  and g_33057_(_22677_, _22680_, _22681_);
  xor g_33058_(_22677_, _22680_, _22682_);
  xor g_33059_(_22675_, _22680_, _22683_);
  and g_33060_(_22673_, _22682_, _22684_);
  or g_33061_(_22674_, _22683_, _22685_);
  or g_33062_(_18601_, _18741_, _22686_);
  not g_33063_(_22686_, _22688_);
  and g_33064_(_22433_, _22686_, _22689_);
  or g_33065_(_22432_, _22688_, _22690_);
  and g_33066_(_22542_, _22608_, _22691_);
  or g_33067_(_22541_, _22607_, _22692_);
  and g_33068_(_22547_, _22607_, _22693_);
  or g_33069_(_22546_, _22608_, _22694_);
  and g_33070_(_22692_, _22694_, _22695_);
  or g_33071_(_22691_, _22693_, _22696_);
  and g_33072_(_22690_, _22695_, _22697_);
  or g_33073_(_22689_, _22696_, _22699_);
  xor g_33074_(out[197], _22432_, _22700_);
  xor g_33075_(_18881_, _22432_, _22701_);
  and g_33076_(_22551_, _22608_, _22702_);
  or g_33077_(_22550_, _22607_, _22703_);
  and g_33078_(_22553_, _22607_, _22704_);
  or g_33079_(_22552_, _22608_, _22705_);
  and g_33080_(_22703_, _22705_, _22706_);
  or g_33081_(_22702_, _22704_, _22707_);
  and g_33082_(_22701_, _22706_, _22708_);
  or g_33083_(_22700_, _22707_, _22710_);
  and g_33084_(_22699_, _22710_, _22711_);
  or g_33085_(_22697_, _22708_, _22712_);
  and g_33086_(_22700_, _22707_, _22713_);
  or g_33087_(_22701_, _22706_, _22714_);
  and g_33088_(_22689_, _22696_, _22715_);
  or g_33089_(_22690_, _22695_, _22716_);
  and g_33090_(_22714_, _22716_, _22717_);
  or g_33091_(_22713_, _22715_, _22718_);
  and g_33092_(_22711_, _22717_, _22719_);
  or g_33093_(_22712_, _22718_, _22721_);
  and g_33094_(_22684_, _22719_, _22722_);
  or g_33095_(_22685_, _22721_, _22723_);
  and g_33096_(_22663_, _22722_, _22724_);
  or g_33097_(_22664_, _22723_, _22725_);
  xor g_33098_(out[195], _18741_, _22726_);
  xor g_33099_(_18936_, _18741_, _22727_);
  and g_33100_(_22576_, _22607_, _22728_);
  and g_33101_(_22574_, _22608_, _22729_);
  or g_33102_(_22728_, _22729_, _22730_);
  not g_33103_(_22730_, _22732_);
  or g_33104_(_22727_, _22730_, _22733_);
  and g_33105_(_18468_, _22608_, _22734_);
  and g_33106_(_18465_, _22607_, _22735_);
  or g_33107_(_22734_, _22735_, _22736_);
  not g_33108_(_22736_, _22737_);
  or g_33109_(_18743_, _22736_, _22738_);
  and g_33110_(_22733_, _22738_, _22739_);
  and g_33111_(_22727_, _22730_, _22740_);
  or g_33112_(_22726_, _22732_, _22741_);
  or g_33113_(_18742_, _22737_, _22743_);
  and g_33114_(_22741_, _22743_, _22744_);
  xor g_33115_(_22726_, _22730_, _22745_);
  xor g_33116_(_18742_, _22736_, _22746_);
  and g_33117_(_22739_, _22744_, _22747_);
  or g_33118_(_22745_, _22746_, _22748_);
  or g_33119_(_18771_, _22608_, _22749_);
  or g_33120_(_18650_, _22607_, _22750_);
  and g_33121_(_22749_, _22750_, _22751_);
  and g_33122_(out[193], _22751_, _22752_);
  not g_33123_(_22752_, _22754_);
  and g_33124_(_18584_, _22608_, _22755_);
  or g_33125_(out[160], _22607_, _22756_);
  or g_33126_(out[176], _22608_, _22757_);
  not g_33127_(_22757_, _22758_);
  and g_33128_(_22756_, _22757_, _22759_);
  or g_33129_(_22755_, _22758_, _22760_);
  and g_33130_(out[192], _22760_, _22761_);
  or g_33131_(_18914_, _22759_, _22762_);
  xor g_33132_(out[193], _22751_, _22763_);
  xor g_33133_(_18903_, _22751_, _22765_);
  and g_33134_(_22762_, _22763_, _22766_);
  or g_33135_(_22761_, _22765_, _22767_);
  and g_33136_(_22754_, _22767_, _22768_);
  or g_33137_(_22752_, _22766_, _22769_);
  and g_33138_(_22747_, _22769_, _22770_);
  or g_33139_(_22748_, _22768_, _22771_);
  or g_33140_(_22739_, _22740_, _22772_);
  not g_33141_(_22772_, _22773_);
  and g_33142_(_22771_, _22772_, _22774_);
  or g_33143_(_22770_, _22773_, _22776_);
  and g_33144_(_22724_, _22776_, _22777_);
  or g_33145_(_22725_, _22774_, _22778_);
  and g_33146_(_22684_, _22712_, _22779_);
  or g_33147_(_22685_, _22711_, _22780_);
  and g_33148_(_22714_, _22779_, _22781_);
  or g_33149_(_22713_, _22780_, _22782_);
  and g_33150_(_22672_, _22681_, _22783_);
  or g_33151_(_22671_, _22783_, _22784_);
  not g_33152_(_22784_, _22785_);
  and g_33153_(_22782_, _22785_, _22787_);
  or g_33154_(_22781_, _22784_, _22788_);
  and g_33155_(_22663_, _22788_, _22789_);
  or g_33156_(_22664_, _22787_, _22790_);
  and g_33157_(_22641_, _22658_, _22791_);
  or g_33158_(_22642_, _22657_, _22792_);
  and g_33159_(_22619_, _22624_, _22793_);
  or g_33160_(_22618_, _22623_, _22794_);
  and g_33161_(_22792_, _22794_, _22795_);
  or g_33162_(_22791_, _22793_, _22796_);
  and g_33163_(_22790_, _22795_, _22798_);
  or g_33164_(_22789_, _22796_, _22799_);
  and g_33165_(_22778_, _22798_, _22800_);
  or g_33166_(_22777_, _22799_, _22801_);
  and g_33167_(_18914_, _22759_, _22802_);
  or g_33168_(out[192], _22760_, _22803_);
  and g_33169_(_22747_, _22803_, _22804_);
  or g_33170_(_22748_, _22802_, _22805_);
  and g_33171_(_22766_, _22804_, _22806_);
  or g_33172_(_22767_, _22805_, _22807_);
  and g_33173_(_22724_, _22806_, _22809_);
  or g_33174_(_22725_, _22807_, _22810_);
  and g_33175_(_22801_, _22810_, _22811_);
  or g_33176_(_22800_, _22809_, _22812_);
  and g_33177_(_22442_, _22811_, _22813_);
  or g_33178_(_22443_, _22812_, _22814_);
  and g_33179_(_22615_, _22812_, _22815_);
  or g_33180_(_22614_, _22811_, _22816_);
  and g_33181_(_22814_, _22816_, _22817_);
  or g_33182_(_22813_, _22815_, _22818_);
  or g_33183_(out[211], _18849_, _22820_);
  not g_33184_(_22820_, _22821_);
  and g_33185_(out[212], _22820_, _22822_);
  or g_33186_(_19002_, _22821_, _22823_);
  and g_33187_(out[213], _22822_, _22824_);
  and g_33188_(out[214], _22824_, _22825_);
  xor g_33189_(out[214], _22824_, _22826_);
  xor g_33190_(_18980_, _22824_, _22827_);
  or g_33191_(_22675_, _22812_, _22828_);
  or g_33192_(_22680_, _22811_, _22829_);
  and g_33193_(_22828_, _22829_, _22831_);
  and g_33194_(_22827_, _22831_, _22832_);
  xor g_33195_(out[213], _22822_, _22833_);
  xor g_33196_(_18991_, _22822_, _22834_);
  or g_33197_(_22700_, _22812_, _22835_);
  or g_33198_(_22706_, _22811_, _22836_);
  and g_33199_(_22835_, _22836_, _22837_);
  or g_33200_(_22834_, _22837_, _22838_);
  not g_33201_(_22838_, _22839_);
  or g_33202_(out[215], _22825_, _22840_);
  xor g_33203_(out[215], _22825_, _22842_);
  xor g_33204_(_18969_, _22825_, _22843_);
  or g_33205_(_22667_, _22812_, _22844_);
  or g_33206_(_22670_, _22811_, _22845_);
  and g_33207_(_22844_, _22845_, _22846_);
  and g_33208_(_22842_, _22846_, _22847_);
  or g_33209_(_22842_, _22846_, _22848_);
  xor g_33210_(_22842_, _22846_, _22849_);
  xor g_33211_(_22843_, _22846_, _22850_);
  xor g_33212_(_22827_, _22831_, _22851_);
  xor g_33213_(_22826_, _22831_, _22853_);
  and g_33214_(_22849_, _22851_, _22854_);
  or g_33215_(_22850_, _22853_, _22855_);
  and g_33216_(_22838_, _22854_, _22856_);
  or g_33217_(_22839_, _22855_, _22857_);
  or g_33218_(_18849_, _18897_, _22858_);
  not g_33219_(_22858_, _22859_);
  and g_33220_(_22823_, _22858_, _22860_);
  or g_33221_(_22822_, _22859_, _22861_);
  or g_33222_(_22695_, _22811_, _22862_);
  or g_33223_(_22689_, _22812_, _22864_);
  and g_33224_(_22862_, _22864_, _22865_);
  and g_33225_(_22861_, _22865_, _22866_);
  not g_33226_(_22866_, _22867_);
  and g_33227_(_22834_, _22837_, _22868_);
  not g_33228_(_22868_, _22869_);
  and g_33229_(_22867_, _22869_, _22870_);
  or g_33230_(_22866_, _22868_, _22871_);
  or g_33231_(_22861_, _22865_, _22872_);
  not g_33232_(_22872_, _22873_);
  and g_33233_(_22870_, _22872_, _22875_);
  or g_33234_(_22871_, _22873_, _22876_);
  and g_33235_(_22856_, _22875_, _22877_);
  or g_33236_(_22857_, _22876_, _22878_);
  and g_33237_(out[216], _22840_, _22879_);
  or g_33238_(out[217], _22879_, _22880_);
  not g_33239_(_22880_, _22881_);
  or g_33240_(out[218], _22880_, _22882_);
  xor g_33241_(out[218], _22880_, _22883_);
  xor g_33242_(_19079_, _22880_, _22884_);
  and g_33243_(_22817_, _22883_, _22886_);
  or g_33244_(_22818_, _22884_, _22887_);
  and g_33245_(_22469_, _22471_, _22888_);
  or g_33246_(_22470_, _22472_, _22889_);
  xor g_33247_(out[219], _22882_, _22890_);
  xor g_33248_(_18958_, _22882_, _22891_);
  and g_33249_(_22888_, _22891_, _22892_);
  or g_33250_(_22889_, _22890_, _22893_);
  and g_33251_(_22887_, _22893_, _22894_);
  or g_33252_(_22886_, _22892_, _22895_);
  and g_33253_(_22889_, _22890_, _22897_);
  or g_33254_(_22888_, _22891_, _22898_);
  and g_33255_(_22818_, _22884_, _22899_);
  or g_33256_(_22817_, _22883_, _22900_);
  and g_33257_(_22898_, _22900_, _22901_);
  or g_33258_(_22897_, _22899_, _22902_);
  and g_33259_(_22894_, _22901_, _22903_);
  or g_33260_(_22895_, _22902_, _22904_);
  xor g_33261_(out[216], _22840_, _22905_);
  xor g_33262_(_19057_, _22840_, _22906_);
  or g_33263_(_22646_, _22812_, _22908_);
  or g_33264_(_22652_, _22811_, _22909_);
  and g_33265_(_22908_, _22909_, _22910_);
  not g_33266_(_22910_, _22911_);
  or g_33267_(_22906_, _22910_, _22912_);
  not g_33268_(_22912_, _22913_);
  or g_33269_(_22626_, _22812_, _22914_);
  or g_33270_(_22634_, _22811_, _22915_);
  and g_33271_(_22914_, _22915_, _22916_);
  not g_33272_(_22916_, _22917_);
  and g_33273_(out[217], _22879_, _22919_);
  xor g_33274_(out[217], _22879_, _22920_);
  or g_33275_(_22881_, _22919_, _22921_);
  and g_33276_(_22916_, _22921_, _22922_);
  or g_33277_(_22917_, _22920_, _22923_);
  and g_33278_(_22912_, _22923_, _22924_);
  or g_33279_(_22913_, _22922_, _22925_);
  or g_33280_(_22916_, _22921_, _22926_);
  not g_33281_(_22926_, _22927_);
  and g_33282_(_22906_, _22910_, _22928_);
  or g_33283_(_22905_, _22911_, _22930_);
  and g_33284_(_22926_, _22930_, _22931_);
  or g_33285_(_22927_, _22928_, _22932_);
  and g_33286_(_22924_, _22931_, _22933_);
  or g_33287_(_22925_, _22932_, _22934_);
  and g_33288_(_22903_, _22933_, _22935_);
  or g_33289_(_22904_, _22934_, _22936_);
  or g_33290_(_18903_, _22812_, _22937_);
  or g_33291_(_22751_, _22811_, _22938_);
  and g_33292_(_22937_, _22938_, _22939_);
  and g_33293_(out[192], _22811_, _22941_);
  or g_33294_(_18914_, _22812_, _22942_);
  and g_33295_(_22759_, _22812_, _22943_);
  or g_33296_(_22760_, _22811_, _22944_);
  and g_33297_(_22942_, _22944_, _22945_);
  or g_33298_(_22941_, _22943_, _22946_);
  and g_33299_(out[208], _22945_, _22947_);
  or g_33300_(_19024_, _22946_, _22948_);
  and g_33301_(out[209], _22939_, _22949_);
  not g_33302_(_22949_, _22950_);
  xor g_33303_(out[209], _22939_, _22952_);
  xor g_33304_(_19013_, _22939_, _22953_);
  and g_33305_(_22948_, _22952_, _22954_);
  or g_33306_(_22947_, _22953_, _22955_);
  or g_33307_(_22737_, _22811_, _22956_);
  or g_33308_(_18743_, _22812_, _22957_);
  and g_33309_(_22956_, _22957_, _22958_);
  not g_33310_(_22958_, _22959_);
  and g_33311_(_18850_, _22958_, _22960_);
  not g_33312_(_22960_, _22961_);
  xor g_33313_(out[211], _18849_, _22963_);
  xor g_33314_(_19046_, _18849_, _22964_);
  or g_33315_(_22727_, _22812_, _22965_);
  or g_33316_(_22732_, _22811_, _22966_);
  and g_33317_(_22965_, _22966_, _22967_);
  not g_33318_(_22967_, _22968_);
  and g_33319_(_22963_, _22967_, _22969_);
  not g_33320_(_22969_, _22970_);
  and g_33321_(_22961_, _22970_, _22971_);
  or g_33322_(_22960_, _22969_, _22972_);
  and g_33323_(_22964_, _22968_, _22974_);
  or g_33324_(_22963_, _22967_, _22975_);
  and g_33325_(_18851_, _22959_, _22976_);
  or g_33326_(_18850_, _22958_, _22977_);
  and g_33327_(_19024_, _22946_, _22978_);
  or g_33328_(_22972_, _22976_, _22979_);
  or g_33329_(_22974_, _22978_, _22980_);
  or g_33330_(_22955_, _22980_, _22981_);
  or g_33331_(_22979_, _22981_, _22982_);
  not g_33332_(_22982_, _22983_);
  and g_33333_(_22935_, _22983_, _22985_);
  or g_33334_(_22936_, _22982_, _22986_);
  and g_33335_(_22877_, _22985_, _22987_);
  or g_33336_(_22878_, _22986_, _22988_);
  and g_33337_(_22950_, _22955_, _22989_);
  or g_33338_(_22949_, _22954_, _22990_);
  and g_33339_(_22977_, _22990_, _22991_);
  or g_33340_(_22976_, _22989_, _22992_);
  and g_33341_(_22971_, _22992_, _22993_);
  or g_33342_(_22972_, _22991_, _22994_);
  or g_33343_(_22878_, _22974_, _22996_);
  and g_33344_(_22877_, _22994_, _22997_);
  and g_33345_(_22975_, _22997_, _22998_);
  or g_33346_(_22993_, _22996_, _22999_);
  and g_33347_(_22856_, _22871_, _23000_);
  and g_33348_(_22832_, _22848_, _23001_);
  or g_33349_(_22847_, _23001_, _23002_);
  or g_33350_(_23000_, _23002_, _23003_);
  not g_33351_(_23003_, _23004_);
  and g_33352_(_22999_, _23004_, _23005_);
  or g_33353_(_22998_, _23003_, _23007_);
  and g_33354_(_22935_, _23007_, _23008_);
  or g_33355_(_22936_, _23005_, _23009_);
  and g_33356_(_22895_, _22898_, _23010_);
  or g_33357_(_22894_, _22897_, _23011_);
  and g_33358_(_22903_, _22932_, _23012_);
  or g_33359_(_22904_, _22931_, _23013_);
  and g_33360_(_22923_, _23012_, _23014_);
  or g_33361_(_22922_, _23013_, _23015_);
  and g_33362_(_23011_, _23015_, _23016_);
  or g_33363_(_23010_, _23014_, _23018_);
  and g_33364_(_23009_, _23016_, _23019_);
  or g_33365_(_23008_, _23018_, _23020_);
  and g_33366_(_22988_, _23020_, _23021_);
  or g_33367_(_22987_, _23019_, _23022_);
  and g_33368_(_22818_, _23022_, _23023_);
  or g_33369_(_22817_, _23021_, _23024_);
  and g_33370_(_22883_, _23021_, _23025_);
  or g_33371_(_22884_, _23022_, _23026_);
  and g_33372_(_23024_, _23026_, _23027_);
  or g_33373_(_23023_, _23025_, _23029_);
  and g_33374_(_22888_, _22890_, _23030_);
  or g_33375_(_22889_, _22891_, _23031_);
  or g_33376_(out[227], _19229_, _23032_);
  not g_33377_(_23032_, _23033_);
  and g_33378_(out[228], _23032_, _23034_);
  or g_33379_(_19134_, _23033_, _23035_);
  and g_33380_(out[229], _23034_, _23036_);
  and g_33381_(out[230], _23036_, _23037_);
  or g_33382_(out[231], _23037_, _23038_);
  and g_33383_(out[232], _23038_, _23040_);
  or g_33384_(out[233], _23040_, _23041_);
  not g_33385_(_23041_, _23042_);
  or g_33386_(out[234], _23041_, _23043_);
  xor g_33387_(out[235], _23043_, _23044_);
  xor g_33388_(_19090_, _23043_, _23045_);
  and g_33389_(_23030_, _23045_, _23046_);
  or g_33390_(_23031_, _23044_, _23047_);
  xor g_33391_(out[234], _23041_, _23048_);
  xor g_33392_(_19211_, _23041_, _23049_);
  and g_33393_(_23027_, _23048_, _23051_);
  or g_33394_(_23029_, _23049_, _23052_);
  and g_33395_(_23047_, _23052_, _23053_);
  or g_33396_(_23046_, _23051_, _23054_);
  and g_33397_(_23031_, _23044_, _23055_);
  or g_33398_(_23030_, _23045_, _23056_);
  and g_33399_(_23029_, _23049_, _23057_);
  or g_33400_(_23027_, _23048_, _23058_);
  and g_33401_(_23056_, _23058_, _23059_);
  or g_33402_(_23055_, _23057_, _23060_);
  or g_33403_(_22916_, _23021_, _23062_);
  not g_33404_(_23062_, _23063_);
  and g_33405_(_22921_, _23021_, _23064_);
  not g_33406_(_23064_, _23065_);
  and g_33407_(_23062_, _23065_, _23066_);
  or g_33408_(_23063_, _23064_, _23067_);
  and g_33409_(out[233], _23040_, _23068_);
  xor g_33410_(out[233], _23040_, _23069_);
  or g_33411_(_23042_, _23068_, _23070_);
  and g_33412_(_23066_, _23070_, _23071_);
  or g_33413_(_23067_, _23069_, _23073_);
  and g_33414_(_23059_, _23073_, _23074_);
  or g_33415_(_23060_, _23071_, _23075_);
  and g_33416_(_23053_, _23074_, _23076_);
  or g_33417_(_23054_, _23075_, _23077_);
  xor g_33418_(out[232], _23038_, _23078_);
  xor g_33419_(_19189_, _23038_, _23079_);
  or g_33420_(_22910_, _23021_, _23080_);
  not g_33421_(_23080_, _23081_);
  and g_33422_(_22906_, _23021_, _23082_);
  not g_33423_(_23082_, _23084_);
  and g_33424_(_23080_, _23084_, _23085_);
  or g_33425_(_23081_, _23082_, _23086_);
  or g_33426_(_23079_, _23085_, _23087_);
  not g_33427_(_23087_, _23088_);
  and g_33428_(_23067_, _23069_, _23089_);
  or g_33429_(_23066_, _23070_, _23090_);
  and g_33430_(_23079_, _23085_, _23091_);
  or g_33431_(_23078_, _23086_, _23092_);
  and g_33432_(_23090_, _23092_, _23093_);
  or g_33433_(_23089_, _23091_, _23095_);
  and g_33434_(_23087_, _23093_, _23096_);
  or g_33435_(_23088_, _23095_, _23097_);
  and g_33436_(_23076_, _23096_, _23098_);
  or g_33437_(_23077_, _23097_, _23099_);
  xor g_33438_(out[231], _23037_, _23100_);
  xor g_33439_(_19101_, _23037_, _23101_);
  or g_33440_(_22843_, _23022_, _23102_);
  or g_33441_(_22846_, _23021_, _23103_);
  and g_33442_(_23102_, _23103_, _23104_);
  or g_33443_(_23100_, _23104_, _23106_);
  xor g_33444_(out[230], _23036_, _23107_);
  xor g_33445_(_19112_, _23036_, _23108_);
  or g_33446_(_22826_, _23022_, _23109_);
  or g_33447_(_22831_, _23021_, _23110_);
  and g_33448_(_23109_, _23110_, _23111_);
  and g_33449_(_23108_, _23111_, _23112_);
  and g_33450_(_23100_, _23104_, _23113_);
  xor g_33451_(_23100_, _23104_, _23114_);
  xor g_33452_(_23101_, _23104_, _23115_);
  xor g_33453_(_23108_, _23111_, _23117_);
  xor g_33454_(_23107_, _23111_, _23118_);
  and g_33455_(_23114_, _23117_, _23119_);
  or g_33456_(_23115_, _23118_, _23120_);
  or g_33457_(_19082_, _19229_, _23121_);
  not g_33458_(_23121_, _23122_);
  and g_33459_(_23035_, _23121_, _23123_);
  or g_33460_(_23034_, _23122_, _23124_);
  or g_33461_(_22865_, _23021_, _23125_);
  or g_33462_(_22860_, _23022_, _23126_);
  and g_33463_(_23125_, _23126_, _23128_);
  and g_33464_(_23124_, _23128_, _23129_);
  not g_33465_(_23129_, _23130_);
  xor g_33466_(out[229], _23034_, _23131_);
  xor g_33467_(_19123_, _23034_, _23132_);
  or g_33468_(_22833_, _23022_, _23133_);
  or g_33469_(_22837_, _23021_, _23134_);
  and g_33470_(_23133_, _23134_, _23135_);
  not g_33471_(_23135_, _23136_);
  and g_33472_(_23132_, _23135_, _23137_);
  or g_33473_(_23131_, _23136_, _23139_);
  and g_33474_(_23130_, _23139_, _23140_);
  or g_33475_(_23129_, _23137_, _23141_);
  or g_33476_(_23132_, _23135_, _23142_);
  or g_33477_(_23124_, _23128_, _23143_);
  and g_33478_(_23142_, _23143_, _23144_);
  not g_33479_(_23144_, _23145_);
  and g_33480_(_23140_, _23144_, _23146_);
  or g_33481_(_23141_, _23145_, _23147_);
  and g_33482_(_23119_, _23146_, _23148_);
  or g_33483_(_23120_, _23147_, _23150_);
  and g_33484_(_23098_, _23148_, _23151_);
  or g_33485_(_23099_, _23150_, _23152_);
  xor g_33486_(out[227], _19229_, _23153_);
  xor g_33487_(_19178_, _19229_, _23154_);
  or g_33488_(_22964_, _23022_, _23155_);
  or g_33489_(_22967_, _23021_, _23156_);
  and g_33490_(_23155_, _23156_, _23157_);
  and g_33491_(_23153_, _23157_, _23158_);
  or g_33492_(_22958_, _23021_, _23159_);
  or g_33493_(_18851_, _23022_, _23161_);
  and g_33494_(_23159_, _23161_, _23162_);
  or g_33495_(_23153_, _23157_, _23163_);
  and g_33496_(_19230_, _23162_, _23164_);
  xor g_33497_(_23153_, _23157_, _23165_);
  xor g_33498_(_23154_, _23157_, _23166_);
  xor g_33499_(_19230_, _23162_, _23167_);
  xor g_33500_(_19231_, _23162_, _23168_);
  and g_33501_(_23165_, _23167_, _23169_);
  or g_33502_(_23166_, _23168_, _23170_);
  or g_33503_(_19013_, _23022_, _23172_);
  or g_33504_(_22939_, _23021_, _23173_);
  and g_33505_(_23172_, _23173_, _23174_);
  and g_33506_(out[225], _23174_, _23175_);
  not g_33507_(_23175_, _23176_);
  or g_33508_(_19024_, _23022_, _23177_);
  or g_33509_(_22945_, _23021_, _23178_);
  and g_33510_(_23177_, _23178_, _23179_);
  and g_33511_(out[224], _23179_, _23180_);
  not g_33512_(_23180_, _23181_);
  xor g_33513_(out[225], _23174_, _23183_);
  xor g_33514_(_19145_, _23174_, _23184_);
  and g_33515_(_23181_, _23183_, _23185_);
  or g_33516_(_23180_, _23184_, _23186_);
  and g_33517_(_23176_, _23186_, _23187_);
  or g_33518_(_23175_, _23185_, _23188_);
  and g_33519_(_23169_, _23188_, _23189_);
  or g_33520_(_23170_, _23187_, _23190_);
  and g_33521_(_23163_, _23164_, _23191_);
  or g_33522_(_23158_, _23191_, _23192_);
  not g_33523_(_23192_, _23194_);
  and g_33524_(_23190_, _23194_, _23195_);
  or g_33525_(_23189_, _23192_, _23196_);
  and g_33526_(_23151_, _23196_, _23197_);
  or g_33527_(_23152_, _23195_, _23198_);
  and g_33528_(_23119_, _23141_, _23199_);
  and g_33529_(_23142_, _23199_, _23200_);
  and g_33530_(_23106_, _23112_, _23201_);
  or g_33531_(_23113_, _23201_, _23202_);
  or g_33532_(_23200_, _23202_, _23203_);
  not g_33533_(_23203_, _23205_);
  and g_33534_(_23098_, _23203_, _23206_);
  or g_33535_(_23099_, _23205_, _23207_);
  or g_33536_(_23077_, _23093_, _23208_);
  not g_33537_(_23208_, _23209_);
  and g_33538_(_23054_, _23056_, _23210_);
  or g_33539_(_23053_, _23055_, _23211_);
  and g_33540_(_23208_, _23211_, _23212_);
  or g_33541_(_23209_, _23210_, _23213_);
  and g_33542_(_23207_, _23212_, _23214_);
  or g_33543_(_23206_, _23213_, _23216_);
  and g_33544_(_23198_, _23214_, _23217_);
  or g_33545_(_23197_, _23216_, _23218_);
  or g_33546_(out[224], _23179_, _23219_);
  and g_33547_(_23169_, _23219_, _23220_);
  not g_33548_(_23220_, _23221_);
  and g_33549_(_23185_, _23220_, _23222_);
  or g_33550_(_23186_, _23221_, _23223_);
  and g_33551_(_23151_, _23222_, _23224_);
  or g_33552_(_23152_, _23223_, _23225_);
  and g_33553_(_23218_, _23225_, _23227_);
  or g_33554_(_23217_, _23224_, _23228_);
  and g_33555_(_23029_, _23228_, _23229_);
  or g_33556_(_23027_, _23227_, _23230_);
  and g_33557_(_23048_, _23227_, _23231_);
  or g_33558_(_23049_, _23228_, _23232_);
  and g_33559_(_23230_, _23232_, _23233_);
  or g_33560_(_23229_, _23231_, _23234_);
  or g_33561_(out[243], _19441_, _23235_);
  not g_33562_(_23235_, _23236_);
  and g_33563_(out[244], _23235_, _23238_);
  or g_33564_(_19266_, _23236_, _23239_);
  and g_33565_(out[245], _23238_, _23240_);
  and g_33566_(out[246], _23240_, _23241_);
  or g_33567_(out[247], _23241_, _23242_);
  and g_33568_(out[248], _23242_, _23243_);
  or g_33569_(out[249], _23243_, _23244_);
  not g_33570_(_23244_, _23245_);
  or g_33571_(out[250], _23244_, _23246_);
  xor g_33572_(out[250], _23244_, _23247_);
  xor g_33573_(_19343_, _23244_, _23249_);
  and g_33574_(_23233_, _23247_, _23250_);
  or g_33575_(_23234_, _23249_, _23251_);
  and g_33576_(_23030_, _23044_, _23252_);
  or g_33577_(_23031_, _23045_, _23253_);
  xor g_33578_(out[251], _23246_, _23254_);
  xor g_33579_(_19222_, _23246_, _23255_);
  and g_33580_(_23252_, _23255_, _23256_);
  or g_33581_(_23253_, _23254_, _23257_);
  and g_33582_(_23251_, _23257_, _23258_);
  or g_33583_(_23250_, _23256_, _23260_);
  and g_33584_(_23253_, _23254_, _23261_);
  or g_33585_(_23252_, _23255_, _23262_);
  and g_33586_(_23234_, _23249_, _23263_);
  or g_33587_(_23233_, _23247_, _23264_);
  and g_33588_(_23262_, _23264_, _23265_);
  or g_33589_(_23261_, _23263_, _23266_);
  and g_33590_(_23258_, _23265_, _23267_);
  or g_33591_(_23260_, _23266_, _23268_);
  xor g_33592_(out[248], _23242_, _23269_);
  xor g_33593_(_19321_, _23242_, _23271_);
  and g_33594_(_23079_, _23227_, _23272_);
  not g_33595_(_23272_, _23273_);
  or g_33596_(_23085_, _23227_, _23274_);
  not g_33597_(_23274_, _23275_);
  and g_33598_(_23273_, _23274_, _23276_);
  or g_33599_(_23272_, _23275_, _23277_);
  and g_33600_(_23269_, _23277_, _23278_);
  or g_33601_(_23271_, _23276_, _23279_);
  and g_33602_(out[249], _23243_, _23280_);
  xor g_33603_(out[249], _23243_, _23282_);
  or g_33604_(_23245_, _23280_, _23283_);
  or g_33605_(_23066_, _23227_, _23284_);
  not g_33606_(_23284_, _23285_);
  and g_33607_(_23070_, _23227_, _23286_);
  not g_33608_(_23286_, _23287_);
  and g_33609_(_23284_, _23287_, _23288_);
  or g_33610_(_23285_, _23286_, _23289_);
  and g_33611_(_23283_, _23288_, _23290_);
  or g_33612_(_23282_, _23289_, _23291_);
  and g_33613_(_23279_, _23291_, _23293_);
  or g_33614_(_23278_, _23290_, _23294_);
  and g_33615_(_23282_, _23289_, _23295_);
  or g_33616_(_23283_, _23288_, _23296_);
  and g_33617_(_23271_, _23276_, _23297_);
  or g_33618_(_23269_, _23277_, _23298_);
  and g_33619_(_23296_, _23298_, _23299_);
  or g_33620_(_23295_, _23297_, _23300_);
  and g_33621_(_23293_, _23299_, _23301_);
  or g_33622_(_23294_, _23300_, _23302_);
  and g_33623_(_23267_, _23301_, _23304_);
  or g_33624_(_23268_, _23302_, _23305_);
  xor g_33625_(out[246], _23240_, _23306_);
  xor g_33626_(_19244_, _23240_, _23307_);
  or g_33627_(_23107_, _23228_, _23308_);
  or g_33628_(_23111_, _23227_, _23309_);
  and g_33629_(_23308_, _23309_, _23310_);
  not g_33630_(_23310_, _23311_);
  and g_33631_(_23307_, _23310_, _23312_);
  or g_33632_(_23306_, _23311_, _23313_);
  xor g_33633_(out[247], _23241_, _23315_);
  xor g_33634_(_19233_, _23241_, _23316_);
  and g_33635_(_23100_, _23227_, _23317_);
  not g_33636_(_23317_, _23318_);
  or g_33637_(_23104_, _23227_, _23319_);
  not g_33638_(_23319_, _23320_);
  and g_33639_(_23318_, _23319_, _23321_);
  or g_33640_(_23317_, _23320_, _23322_);
  and g_33641_(_23315_, _23321_, _23323_);
  or g_33642_(_23316_, _23322_, _23324_);
  and g_33643_(_23313_, _23324_, _23326_);
  or g_33644_(_23312_, _23323_, _23327_);
  and g_33645_(_23306_, _23311_, _23328_);
  or g_33646_(_23307_, _23310_, _23329_);
  and g_33647_(_23316_, _23322_, _23330_);
  or g_33648_(_23315_, _23321_, _23331_);
  xor g_33649_(out[245], _23238_, _23332_);
  xor g_33650_(_19255_, _23238_, _23333_);
  and g_33651_(_23132_, _23227_, _23334_);
  not g_33652_(_23334_, _23335_);
  or g_33653_(_23135_, _23227_, _23337_);
  not g_33654_(_23337_, _23338_);
  and g_33655_(_23335_, _23337_, _23339_);
  or g_33656_(_23334_, _23338_, _23340_);
  and g_33657_(_23332_, _23340_, _23341_);
  or g_33658_(_23333_, _23339_, _23342_);
  and g_33659_(_23331_, _23342_, _23343_);
  or g_33660_(_23330_, _23341_, _23344_);
  and g_33661_(_23329_, _23343_, _23345_);
  or g_33662_(_23328_, _23344_, _23346_);
  and g_33663_(_23326_, _23345_, _23348_);
  or g_33664_(_23327_, _23346_, _23349_);
  and g_33665_(_23304_, _23348_, _23350_);
  or g_33666_(_23305_, _23349_, _23351_);
  or g_33667_(_19318_, _19441_, _23352_);
  not g_33668_(_23352_, _23353_);
  and g_33669_(_23239_, _23352_, _23354_);
  or g_33670_(_23238_, _23353_, _23355_);
  or g_33671_(_23128_, _23227_, _23356_);
  not g_33672_(_23356_, _23357_);
  and g_33673_(_23124_, _23227_, _23359_);
  not g_33674_(_23359_, _23360_);
  and g_33675_(_23356_, _23360_, _23361_);
  or g_33676_(_23357_, _23359_, _23362_);
  and g_33677_(_23355_, _23361_, _23363_);
  or g_33678_(_23354_, _23362_, _23364_);
  and g_33679_(_23333_, _23339_, _23365_);
  or g_33680_(_23332_, _23340_, _23366_);
  and g_33681_(_23364_, _23366_, _23367_);
  or g_33682_(_23363_, _23365_, _23368_);
  and g_33683_(_23354_, _23362_, _23370_);
  or g_33684_(_23355_, _23361_, _23371_);
  and g_33685_(_23367_, _23371_, _23372_);
  or g_33686_(_23368_, _23370_, _23373_);
  and g_33687_(_23350_, _23372_, _23374_);
  or g_33688_(_23351_, _23373_, _23375_);
  xor g_33689_(out[243], _19441_, _23376_);
  xor g_33690_(_19310_, _19441_, _23377_);
  and g_33691_(_23154_, _23227_, _23378_);
  and g_33692_(_23157_, _23228_, _23379_);
  or g_33693_(_23378_, _23379_, _23381_);
  and g_33694_(_23376_, _23381_, _23382_);
  and g_33695_(_19231_, _23227_, _23383_);
  and g_33696_(_23162_, _23228_, _23384_);
  or g_33697_(_23383_, _23384_, _23385_);
  and g_33698_(_19443_, _23385_, _23386_);
  or g_33699_(_23382_, _23386_, _23387_);
  or g_33700_(_23376_, _23381_, _23388_);
  xor g_33701_(_23376_, _23381_, _23389_);
  xor g_33702_(_23377_, _23381_, _23390_);
  xor g_33703_(_19443_, _23385_, _23392_);
  xor g_33704_(_19444_, _23385_, _23393_);
  and g_33705_(_23389_, _23392_, _23394_);
  or g_33706_(_23390_, _23393_, _23395_);
  and g_33707_(out[224], _23227_, _23396_);
  not g_33708_(_23396_, _23397_);
  or g_33709_(_23179_, _23227_, _23398_);
  not g_33710_(_23398_, _23399_);
  and g_33711_(_23397_, _23398_, _23400_);
  or g_33712_(_23396_, _23399_, _23401_);
  and g_33713_(out[240], _23400_, _23403_);
  or g_33714_(_19288_, _23401_, _23404_);
  or g_33715_(_19145_, _23228_, _23405_);
  or g_33716_(_23174_, _23227_, _23406_);
  and g_33717_(_23405_, _23406_, _23407_);
  and g_33718_(out[241], _23407_, _23408_);
  xor g_33719_(out[241], _23407_, _23409_);
  xor g_33720_(_19277_, _23407_, _23410_);
  and g_33721_(_23404_, _23409_, _23411_);
  or g_33722_(_23403_, _23410_, _23412_);
  and g_33723_(_23394_, _23411_, _23414_);
  or g_33724_(_23395_, _23412_, _23415_);
  and g_33725_(_19288_, _23401_, _23416_);
  or g_33726_(out[240], _23400_, _23417_);
  and g_33727_(_23414_, _23417_, _23418_);
  or g_33728_(_23415_, _23416_, _23419_);
  and g_33729_(_23374_, _23418_, _23420_);
  or g_33730_(_23375_, _23419_, _23421_);
  and g_33731_(_23394_, _23408_, _23422_);
  and g_33732_(_23387_, _23388_, _23423_);
  or g_33733_(_23422_, _23423_, _23425_);
  not g_33734_(_23425_, _23426_);
  and g_33735_(_23415_, _23426_, _23427_);
  or g_33736_(_23414_, _23425_, _23428_);
  and g_33737_(_23374_, _23428_, _23429_);
  or g_33738_(_23375_, _23427_, _23430_);
  and g_33739_(_23350_, _23368_, _23431_);
  or g_33740_(_23351_, _23367_, _23432_);
  and g_33741_(_23327_, _23331_, _23433_);
  or g_33742_(_23326_, _23330_, _23434_);
  and g_33743_(_23304_, _23433_, _23436_);
  or g_33744_(_23305_, _23434_, _23437_);
  and g_33745_(_23291_, _23300_, _23438_);
  or g_33746_(_23290_, _23299_, _23439_);
  and g_33747_(_23267_, _23438_, _23440_);
  or g_33748_(_23268_, _23439_, _23441_);
  and g_33749_(_23260_, _23262_, _23442_);
  or g_33750_(_23258_, _23261_, _23443_);
  and g_33751_(_23441_, _23443_, _23444_);
  or g_33752_(_23440_, _23442_, _23445_);
  and g_33753_(_23437_, _23444_, _23447_);
  or g_33754_(_23436_, _23445_, _23448_);
  and g_33755_(_23432_, _23447_, _23449_);
  or g_33756_(_23431_, _23448_, _23450_);
  and g_33757_(_23430_, _23449_, _23451_);
  or g_33758_(_23429_, _23450_, _23452_);
  and g_33759_(_23421_, _23452_, _23453_);
  or g_33760_(_23420_, _23451_, _23454_);
  or g_33761_(_23233_, _23453_, _23455_);
  or g_33762_(_23249_, _23454_, _23456_);
  and g_33763_(_23455_, _23456_, _23458_);
  not g_33764_(_23458_, _23459_);
  or g_33765_(out[259], _19672_, _23460_);
  not g_33766_(_23460_, _23461_);
  and g_33767_(out[260], _23460_, _23462_);
  or g_33768_(_19398_, _23461_, _23463_);
  or g_33769_(_19528_, _19672_, _23464_);
  not g_33770_(_23464_, _23465_);
  and g_33771_(_23463_, _23464_, _23466_);
  or g_33772_(_23462_, _23465_, _23467_);
  or g_33773_(_23361_, _23453_, _23469_);
  or g_33774_(_23354_, _23454_, _23470_);
  and g_33775_(_23469_, _23470_, _23471_);
  not g_33776_(_23471_, _23472_);
  and g_33777_(_23467_, _23471_, _23473_);
  not g_33778_(_23473_, _23474_);
  and g_33779_(out[261], _23462_, _23475_);
  xor g_33780_(out[261], _23462_, _23476_);
  xor g_33781_(_19387_, _23462_, _23477_);
  or g_33782_(_23332_, _23454_, _23478_);
  or g_33783_(_23339_, _23453_, _23480_);
  and g_33784_(_23478_, _23480_, _23481_);
  and g_33785_(_23477_, _23481_, _23482_);
  not g_33786_(_23482_, _23483_);
  and g_33787_(_23474_, _23483_, _23484_);
  or g_33788_(_23473_, _23482_, _23485_);
  and g_33789_(_23466_, _23472_, _23486_);
  or g_33790_(_23467_, _23471_, _23487_);
  or g_33791_(_23385_, _23453_, _23488_);
  or g_33792_(_19444_, _23454_, _23489_);
  and g_33793_(_23488_, _23489_, _23491_);
  xor g_33794_(out[259], _19672_, _23492_);
  xor g_33795_(_19442_, _19672_, _23493_);
  or g_33796_(_23377_, _23454_, _23494_);
  or g_33797_(_23381_, _23453_, _23495_);
  and g_33798_(_23494_, _23495_, _23496_);
  and g_33799_(_23492_, _23496_, _23497_);
  and g_33800_(_19674_, _23491_, _23498_);
  or g_33801_(_23492_, _23496_, _23499_);
  xor g_33802_(_19674_, _23491_, _23500_);
  xor g_33803_(_19675_, _23491_, _23502_);
  xor g_33804_(_23492_, _23496_, _23503_);
  xor g_33805_(_23493_, _23496_, _23504_);
  and g_33806_(_23500_, _23503_, _23505_);
  or g_33807_(_23502_, _23504_, _23506_);
  or g_33808_(_19277_, _23454_, _23507_);
  or g_33809_(_23407_, _23453_, _23508_);
  and g_33810_(_23507_, _23508_, _23509_);
  and g_33811_(out[257], _23509_, _23510_);
  not g_33812_(_23510_, _23511_);
  and g_33813_(out[240], _23453_, _23513_);
  or g_33814_(_19288_, _23454_, _23514_);
  and g_33815_(_23401_, _23454_, _23515_);
  or g_33816_(_23400_, _23453_, _23516_);
  and g_33817_(_23514_, _23516_, _23517_);
  or g_33818_(_23513_, _23515_, _23518_);
  and g_33819_(out[256], _23517_, _23519_);
  or g_33820_(_19420_, _23518_, _23520_);
  xor g_33821_(out[257], _23509_, _23521_);
  xor g_33822_(_19409_, _23509_, _23522_);
  and g_33823_(_23520_, _23521_, _23524_);
  or g_33824_(_23519_, _23522_, _23525_);
  and g_33825_(_23511_, _23525_, _23526_);
  or g_33826_(_23510_, _23524_, _23527_);
  and g_33827_(_23505_, _23527_, _23528_);
  or g_33828_(_23506_, _23526_, _23529_);
  or g_33829_(_23497_, _23498_, _23530_);
  and g_33830_(_23499_, _23530_, _23531_);
  not g_33831_(_23531_, _23532_);
  and g_33832_(_23529_, _23532_, _23533_);
  or g_33833_(_23528_, _23531_, _23535_);
  and g_33834_(_23487_, _23535_, _23536_);
  or g_33835_(_23486_, _23533_, _23537_);
  and g_33836_(_23484_, _23537_, _23538_);
  or g_33837_(_23485_, _23536_, _23539_);
  and g_33838_(out[262], _23475_, _23540_);
  or g_33839_(out[263], _23540_, _23541_);
  and g_33840_(out[264], _23541_, _23542_);
  or g_33841_(out[265], _23542_, _23543_);
  or g_33842_(out[266], _23543_, _23544_);
  xor g_33843_(out[266], _23543_, _23546_);
  and g_33844_(_23458_, _23546_, _23547_);
  and g_33845_(_23252_, _23254_, _23548_);
  or g_33846_(_23253_, _23255_, _23549_);
  xor g_33847_(out[267], _23544_, _23550_);
  xor g_33848_(_19354_, _23544_, _23551_);
  and g_33849_(_23548_, _23551_, _23552_);
  or g_33850_(_23548_, _23551_, _23553_);
  xor g_33851_(_23549_, _23550_, _23554_);
  xor g_33852_(_23548_, _23550_, _23555_);
  xor g_33853_(_23458_, _23546_, _23557_);
  xor g_33854_(_23459_, _23546_, _23558_);
  and g_33855_(_23554_, _23557_, _23559_);
  or g_33856_(_23555_, _23558_, _23560_);
  or g_33857_(_23288_, _23453_, _23561_);
  or g_33858_(_23282_, _23454_, _23562_);
  and g_33859_(_23561_, _23562_, _23563_);
  not g_33860_(_23563_, _23564_);
  and g_33861_(out[265], _23542_, _23565_);
  xor g_33862_(out[265], _23542_, _23566_);
  xor g_33863_(_19464_, _23542_, _23568_);
  or g_33864_(_23563_, _23568_, _23569_);
  not g_33865_(_23569_, _23570_);
  xor g_33866_(out[264], _23541_, _23571_);
  xor g_33867_(_19453_, _23541_, _23572_);
  or g_33868_(_23269_, _23454_, _23573_);
  or g_33869_(_23276_, _23453_, _23574_);
  and g_33870_(_23573_, _23574_, _23575_);
  not g_33871_(_23575_, _23576_);
  and g_33872_(_23572_, _23575_, _23577_);
  or g_33873_(_23570_, _23577_, _23579_);
  and g_33874_(_23563_, _23568_, _23580_);
  or g_33875_(_23564_, _23566_, _23581_);
  and g_33876_(_23571_, _23576_, _23582_);
  or g_33877_(_23580_, _23582_, _23583_);
  or g_33878_(_23579_, _23583_, _23584_);
  xor g_33879_(_23572_, _23575_, _23585_);
  and g_33880_(_23569_, _23581_, _23586_);
  and g_33881_(_23559_, _23586_, _23587_);
  and g_33882_(_23585_, _23587_, _23588_);
  or g_33883_(_23560_, _23584_, _23590_);
  or g_33884_(_23477_, _23481_, _23591_);
  not g_33885_(_23591_, _23592_);
  xor g_33886_(out[262], _23475_, _23593_);
  not g_33887_(_23593_, _23594_);
  or g_33888_(_23306_, _23454_, _23595_);
  or g_33889_(_23310_, _23453_, _23596_);
  and g_33890_(_23595_, _23596_, _23597_);
  xor g_33891_(out[263], _23540_, _23598_);
  xor g_33892_(_19365_, _23540_, _23599_);
  and g_33893_(_23315_, _23453_, _23601_);
  not g_33894_(_23601_, _23602_);
  and g_33895_(_23322_, _23454_, _23603_);
  or g_33896_(_23321_, _23453_, _23604_);
  and g_33897_(_23602_, _23604_, _23605_);
  or g_33898_(_23601_, _23603_, _23606_);
  and g_33899_(_23598_, _23605_, _23607_);
  or g_33900_(_23598_, _23605_, _23608_);
  and g_33901_(_23594_, _23597_, _23609_);
  xor g_33902_(_23599_, _23606_, _23610_);
  xor g_33903_(_23598_, _23606_, _23612_);
  xor g_33904_(_23594_, _23597_, _23613_);
  xor g_33905_(_23593_, _23597_, _23614_);
  and g_33906_(_23591_, _23613_, _23615_);
  or g_33907_(_23592_, _23614_, _23616_);
  and g_33908_(_23588_, _23615_, _23617_);
  or g_33909_(_23590_, _23616_, _23618_);
  and g_33910_(_23610_, _23617_, _23619_);
  or g_33911_(_23612_, _23618_, _23620_);
  and g_33912_(_23539_, _23619_, _23621_);
  or g_33913_(_23538_, _23620_, _23623_);
  and g_33914_(_23608_, _23609_, _23624_);
  or g_33915_(_23607_, _23624_, _23625_);
  and g_33916_(_23588_, _23625_, _23626_);
  and g_33917_(_23559_, _23579_, _23627_);
  and g_33918_(_23581_, _23627_, _23628_);
  and g_33919_(_23547_, _23553_, _23629_);
  or g_33920_(_23552_, _23629_, _23630_);
  or g_33921_(_23628_, _23630_, _23631_);
  or g_33922_(_23626_, _23631_, _23632_);
  not g_33923_(_23632_, _23634_);
  and g_33924_(_23623_, _23634_, _23635_);
  or g_33925_(_23621_, _23632_, _23636_);
  or g_33926_(out[256], _23517_, _23637_);
  and g_33927_(_23487_, _23637_, _23638_);
  and g_33928_(_23505_, _23638_, _23639_);
  and g_33929_(_23484_, _23639_, _23640_);
  and g_33930_(_23524_, _23640_, _23641_);
  and g_33931_(_23619_, _23641_, _23642_);
  not g_33932_(_23642_, _23643_);
  and g_33933_(_23636_, _23643_, _23645_);
  or g_33934_(_23635_, _23642_, _23646_);
  or g_33935_(_23458_, _23645_, _23647_);
  not g_33936_(_23647_, _23648_);
  and g_33937_(_23546_, _23645_, _23649_);
  not g_33938_(_23649_, _23650_);
  and g_33939_(_23647_, _23650_, _23651_);
  or g_33940_(_23648_, _23649_, _23652_);
  or g_33941_(out[275], _19885_, _23653_);
  not g_33942_(_23653_, _23654_);
  and g_33943_(out[276], _23653_, _23656_);
  or g_33944_(_19530_, _23654_, _23657_);
  and g_33945_(out[277], _23656_, _23658_);
  and g_33946_(out[278], _23658_, _23659_);
  or g_33947_(out[279], _23659_, _23660_);
  and g_33948_(out[280], _23660_, _23661_);
  or g_33949_(out[281], _23661_, _23662_);
  not g_33950_(_23662_, _23663_);
  or g_33951_(out[282], _23662_, _23664_);
  xor g_33952_(out[282], _23662_, _23665_);
  xor g_33953_(_19607_, _23662_, _23667_);
  and g_33954_(_23651_, _23665_, _23668_);
  or g_33955_(_23652_, _23667_, _23669_);
  and g_33956_(_23548_, _23550_, _23670_);
  or g_33957_(_23549_, _23551_, _23671_);
  xor g_33958_(out[283], _23664_, _23672_);
  xor g_33959_(_19486_, _23664_, _23673_);
  and g_33960_(_23670_, _23673_, _23674_);
  or g_33961_(_23671_, _23672_, _23675_);
  and g_33962_(_23669_, _23675_, _23676_);
  or g_33963_(_23668_, _23674_, _23678_);
  and g_33964_(_23652_, _23667_, _23679_);
  or g_33965_(_23651_, _23665_, _23680_);
  and g_33966_(_23671_, _23672_, _23681_);
  or g_33967_(_23670_, _23673_, _23682_);
  or g_33968_(_23563_, _23645_, _23683_);
  not g_33969_(_23683_, _23684_);
  and g_33970_(_23568_, _23645_, _23685_);
  not g_33971_(_23685_, _23686_);
  and g_33972_(_23683_, _23686_, _23687_);
  or g_33973_(_23684_, _23685_, _23689_);
  and g_33974_(out[281], _23661_, _23690_);
  xor g_33975_(out[281], _23661_, _23691_);
  or g_33976_(_23663_, _23690_, _23692_);
  and g_33977_(_23687_, _23692_, _23693_);
  or g_33978_(_23689_, _23691_, _23694_);
  and g_33979_(_23682_, _23694_, _23695_);
  or g_33980_(_23681_, _23693_, _23696_);
  and g_33981_(_23680_, _23695_, _23697_);
  or g_33982_(_23679_, _23696_, _23698_);
  and g_33983_(_23676_, _23697_, _23700_);
  or g_33984_(_23678_, _23698_, _23701_);
  xor g_33985_(out[280], _23660_, _23702_);
  xor g_33986_(_19585_, _23660_, _23703_);
  and g_33987_(_23572_, _23645_, _23704_);
  not g_33988_(_23704_, _23705_);
  or g_33989_(_23575_, _23645_, _23706_);
  not g_33990_(_23706_, _23707_);
  and g_33991_(_23705_, _23706_, _23708_);
  or g_33992_(_23704_, _23707_, _23709_);
  and g_33993_(_23702_, _23709_, _23711_);
  or g_33994_(_23703_, _23708_, _23712_);
  and g_33995_(_23689_, _23691_, _23713_);
  or g_33996_(_23687_, _23692_, _23714_);
  and g_33997_(_23703_, _23708_, _23715_);
  or g_33998_(_23702_, _23709_, _23716_);
  and g_33999_(_23714_, _23716_, _23717_);
  or g_34000_(_23713_, _23715_, _23718_);
  and g_34001_(_23712_, _23717_, _23719_);
  or g_34002_(_23711_, _23718_, _23720_);
  and g_34003_(_23700_, _23719_, _23722_);
  or g_34004_(_23701_, _23720_, _23723_);
  and g_34005_(_23594_, _23645_, _23724_);
  or g_34006_(_23597_, _23645_, _23725_);
  not g_34007_(_23725_, _23726_);
  or g_34008_(_23724_, _23726_, _23727_);
  xor g_34009_(out[278], _23658_, _23728_);
  not g_34010_(_23728_, _23729_);
  or g_34011_(_23727_, _23728_, _23730_);
  xor g_34012_(out[279], _23659_, _23731_);
  xor g_34013_(_19497_, _23659_, _23733_);
  and g_34014_(_23598_, _23645_, _23734_);
  and g_34015_(_23606_, _23646_, _23735_);
  or g_34016_(_23734_, _23735_, _23736_);
  and g_34017_(_23733_, _23736_, _23737_);
  or g_34018_(_23733_, _23736_, _23738_);
  xor g_34019_(_23733_, _23736_, _23739_);
  xor g_34020_(_23731_, _23736_, _23740_);
  xor g_34021_(_23727_, _23728_, _23741_);
  xor g_34022_(_23727_, _23729_, _23742_);
  and g_34023_(_23739_, _23741_, _23744_);
  or g_34024_(_23740_, _23742_, _23745_);
  or g_34025_(_19748_, _19885_, _23746_);
  not g_34026_(_23746_, _23747_);
  and g_34027_(_23657_, _23746_, _23748_);
  or g_34028_(_23656_, _23747_, _23749_);
  or g_34029_(_23471_, _23645_, _23750_);
  not g_34030_(_23750_, _23751_);
  and g_34031_(_23467_, _23645_, _23752_);
  not g_34032_(_23752_, _23753_);
  and g_34033_(_23750_, _23753_, _23755_);
  or g_34034_(_23751_, _23752_, _23756_);
  and g_34035_(_23749_, _23755_, _23757_);
  or g_34036_(_23748_, _23756_, _23758_);
  xor g_34037_(out[277], _23656_, _23759_);
  xor g_34038_(_19519_, _23656_, _23760_);
  and g_34039_(_23477_, _23645_, _23761_);
  not g_34040_(_23761_, _23762_);
  or g_34041_(_23481_, _23645_, _23763_);
  not g_34042_(_23763_, _23764_);
  and g_34043_(_23762_, _23763_, _23766_);
  or g_34044_(_23761_, _23764_, _23767_);
  and g_34045_(_23760_, _23766_, _23768_);
  or g_34046_(_23759_, _23767_, _23769_);
  and g_34047_(_23758_, _23769_, _23770_);
  or g_34048_(_23757_, _23768_, _23771_);
  and g_34049_(_23759_, _23767_, _23772_);
  or g_34050_(_23760_, _23766_, _23773_);
  and g_34051_(_23748_, _23756_, _23774_);
  or g_34052_(_23749_, _23755_, _23775_);
  and g_34053_(_23773_, _23775_, _23777_);
  or g_34054_(_23772_, _23774_, _23778_);
  and g_34055_(_23770_, _23777_, _23779_);
  or g_34056_(_23771_, _23778_, _23780_);
  and g_34057_(_23744_, _23779_, _23781_);
  or g_34058_(_23745_, _23780_, _23782_);
  and g_34059_(_23722_, _23781_, _23783_);
  or g_34060_(_23723_, _23782_, _23784_);
  xor g_34061_(out[275], _19885_, _23785_);
  xor g_34062_(_19574_, _19885_, _23786_);
  or g_34063_(_23496_, _23645_, _23788_);
  not g_34064_(_23788_, _23789_);
  and g_34065_(_23492_, _23645_, _23790_);
  not g_34066_(_23790_, _23791_);
  and g_34067_(_23788_, _23791_, _23792_);
  or g_34068_(_23789_, _23790_, _23793_);
  and g_34069_(_23785_, _23792_, _23794_);
  or g_34070_(_23491_, _23645_, _23795_);
  not g_34071_(_23795_, _23796_);
  and g_34072_(_19674_, _23645_, _23797_);
  not g_34073_(_23797_, _23799_);
  and g_34074_(_23795_, _23799_, _23800_);
  or g_34075_(_23796_, _23797_, _23801_);
  and g_34076_(_19886_, _23800_, _23802_);
  or g_34077_(_23794_, _23802_, _23803_);
  and g_34078_(_23786_, _23793_, _23804_);
  or g_34079_(_23785_, _23792_, _23805_);
  and g_34080_(_19887_, _23801_, _23806_);
  or g_34081_(_23804_, _23806_, _23807_);
  xor g_34082_(_23785_, _23792_, _23808_);
  xor g_34083_(_19886_, _23800_, _23810_);
  and g_34084_(_23808_, _23810_, _23811_);
  or g_34085_(_23803_, _23807_, _23812_);
  or g_34086_(_19409_, _23646_, _23813_);
  or g_34087_(_23509_, _23645_, _23814_);
  and g_34088_(_23813_, _23814_, _23815_);
  and g_34089_(out[273], _23815_, _23816_);
  and g_34090_(out[256], _23645_, _23817_);
  not g_34091_(_23817_, _23818_);
  or g_34092_(_23517_, _23645_, _23819_);
  not g_34093_(_23819_, _23821_);
  and g_34094_(_23818_, _23819_, _23822_);
  or g_34095_(_23817_, _23821_, _23823_);
  and g_34096_(out[272], _23822_, _23824_);
  or g_34097_(_19552_, _23823_, _23825_);
  xor g_34098_(out[273], _23815_, _23826_);
  xor g_34099_(_19541_, _23815_, _23827_);
  and g_34100_(_23825_, _23826_, _23828_);
  or g_34101_(_23824_, _23827_, _23829_);
  or g_34102_(_23816_, _23828_, _23830_);
  and g_34103_(_23811_, _23830_, _23832_);
  and g_34104_(_23803_, _23805_, _23833_);
  or g_34105_(_23832_, _23833_, _23834_);
  not g_34106_(_23834_, _23835_);
  and g_34107_(_23783_, _23834_, _23836_);
  or g_34108_(_23784_, _23835_, _23837_);
  and g_34109_(_23744_, _23771_, _23838_);
  or g_34110_(_23745_, _23770_, _23839_);
  and g_34111_(_23773_, _23838_, _23840_);
  or g_34112_(_23772_, _23839_, _23841_);
  or g_34113_(_23730_, _23737_, _23843_);
  and g_34114_(_23738_, _23843_, _23844_);
  not g_34115_(_23844_, _23845_);
  and g_34116_(_23841_, _23844_, _23846_);
  or g_34117_(_23840_, _23845_, _23847_);
  and g_34118_(_23722_, _23847_, _23848_);
  or g_34119_(_23723_, _23846_, _23849_);
  and g_34120_(_23700_, _23718_, _23850_);
  or g_34121_(_23701_, _23717_, _23851_);
  and g_34122_(_23678_, _23682_, _23852_);
  or g_34123_(_23676_, _23681_, _23854_);
  and g_34124_(_23851_, _23854_, _23855_);
  or g_34125_(_23850_, _23852_, _23856_);
  and g_34126_(_23849_, _23855_, _23857_);
  or g_34127_(_23848_, _23856_, _23858_);
  and g_34128_(_23837_, _23857_, _23859_);
  or g_34129_(_23836_, _23858_, _23860_);
  and g_34130_(_19552_, _23823_, _23861_);
  or g_34131_(out[272], _23822_, _23862_);
  and g_34132_(_23811_, _23862_, _23863_);
  or g_34133_(_23812_, _23861_, _23865_);
  and g_34134_(_23828_, _23863_, _23866_);
  or g_34135_(_23829_, _23865_, _23867_);
  and g_34136_(_23783_, _23866_, _23868_);
  or g_34137_(_23784_, _23867_, _23869_);
  and g_34138_(_23860_, _23869_, _23870_);
  or g_34139_(_23859_, _23868_, _23871_);
  and g_34140_(_23652_, _23871_, _23872_);
  or g_34141_(_23651_, _23870_, _23873_);
  and g_34142_(_23665_, _23870_, _23874_);
  or g_34143_(_23667_, _23871_, _23876_);
  and g_34144_(_23873_, _23876_, _23877_);
  or g_34145_(_23872_, _23874_, _23878_);
  and g_34146_(_22428_, _23877_, _23879_);
  or g_34147_(_22429_, _23878_, _23880_);
  and g_34148_(_23670_, _23672_, _23881_);
  or g_34149_(_23671_, _23673_, _23882_);
  xor g_34150_(out[299], _22427_, _23883_);
  xor g_34151_(_19618_, _22427_, _23884_);
  and g_34152_(_23881_, _23884_, _23885_);
  or g_34153_(_23882_, _23883_, _23887_);
  and g_34154_(_23880_, _23887_, _23888_);
  or g_34155_(_23879_, _23885_, _23889_);
  and g_34156_(_22429_, _23878_, _23890_);
  or g_34157_(_22428_, _23877_, _23891_);
  and g_34158_(_23882_, _23883_, _23892_);
  or g_34159_(_23881_, _23884_, _23893_);
  and g_34160_(out[297], _22424_, _23894_);
  xor g_34161_(out[297], _22424_, _23895_);
  or g_34162_(_22426_, _23894_, _23896_);
  and g_34163_(_23689_, _23871_, _23898_);
  or g_34164_(_23687_, _23870_, _23899_);
  and g_34165_(_23692_, _23870_, _23900_);
  or g_34166_(_23691_, _23871_, _23901_);
  and g_34167_(_23899_, _23901_, _23902_);
  or g_34168_(_23898_, _23900_, _23903_);
  and g_34169_(_23896_, _23902_, _23904_);
  or g_34170_(_23895_, _23903_, _23905_);
  xor g_34171_(out[296], _22422_, _23906_);
  xor g_34172_(_19706_, _22422_, _23907_);
  and g_34173_(_23703_, _23870_, _23909_);
  or g_34174_(_23702_, _23871_, _23910_);
  and g_34175_(_23709_, _23871_, _23911_);
  or g_34176_(_23708_, _23870_, _23912_);
  and g_34177_(_23910_, _23912_, _23913_);
  or g_34178_(_23909_, _23911_, _23914_);
  or g_34179_(_23907_, _23913_, _23915_);
  or g_34180_(_23896_, _23902_, _23916_);
  and g_34181_(_23915_, _23916_, _23917_);
  or g_34182_(_23906_, _23914_, _23918_);
  xor g_34183_(_23906_, _23913_, _23920_);
  and g_34184_(_23891_, _23893_, _23921_);
  or g_34185_(_23890_, _23892_, _23922_);
  and g_34186_(_23888_, _23921_, _23923_);
  or g_34187_(_23889_, _23922_, _23924_);
  xor g_34188_(_23895_, _23902_, _23925_);
  or g_34189_(_23924_, _23925_, _23926_);
  and g_34190_(_23905_, _23918_, _23927_);
  and g_34191_(_23917_, _23927_, _23928_);
  and g_34192_(_23923_, _23928_, _23929_);
  or g_34193_(_23920_, _23926_, _23931_);
  and g_34194_(_23729_, _23870_, _23932_);
  and g_34195_(_23727_, _23871_, _23933_);
  or g_34196_(_23932_, _23933_, _23934_);
  or g_34197_(_22420_, _23934_, _23935_);
  xor g_34198_(out[295], _22419_, _23936_);
  xor g_34199_(_19629_, _22419_, _23937_);
  and g_34200_(_23731_, _23870_, _23938_);
  and g_34201_(_23736_, _23871_, _23939_);
  or g_34202_(_23938_, _23939_, _23940_);
  and g_34203_(_23937_, _23940_, _23942_);
  or g_34204_(_23937_, _23940_, _23943_);
  xor g_34205_(_22420_, _23934_, _23944_);
  and g_34206_(_23943_, _23944_, _23945_);
  not g_34207_(_23945_, _23946_);
  xor g_34208_(_23937_, _23940_, _23947_);
  and g_34209_(_23944_, _23947_, _23948_);
  or g_34210_(_23942_, _23946_, _23949_);
  or g_34211_(_19983_, _20106_, _23950_);
  not g_34212_(_23950_, _23951_);
  and g_34213_(_22417_, _23950_, _23953_);
  or g_34214_(_22416_, _23951_, _23954_);
  or g_34215_(_23755_, _23870_, _23955_);
  or g_34216_(_23748_, _23871_, _23956_);
  and g_34217_(_23955_, _23956_, _23957_);
  and g_34218_(_23954_, _23957_, _23958_);
  xor g_34219_(out[293], _22416_, _23959_);
  xor g_34220_(_19651_, _22416_, _23960_);
  and g_34221_(_23760_, _23870_, _23961_);
  or g_34222_(_23759_, _23871_, _23962_);
  and g_34223_(_23767_, _23871_, _23964_);
  or g_34224_(_23766_, _23870_, _23965_);
  and g_34225_(_23962_, _23965_, _23966_);
  or g_34226_(_23961_, _23964_, _23967_);
  and g_34227_(_23960_, _23966_, _23968_);
  or g_34228_(_23958_, _23968_, _23969_);
  or g_34229_(_23960_, _23966_, _23970_);
  or g_34230_(_23954_, _23957_, _23971_);
  and g_34231_(_23970_, _23971_, _23972_);
  not g_34232_(_23972_, _23973_);
  or g_34233_(_23969_, _23973_, _23975_);
  or g_34234_(_23931_, _23975_, _23976_);
  or g_34235_(_23949_, _23976_, _23977_);
  xor g_34236_(out[291], _20106_, _23978_);
  xor g_34237_(_19695_, _20106_, _23979_);
  and g_34238_(_23785_, _23870_, _23980_);
  and g_34239_(_23793_, _23871_, _23981_);
  or g_34240_(_23980_, _23981_, _23982_);
  or g_34241_(_23979_, _23982_, _23983_);
  and g_34242_(_23801_, _23871_, _23984_);
  and g_34243_(_19886_, _23870_, _23986_);
  or g_34244_(_23984_, _23986_, _23987_);
  and g_34245_(_23979_, _23982_, _23988_);
  or g_34246_(_20108_, _23987_, _23989_);
  xor g_34247_(_20108_, _23987_, _23990_);
  xor g_34248_(_20107_, _23987_, _23991_);
  xor g_34249_(_23979_, _23982_, _23992_);
  xor g_34250_(_23978_, _23982_, _23993_);
  and g_34251_(_23990_, _23992_, _23994_);
  or g_34252_(_23991_, _23993_, _23995_);
  or g_34253_(_19541_, _23871_, _23997_);
  or g_34254_(_23815_, _23870_, _23998_);
  and g_34255_(_23997_, _23998_, _23999_);
  and g_34256_(out[289], _23999_, _24000_);
  or g_34257_(_19552_, _23871_, _24001_);
  or g_34258_(_23822_, _23870_, _24002_);
  and g_34259_(_24001_, _24002_, _24003_);
  and g_34260_(out[288], _24003_, _24004_);
  not g_34261_(_24004_, _24005_);
  xor g_34262_(out[289], _23999_, _24006_);
  xor g_34263_(_19673_, _23999_, _24008_);
  and g_34264_(_24005_, _24006_, _24009_);
  or g_34265_(_24004_, _24008_, _24010_);
  and g_34266_(_23994_, _24009_, _24011_);
  or g_34267_(_23995_, _24010_, _24012_);
  or g_34268_(_23988_, _23989_, _24013_);
  and g_34269_(_23983_, _24013_, _24014_);
  and g_34270_(_23994_, _24000_, _24015_);
  not g_34271_(_24015_, _24016_);
  and g_34272_(_24012_, _24014_, _24017_);
  and g_34273_(_24016_, _24017_, _24019_);
  or g_34274_(_23977_, _24019_, _24020_);
  and g_34275_(_23948_, _23969_, _24021_);
  and g_34276_(_23970_, _24021_, _24022_);
  or g_34277_(_23935_, _23942_, _24023_);
  and g_34278_(_23943_, _24023_, _24024_);
  not g_34279_(_24024_, _24025_);
  or g_34280_(_24022_, _24025_, _24026_);
  and g_34281_(_23929_, _24026_, _24027_);
  not g_34282_(_24027_, _24028_);
  or g_34283_(_23904_, _23918_, _24030_);
  and g_34284_(_23916_, _24030_, _24031_);
  or g_34285_(_23924_, _24031_, _24032_);
  and g_34286_(_23889_, _23893_, _24033_);
  or g_34287_(_23888_, _23892_, _24034_);
  and g_34288_(_24020_, _24032_, _24035_);
  not g_34289_(_24035_, _24036_);
  and g_34290_(_24028_, _24034_, _24037_);
  or g_34291_(_24027_, _24033_, _24038_);
  and g_34292_(_24035_, _24037_, _24039_);
  or g_34293_(_24036_, _24038_, _24041_);
  or g_34294_(out[288], _24003_, _24042_);
  not g_34295_(_24042_, _24043_);
  or g_34296_(_23977_, _24043_, _24044_);
  not g_34297_(_24044_, _24045_);
  and g_34298_(_24011_, _24045_, _24046_);
  or g_34299_(_24012_, _24044_, _24047_);
  and g_34300_(_24041_, _24047_, _24048_);
  or g_34301_(_24039_, _24046_, _24049_);
  and g_34302_(_22421_, _24048_, _24050_);
  and g_34303_(_23934_, _24049_, _24052_);
  or g_34304_(_24050_, _24052_, _24053_);
  or g_34305_(_22411_, _24053_, _24054_);
  or g_34306_(out[311], _22410_, _24055_);
  xor g_34307_(out[311], _22410_, _24056_);
  xor g_34308_(_19750_, _22410_, _24057_);
  or g_34309_(_23937_, _24049_, _24058_);
  not g_34310_(_24058_, _24059_);
  and g_34311_(_23940_, _24049_, _24060_);
  not g_34312_(_24060_, _24061_);
  and g_34313_(_24058_, _24061_, _24063_);
  or g_34314_(_24059_, _24060_, _24064_);
  and g_34315_(_24057_, _24064_, _24065_);
  or g_34316_(_24057_, _24064_, _24066_);
  xor g_34317_(out[309], _22407_, _24067_);
  xor g_34318_(_19783_, _22407_, _24068_);
  and g_34319_(_23967_, _24049_, _24069_);
  not g_34320_(_24069_, _24070_);
  or g_34321_(_23959_, _24049_, _24071_);
  not g_34322_(_24071_, _24072_);
  and g_34323_(_24070_, _24071_, _24074_);
  or g_34324_(_24069_, _24072_, _24075_);
  and g_34325_(_24067_, _24075_, _24076_);
  xor g_34326_(_22413_, _24053_, _24077_);
  xor g_34327_(_24057_, _24063_, _24078_);
  or g_34328_(_24077_, _24078_, _24079_);
  or g_34329_(_24076_, _24079_, _24080_);
  and g_34330_(out[312], _24055_, _24081_);
  or g_34331_(out[313], _24081_, _24082_);
  not g_34332_(_24082_, _24083_);
  or g_34333_(out[314], _24082_, _24085_);
  xor g_34334_(out[314], _24082_, _24086_);
  xor g_34335_(_19849_, _24082_, _24087_);
  or g_34336_(_22429_, _24049_, _24088_);
  not g_34337_(_24088_, _24089_);
  and g_34338_(_23878_, _24049_, _24090_);
  or g_34339_(_23877_, _24048_, _24091_);
  and g_34340_(_24088_, _24091_, _24092_);
  or g_34341_(_24089_, _24090_, _24093_);
  and g_34342_(_24086_, _24092_, _24094_);
  or g_34343_(_24087_, _24093_, _24096_);
  and g_34344_(_23881_, _23883_, _24097_);
  or g_34345_(_23882_, _23884_, _24098_);
  xor g_34346_(out[315], _24085_, _24099_);
  xor g_34347_(_19739_, _24085_, _24100_);
  and g_34348_(_24097_, _24100_, _24101_);
  or g_34349_(_24098_, _24099_, _24102_);
  and g_34350_(_24096_, _24102_, _24103_);
  or g_34351_(_24094_, _24101_, _24104_);
  and g_34352_(_24098_, _24099_, _24105_);
  and g_34353_(_24087_, _24093_, _24107_);
  or g_34354_(_24105_, _24107_, _24108_);
  or g_34355_(_24104_, _24108_, _24109_);
  and g_34356_(_23914_, _24049_, _24110_);
  not g_34357_(_24110_, _24111_);
  or g_34358_(_23906_, _24049_, _24112_);
  not g_34359_(_24112_, _24113_);
  and g_34360_(_24111_, _24112_, _24114_);
  or g_34361_(_24110_, _24113_, _24115_);
  xor g_34362_(out[312], _24055_, _24116_);
  xor g_34363_(_19827_, _24055_, _24118_);
  and g_34364_(_24114_, _24118_, _24119_);
  or g_34365_(_24115_, _24116_, _24120_);
  and g_34366_(out[313], _24081_, _24121_);
  xor g_34367_(out[313], _24081_, _24122_);
  or g_34368_(_24083_, _24121_, _24123_);
  or g_34369_(_23902_, _24048_, _24124_);
  or g_34370_(_23895_, _24049_, _24125_);
  and g_34371_(_24124_, _24125_, _24126_);
  not g_34372_(_24126_, _24127_);
  and g_34373_(_24122_, _24127_, _24129_);
  or g_34374_(_24123_, _24126_, _24130_);
  and g_34375_(_24120_, _24130_, _24131_);
  or g_34376_(_24119_, _24129_, _24132_);
  and g_34377_(_24123_, _24126_, _24133_);
  and g_34378_(_24115_, _24116_, _24134_);
  or g_34379_(_24133_, _24134_, _24135_);
  or g_34380_(_24132_, _24135_, _24136_);
  or g_34381_(_24109_, _24136_, _24137_);
  or g_34382_(_18408_, _20292_, _24138_);
  not g_34383_(_24138_, _24140_);
  and g_34384_(_22408_, _24138_, _24141_);
  or g_34385_(_22407_, _24140_, _24142_);
  or g_34386_(_23957_, _24048_, _24143_);
  or g_34387_(_23953_, _24049_, _24144_);
  and g_34388_(_24143_, _24144_, _24145_);
  not g_34389_(_24145_, _24146_);
  and g_34390_(_24142_, _24145_, _24147_);
  or g_34391_(_24141_, _24146_, _24148_);
  and g_34392_(_24068_, _24074_, _24149_);
  or g_34393_(_24067_, _24075_, _24151_);
  and g_34394_(_24148_, _24151_, _24152_);
  or g_34395_(_24147_, _24149_, _24153_);
  and g_34396_(_24141_, _24146_, _24154_);
  or g_34397_(_24142_, _24145_, _24155_);
  and g_34398_(_24152_, _24155_, _24156_);
  or g_34399_(_24153_, _24154_, _24157_);
  or g_34400_(_24080_, _24137_, _24158_);
  not g_34401_(_24158_, _24159_);
  and g_34402_(_24156_, _24159_, _24160_);
  or g_34403_(_24157_, _24158_, _24162_);
  xor g_34404_(out[307], _20292_, _24163_);
  not g_34405_(_24163_, _24164_);
  or g_34406_(_23979_, _24049_, _24165_);
  and g_34407_(_23982_, _24049_, _24166_);
  not g_34408_(_24166_, _24167_);
  and g_34409_(_24165_, _24167_, _24168_);
  and g_34410_(_24163_, _24168_, _24169_);
  and g_34411_(_23987_, _24049_, _24170_);
  not g_34412_(_24170_, _24171_);
  or g_34413_(_20108_, _24049_, _24173_);
  and g_34414_(_24171_, _24173_, _24174_);
  and g_34415_(_20293_, _24174_, _24175_);
  or g_34416_(_24169_, _24175_, _24176_);
  or g_34417_(_24163_, _24168_, _24177_);
  xor g_34418_(_24163_, _24168_, _24178_);
  xor g_34419_(_20293_, _24174_, _24179_);
  and g_34420_(_24178_, _24179_, _24180_);
  or g_34421_(_19673_, _24049_, _24181_);
  or g_34422_(_23999_, _24048_, _24182_);
  and g_34423_(_24181_, _24182_, _24184_);
  and g_34424_(out[305], _24184_, _24185_);
  and g_34425_(_24003_, _24049_, _24186_);
  not g_34426_(_24186_, _24187_);
  or g_34427_(out[288], _24049_, _24188_);
  and g_34428_(_24187_, _24188_, _24189_);
  not g_34429_(_24189_, _24190_);
  or g_34430_(_18562_, _24189_, _24191_);
  xor g_34431_(out[305], _24184_, _24192_);
  and g_34432_(_24191_, _24192_, _24193_);
  or g_34433_(_24185_, _24193_, _24195_);
  and g_34434_(_24180_, _24195_, _24196_);
  and g_34435_(_24176_, _24177_, _24197_);
  or g_34436_(_24196_, _24197_, _24198_);
  not g_34437_(_24198_, _24199_);
  or g_34438_(_24162_, _24199_, _24200_);
  or g_34439_(_24080_, _24152_, _24201_);
  or g_34440_(_24054_, _24065_, _24202_);
  and g_34441_(_24066_, _24202_, _24203_);
  and g_34442_(_24201_, _24203_, _24204_);
  or g_34443_(_24137_, _24204_, _24206_);
  or g_34444_(_24131_, _24133_, _24207_);
  or g_34445_(_24109_, _24207_, _24208_);
  or g_34446_(_24103_, _24105_, _24209_);
  and g_34447_(_24208_, _24209_, _24210_);
  and g_34448_(_24206_, _24210_, _24211_);
  and g_34449_(_24200_, _24211_, _24212_);
  or g_34450_(out[304], _24190_, _24213_);
  and g_34451_(_24180_, _24213_, _24214_);
  and g_34452_(_24193_, _24214_, _24215_);
  and g_34453_(_24160_, _24215_, _24217_);
  or g_34454_(_24212_, _24217_, _24218_);
  not g_34455_(_24218_, _24219_);
  and g_34456_(_24184_, _24218_, _24220_);
  not g_34457_(_24220_, _24221_);
  or g_34458_(out[305], _24218_, _24222_);
  not g_34459_(_24222_, _24223_);
  or g_34460_(_24220_, _24223_, _24224_);
  and g_34461_(_24221_, _24222_, _24225_);
  and g_34462_(_22403_, _24225_, _24226_);
  or g_34463_(_22404_, _24224_, _24228_);
  and g_34464_(_24146_, _24218_, _24229_);
  or g_34465_(_24145_, _24219_, _24230_);
  and g_34466_(_24142_, _24219_, _24231_);
  or g_34467_(_24141_, _24218_, _24232_);
  and g_34468_(_24230_, _24232_, _24233_);
  or g_34469_(_24229_, _24231_, _24234_);
  or g_34470_(_22358_, _22396_, _24235_);
  or g_34471_(_22364_, _22397_, _24236_);
  and g_34472_(_24235_, _24236_, _24237_);
  and g_34473_(_22233_, _22396_, _24239_);
  not g_34474_(_24239_, _24240_);
  and g_34475_(_18337_, _22397_, _24241_);
  or g_34476_(_18338_, _22396_, _24242_);
  and g_34477_(_24240_, _24242_, _24243_);
  or g_34478_(_24239_, _24241_, _24244_);
  or g_34479_(_20293_, _24218_, _24245_);
  not g_34480_(_24245_, _24246_);
  and g_34481_(_24174_, _24218_, _24247_);
  not g_34482_(_24247_, _24248_);
  or g_34483_(_24246_, _24247_, _24250_);
  and g_34484_(_24245_, _24248_, _24251_);
  and g_34485_(_24243_, _24251_, _24252_);
  or g_34486_(_24244_, _24250_, _24253_);
  and g_34487_(_22267_, _22397_, _24254_);
  and g_34488_(_22272_, _22396_, _24255_);
  or g_34489_(_24254_, _24255_, _24256_);
  and g_34490_(_24056_, _24219_, _24257_);
  or g_34491_(_24057_, _24218_, _24258_);
  and g_34492_(_24064_, _24218_, _24259_);
  or g_34493_(_24063_, _24219_, _24261_);
  and g_34494_(_24258_, _24261_, _24262_);
  or g_34495_(_24257_, _24259_, _24263_);
  xor g_34496_(_24256_, _24263_, _24264_);
  xor g_34497_(_24256_, _24262_, _24265_);
  and g_34498_(_22297_, _22303_, _24266_);
  and g_34499_(_24097_, _24099_, _24267_);
  or g_34500_(_24098_, _24100_, _24268_);
  xor g_34501_(_24266_, _24268_, _24269_);
  xor g_34502_(_24266_, _24267_, _24270_);
  or g_34503_(_22282_, _22396_, _24272_);
  not g_34504_(_24272_, _24273_);
  and g_34505_(_22289_, _22396_, _24274_);
  or g_34506_(_22288_, _22397_, _24275_);
  and g_34507_(_24272_, _24275_, _24276_);
  or g_34508_(_24273_, _24274_, _24277_);
  or g_34509_(_24067_, _24218_, _24278_);
  not g_34510_(_24278_, _24279_);
  and g_34511_(_24075_, _24218_, _24280_);
  or g_34512_(_24074_, _24219_, _24281_);
  and g_34513_(_24278_, _24281_, _24283_);
  or g_34514_(_24279_, _24280_, _24284_);
  and g_34515_(_24277_, _24283_, _24285_);
  or g_34516_(_24276_, _24284_, _24286_);
  or g_34517_(_22327_, _22396_, _24287_);
  not g_34518_(_24287_, _24288_);
  and g_34519_(_22334_, _22396_, _24289_);
  or g_34520_(_22333_, _22397_, _24290_);
  and g_34521_(_24287_, _24290_, _24291_);
  or g_34522_(_24288_, _24289_, _24292_);
  or g_34523_(_24116_, _24218_, _24294_);
  not g_34524_(_24294_, _24295_);
  and g_34525_(_24115_, _24218_, _24296_);
  or g_34526_(_24114_, _24219_, _24297_);
  and g_34527_(_24294_, _24297_, _24298_);
  or g_34528_(_24295_, _24296_, _24299_);
  and g_34529_(_24292_, _24298_, _24300_);
  or g_34530_(_24291_, _24299_, _24301_);
  or g_34531_(_22250_, _22397_, _24302_);
  or g_34532_(out[144], _22396_, _24303_);
  and g_34533_(_24302_, _24303_, _24305_);
  or g_34534_(_24189_, _24219_, _24306_);
  or g_34535_(out[304], _24218_, _24307_);
  and g_34536_(_24306_, _24307_, _24308_);
  or g_34537_(_22344_, _22397_, _24309_);
  or g_34538_(_22340_, _22396_, _24310_);
  and g_34539_(_24309_, _24310_, _24311_);
  and g_34540_(_24127_, _24218_, _24312_);
  or g_34541_(_24126_, _24219_, _24313_);
  and g_34542_(_24123_, _24219_, _24314_);
  or g_34543_(_24122_, _24218_, _24316_);
  and g_34544_(_24313_, _24316_, _24317_);
  or g_34545_(_24312_, _24314_, _24318_);
  and g_34546_(_22311_, _22396_, _24319_);
  and g_34547_(_22307_, _22397_, _24320_);
  or g_34548_(_24319_, _24320_, _24321_);
  and g_34549_(_24086_, _24219_, _24322_);
  or g_34550_(_24087_, _24218_, _24323_);
  and g_34551_(_24093_, _24218_, _24324_);
  not g_34552_(_24324_, _24325_);
  and g_34553_(_24323_, _24325_, _24327_);
  or g_34554_(_24322_, _24324_, _24328_);
  xor g_34555_(_24321_, _24327_, _24329_);
  xor g_34556_(_24321_, _24328_, _24330_);
  and g_34557_(_24291_, _24299_, _24331_);
  or g_34558_(_24292_, _24298_, _24332_);
  and g_34559_(_24276_, _24284_, _24333_);
  or g_34560_(_24277_, _24283_, _24334_);
  and g_34561_(_22404_, _24224_, _24335_);
  or g_34562_(_22403_, _24225_, _24336_);
  and g_34563_(_22229_, _22396_, _24338_);
  or g_34564_(_22228_, _22397_, _24339_);
  and g_34565_(_20525_, _22397_, _24340_);
  or g_34566_(_20526_, _22396_, _24341_);
  and g_34567_(_24339_, _24341_, _24342_);
  or g_34568_(_24338_, _24340_, _24343_);
  and g_34569_(_24168_, _24218_, _24344_);
  not g_34570_(_24344_, _24345_);
  or g_34571_(_24163_, _24218_, _24346_);
  not g_34572_(_24346_, _24347_);
  or g_34573_(_24344_, _24347_, _24349_);
  and g_34574_(_24345_, _24346_, _24350_);
  and g_34575_(_24342_, _24350_, _24351_);
  or g_34576_(_24343_, _24349_, _24352_);
  or g_34577_(_22274_, _22396_, _24353_);
  not g_34578_(_24353_, _24354_);
  and g_34579_(_22278_, _22396_, _24355_);
  not g_34580_(_24355_, _24356_);
  and g_34581_(_24353_, _24356_, _24357_);
  or g_34582_(_24354_, _24355_, _24358_);
  or g_34583_(_22411_, _24218_, _24360_);
  not g_34584_(_24360_, _24361_);
  and g_34585_(_24053_, _24218_, _24362_);
  not g_34586_(_24362_, _24363_);
  and g_34587_(_24360_, _24363_, _24364_);
  or g_34588_(_24361_, _24362_, _24365_);
  and g_34589_(_24358_, _24364_, _24366_);
  or g_34590_(_24357_, _24365_, _24367_);
  and g_34591_(_24343_, _24349_, _24368_);
  or g_34592_(_24342_, _24350_, _24369_);
  and g_34593_(_24244_, _24250_, _24371_);
  or g_34594_(_24243_, _24251_, _24372_);
  and g_34595_(_24357_, _24365_, _24373_);
  xor g_34596_(_24233_, _24237_, _24374_);
  xor g_34597_(_24234_, _24237_, _24375_);
  and g_34598_(_24329_, _24374_, _24376_);
  or g_34599_(_24330_, _24375_, _24377_);
  and g_34600_(_24301_, _24376_, _24378_);
  or g_34601_(_24300_, _24377_, _24379_);
  and g_34602_(_24228_, _24286_, _24380_);
  or g_34603_(_24226_, _24285_, _24382_);
  and g_34604_(_24265_, _24380_, _24383_);
  or g_34605_(_24264_, _24382_, _24384_);
  xor g_34606_(_24305_, _24308_, _24385_);
  or g_34607_(_24373_, _24385_, _24386_);
  not g_34608_(_24386_, _24387_);
  and g_34609_(_24383_, _24387_, _24388_);
  or g_34610_(_24384_, _24386_, _24389_);
  and g_34611_(_24378_, _24388_, _24390_);
  or g_34612_(_24379_, _24389_, _24391_);
  and g_34613_(_24269_, _24352_, _24393_);
  or g_34614_(_24270_, _24351_, _24394_);
  and g_34615_(_24336_, _24393_, _24395_);
  or g_34616_(_24335_, _24394_, _24396_);
  xor g_34617_(_24311_, _24318_, _24397_);
  xor g_34618_(_24311_, _24317_, _24398_);
  and g_34619_(_24367_, _24369_, _24399_);
  or g_34620_(_24366_, _24368_, _24400_);
  and g_34621_(_24397_, _24399_, _24401_);
  or g_34622_(_24398_, _24400_, _24402_);
  and g_34623_(_24334_, _24372_, _24404_);
  or g_34624_(_24333_, _24371_, _24405_);
  and g_34625_(_24253_, _24332_, _24406_);
  or g_34626_(_24252_, _24331_, _24407_);
  and g_34627_(_24404_, _24406_, _24408_);
  or g_34628_(_24405_, _24407_, _24409_);
  and g_34629_(_24401_, _24408_, _24410_);
  or g_34630_(_24402_, _24409_, _24411_);
  and g_34631_(_24395_, _24410_, _24412_);
  or g_34632_(_24396_, _24411_, _24413_);
  and g_34633_(_24390_, _24412_, _24415_);
  or g_34634_(_24391_, _24413_, _24416_);
  or g_34635_(out[5], _23050_, _24417_);
  or g_34636_(out[6], _24417_, _24418_);
  or g_34637_(out[7], _24418_, _24419_);
  or g_34638_(out[8], _24419_, _24420_);
  and g_34639_(out[9], _24420_, _24421_);
  or g_34640_(out[10], _24421_, _24422_);
  xor g_34641_(out[11], _24422_, _24423_);
  xor g_34642_(_19871_, _24422_, _24424_);
  or g_34643_(out[21], _23138_, _24426_);
  or g_34644_(out[22], _24426_, _24427_);
  or g_34645_(out[23], _24427_, _24428_);
  or g_34646_(out[24], _24428_, _24429_);
  and g_34647_(out[25], _24429_, _24430_);
  or g_34648_(out[26], _24430_, _24431_);
  xor g_34649_(out[27], _24431_, _24432_);
  xor g_34650_(_20003_, _24431_, _24433_);
  and g_34651_(_24424_, _24432_, _24434_);
  or g_34652_(_24423_, _24433_, _24435_);
  xor g_34653_(out[9], _24420_, _24437_);
  xor g_34654_(_19981_, _24420_, _24438_);
  xor g_34655_(out[25], _24429_, _24439_);
  xor g_34656_(_20113_, _24429_, _24440_);
  and g_34657_(_24437_, _24440_, _24441_);
  or g_34658_(_24438_, _24439_, _24442_);
  xor g_34659_(out[8], _24419_, _24443_);
  xor g_34660_(_19970_, _24419_, _24444_);
  xor g_34661_(out[24], _24428_, _24445_);
  xor g_34662_(_20102_, _24428_, _24446_);
  and g_34663_(_24443_, _24446_, _24448_);
  or g_34664_(_24444_, _24445_, _24449_);
  xor g_34665_(out[7], _24418_, _24450_);
  xor g_34666_(_19893_, _24418_, _24451_);
  xor g_34667_(out[23], _24427_, _24452_);
  xor g_34668_(_20014_, _24427_, _24453_);
  and g_34669_(_24450_, _24453_, _24454_);
  or g_34670_(_24451_, _24452_, _24455_);
  and g_34671_(_19959_, out[19], _24456_);
  or g_34672_(out[3], _20091_, _24457_);
  and g_34673_(out[2], _20080_, _24459_);
  or g_34674_(_19948_, out[18], _24460_);
  and g_34675_(_22599_, _24460_, _24461_);
  or g_34676_(_22588_, _24459_, _24462_);
  and g_34677_(_22786_, _24461_, _24463_);
  or g_34678_(_22775_, _24462_, _24464_);
  and g_34679_(_19948_, out[18], _24465_);
  or g_34680_(out[2], _20080_, _24466_);
  and g_34681_(out[3], _20091_, _24467_);
  or g_34682_(_19959_, out[19], _24468_);
  and g_34683_(_24466_, _24468_, _24470_);
  or g_34684_(_24465_, _24467_, _24471_);
  and g_34685_(_24464_, _24470_, _24472_);
  or g_34686_(_24463_, _24471_, _24473_);
  and g_34687_(_24457_, _24473_, _24474_);
  or g_34688_(_24456_, _24472_, _24475_);
  xor g_34689_(out[4], out[3], _24476_);
  xor g_34690_(_19915_, out[3], _24477_);
  xor g_34691_(out[20], out[19], _24478_);
  xor g_34692_(_20047_, out[19], _24479_);
  and g_34693_(_24477_, _24478_, _24481_);
  or g_34694_(_24476_, _24479_, _24482_);
  and g_34695_(_24475_, _24482_, _24483_);
  or g_34696_(_24474_, _24481_, _24484_);
  and g_34697_(_22830_, _24483_, _24485_);
  or g_34698_(_22819_, _24484_, _24486_);
  xor g_34699_(out[5], _23050_, _24487_);
  xor g_34700_(_19904_, _23050_, _24488_);
  xor g_34701_(out[21], _23138_, _24489_);
  xor g_34702_(_20036_, _23138_, _24490_);
  and g_34703_(_24488_, _24489_, _24492_);
  or g_34704_(_24487_, _24490_, _24493_);
  and g_34705_(_24476_, _24479_, _24494_);
  or g_34706_(_24477_, _24478_, _24495_);
  and g_34707_(_24493_, _24495_, _24496_);
  or g_34708_(_24492_, _24494_, _24497_);
  and g_34709_(_24486_, _24496_, _24498_);
  or g_34710_(_24485_, _24497_, _24499_);
  xor g_34711_(out[6], _24417_, _24500_);
  xor g_34712_(_19882_, _24417_, _24501_);
  xor g_34713_(out[22], _24426_, _24503_);
  xor g_34714_(_20025_, _24426_, _24504_);
  and g_34715_(_24500_, _24504_, _24505_);
  or g_34716_(_24501_, _24503_, _24506_);
  and g_34717_(_24487_, _24490_, _24507_);
  or g_34718_(_24488_, _24489_, _24508_);
  and g_34719_(_24506_, _24508_, _24509_);
  or g_34720_(_24505_, _24507_, _24510_);
  and g_34721_(_24499_, _24509_, _24511_);
  or g_34722_(_24498_, _24510_, _24512_);
  and g_34723_(_24451_, _24452_, _24514_);
  or g_34724_(_24450_, _24453_, _24515_);
  and g_34725_(_24501_, _24503_, _24516_);
  or g_34726_(_24500_, _24504_, _24517_);
  and g_34727_(_24515_, _24517_, _24518_);
  or g_34728_(_24514_, _24516_, _24519_);
  and g_34729_(_24512_, _24518_, _24520_);
  or g_34730_(_24511_, _24519_, _24521_);
  and g_34731_(_24455_, _24521_, _24522_);
  or g_34732_(_24454_, _24520_, _24523_);
  and g_34733_(_24444_, _24445_, _24525_);
  or g_34734_(_24443_, _24446_, _24526_);
  and g_34735_(_24449_, _24522_, _24527_);
  or g_34736_(_24448_, _24523_, _24528_);
  and g_34737_(_24442_, _24526_, _24529_);
  or g_34738_(_24441_, _24525_, _24530_);
  and g_34739_(_24528_, _24529_, _24531_);
  or g_34740_(_24527_, _24530_, _24532_);
  xor g_34741_(out[10], _24421_, _24533_);
  xor g_34742_(_19992_, _24421_, _24534_);
  xor g_34743_(out[26], _24430_, _24536_);
  xor g_34744_(_20124_, _24430_, _24537_);
  and g_34745_(_24533_, _24537_, _24538_);
  or g_34746_(_24534_, _24536_, _24539_);
  and g_34747_(_24438_, _24439_, _24540_);
  or g_34748_(_24437_, _24440_, _24541_);
  and g_34749_(_24539_, _24541_, _24542_);
  or g_34750_(_24538_, _24540_, _24543_);
  and g_34751_(_24532_, _24542_, _24544_);
  or g_34752_(_24531_, _24543_, _24545_);
  and g_34753_(_24423_, _24433_, _24547_);
  or g_34754_(_24424_, _24432_, _24548_);
  and g_34755_(_24534_, _24536_, _24549_);
  or g_34756_(_24533_, _24537_, _24550_);
  and g_34757_(_24548_, _24550_, _24551_);
  or g_34758_(_24547_, _24549_, _24552_);
  and g_34759_(_24545_, _24551_, _24553_);
  or g_34760_(_24544_, _24552_, _24554_);
  and g_34761_(_24435_, _24554_, _24555_);
  or g_34762_(_24434_, _24553_, _24556_);
  and g_34763_(_19937_, _24556_, _24558_);
  or g_34764_(out[0], _24555_, _24559_);
  and g_34765_(_20069_, _24555_, _24560_);
  or g_34766_(out[16], _24556_, _24561_);
  and g_34767_(_24559_, _24561_, _24562_);
  or g_34768_(_24558_, _24560_, _24563_);
  and g_34769_(_24536_, _24555_, _24564_);
  or g_34770_(_24537_, _24556_, _24565_);
  and g_34771_(_24533_, _24556_, _24566_);
  or g_34772_(_24534_, _24555_, _24567_);
  and g_34773_(_24565_, _24567_, _24569_);
  or g_34774_(_24564_, _24566_, _24570_);
  and g_34775_(out[36], out[35], _24571_);
  or g_34776_(out[37], _24571_, _24572_);
  or g_34777_(out[38], _24572_, _24573_);
  or g_34778_(out[39], _24573_, _24574_);
  or g_34779_(out[40], _24574_, _24575_);
  and g_34780_(out[41], _24575_, _24576_);
  or g_34781_(out[42], _24576_, _24577_);
  xor g_34782_(out[42], _24576_, _24578_);
  not g_34783_(_24578_, _24580_);
  or g_34784_(_24570_, _24580_, _24581_);
  and g_34785_(_24423_, _24432_, _24582_);
  or g_34786_(_24424_, _24433_, _24583_);
  xor g_34787_(out[43], _24577_, _24584_);
  xor g_34788_(_20135_, _24577_, _24585_);
  or g_34789_(_24583_, _24584_, _24586_);
  and g_34790_(_24581_, _24586_, _24587_);
  not g_34791_(_24587_, _24588_);
  and g_34792_(_24570_, _24580_, _24589_);
  or g_34793_(_24569_, _24578_, _24591_);
  or g_34794_(_24582_, _24585_, _24592_);
  not g_34795_(_24592_, _24593_);
  and g_34796_(_24591_, _24592_, _24594_);
  or g_34797_(_24589_, _24593_, _24595_);
  and g_34798_(_24587_, _24594_, _24596_);
  or g_34799_(_24588_, _24595_, _24597_);
  xor g_34800_(out[40], _24574_, _24598_);
  xor g_34801_(_20234_, _24574_, _24599_);
  and g_34802_(_24446_, _24555_, _24600_);
  or g_34803_(_24445_, _24556_, _24602_);
  and g_34804_(_24444_, _24556_, _24603_);
  or g_34805_(_24443_, _24555_, _24604_);
  and g_34806_(_24602_, _24604_, _24605_);
  or g_34807_(_24600_, _24603_, _24606_);
  and g_34808_(_24598_, _24606_, _24607_);
  or g_34809_(_24599_, _24605_, _24608_);
  xor g_34810_(out[41], _24575_, _24609_);
  xor g_34811_(_20245_, _24575_, _24610_);
  and g_34812_(_24439_, _24555_, _24611_);
  or g_34813_(_24440_, _24556_, _24613_);
  and g_34814_(_24437_, _24556_, _24614_);
  or g_34815_(_24438_, _24555_, _24615_);
  and g_34816_(_24613_, _24615_, _24616_);
  or g_34817_(_24611_, _24614_, _24617_);
  and g_34818_(_24610_, _24617_, _24618_);
  or g_34819_(_24609_, _24616_, _24619_);
  and g_34820_(_24608_, _24619_, _24620_);
  or g_34821_(_24607_, _24618_, _24621_);
  and g_34822_(_24599_, _24605_, _24622_);
  or g_34823_(_24598_, _24606_, _24624_);
  and g_34824_(_24609_, _24616_, _24625_);
  or g_34825_(_24610_, _24617_, _24626_);
  and g_34826_(_24624_, _24626_, _24627_);
  or g_34827_(_24622_, _24625_, _24628_);
  and g_34828_(_24620_, _24627_, _24629_);
  or g_34829_(_24621_, _24628_, _24630_);
  and g_34830_(_24596_, _24629_, _24631_);
  or g_34831_(_24597_, _24630_, _24632_);
  xor g_34832_(out[38], _24572_, _24633_);
  xor g_34833_(_20157_, _24572_, _24635_);
  and g_34834_(_24503_, _24555_, _24636_);
  or g_34835_(_24504_, _24556_, _24637_);
  and g_34836_(_24500_, _24556_, _24638_);
  or g_34837_(_24501_, _24555_, _24639_);
  and g_34838_(_24637_, _24639_, _24640_);
  or g_34839_(_24636_, _24638_, _24641_);
  and g_34840_(_24633_, _24640_, _24642_);
  or g_34841_(_24635_, _24641_, _24643_);
  xor g_34842_(out[39], _24573_, _24644_);
  xor g_34843_(_20146_, _24573_, _24646_);
  and g_34844_(_24453_, _24555_, _24647_);
  or g_34845_(_24452_, _24556_, _24648_);
  and g_34846_(_24451_, _24556_, _24649_);
  or g_34847_(_24450_, _24555_, _24650_);
  and g_34848_(_24648_, _24650_, _24651_);
  or g_34849_(_24647_, _24649_, _24652_);
  and g_34850_(_24644_, _24652_, _24653_);
  or g_34851_(_24646_, _24651_, _24654_);
  and g_34852_(_24643_, _24654_, _24655_);
  or g_34853_(_24642_, _24653_, _24657_);
  and g_34854_(_24646_, _24651_, _24658_);
  or g_34855_(_24644_, _24652_, _24659_);
  and g_34856_(_24635_, _24641_, _24660_);
  or g_34857_(_24633_, _24640_, _24661_);
  and g_34858_(_24659_, _24661_, _24662_);
  or g_34859_(_24658_, _24660_, _24663_);
  and g_34860_(_24655_, _24662_, _24664_);
  or g_34861_(_24657_, _24663_, _24665_);
  xor g_34862_(out[37], _24571_, _24666_);
  xor g_34863_(_20168_, _24571_, _24668_);
  and g_34864_(_24490_, _24555_, _24669_);
  or g_34865_(_24489_, _24556_, _24670_);
  and g_34866_(_24488_, _24556_, _24671_);
  or g_34867_(_24487_, _24555_, _24672_);
  and g_34868_(_24670_, _24672_, _24673_);
  or g_34869_(_24669_, _24671_, _24674_);
  and g_34870_(_24666_, _24674_, _24675_);
  or g_34871_(_24668_, _24673_, _24676_);
  xor g_34872_(out[36], out[35], _24677_);
  xor g_34873_(_20179_, out[35], _24679_);
  and g_34874_(_24478_, _24555_, _24680_);
  or g_34875_(_24479_, _24556_, _24681_);
  and g_34876_(_24476_, _24556_, _24682_);
  or g_34877_(_24477_, _24555_, _24683_);
  and g_34878_(_24681_, _24683_, _24684_);
  or g_34879_(_24680_, _24682_, _24685_);
  and g_34880_(_24679_, _24685_, _24686_);
  or g_34881_(_24677_, _24684_, _24687_);
  and g_34882_(_24676_, _24687_, _24688_);
  or g_34883_(_24675_, _24686_, _24690_);
  and g_34884_(_24677_, _24684_, _24691_);
  or g_34885_(_24679_, _24685_, _24692_);
  and g_34886_(_24668_, _24673_, _24693_);
  or g_34887_(_24666_, _24674_, _24694_);
  and g_34888_(_24692_, _24694_, _24695_);
  or g_34889_(_24691_, _24693_, _24696_);
  and g_34890_(_24688_, _24695_, _24697_);
  or g_34891_(_24690_, _24696_, _24698_);
  and g_34892_(_24664_, _24697_, _24699_);
  or g_34893_(_24665_, _24698_, _24701_);
  and g_34894_(_24631_, _24699_, _24702_);
  or g_34895_(_24632_, _24701_, _24703_);
  and g_34896_(out[19], _24555_, _24704_);
  or g_34897_(_20091_, _24556_, _24705_);
  and g_34898_(out[3], _24556_, _24706_);
  or g_34899_(_19959_, _24555_, _24707_);
  and g_34900_(_24705_, _24707_, _24708_);
  or g_34901_(_24704_, _24706_, _24709_);
  or g_34902_(_20223_, _24709_, _24710_);
  not g_34903_(_24710_, _24712_);
  and g_34904_(_19948_, _24556_, _24713_);
  or g_34905_(out[2], _24555_, _24714_);
  and g_34906_(_20080_, _24555_, _24715_);
  or g_34907_(out[18], _24556_, _24716_);
  and g_34908_(_24714_, _24716_, _24717_);
  or g_34909_(_24713_, _24715_, _24718_);
  and g_34910_(out[34], _24718_, _24719_);
  or g_34911_(_20212_, _24717_, _24720_);
  and g_34912_(_24710_, _24720_, _24721_);
  or g_34913_(_24712_, _24719_, _24723_);
  or g_34914_(out[35], _24708_, _24724_);
  not g_34915_(_24724_, _24725_);
  and g_34916_(_20212_, _24717_, _24726_);
  or g_34917_(out[34], _24718_, _24727_);
  and g_34918_(_24724_, _24727_, _24728_);
  or g_34919_(_24725_, _24726_, _24729_);
  and g_34920_(_24721_, _24728_, _24730_);
  or g_34921_(_24723_, _24729_, _24731_);
  and g_34922_(_20201_, _24562_, _24732_);
  or g_34923_(out[32], _24563_, _24734_);
  or g_34924_(out[1], _24555_, _24735_);
  or g_34925_(out[17], _24556_, _24736_);
  and g_34926_(_24735_, _24736_, _24737_);
  not g_34927_(_24737_, _24738_);
  and g_34928_(out[32], _24563_, _24739_);
  or g_34929_(_20201_, _24562_, _24740_);
  and g_34930_(_20190_, _24737_, _24741_);
  or g_34931_(out[33], _24738_, _24742_);
  xor g_34932_(_20190_, _24737_, _24743_);
  xor g_34933_(out[33], _24737_, _24745_);
  and g_34934_(_24740_, _24743_, _24746_);
  or g_34935_(_24739_, _24745_, _24747_);
  and g_34936_(_24734_, _24746_, _24748_);
  or g_34937_(_24732_, _24747_, _24749_);
  and g_34938_(_24730_, _24748_, _24750_);
  or g_34939_(_24731_, _24749_, _24751_);
  and g_34940_(_24702_, _24750_, _24752_);
  or g_34941_(_24703_, _24751_, _24753_);
  and g_34942_(_24742_, _24747_, _24754_);
  or g_34943_(_24741_, _24746_, _24756_);
  and g_34944_(_24730_, _24756_, _24757_);
  or g_34945_(_24731_, _24754_, _24758_);
  and g_34946_(_24724_, _24726_, _24759_);
  or g_34947_(_24725_, _24727_, _24760_);
  and g_34948_(_24710_, _24760_, _24761_);
  or g_34949_(_24712_, _24759_, _24762_);
  and g_34950_(_24758_, _24761_, _24763_);
  or g_34951_(_24757_, _24762_, _24764_);
  and g_34952_(_24702_, _24764_, _24765_);
  or g_34953_(_24703_, _24763_, _24767_);
  and g_34954_(_24657_, _24659_, _24768_);
  or g_34955_(_24655_, _24658_, _24769_);
  and g_34956_(_24690_, _24694_, _24770_);
  or g_34957_(_24688_, _24693_, _24771_);
  and g_34958_(_24664_, _24770_, _24772_);
  or g_34959_(_24665_, _24771_, _24773_);
  and g_34960_(_24769_, _24773_, _24774_);
  or g_34961_(_24768_, _24772_, _24775_);
  and g_34962_(_24631_, _24775_, _24776_);
  or g_34963_(_24632_, _24774_, _24778_);
  and g_34964_(_24621_, _24626_, _24779_);
  or g_34965_(_24620_, _24625_, _24780_);
  and g_34966_(_24596_, _24779_, _24781_);
  or g_34967_(_24597_, _24780_, _24782_);
  and g_34968_(_24588_, _24592_, _24783_);
  or g_34969_(_24587_, _24593_, _24784_);
  and g_34970_(_24782_, _24784_, _24785_);
  or g_34971_(_24781_, _24783_, _24786_);
  and g_34972_(_24767_, _24785_, _24787_);
  or g_34973_(_24765_, _24786_, _24789_);
  and g_34974_(_24778_, _24787_, _24790_);
  or g_34975_(_24776_, _24789_, _24791_);
  and g_34976_(_24753_, _24791_, _24792_);
  or g_34977_(_24752_, _24790_, _24793_);
  and g_34978_(_24563_, _24793_, _24794_);
  or g_34979_(_24562_, _24792_, _24795_);
  and g_34980_(_20201_, _24792_, _24796_);
  or g_34981_(out[32], _24793_, _24797_);
  and g_34982_(_24795_, _24797_, _24798_);
  or g_34983_(_24794_, _24796_, _24800_);
  and g_34984_(_24582_, _24584_, _24801_);
  or g_34985_(_24583_, _24585_, _24802_);
  and g_34986_(out[52], out[51], _24803_);
  or g_34987_(out[53], _24803_, _24804_);
  or g_34988_(out[54], _24804_, _24805_);
  or g_34989_(out[55], _24805_, _24806_);
  or g_34990_(out[56], _24806_, _24807_);
  and g_34991_(out[57], _24807_, _24808_);
  or g_34992_(out[58], _24808_, _24809_);
  xor g_34993_(out[59], _24809_, _24811_);
  xor g_34994_(_20267_, _24809_, _24812_);
  and g_34995_(_24801_, _24812_, _24813_);
  or g_34996_(_24802_, _24811_, _24814_);
  and g_34997_(_24578_, _24792_, _24815_);
  or g_34998_(_24580_, _24793_, _24816_);
  and g_34999_(_24570_, _24793_, _24817_);
  not g_35000_(_24817_, _24818_);
  and g_35001_(_24816_, _24818_, _24819_);
  or g_35002_(_24815_, _24817_, _24820_);
  xor g_35003_(out[58], _24808_, _24822_);
  xor g_35004_(_20388_, _24808_, _24823_);
  and g_35005_(_24819_, _24822_, _24824_);
  or g_35006_(_24820_, _24823_, _24825_);
  and g_35007_(_24814_, _24825_, _24826_);
  or g_35008_(_24813_, _24824_, _24827_);
  xor g_35009_(out[57], _24807_, _24828_);
  xor g_35010_(_20377_, _24807_, _24829_);
  and g_35011_(_24609_, _24792_, _24830_);
  or g_35012_(_24610_, _24793_, _24831_);
  and g_35013_(_24617_, _24793_, _24833_);
  not g_35014_(_24833_, _24834_);
  and g_35015_(_24831_, _24834_, _24835_);
  or g_35016_(_24830_, _24833_, _24836_);
  and g_35017_(_24828_, _24835_, _24837_);
  or g_35018_(_24829_, _24836_, _24838_);
  and g_35019_(_24820_, _24823_, _24839_);
  or g_35020_(_24819_, _24822_, _24840_);
  and g_35021_(_24802_, _24811_, _24841_);
  or g_35022_(_24801_, _24812_, _24842_);
  and g_35023_(_24840_, _24842_, _24844_);
  or g_35024_(_24839_, _24841_, _24845_);
  and g_35025_(_24838_, _24844_, _24846_);
  or g_35026_(_24837_, _24845_, _24847_);
  and g_35027_(_24826_, _24846_, _24848_);
  or g_35028_(_24827_, _24847_, _24849_);
  and g_35029_(_24829_, _24836_, _24850_);
  or g_35030_(_24828_, _24835_, _24851_);
  xor g_35031_(out[56], _24806_, _24852_);
  xor g_35032_(_20366_, _24806_, _24853_);
  or g_35033_(_24598_, _24793_, _24855_);
  not g_35034_(_24855_, _24856_);
  and g_35035_(_24606_, _24793_, _24857_);
  or g_35036_(_24605_, _24792_, _24858_);
  and g_35037_(_24855_, _24858_, _24859_);
  or g_35038_(_24856_, _24857_, _24860_);
  and g_35039_(_24852_, _24860_, _24861_);
  or g_35040_(_24853_, _24859_, _24862_);
  and g_35041_(_24851_, _24862_, _24863_);
  or g_35042_(_24850_, _24861_, _24864_);
  and g_35043_(_24853_, _24859_, _24866_);
  or g_35044_(_24852_, _24860_, _24867_);
  and g_35045_(_24863_, _24867_, _24868_);
  or g_35046_(_24864_, _24866_, _24869_);
  and g_35047_(_24848_, _24868_, _24870_);
  or g_35048_(_24849_, _24869_, _24871_);
  xor g_35049_(out[54], _24804_, _24872_);
  xor g_35050_(_20289_, _24804_, _24873_);
  and g_35051_(_24633_, _24792_, _24874_);
  or g_35052_(_24635_, _24793_, _24875_);
  and g_35053_(_24641_, _24793_, _24877_);
  not g_35054_(_24877_, _24878_);
  and g_35055_(_24875_, _24878_, _24879_);
  or g_35056_(_24874_, _24877_, _24880_);
  and g_35057_(_24872_, _24879_, _24881_);
  or g_35058_(_24873_, _24880_, _24882_);
  xor g_35059_(out[55], _24805_, _24883_);
  xor g_35060_(_20278_, _24805_, _24884_);
  and g_35061_(_24646_, _24792_, _24885_);
  or g_35062_(_24644_, _24793_, _24886_);
  and g_35063_(_24652_, _24793_, _24888_);
  or g_35064_(_24651_, _24792_, _24889_);
  and g_35065_(_24886_, _24889_, _24890_);
  or g_35066_(_24885_, _24888_, _24891_);
  and g_35067_(_24883_, _24891_, _24892_);
  or g_35068_(_24884_, _24890_, _24893_);
  and g_35069_(_24882_, _24893_, _24894_);
  or g_35070_(_24881_, _24892_, _24895_);
  and g_35071_(_24873_, _24880_, _24896_);
  or g_35072_(_24872_, _24879_, _24897_);
  xor g_35073_(out[53], _24803_, _24899_);
  xor g_35074_(_20300_, _24803_, _24900_);
  and g_35075_(_24668_, _24792_, _24901_);
  or g_35076_(_24666_, _24793_, _24902_);
  and g_35077_(_24674_, _24793_, _24903_);
  or g_35078_(_24673_, _24792_, _24904_);
  and g_35079_(_24902_, _24904_, _24905_);
  or g_35080_(_24901_, _24903_, _24906_);
  and g_35081_(_24900_, _24905_, _24907_);
  or g_35082_(_24899_, _24906_, _24908_);
  and g_35083_(_24884_, _24890_, _24910_);
  or g_35084_(_24883_, _24891_, _24911_);
  and g_35085_(_24908_, _24911_, _24912_);
  or g_35086_(_24907_, _24910_, _24913_);
  and g_35087_(_24897_, _24912_, _24914_);
  or g_35088_(_24896_, _24913_, _24915_);
  and g_35089_(_24894_, _24914_, _24916_);
  or g_35090_(_24895_, _24915_, _24917_);
  and g_35091_(_24899_, _24906_, _24918_);
  or g_35092_(_24900_, _24905_, _24919_);
  xor g_35093_(out[52], out[51], _24921_);
  xor g_35094_(_20311_, out[51], _24922_);
  and g_35095_(_24677_, _24792_, _24923_);
  or g_35096_(_24679_, _24793_, _24924_);
  and g_35097_(_24685_, _24793_, _24925_);
  not g_35098_(_24925_, _24926_);
  and g_35099_(_24924_, _24926_, _24927_);
  or g_35100_(_24923_, _24925_, _24928_);
  and g_35101_(_24922_, _24928_, _24929_);
  or g_35102_(_24921_, _24927_, _24930_);
  and g_35103_(_24919_, _24930_, _24932_);
  or g_35104_(_24918_, _24929_, _24933_);
  and g_35105_(_24921_, _24927_, _24934_);
  or g_35106_(_24922_, _24928_, _24935_);
  and g_35107_(_24932_, _24935_, _24936_);
  or g_35108_(_24933_, _24934_, _24937_);
  and g_35109_(_24916_, _24936_, _24938_);
  or g_35110_(_24917_, _24937_, _24939_);
  and g_35111_(out[35], _24792_, _24940_);
  or g_35112_(_20223_, _24793_, _24941_);
  and g_35113_(_24709_, _24793_, _24943_);
  or g_35114_(_24708_, _24792_, _24944_);
  and g_35115_(_24941_, _24944_, _24945_);
  or g_35116_(_24940_, _24943_, _24946_);
  or g_35117_(_20355_, _24946_, _24947_);
  not g_35118_(_24947_, _24948_);
  or g_35119_(_24717_, _24792_, _24949_);
  or g_35120_(out[34], _24793_, _24950_);
  and g_35121_(_24949_, _24950_, _24951_);
  not g_35122_(_24951_, _24952_);
  or g_35123_(out[51], _24945_, _24954_);
  and g_35124_(_20344_, _24951_, _24955_);
  and g_35125_(_24947_, _24954_, _24956_);
  xor g_35126_(_20355_, _24945_, _24957_);
  xor g_35127_(_20344_, _24951_, _24958_);
  xor g_35128_(out[50], _24951_, _24959_);
  and g_35129_(_24956_, _24958_, _24960_);
  or g_35130_(_24957_, _24959_, _24961_);
  and g_35131_(_24738_, _24793_, _24962_);
  or g_35132_(_24737_, _24792_, _24963_);
  and g_35133_(_20190_, _24792_, _24965_);
  or g_35134_(out[33], _24793_, _24966_);
  and g_35135_(_24963_, _24966_, _24967_);
  or g_35136_(_24962_, _24965_, _24968_);
  and g_35137_(_20322_, _24967_, _24969_);
  or g_35138_(out[49], _24968_, _24970_);
  and g_35139_(out[48], _24800_, _24971_);
  or g_35140_(_20333_, _24798_, _24972_);
  and g_35141_(out[49], _24968_, _24973_);
  or g_35142_(_20322_, _24967_, _24974_);
  and g_35143_(_24972_, _24974_, _24976_);
  or g_35144_(_24971_, _24973_, _24977_);
  and g_35145_(_24970_, _24977_, _24978_);
  or g_35146_(_24969_, _24976_, _24979_);
  and g_35147_(_24960_, _24979_, _24980_);
  or g_35148_(_24961_, _24978_, _24981_);
  and g_35149_(_24954_, _24955_, _24982_);
  not g_35150_(_24982_, _24983_);
  and g_35151_(_24947_, _24983_, _24984_);
  or g_35152_(_24948_, _24982_, _24985_);
  and g_35153_(_24981_, _24984_, _24987_);
  or g_35154_(_24980_, _24985_, _24988_);
  and g_35155_(_24938_, _24988_, _24989_);
  or g_35156_(_24939_, _24987_, _24990_);
  and g_35157_(_24916_, _24933_, _24991_);
  or g_35158_(_24917_, _24932_, _24992_);
  or g_35159_(_24894_, _24910_, _24993_);
  and g_35160_(_24895_, _24911_, _24994_);
  and g_35161_(_24992_, _24993_, _24995_);
  or g_35162_(_24991_, _24994_, _24996_);
  and g_35163_(_24990_, _24995_, _24998_);
  or g_35164_(_24989_, _24996_, _24999_);
  and g_35165_(_24870_, _24999_, _25000_);
  or g_35166_(_24871_, _24998_, _25001_);
  and g_35167_(_24848_, _24864_, _25002_);
  or g_35168_(_24849_, _24863_, _25003_);
  and g_35169_(_24827_, _24842_, _25004_);
  or g_35170_(_24826_, _24841_, _25005_);
  and g_35171_(_25003_, _25005_, _25006_);
  or g_35172_(_25002_, _25004_, _25007_);
  and g_35173_(_25001_, _25006_, _25009_);
  or g_35174_(_25000_, _25007_, _25010_);
  and g_35175_(_20333_, _24798_, _25011_);
  or g_35176_(out[48], _24800_, _25012_);
  and g_35177_(_24970_, _25012_, _25013_);
  or g_35178_(_24969_, _25011_, _25014_);
  and g_35179_(_24976_, _25013_, _25015_);
  or g_35180_(_24977_, _25014_, _25016_);
  and g_35181_(_24960_, _25015_, _25017_);
  or g_35182_(_24961_, _25016_, _25018_);
  and g_35183_(_24938_, _25017_, _25020_);
  or g_35184_(_24939_, _25018_, _25021_);
  and g_35185_(_24870_, _25020_, _25022_);
  or g_35186_(_24871_, _25021_, _25023_);
  and g_35187_(_25010_, _25023_, _25024_);
  or g_35188_(_25009_, _25022_, _25025_);
  and g_35189_(_24800_, _25025_, _25026_);
  or g_35190_(_24798_, _25024_, _25027_);
  or g_35191_(out[48], _25025_, _25028_);
  not g_35192_(_25028_, _25029_);
  and g_35193_(_25027_, _25028_, _25031_);
  or g_35194_(_25026_, _25029_, _25032_);
  and g_35195_(_24820_, _25025_, _25033_);
  not g_35196_(_25033_, _25034_);
  and g_35197_(_24822_, _25024_, _25035_);
  or g_35198_(_24823_, _25025_, _25036_);
  and g_35199_(_25034_, _25036_, _25037_);
  or g_35200_(_25033_, _25035_, _25038_);
  and g_35201_(out[68], out[67], _25039_);
  or g_35202_(out[69], _25039_, _25040_);
  or g_35203_(out[70], _25040_, _25042_);
  or g_35204_(out[71], _25042_, _25043_);
  or g_35205_(out[72], _25043_, _25044_);
  and g_35206_(out[73], _25044_, _25045_);
  or g_35207_(out[74], _25045_, _25046_);
  xor g_35208_(out[74], _25045_, _25047_);
  xor g_35209_(_20520_, _25045_, _25048_);
  and g_35210_(_25037_, _25047_, _25049_);
  or g_35211_(_25038_, _25048_, _25050_);
  and g_35212_(_24801_, _24811_, _25051_);
  or g_35213_(_24802_, _24812_, _25053_);
  xor g_35214_(out[75], _25046_, _25054_);
  xor g_35215_(_20399_, _25046_, _25055_);
  and g_35216_(_25051_, _25055_, _25056_);
  or g_35217_(_25053_, _25054_, _25057_);
  and g_35218_(_25050_, _25057_, _25058_);
  or g_35219_(_25049_, _25056_, _25059_);
  and g_35220_(_25038_, _25048_, _25060_);
  or g_35221_(_25037_, _25047_, _25061_);
  and g_35222_(_25053_, _25054_, _25062_);
  or g_35223_(_25051_, _25055_, _25064_);
  or g_35224_(_25060_, _25062_, _25065_);
  and g_35225_(_25058_, _25064_, _25066_);
  and g_35226_(_25061_, _25066_, _25067_);
  or g_35227_(_25059_, _25065_, _25068_);
  xor g_35228_(out[72], _25043_, _25069_);
  not g_35229_(_25069_, _25070_);
  and g_35230_(_24860_, _25025_, _25071_);
  or g_35231_(_24859_, _25024_, _25072_);
  or g_35232_(_24852_, _25025_, _25073_);
  not g_35233_(_25073_, _25075_);
  and g_35234_(_25072_, _25073_, _25076_);
  or g_35235_(_25071_, _25075_, _25077_);
  and g_35236_(_25069_, _25077_, _25078_);
  or g_35237_(_25070_, _25076_, _25079_);
  xor g_35238_(out[73], _25044_, _25080_);
  xor g_35239_(_20509_, _25044_, _25081_);
  and g_35240_(_24836_, _25025_, _25082_);
  not g_35241_(_25082_, _25083_);
  and g_35242_(_24828_, _25024_, _25084_);
  or g_35243_(_24829_, _25025_, _25086_);
  and g_35244_(_25083_, _25086_, _25087_);
  or g_35245_(_25082_, _25084_, _25088_);
  and g_35246_(_25081_, _25088_, _25089_);
  or g_35247_(_25080_, _25087_, _25090_);
  and g_35248_(_25079_, _25090_, _25091_);
  or g_35249_(_25078_, _25089_, _25092_);
  and g_35250_(_25080_, _25087_, _25093_);
  or g_35251_(_25081_, _25088_, _25094_);
  or g_35252_(_25069_, _25077_, _25095_);
  and g_35253_(_25091_, _25094_, _25097_);
  or g_35254_(_25092_, _25093_, _25098_);
  and g_35255_(_25067_, _25095_, _25099_);
  not g_35256_(_25099_, _25100_);
  and g_35257_(_25097_, _25099_, _25101_);
  or g_35258_(_25098_, _25100_, _25102_);
  and g_35259_(_24891_, _25025_, _25103_);
  or g_35260_(_24890_, _25024_, _25104_);
  or g_35261_(_24883_, _25025_, _25105_);
  not g_35262_(_25105_, _25106_);
  and g_35263_(_25104_, _25105_, _25108_);
  or g_35264_(_25103_, _25106_, _25109_);
  xor g_35265_(out[71], _25042_, _25110_);
  xor g_35266_(_20410_, _25042_, _25111_);
  and g_35267_(_25109_, _25110_, _25112_);
  or g_35268_(_25108_, _25111_, _25113_);
  xor g_35269_(out[70], _25040_, _25114_);
  xor g_35270_(_20421_, _25040_, _25115_);
  and g_35271_(_24880_, _25025_, _25116_);
  not g_35272_(_25116_, _25117_);
  and g_35273_(_24872_, _25024_, _25119_);
  or g_35274_(_24873_, _25025_, _25120_);
  and g_35275_(_25117_, _25120_, _25121_);
  or g_35276_(_25116_, _25119_, _25122_);
  and g_35277_(_25114_, _25121_, _25123_);
  or g_35278_(_25115_, _25122_, _25124_);
  and g_35279_(_25113_, _25124_, _25125_);
  or g_35280_(_25112_, _25123_, _25126_);
  and g_35281_(_25108_, _25111_, _25127_);
  or g_35282_(_25109_, _25110_, _25128_);
  and g_35283_(_25126_, _25128_, _25130_);
  or g_35284_(_25125_, _25127_, _25131_);
  xor g_35285_(out[69], _25039_, _25132_);
  xor g_35286_(_20432_, _25039_, _25133_);
  and g_35287_(_24906_, _25025_, _25134_);
  or g_35288_(_24905_, _25024_, _25135_);
  or g_35289_(_24899_, _25025_, _25136_);
  not g_35290_(_25136_, _25137_);
  and g_35291_(_25135_, _25136_, _25138_);
  or g_35292_(_25134_, _25137_, _25139_);
  and g_35293_(_25132_, _25139_, _25141_);
  or g_35294_(_25133_, _25138_, _25142_);
  xor g_35295_(out[68], out[67], _25143_);
  xor g_35296_(_20443_, out[67], _25144_);
  and g_35297_(_24921_, _25024_, _25145_);
  or g_35298_(_24922_, _25025_, _25146_);
  and g_35299_(_24928_, _25025_, _25147_);
  not g_35300_(_25147_, _25148_);
  and g_35301_(_25146_, _25148_, _25149_);
  or g_35302_(_25145_, _25147_, _25150_);
  and g_35303_(_25143_, _25149_, _25152_);
  or g_35304_(_25144_, _25150_, _25153_);
  and g_35305_(out[51], _25024_, _25154_);
  or g_35306_(_20355_, _25025_, _25155_);
  and g_35307_(_24946_, _25025_, _25156_);
  or g_35308_(_24945_, _25024_, _25157_);
  and g_35309_(_25155_, _25157_, _25158_);
  or g_35310_(_25154_, _25156_, _25159_);
  and g_35311_(_20487_, _25159_, _25160_);
  or g_35312_(out[67], _25158_, _25161_);
  and g_35313_(_24952_, _25025_, _25163_);
  or g_35314_(_24951_, _25024_, _25164_);
  and g_35315_(_20344_, _25024_, _25165_);
  or g_35316_(out[50], _25025_, _25166_);
  and g_35317_(_25164_, _25166_, _25167_);
  or g_35318_(_25163_, _25165_, _25168_);
  and g_35319_(out[66], _25168_, _25169_);
  or g_35320_(_20476_, _25167_, _25170_);
  and g_35321_(_25161_, _25170_, _25171_);
  or g_35322_(_25160_, _25169_, _25172_);
  and g_35323_(_20476_, _25167_, _25174_);
  or g_35324_(out[66], _25168_, _25175_);
  and g_35325_(_24968_, _25025_, _25176_);
  or g_35326_(_24967_, _25024_, _25177_);
  and g_35327_(_20322_, _25024_, _25178_);
  or g_35328_(out[49], _25025_, _25179_);
  and g_35329_(_25177_, _25179_, _25180_);
  or g_35330_(_25176_, _25178_, _25181_);
  and g_35331_(_20454_, _25180_, _25182_);
  or g_35332_(out[65], _25181_, _25183_);
  and g_35333_(_25175_, _25183_, _25185_);
  or g_35334_(_25174_, _25182_, _25186_);
  or g_35335_(_25172_, _25185_, _25187_);
  and g_35336_(_25144_, _25150_, _25188_);
  or g_35337_(_25143_, _25149_, _25189_);
  or g_35338_(_20487_, _25159_, _25190_);
  not g_35339_(_25190_, _25191_);
  and g_35340_(_25189_, _25190_, _25192_);
  or g_35341_(_25188_, _25191_, _25193_);
  and g_35342_(out[65], _25181_, _25194_);
  or g_35343_(_20454_, _25180_, _25196_);
  and g_35344_(out[64], _25032_, _25197_);
  or g_35345_(_20465_, _25031_, _25198_);
  and g_35346_(_25196_, _25198_, _25199_);
  or g_35347_(_25194_, _25197_, _25200_);
  or g_35348_(_25172_, _25200_, _25201_);
  and g_35349_(_25187_, _25192_, _25202_);
  or g_35350_(_25186_, _25199_, _25203_);
  and g_35351_(_25171_, _25203_, _25204_);
  and g_35352_(_25201_, _25202_, _25205_);
  or g_35353_(_25193_, _25204_, _25207_);
  and g_35354_(_25153_, _25207_, _25208_);
  or g_35355_(_25152_, _25205_, _25209_);
  and g_35356_(_25142_, _25209_, _25210_);
  or g_35357_(_25141_, _25208_, _25211_);
  and g_35358_(_25133_, _25138_, _25212_);
  or g_35359_(_25132_, _25139_, _25213_);
  and g_35360_(_25115_, _25122_, _25214_);
  or g_35361_(_25114_, _25121_, _25215_);
  or g_35362_(_25127_, _25214_, _25216_);
  and g_35363_(_25125_, _25128_, _25218_);
  and g_35364_(_25215_, _25218_, _25219_);
  or g_35365_(_25126_, _25216_, _25220_);
  and g_35366_(_25213_, _25219_, _25221_);
  or g_35367_(_25212_, _25220_, _25222_);
  and g_35368_(_25211_, _25221_, _25223_);
  or g_35369_(_25210_, _25222_, _25224_);
  and g_35370_(_25131_, _25224_, _25225_);
  or g_35371_(_25130_, _25223_, _25226_);
  and g_35372_(_25101_, _25226_, _25227_);
  or g_35373_(_25102_, _25225_, _25229_);
  and g_35374_(_25059_, _25064_, _25230_);
  or g_35375_(_25058_, _25062_, _25231_);
  and g_35376_(_25092_, _25094_, _25232_);
  or g_35377_(_25091_, _25093_, _25233_);
  and g_35378_(_25067_, _25232_, _25234_);
  or g_35379_(_25068_, _25233_, _25235_);
  and g_35380_(_25231_, _25235_, _25236_);
  or g_35381_(_25230_, _25234_, _25237_);
  and g_35382_(_25229_, _25236_, _25238_);
  or g_35383_(_25227_, _25237_, _25240_);
  and g_35384_(_20465_, _25031_, _25241_);
  or g_35385_(_25212_, _25241_, _25242_);
  or g_35386_(_25186_, _25242_, _25243_);
  or g_35387_(_25201_, _25243_, _25244_);
  not g_35388_(_25244_, _25245_);
  and g_35389_(_25142_, _25192_, _25246_);
  or g_35390_(_25141_, _25193_, _25247_);
  and g_35391_(_25153_, _25246_, _25248_);
  or g_35392_(_25152_, _25247_, _25249_);
  and g_35393_(_25245_, _25248_, _25251_);
  or g_35394_(_25244_, _25249_, _25252_);
  and g_35395_(_25101_, _25251_, _25253_);
  or g_35396_(_25102_, _25252_, _25254_);
  and g_35397_(_25219_, _25253_, _25255_);
  or g_35398_(_25220_, _25254_, _25256_);
  and g_35399_(_25240_, _25256_, _25257_);
  or g_35400_(_25238_, _25255_, _25258_);
  and g_35401_(_25032_, _25258_, _25259_);
  not g_35402_(_25259_, _25260_);
  or g_35403_(out[64], _25258_, _25262_);
  not g_35404_(_25262_, _25263_);
  and g_35405_(_25260_, _25262_, _25264_);
  or g_35406_(_25259_, _25263_, _25265_);
  and g_35407_(_25038_, _25258_, _25266_);
  not g_35408_(_25266_, _25267_);
  or g_35409_(_25048_, _25258_, _25268_);
  not g_35410_(_25268_, _25269_);
  and g_35411_(_25267_, _25268_, _25270_);
  or g_35412_(_25266_, _25269_, _25271_);
  and g_35413_(out[84], out[83], _25273_);
  or g_35414_(out[85], _25273_, _25274_);
  or g_35415_(out[86], _25274_, _25275_);
  or g_35416_(out[87], _25275_, _25276_);
  or g_35417_(out[88], _25276_, _25277_);
  and g_35418_(out[89], _25277_, _25278_);
  or g_35419_(out[90], _25278_, _25279_);
  xor g_35420_(out[90], _25278_, _25280_);
  xor g_35421_(_20652_, _25278_, _25281_);
  and g_35422_(_25270_, _25280_, _25282_);
  or g_35423_(_25271_, _25281_, _25284_);
  and g_35424_(_25051_, _25054_, _25285_);
  or g_35425_(_25053_, _25055_, _25286_);
  xor g_35426_(out[91], _25279_, _25287_);
  xor g_35427_(_20531_, _25279_, _25288_);
  and g_35428_(_25285_, _25288_, _25289_);
  or g_35429_(_25286_, _25287_, _25290_);
  and g_35430_(_25284_, _25290_, _25291_);
  or g_35431_(_25282_, _25289_, _25292_);
  and g_35432_(_25286_, _25287_, _25293_);
  or g_35433_(_25285_, _25288_, _25295_);
  and g_35434_(_25271_, _25281_, _25296_);
  or g_35435_(_25270_, _25280_, _25297_);
  and g_35436_(_25295_, _25297_, _25298_);
  or g_35437_(_25293_, _25296_, _25299_);
  xor g_35438_(out[89], _25277_, _25300_);
  xor g_35439_(_20641_, _25277_, _25301_);
  and g_35440_(_25088_, _25258_, _25302_);
  not g_35441_(_25302_, _25303_);
  or g_35442_(_25081_, _25258_, _25304_);
  not g_35443_(_25304_, _25306_);
  and g_35444_(_25303_, _25304_, _25307_);
  or g_35445_(_25302_, _25306_, _25308_);
  and g_35446_(_25300_, _25307_, _25309_);
  or g_35447_(_25301_, _25308_, _25310_);
  and g_35448_(_25291_, _25298_, _25311_);
  or g_35449_(_25292_, _25299_, _25312_);
  and g_35450_(_25310_, _25311_, _25313_);
  or g_35451_(_25309_, _25312_, _25314_);
  and g_35452_(_25301_, _25308_, _25315_);
  or g_35453_(_25300_, _25307_, _25317_);
  xor g_35454_(out[88], _25276_, _25318_);
  xor g_35455_(_20630_, _25276_, _25319_);
  and g_35456_(_25077_, _25258_, _25320_);
  not g_35457_(_25320_, _25321_);
  or g_35458_(_25069_, _25258_, _25322_);
  not g_35459_(_25322_, _25323_);
  and g_35460_(_25321_, _25322_, _25324_);
  or g_35461_(_25320_, _25323_, _25325_);
  and g_35462_(_25318_, _25325_, _25326_);
  or g_35463_(_25319_, _25324_, _25328_);
  and g_35464_(_25317_, _25328_, _25329_);
  or g_35465_(_25315_, _25326_, _25330_);
  and g_35466_(_25319_, _25324_, _25331_);
  or g_35467_(_25318_, _25325_, _25332_);
  and g_35468_(_25329_, _25332_, _25333_);
  or g_35469_(_25330_, _25331_, _25334_);
  and g_35470_(_25313_, _25333_, _25335_);
  or g_35471_(_25314_, _25334_, _25336_);
  xor g_35472_(out[86], _25274_, _25337_);
  xor g_35473_(_20553_, _25274_, _25339_);
  and g_35474_(_25122_, _25258_, _25340_);
  or g_35475_(_25121_, _25257_, _25341_);
  and g_35476_(_25114_, _25257_, _25342_);
  or g_35477_(_25115_, _25258_, _25343_);
  and g_35478_(_25341_, _25343_, _25344_);
  or g_35479_(_25340_, _25342_, _25345_);
  and g_35480_(_25337_, _25344_, _25346_);
  or g_35481_(_25339_, _25345_, _25347_);
  and g_35482_(_25109_, _25258_, _25348_);
  or g_35483_(_25108_, _25257_, _25350_);
  and g_35484_(_25111_, _25257_, _25351_);
  or g_35485_(_25110_, _25258_, _25352_);
  and g_35486_(_25350_, _25352_, _25353_);
  or g_35487_(_25348_, _25351_, _25354_);
  xor g_35488_(out[87], _25275_, _25355_);
  xor g_35489_(_20542_, _25275_, _25356_);
  and g_35490_(_25354_, _25355_, _25357_);
  or g_35491_(_25353_, _25356_, _25358_);
  and g_35492_(_25347_, _25358_, _25359_);
  or g_35493_(_25346_, _25357_, _25361_);
  and g_35494_(_25339_, _25345_, _25362_);
  or g_35495_(_25337_, _25344_, _25363_);
  and g_35496_(_25353_, _25356_, _25364_);
  or g_35497_(_25354_, _25355_, _25365_);
  xor g_35498_(out[85], _25273_, _25366_);
  xor g_35499_(_20564_, _25273_, _25367_);
  and g_35500_(_25139_, _25258_, _25368_);
  not g_35501_(_25368_, _25369_);
  or g_35502_(_25132_, _25258_, _25370_);
  not g_35503_(_25370_, _25372_);
  and g_35504_(_25369_, _25370_, _25373_);
  or g_35505_(_25368_, _25372_, _25374_);
  and g_35506_(_25367_, _25373_, _25375_);
  or g_35507_(_25366_, _25374_, _25376_);
  xor g_35508_(out[84], out[83], _25377_);
  xor g_35509_(_20575_, out[83], _25378_);
  or g_35510_(_25144_, _25258_, _25379_);
  not g_35511_(_25379_, _25380_);
  and g_35512_(_25150_, _25258_, _25381_);
  not g_35513_(_25381_, _25383_);
  and g_35514_(_25379_, _25383_, _25384_);
  or g_35515_(_25380_, _25381_, _25385_);
  and g_35516_(_25377_, _25384_, _25386_);
  or g_35517_(_25378_, _25385_, _25387_);
  and g_35518_(_25366_, _25374_, _25388_);
  or g_35519_(_25367_, _25373_, _25389_);
  and g_35520_(_25378_, _25385_, _25390_);
  or g_35521_(_25377_, _25384_, _25391_);
  and g_35522_(_25389_, _25391_, _25392_);
  or g_35523_(_25388_, _25390_, _25394_);
  and g_35524_(_25376_, _25392_, _25395_);
  or g_35525_(_25375_, _25394_, _25396_);
  and g_35526_(_25359_, _25363_, _25397_);
  or g_35527_(_25361_, _25362_, _25398_);
  and g_35528_(_25365_, _25397_, _25399_);
  or g_35529_(_25364_, _25398_, _25400_);
  and g_35530_(_25387_, _25395_, _25401_);
  or g_35531_(_25386_, _25396_, _25402_);
  and g_35532_(_25399_, _25401_, _25403_);
  or g_35533_(_25400_, _25402_, _25405_);
  or g_35534_(_20487_, _25258_, _25406_);
  not g_35535_(_25406_, _25407_);
  and g_35536_(_25159_, _25258_, _25408_);
  not g_35537_(_25408_, _25409_);
  and g_35538_(_25406_, _25409_, _25410_);
  or g_35539_(_25407_, _25408_, _25411_);
  and g_35540_(out[83], _25410_, _25412_);
  or g_35541_(_20619_, _25411_, _25413_);
  or g_35542_(_25167_, _25257_, _25414_);
  not g_35543_(_25414_, _25416_);
  or g_35544_(out[66], _25258_, _25417_);
  not g_35545_(_25417_, _25418_);
  and g_35546_(_25414_, _25417_, _25419_);
  or g_35547_(_25416_, _25418_, _25420_);
  and g_35548_(out[82], _25420_, _25421_);
  or g_35549_(_20608_, _25419_, _25422_);
  and g_35550_(_25413_, _25422_, _25423_);
  or g_35551_(_25412_, _25421_, _25424_);
  and g_35552_(_20619_, _25411_, _25425_);
  or g_35553_(out[83], _25410_, _25427_);
  and g_35554_(_20608_, _25419_, _25428_);
  or g_35555_(out[82], _25420_, _25429_);
  and g_35556_(_25427_, _25429_, _25430_);
  or g_35557_(_25425_, _25428_, _25431_);
  and g_35558_(_25423_, _25430_, _25432_);
  or g_35559_(_25424_, _25431_, _25433_);
  and g_35560_(_25181_, _25258_, _25434_);
  not g_35561_(_25434_, _25435_);
  or g_35562_(out[65], _25258_, _25436_);
  not g_35563_(_25436_, _25438_);
  and g_35564_(_25435_, _25436_, _25439_);
  or g_35565_(_25434_, _25438_, _25440_);
  and g_35566_(_20586_, _25439_, _25441_);
  or g_35567_(out[81], _25440_, _25442_);
  and g_35568_(out[80], _25265_, _25443_);
  or g_35569_(_20597_, _25264_, _25444_);
  xor g_35570_(_20586_, _25439_, _25445_);
  xor g_35571_(out[81], _25439_, _25446_);
  and g_35572_(_25444_, _25445_, _25447_);
  or g_35573_(_25443_, _25446_, _25449_);
  and g_35574_(_25442_, _25449_, _25450_);
  or g_35575_(_25441_, _25447_, _25451_);
  and g_35576_(_25432_, _25451_, _25452_);
  or g_35577_(_25433_, _25450_, _25453_);
  and g_35578_(_25427_, _25428_, _25454_);
  or g_35579_(_25425_, _25429_, _25455_);
  and g_35580_(_25413_, _25455_, _25456_);
  or g_35581_(_25412_, _25454_, _25457_);
  and g_35582_(_25453_, _25456_, _25458_);
  or g_35583_(_25452_, _25457_, _25460_);
  and g_35584_(_25403_, _25460_, _25461_);
  or g_35585_(_25405_, _25458_, _25462_);
  and g_35586_(_25394_, _25399_, _25463_);
  or g_35587_(_25392_, _25400_, _25464_);
  and g_35588_(_25376_, _25463_, _25465_);
  or g_35589_(_25375_, _25464_, _25466_);
  and g_35590_(_25361_, _25365_, _25467_);
  or g_35591_(_25359_, _25364_, _25468_);
  and g_35592_(_25466_, _25468_, _25469_);
  or g_35593_(_25465_, _25467_, _25471_);
  and g_35594_(_25462_, _25469_, _25472_);
  or g_35595_(_25461_, _25471_, _25473_);
  and g_35596_(_25335_, _25473_, _25474_);
  or g_35597_(_25336_, _25472_, _25475_);
  and g_35598_(_25313_, _25330_, _25476_);
  or g_35599_(_25314_, _25329_, _25477_);
  and g_35600_(_25292_, _25295_, _25478_);
  or g_35601_(_25291_, _25293_, _25479_);
  and g_35602_(_25477_, _25479_, _25480_);
  or g_35603_(_25476_, _25478_, _25482_);
  and g_35604_(_25475_, _25480_, _25483_);
  or g_35605_(_25474_, _25482_, _25484_);
  and g_35606_(_20597_, _25264_, _25485_);
  or g_35607_(out[80], _25265_, _25486_);
  and g_35608_(_25432_, _25447_, _25487_);
  or g_35609_(_25433_, _25449_, _25488_);
  and g_35610_(_25486_, _25487_, _25489_);
  or g_35611_(_25485_, _25488_, _25490_);
  and g_35612_(_25335_, _25489_, _25491_);
  or g_35613_(_25336_, _25490_, _25493_);
  and g_35614_(_25403_, _25491_, _25494_);
  or g_35615_(_25405_, _25493_, _25495_);
  and g_35616_(_25484_, _25495_, _25496_);
  or g_35617_(_25483_, _25494_, _25497_);
  and g_35618_(_25265_, _25497_, _25498_);
  and g_35619_(_20597_, _25496_, _25499_);
  or g_35620_(_25498_, _25499_, _25500_);
  and g_35621_(out[83], _25496_, _25501_);
  and g_35622_(_25411_, _25497_, _25502_);
  or g_35623_(_25501_, _25502_, _25504_);
  not g_35624_(_25504_, _25505_);
  or g_35625_(_20751_, _25504_, _25506_);
  and g_35626_(_25420_, _25497_, _25507_);
  and g_35627_(_20608_, _25496_, _25508_);
  or g_35628_(_25507_, _25508_, _25509_);
  not g_35629_(_25509_, _25510_);
  and g_35630_(out[98], _25509_, _25511_);
  or g_35631_(_20740_, _25510_, _25512_);
  and g_35632_(out[96], _25500_, _25513_);
  not g_35633_(_25513_, _25515_);
  and g_35634_(_25440_, _25497_, _25516_);
  and g_35635_(_20586_, _25496_, _25517_);
  or g_35636_(_25516_, _25517_, _25518_);
  and g_35637_(out[97], _25518_, _25519_);
  not g_35638_(_25519_, _25520_);
  and g_35639_(_25515_, _25520_, _25521_);
  or g_35640_(_25513_, _25519_, _25522_);
  or g_35641_(out[97], _25518_, _25523_);
  or g_35642_(out[98], _25509_, _25524_);
  and g_35643_(_25523_, _25524_, _25526_);
  and g_35644_(_25522_, _25526_, _25527_);
  or g_35645_(_25511_, _25527_, _25528_);
  and g_35646_(_25506_, _25528_, _25529_);
  and g_35647_(out[100], out[99], _25530_);
  xor g_35648_(_20707_, out[99], _25531_);
  and g_35649_(_25377_, _25496_, _25532_);
  and g_35650_(_25385_, _25497_, _25533_);
  or g_35651_(_25532_, _25533_, _25534_);
  or g_35652_(_25531_, _25534_, _25535_);
  not g_35653_(_25535_, _25537_);
  and g_35654_(_20751_, _25504_, _25538_);
  or g_35655_(out[99], _25505_, _25539_);
  and g_35656_(_25535_, _25539_, _25540_);
  or g_35657_(_25537_, _25538_, _25541_);
  or g_35658_(_25529_, _25541_, _25542_);
  or g_35659_(out[101], _25530_, _25543_);
  or g_35660_(out[102], _25543_, _25544_);
  xor g_35661_(out[102], _25543_, _25545_);
  xor g_35662_(_20685_, _25543_, _25546_);
  and g_35663_(_25345_, _25497_, _25548_);
  or g_35664_(_25344_, _25496_, _25549_);
  and g_35665_(_25337_, _25496_, _25550_);
  or g_35666_(_25339_, _25497_, _25551_);
  and g_35667_(_25549_, _25551_, _25552_);
  or g_35668_(_25548_, _25550_, _25553_);
  or g_35669_(_25546_, _25553_, _25554_);
  or g_35670_(out[103], _25544_, _25555_);
  xor g_35671_(out[103], _25544_, _25556_);
  xor g_35672_(_20674_, _25544_, _25557_);
  and g_35673_(_25354_, _25497_, _25559_);
  or g_35674_(_25353_, _25496_, _25560_);
  and g_35675_(_25356_, _25496_, _25561_);
  or g_35676_(_25355_, _25497_, _25562_);
  and g_35677_(_25560_, _25562_, _25563_);
  or g_35678_(_25559_, _25561_, _25564_);
  or g_35679_(_25557_, _25563_, _25565_);
  and g_35680_(_25554_, _25565_, _25566_);
  and g_35681_(_25531_, _25534_, _25567_);
  xor g_35682_(out[101], _25530_, _25568_);
  and g_35683_(_25374_, _25497_, _25570_);
  and g_35684_(_25367_, _25496_, _25571_);
  or g_35685_(_25570_, _25571_, _25572_);
  and g_35686_(_25568_, _25572_, _25573_);
  or g_35687_(_25567_, _25573_, _25574_);
  not g_35688_(_25574_, _25575_);
  and g_35689_(_25566_, _25575_, _25576_);
  and g_35690_(_25542_, _25576_, _25577_);
  or g_35691_(out[104], _25555_, _25578_);
  and g_35692_(out[105], _25578_, _25579_);
  or g_35693_(out[106], _25579_, _25581_);
  xor g_35694_(out[106], _25579_, _25582_);
  xor g_35695_(_20784_, _25579_, _25583_);
  and g_35696_(_25271_, _25497_, _25584_);
  and g_35697_(_25280_, _25496_, _25585_);
  or g_35698_(_25584_, _25585_, _25586_);
  not g_35699_(_25586_, _25587_);
  and g_35700_(_25582_, _25587_, _25588_);
  or g_35701_(_25583_, _25586_, _25589_);
  and g_35702_(_25285_, _25287_, _25590_);
  or g_35703_(_25286_, _25288_, _25592_);
  xor g_35704_(out[107], _25581_, _25593_);
  xor g_35705_(_20663_, _25581_, _25594_);
  and g_35706_(_25590_, _25594_, _25595_);
  or g_35707_(_25592_, _25593_, _25596_);
  and g_35708_(_25592_, _25593_, _25597_);
  or g_35709_(_25590_, _25594_, _25598_);
  and g_35710_(_25583_, _25586_, _25599_);
  not g_35711_(_25599_, _25600_);
  xor g_35712_(_20773_, _25578_, _25601_);
  and g_35713_(_25308_, _25497_, _25603_);
  and g_35714_(_25300_, _25496_, _25604_);
  or g_35715_(_25603_, _25604_, _25605_);
  or g_35716_(_25601_, _25605_, _25606_);
  xor g_35717_(out[104], _25555_, _25607_);
  and g_35718_(_25325_, _25497_, _25608_);
  and g_35719_(_25319_, _25496_, _25609_);
  or g_35720_(_25608_, _25609_, _25610_);
  and g_35721_(_25607_, _25610_, _25611_);
  not g_35722_(_25611_, _25612_);
  and g_35723_(_25601_, _25605_, _25614_);
  not g_35724_(_25614_, _25615_);
  and g_35725_(_25612_, _25615_, _25616_);
  or g_35726_(_25611_, _25614_, _25617_);
  or g_35727_(_25607_, _25610_, _25618_);
  and g_35728_(_25596_, _25600_, _25619_);
  or g_35729_(_25595_, _25599_, _25620_);
  and g_35730_(_25589_, _25598_, _25621_);
  or g_35731_(_25588_, _25597_, _25622_);
  and g_35732_(_25619_, _25621_, _25623_);
  or g_35733_(_25620_, _25622_, _25625_);
  and g_35734_(_25606_, _25618_, _25626_);
  not g_35735_(_25626_, _25627_);
  and g_35736_(_25616_, _25626_, _25628_);
  or g_35737_(_25617_, _25627_, _25629_);
  and g_35738_(_25623_, _25628_, _25630_);
  or g_35739_(_25625_, _25629_, _25631_);
  and g_35740_(_25557_, _25563_, _25632_);
  or g_35741_(_25556_, _25564_, _25633_);
  and g_35742_(_25546_, _25553_, _25634_);
  or g_35743_(_25545_, _25552_, _25636_);
  or g_35744_(_25568_, _25572_, _25637_);
  not g_35745_(_25637_, _25638_);
  and g_35746_(_25636_, _25637_, _25639_);
  or g_35747_(_25634_, _25638_, _25640_);
  and g_35748_(_25566_, _25640_, _25641_);
  or g_35749_(_25632_, _25641_, _25642_);
  or g_35750_(_25631_, _25642_, _25643_);
  or g_35751_(_25577_, _25643_, _25644_);
  and g_35752_(_25606_, _25617_, _25645_);
  not g_35753_(_25645_, _25647_);
  or g_35754_(_25625_, _25647_, _25648_);
  or g_35755_(_25589_, _25597_, _25649_);
  and g_35756_(_25596_, _25649_, _25650_);
  and g_35757_(_25648_, _25650_, _25651_);
  and g_35758_(_25644_, _25651_, _25652_);
  and g_35759_(_25521_, _25526_, _25653_);
  and g_35760_(_25540_, _25639_, _25654_);
  and g_35761_(_25653_, _25654_, _25655_);
  and g_35762_(_25506_, _25512_, _25656_);
  or g_35763_(out[96], _25500_, _25658_);
  and g_35764_(_25633_, _25658_, _25659_);
  and g_35765_(_25656_, _25659_, _25660_);
  and g_35766_(_25576_, _25660_, _25661_);
  and g_35767_(_25655_, _25661_, _25662_);
  and g_35768_(_25630_, _25662_, _25663_);
  or g_35769_(_25652_, _25663_, _25664_);
  not g_35770_(_25664_, _25665_);
  and g_35771_(_25500_, _25664_, _25666_);
  and g_35772_(_20729_, _25665_, _25667_);
  or g_35773_(_25666_, _25667_, _25669_);
  and g_35774_(out[99], _25665_, _25670_);
  and g_35775_(_25504_, _25664_, _25671_);
  or g_35776_(_25670_, _25671_, _25672_);
  or g_35777_(_20872_, _25672_, _25673_);
  and g_35778_(_25509_, _25664_, _25674_);
  and g_35779_(_20740_, _25665_, _25675_);
  or g_35780_(_25674_, _25675_, _25676_);
  and g_35781_(_20872_, _25672_, _25677_);
  or g_35782_(out[114], _25676_, _25678_);
  xor g_35783_(_20872_, _25672_, _25680_);
  xor g_35784_(out[115], _25672_, _25681_);
  xor g_35785_(out[114], _25676_, _25682_);
  xor g_35786_(_20861_, _25676_, _25683_);
  and g_35787_(_25680_, _25682_, _25684_);
  or g_35788_(_25681_, _25683_, _25685_);
  and g_35789_(_25518_, _25664_, _25686_);
  and g_35790_(_20718_, _25665_, _25687_);
  or g_35791_(_25686_, _25687_, _25688_);
  or g_35792_(out[113], _25688_, _25689_);
  and g_35793_(out[112], _25669_, _25691_);
  not g_35794_(_25691_, _25692_);
  xor g_35795_(out[113], _25688_, _25693_);
  xor g_35796_(_20850_, _25688_, _25694_);
  and g_35797_(_25692_, _25693_, _25695_);
  or g_35798_(_25691_, _25694_, _25696_);
  and g_35799_(_25689_, _25696_, _25697_);
  or g_35800_(_25685_, _25697_, _25698_);
  or g_35801_(_25677_, _25678_, _25699_);
  and g_35802_(_25673_, _25699_, _25700_);
  and g_35803_(_25698_, _25700_, _25702_);
  and g_35804_(_25590_, _25593_, _25703_);
  or g_35805_(_25592_, _25594_, _25704_);
  and g_35806_(out[116], out[115], _25705_);
  or g_35807_(out[117], _25705_, _25706_);
  or g_35808_(out[118], _25706_, _25707_);
  or g_35809_(out[119], _25707_, _25708_);
  or g_35810_(out[120], _25708_, _25709_);
  and g_35811_(out[121], _25709_, _25710_);
  or g_35812_(out[122], _25710_, _25711_);
  xor g_35813_(out[123], _25711_, _25713_);
  xor g_35814_(_20795_, _25711_, _25714_);
  and g_35815_(_25703_, _25714_, _25715_);
  or g_35816_(_25704_, _25713_, _25716_);
  and g_35817_(_25586_, _25664_, _25717_);
  not g_35818_(_25717_, _25718_);
  or g_35819_(_25583_, _25664_, _25719_);
  not g_35820_(_25719_, _25720_);
  and g_35821_(_25718_, _25719_, _25721_);
  or g_35822_(_25717_, _25720_, _25722_);
  xor g_35823_(out[122], _25710_, _25724_);
  not g_35824_(_25724_, _25725_);
  and g_35825_(_25721_, _25724_, _25726_);
  or g_35826_(_25722_, _25725_, _25727_);
  and g_35827_(_25716_, _25727_, _25728_);
  or g_35828_(_25715_, _25726_, _25729_);
  and g_35829_(_25704_, _25713_, _25730_);
  not g_35830_(_25730_, _25731_);
  and g_35831_(_25722_, _25725_, _25732_);
  or g_35832_(_25721_, _25724_, _25733_);
  and g_35833_(_25731_, _25733_, _25735_);
  or g_35834_(_25730_, _25732_, _25736_);
  and g_35835_(_25728_, _25735_, _25737_);
  or g_35836_(_25729_, _25736_, _25738_);
  xor g_35837_(out[121], _25709_, _25739_);
  and g_35838_(_25605_, _25664_, _25740_);
  not g_35839_(_25740_, _25741_);
  or g_35840_(_25601_, _25664_, _25742_);
  not g_35841_(_25742_, _25743_);
  and g_35842_(_25741_, _25742_, _25744_);
  or g_35843_(_25740_, _25743_, _25746_);
  or g_35844_(_25739_, _25744_, _25747_);
  xor g_35845_(out[120], _25708_, _25748_);
  not g_35846_(_25748_, _25749_);
  and g_35847_(_25610_, _25664_, _25750_);
  not g_35848_(_25750_, _25751_);
  or g_35849_(_25607_, _25664_, _25752_);
  not g_35850_(_25752_, _25753_);
  and g_35851_(_25751_, _25752_, _25754_);
  or g_35852_(_25750_, _25753_, _25755_);
  or g_35853_(_25749_, _25754_, _25757_);
  and g_35854_(_25747_, _25757_, _25758_);
  not g_35855_(_25758_, _25759_);
  and g_35856_(_25739_, _25744_, _25760_);
  not g_35857_(_25760_, _25761_);
  and g_35858_(_25749_, _25754_, _25762_);
  or g_35859_(_25748_, _25755_, _25763_);
  and g_35860_(_25761_, _25763_, _25764_);
  or g_35861_(_25760_, _25762_, _25765_);
  and g_35862_(_25758_, _25764_, _25766_);
  or g_35863_(_25759_, _25765_, _25768_);
  and g_35864_(_25737_, _25766_, _25769_);
  or g_35865_(_25738_, _25768_, _25770_);
  xor g_35866_(out[119], _25707_, _25771_);
  not g_35867_(_25771_, _25772_);
  or g_35868_(_25563_, _25665_, _25773_);
  or g_35869_(_25556_, _25664_, _25774_);
  and g_35870_(_25773_, _25774_, _25775_);
  or g_35871_(_25772_, _25775_, _25776_);
  xor g_35872_(out[118], _25706_, _25777_);
  not g_35873_(_25777_, _25779_);
  and g_35874_(_25553_, _25664_, _25780_);
  and g_35875_(_25545_, _25665_, _25781_);
  or g_35876_(_25780_, _25781_, _25782_);
  or g_35877_(_25779_, _25782_, _25783_);
  and g_35878_(_25776_, _25783_, _25784_);
  and g_35879_(_25772_, _25775_, _25785_);
  xor g_35880_(_25771_, _25775_, _25786_);
  xor g_35881_(_25777_, _25782_, _25787_);
  or g_35882_(_25786_, _25787_, _25788_);
  not g_35883_(_25788_, _25790_);
  xor g_35884_(out[116], out[115], _25791_);
  or g_35885_(_25531_, _25664_, _25792_);
  not g_35886_(_25792_, _25793_);
  and g_35887_(_25534_, _25664_, _25794_);
  not g_35888_(_25794_, _25795_);
  and g_35889_(_25792_, _25795_, _25796_);
  or g_35890_(_25793_, _25794_, _25797_);
  or g_35891_(_25791_, _25796_, _25798_);
  xor g_35892_(out[117], _25705_, _25799_);
  xor g_35893_(_20828_, _25705_, _25801_);
  and g_35894_(_25572_, _25664_, _25802_);
  not g_35895_(_25802_, _25803_);
  or g_35896_(_25568_, _25664_, _25804_);
  not g_35897_(_25804_, _25805_);
  and g_35898_(_25803_, _25804_, _25806_);
  or g_35899_(_25802_, _25805_, _25807_);
  or g_35900_(_25801_, _25806_, _25808_);
  and g_35901_(_25798_, _25808_, _25809_);
  not g_35902_(_25809_, _25810_);
  and g_35903_(_25801_, _25806_, _25812_);
  and g_35904_(_25791_, _25796_, _25813_);
  or g_35905_(_25812_, _25813_, _25814_);
  not g_35906_(_25814_, _25815_);
  and g_35907_(_25809_, _25815_, _25816_);
  or g_35908_(_25810_, _25814_, _25817_);
  and g_35909_(_25790_, _25816_, _25818_);
  or g_35910_(_25788_, _25817_, _25819_);
  and g_35911_(_25769_, _25818_, _25820_);
  or g_35912_(_25770_, _25819_, _25821_);
  or g_35913_(_25702_, _25821_, _25823_);
  or g_35914_(_25728_, _25730_, _25824_);
  or g_35915_(_25758_, _25760_, _25825_);
  or g_35916_(_25738_, _25825_, _25826_);
  and g_35917_(_25824_, _25826_, _25827_);
  or g_35918_(_25784_, _25785_, _25828_);
  or g_35919_(_25788_, _25809_, _25829_);
  or g_35920_(_25812_, _25829_, _25830_);
  and g_35921_(_25828_, _25830_, _25831_);
  or g_35922_(_25770_, _25831_, _25832_);
  and g_35923_(_25827_, _25832_, _25834_);
  and g_35924_(_25823_, _25834_, _25835_);
  or g_35925_(out[112], _25669_, _25836_);
  and g_35926_(_25684_, _25836_, _25837_);
  and g_35927_(_25695_, _25837_, _25838_);
  and g_35928_(_25820_, _25838_, _25839_);
  or g_35929_(_25835_, _25839_, _25840_);
  not g_35930_(_25840_, _25841_);
  and g_35931_(_25669_, _25840_, _25842_);
  not g_35932_(_25842_, _25843_);
  or g_35933_(out[112], _25840_, _25845_);
  not g_35934_(_25845_, _25846_);
  and g_35935_(_25843_, _25845_, _25847_);
  or g_35936_(_25842_, _25846_, _25848_);
  and g_35937_(_25724_, _25841_, _25849_);
  or g_35938_(_25725_, _25840_, _25850_);
  and g_35939_(_25722_, _25840_, _25851_);
  or g_35940_(_25721_, _25841_, _25852_);
  and g_35941_(_25850_, _25852_, _25853_);
  or g_35942_(_25849_, _25851_, _25854_);
  and g_35943_(out[132], out[131], _25856_);
  or g_35944_(out[133], _25856_, _25857_);
  or g_35945_(out[134], _25857_, _25858_);
  or g_35946_(out[135], _25858_, _25859_);
  or g_35947_(out[136], _25859_, _25860_);
  and g_35948_(out[137], _25860_, _25861_);
  or g_35949_(out[138], _25861_, _25862_);
  xor g_35950_(out[138], _25861_, _25863_);
  not g_35951_(_25863_, _25864_);
  or g_35952_(_25854_, _25864_, _25865_);
  not g_35953_(_25865_, _25867_);
  and g_35954_(_25703_, _25713_, _25868_);
  not g_35955_(_25868_, _25869_);
  xor g_35956_(out[139], _25862_, _25870_);
  or g_35957_(_25869_, _25870_, _25871_);
  and g_35958_(_25865_, _25871_, _25872_);
  or g_35959_(_25853_, _25863_, _25873_);
  and g_35960_(_25869_, _25870_, _25874_);
  xor g_35961_(out[137], _25860_, _25875_);
  and g_35962_(_25744_, _25840_, _25876_);
  or g_35963_(_25746_, _25841_, _25878_);
  or g_35964_(_25739_, _25840_, _25879_);
  not g_35965_(_25879_, _25880_);
  or g_35966_(_25876_, _25880_, _25881_);
  and g_35967_(_25878_, _25879_, _25882_);
  and g_35968_(_25875_, _25881_, _25883_);
  not g_35969_(_25883_, _25884_);
  xor g_35970_(out[136], _25859_, _25885_);
  not g_35971_(_25885_, _25886_);
  and g_35972_(_25748_, _25841_, _25887_);
  or g_35973_(_25749_, _25840_, _25889_);
  and g_35974_(_25754_, _25840_, _25890_);
  or g_35975_(_25755_, _25841_, _25891_);
  and g_35976_(_25889_, _25891_, _25892_);
  or g_35977_(_25887_, _25890_, _25893_);
  and g_35978_(_25886_, _25893_, _25894_);
  or g_35979_(_25885_, _25892_, _25895_);
  or g_35980_(_25875_, _25881_, _25896_);
  or g_35981_(_25886_, _25893_, _25897_);
  and g_35982_(_25896_, _25897_, _25898_);
  not g_35983_(_25898_, _25900_);
  and g_35984_(_25884_, _25898_, _25901_);
  or g_35985_(_25883_, _25900_, _25902_);
  or g_35986_(_25867_, _25874_, _25903_);
  and g_35987_(_25871_, _25873_, _25904_);
  not g_35988_(_25904_, _25905_);
  or g_35989_(_25903_, _25905_, _25906_);
  not g_35990_(_25906_, _25907_);
  and g_35991_(_25895_, _25907_, _25908_);
  or g_35992_(_25894_, _25906_, _25909_);
  and g_35993_(_25901_, _25908_, _25911_);
  or g_35994_(_25902_, _25909_, _25912_);
  xor g_35995_(out[134], _25857_, _25913_);
  not g_35996_(_25913_, _25914_);
  and g_35997_(_25777_, _25841_, _25915_);
  and g_35998_(_25782_, _25840_, _25916_);
  or g_35999_(_25915_, _25916_, _25917_);
  or g_36000_(_25914_, _25917_, _25918_);
  xor g_36001_(out[135], _25858_, _25919_);
  not g_36002_(_25919_, _25920_);
  or g_36003_(_25771_, _25840_, _25922_);
  or g_36004_(_25775_, _25841_, _25923_);
  and g_36005_(_25922_, _25923_, _25924_);
  or g_36006_(_25920_, _25924_, _25925_);
  and g_36007_(_25918_, _25925_, _25926_);
  not g_36008_(_25926_, _25927_);
  xor g_36009_(out[133], _25856_, _25928_);
  xor g_36010_(_20949_, _25856_, _25929_);
  or g_36011_(_25799_, _25840_, _25930_);
  not g_36012_(_25930_, _25931_);
  and g_36013_(_25807_, _25840_, _25933_);
  or g_36014_(_25806_, _25841_, _25934_);
  and g_36015_(_25930_, _25934_, _25935_);
  or g_36016_(_25931_, _25933_, _25936_);
  and g_36017_(_25929_, _25935_, _25937_);
  and g_36018_(_25914_, _25917_, _25938_);
  and g_36019_(_25920_, _25924_, _25939_);
  or g_36020_(_25938_, _25939_, _25940_);
  or g_36021_(_25937_, _25940_, _25941_);
  or g_36022_(_25927_, _25941_, _25942_);
  not g_36023_(_25942_, _25944_);
  xor g_36024_(out[132], out[131], _25945_);
  not g_36025_(_25945_, _25946_);
  and g_36026_(_25791_, _25841_, _25947_);
  and g_36027_(_25797_, _25840_, _25948_);
  or g_36028_(_25947_, _25948_, _25949_);
  not g_36029_(_25949_, _25950_);
  and g_36030_(_25946_, _25949_, _25951_);
  or g_36031_(_25945_, _25950_, _25952_);
  and g_36032_(_25928_, _25936_, _25953_);
  or g_36033_(_25929_, _25935_, _25955_);
  and g_36034_(_25952_, _25955_, _25956_);
  or g_36035_(_25951_, _25953_, _25957_);
  and g_36036_(_25945_, _25950_, _25958_);
  or g_36037_(_25946_, _25949_, _25959_);
  and g_36038_(_25956_, _25959_, _25960_);
  or g_36039_(_25957_, _25958_, _25961_);
  and g_36040_(_25944_, _25960_, _25962_);
  or g_36041_(_25942_, _25961_, _25963_);
  and g_36042_(out[115], _25841_, _25964_);
  and g_36043_(_25672_, _25840_, _25966_);
  or g_36044_(_25964_, _25966_, _25967_);
  or g_36045_(_21004_, _25967_, _25968_);
  and g_36046_(_21004_, _25967_, _25969_);
  and g_36047_(_25676_, _25840_, _25970_);
  and g_36048_(_20861_, _25841_, _25971_);
  or g_36049_(_25970_, _25971_, _25972_);
  or g_36050_(out[130], _25972_, _25973_);
  or g_36051_(_25969_, _25973_, _25974_);
  and g_36052_(_25968_, _25974_, _25975_);
  xor g_36053_(out[131], _25967_, _25977_);
  xor g_36054_(_20993_, _25972_, _25978_);
  or g_36055_(_25977_, _25978_, _25979_);
  not g_36056_(_25979_, _25980_);
  and g_36057_(_25688_, _25840_, _25981_);
  and g_36058_(_20850_, _25841_, _25982_);
  or g_36059_(_25981_, _25982_, _25983_);
  or g_36060_(out[129], _25983_, _25984_);
  and g_36061_(out[128], _25848_, _25985_);
  or g_36062_(_20982_, _25847_, _25986_);
  xor g_36063_(out[129], _25983_, _25988_);
  xor g_36064_(_20971_, _25983_, _25989_);
  and g_36065_(_25986_, _25988_, _25990_);
  or g_36066_(_25985_, _25989_, _25991_);
  and g_36067_(_25984_, _25991_, _25992_);
  or g_36068_(_25979_, _25992_, _25993_);
  and g_36069_(_25975_, _25993_, _25994_);
  or g_36070_(_25963_, _25994_, _25995_);
  or g_36071_(_25942_, _25956_, _25996_);
  or g_36072_(_25926_, _25939_, _25997_);
  and g_36073_(_25996_, _25997_, _25999_);
  and g_36074_(_25995_, _25999_, _26000_);
  or g_36075_(_25912_, _26000_, _26001_);
  or g_36076_(_25883_, _25898_, _26002_);
  or g_36077_(_25906_, _26002_, _26003_);
  or g_36078_(_25872_, _25874_, _26004_);
  and g_36079_(_26003_, _26004_, _26005_);
  and g_36080_(_26001_, _26005_, _26006_);
  or g_36081_(out[128], _25848_, _26007_);
  and g_36082_(_25980_, _26007_, _26008_);
  and g_36083_(_25990_, _26008_, _26010_);
  and g_36084_(_25911_, _26010_, _26011_);
  and g_36085_(_25962_, _26011_, _26012_);
  or g_36086_(_26006_, _26012_, _26013_);
  not g_36087_(_26013_, _26014_);
  or g_36088_(_25847_, _26014_, _26015_);
  or g_36089_(out[128], _26013_, _26016_);
  and g_36090_(_26015_, _26016_, _26017_);
  not g_36091_(_26017_, _26018_);
  and g_36092_(out[131], _26014_, _26019_);
  and g_36093_(_25967_, _26013_, _26021_);
  or g_36094_(_26019_, _26021_, _26022_);
  or g_36095_(_21136_, _26022_, _26023_);
  and g_36096_(_25972_, _26013_, _26024_);
  not g_36097_(_26024_, _26025_);
  or g_36098_(out[130], _26013_, _26026_);
  not g_36099_(_26026_, _26027_);
  and g_36100_(_26025_, _26026_, _26028_);
  or g_36101_(_26024_, _26027_, _26029_);
  and g_36102_(_21136_, _26022_, _26030_);
  or g_36103_(out[146], _26029_, _26032_);
  xor g_36104_(out[147], _26022_, _26033_);
  xor g_36105_(out[146], _26028_, _26034_);
  or g_36106_(_26033_, _26034_, _26035_);
  and g_36107_(_25983_, _26013_, _26036_);
  and g_36108_(_20971_, _26014_, _26037_);
  or g_36109_(_26036_, _26037_, _26038_);
  not g_36110_(_26038_, _26039_);
  or g_36111_(out[145], _26038_, _26040_);
  and g_36112_(out[144], _26018_, _26041_);
  xor g_36113_(_21103_, _26038_, _26043_);
  or g_36114_(_26041_, _26043_, _26044_);
  and g_36115_(_26040_, _26044_, _26045_);
  or g_36116_(_26035_, _26045_, _26046_);
  or g_36117_(_26030_, _26032_, _26047_);
  and g_36118_(_26023_, _26047_, _26048_);
  and g_36119_(_26046_, _26048_, _26049_);
  not g_36120_(_26049_, _26050_);
  and g_36121_(_25868_, _25870_, _26051_);
  not g_36122_(_26051_, _26052_);
  and g_36123_(out[148], out[147], _26054_);
  or g_36124_(out[149], _26054_, _26055_);
  or g_36125_(out[150], _26055_, _26056_);
  or g_36126_(out[151], _26056_, _26057_);
  or g_36127_(out[152], _26057_, _26058_);
  and g_36128_(out[153], _26058_, _26059_);
  or g_36129_(out[154], _26059_, _26060_);
  xor g_36130_(out[155], _26060_, _26061_);
  not g_36131_(_26061_, _26062_);
  and g_36132_(_26051_, _26062_, _26063_);
  or g_36133_(_26052_, _26061_, _26065_);
  xor g_36134_(out[154], _26059_, _26066_);
  not g_36135_(_26066_, _26067_);
  and g_36136_(_25854_, _26013_, _26068_);
  and g_36137_(_25863_, _26014_, _26069_);
  or g_36138_(_26068_, _26069_, _26070_);
  or g_36139_(_26067_, _26070_, _26071_);
  and g_36140_(_26065_, _26071_, _26072_);
  and g_36141_(_26052_, _26061_, _26073_);
  not g_36142_(_26073_, _26074_);
  and g_36143_(_26067_, _26070_, _26076_);
  or g_36144_(_26073_, _26076_, _26077_);
  not g_36145_(_26077_, _26078_);
  or g_36146_(_26063_, _26076_, _26079_);
  and g_36147_(_26071_, _26074_, _26080_);
  not g_36148_(_26080_, _26081_);
  and g_36149_(_26072_, _26078_, _26082_);
  or g_36150_(_26079_, _26081_, _26083_);
  or g_36151_(_25875_, _26013_, _26084_);
  not g_36152_(_26084_, _26085_);
  and g_36153_(_25881_, _26013_, _26087_);
  or g_36154_(_25882_, _26014_, _26088_);
  or g_36155_(_26085_, _26087_, _26089_);
  and g_36156_(_26084_, _26088_, _26090_);
  xor g_36157_(out[153], _26058_, _26091_);
  xor g_36158_(_21158_, _26058_, _26092_);
  and g_36159_(_26090_, _26092_, _26093_);
  or g_36160_(_26089_, _26091_, _26094_);
  xor g_36161_(out[152], _26057_, _26095_);
  not g_36162_(_26095_, _26096_);
  and g_36163_(_25893_, _26013_, _26098_);
  and g_36164_(_25885_, _26014_, _26099_);
  or g_36165_(_26098_, _26099_, _26100_);
  not g_36166_(_26100_, _26101_);
  and g_36167_(_26095_, _26101_, _26102_);
  or g_36168_(_26096_, _26100_, _26103_);
  and g_36169_(_26094_, _26103_, _26104_);
  or g_36170_(_26093_, _26102_, _26105_);
  and g_36171_(_26089_, _26091_, _26106_);
  or g_36172_(_26090_, _26092_, _26107_);
  or g_36173_(_26095_, _26101_, _26109_);
  and g_36174_(_26107_, _26109_, _26110_);
  and g_36175_(_26104_, _26110_, _26111_);
  and g_36176_(_26082_, _26111_, _26112_);
  not g_36177_(_26112_, _26113_);
  xor g_36178_(out[150], _26055_, _26114_);
  not g_36179_(_26114_, _26115_);
  and g_36180_(_25917_, _26013_, _26116_);
  and g_36181_(_25913_, _26014_, _26117_);
  or g_36182_(_26116_, _26117_, _26118_);
  not g_36183_(_26118_, _26120_);
  and g_36184_(_26114_, _26120_, _26121_);
  or g_36185_(_26115_, _26118_, _26122_);
  xor g_36186_(out[151], _26056_, _26123_);
  not g_36187_(_26123_, _26124_);
  or g_36188_(_25924_, _26014_, _26125_);
  or g_36189_(_25919_, _26013_, _26126_);
  and g_36190_(_26125_, _26126_, _26127_);
  not g_36191_(_26127_, _26128_);
  and g_36192_(_26123_, _26128_, _26129_);
  or g_36193_(_26124_, _26127_, _26131_);
  and g_36194_(_26122_, _26131_, _26132_);
  or g_36195_(_26121_, _26129_, _26133_);
  and g_36196_(_26124_, _26127_, _26134_);
  or g_36197_(_26123_, _26128_, _26135_);
  and g_36198_(_26115_, _26118_, _26136_);
  or g_36199_(_26114_, _26120_, _26137_);
  and g_36200_(_26135_, _26137_, _26138_);
  or g_36201_(_26134_, _26136_, _26139_);
  and g_36202_(_26132_, _26138_, _26140_);
  or g_36203_(_26133_, _26139_, _26142_);
  xor g_36204_(out[149], _26054_, _26143_);
  xor g_36205_(_21092_, _26054_, _26144_);
  or g_36206_(_25935_, _26014_, _26145_);
  or g_36207_(_25928_, _26013_, _26146_);
  and g_36208_(_26145_, _26146_, _26147_);
  not g_36209_(_26147_, _26148_);
  and g_36210_(_26143_, _26148_, _26149_);
  or g_36211_(_26144_, _26147_, _26150_);
  xor g_36212_(out[148], out[147], _26151_);
  not g_36213_(_26151_, _26153_);
  or g_36214_(_25945_, _26013_, _26154_);
  or g_36215_(_25949_, _26014_, _26155_);
  and g_36216_(_26154_, _26155_, _26156_);
  not g_36217_(_26156_, _26157_);
  and g_36218_(_26153_, _26156_, _26158_);
  or g_36219_(_26151_, _26157_, _26159_);
  and g_36220_(_26150_, _26159_, _26160_);
  or g_36221_(_26149_, _26158_, _26161_);
  and g_36222_(_26144_, _26147_, _26162_);
  or g_36223_(_26143_, _26148_, _26164_);
  and g_36224_(_26151_, _26157_, _26165_);
  or g_36225_(_26153_, _26156_, _26166_);
  and g_36226_(_26164_, _26166_, _26167_);
  or g_36227_(_26162_, _26165_, _26168_);
  and g_36228_(_26160_, _26167_, _26169_);
  or g_36229_(_26161_, _26168_, _26170_);
  and g_36230_(_26140_, _26169_, _26171_);
  or g_36231_(_26142_, _26170_, _26172_);
  and g_36232_(_26112_, _26171_, _26173_);
  or g_36233_(_26113_, _26172_, _26175_);
  and g_36234_(_26050_, _26173_, _26176_);
  or g_36235_(_26049_, _26175_, _26177_);
  or g_36236_(_26072_, _26073_, _26178_);
  not g_36237_(_26178_, _26179_);
  and g_36238_(_26105_, _26107_, _26180_);
  or g_36239_(_26104_, _26106_, _26181_);
  and g_36240_(_26082_, _26180_, _26182_);
  or g_36241_(_26083_, _26181_, _26183_);
  and g_36242_(_26178_, _26183_, _26184_);
  or g_36243_(_26179_, _26182_, _26186_);
  and g_36244_(_26133_, _26135_, _26187_);
  or g_36245_(_26132_, _26134_, _26188_);
  and g_36246_(_26161_, _26164_, _26189_);
  or g_36247_(_26160_, _26162_, _26190_);
  and g_36248_(_26140_, _26189_, _26191_);
  or g_36249_(_26142_, _26190_, _26192_);
  and g_36250_(_26188_, _26192_, _26193_);
  or g_36251_(_26187_, _26191_, _26194_);
  and g_36252_(_26112_, _26194_, _26195_);
  or g_36253_(_26113_, _26193_, _26197_);
  and g_36254_(_26184_, _26197_, _26198_);
  or g_36255_(_26186_, _26195_, _26199_);
  and g_36256_(_26177_, _26198_, _26200_);
  or g_36257_(_26176_, _26199_, _26201_);
  and g_36258_(_21114_, _26017_, _26202_);
  or g_36259_(_26035_, _26202_, _26203_);
  or g_36260_(_26044_, _26203_, _26204_);
  not g_36261_(_26204_, _26205_);
  and g_36262_(_26173_, _26205_, _26206_);
  or g_36263_(_26175_, _26204_, _26208_);
  and g_36264_(_26201_, _26208_, _26209_);
  or g_36265_(_26200_, _26206_, _26210_);
  or g_36266_(_26017_, _26209_, _26211_);
  or g_36267_(out[144], _26210_, _26212_);
  and g_36268_(_26211_, _26212_, _26213_);
  and g_36269_(out[164], out[163], _26214_);
  or g_36270_(out[165], _26214_, _26215_);
  or g_36271_(out[166], _26215_, _26216_);
  or g_36272_(out[167], _26216_, _26217_);
  or g_36273_(out[168], _26217_, _26219_);
  and g_36274_(out[169], _26219_, _26220_);
  or g_36275_(out[170], _26220_, _26221_);
  xor g_36276_(out[171], _26221_, _26222_);
  xor g_36277_(_18595_, _26221_, _26223_);
  and g_36278_(out[180], out[179], _26224_);
  or g_36279_(out[181], _26224_, _26225_);
  or g_36280_(out[182], _26225_, _26226_);
  or g_36281_(out[183], _26226_, _26227_);
  or g_36282_(out[184], _26227_, _26228_);
  and g_36283_(out[185], _26228_, _26230_);
  or g_36284_(out[186], _26230_, _26231_);
  xor g_36285_(out[187], _26231_, _26232_);
  xor g_36286_(_18716_, _26231_, _26233_);
  and g_36287_(_26223_, _26232_, _26234_);
  or g_36288_(_26222_, _26233_, _26235_);
  xor g_36289_(out[164], out[163], _26236_);
  xor g_36290_(_18639_, out[163], _26237_);
  xor g_36291_(out[180], out[179], _26238_);
  xor g_36292_(_18760_, out[179], _26239_);
  and g_36293_(_26236_, _26239_, _26241_);
  or g_36294_(_26237_, _26238_, _26242_);
  and g_36295_(_18672_, out[179], _26243_);
  or g_36296_(out[163], _18804_, _26244_);
  and g_36297_(out[163], _18804_, _26245_);
  or g_36298_(_18672_, out[179], _26246_);
  and g_36299_(out[162], _18793_, _26247_);
  or g_36300_(_18661_, out[178], _26248_);
  and g_36301_(_18661_, out[178], _26249_);
  or g_36302_(out[162], _18793_, _26250_);
  and g_36303_(_18485_, _26248_, _26252_);
  or g_36304_(_18484_, _26247_, _26253_);
  and g_36305_(_18489_, _26252_, _26254_);
  or g_36306_(_18488_, _26253_, _26255_);
  and g_36307_(_26246_, _26255_, _26256_);
  or g_36308_(_26245_, _26254_, _26257_);
  and g_36309_(_26250_, _26256_, _26258_);
  or g_36310_(_26249_, _26257_, _26259_);
  and g_36311_(_26244_, _26259_, _26260_);
  or g_36312_(_26243_, _26258_, _26261_);
  and g_36313_(_18511_, _26261_, _26263_);
  or g_36314_(_18510_, _26260_, _26264_);
  and g_36315_(_26242_, _26264_, _26265_);
  or g_36316_(_26241_, _26263_, _26266_);
  xor g_36317_(out[166], _26215_, _26267_);
  xor g_36318_(_18617_, _26215_, _26268_);
  xor g_36319_(out[182], _26225_, _26269_);
  xor g_36320_(_18738_, _26225_, _26270_);
  and g_36321_(_26267_, _26270_, _26271_);
  or g_36322_(_26268_, _26269_, _26272_);
  and g_36323_(_26237_, _26238_, _26274_);
  or g_36324_(_26236_, _26239_, _26275_);
  xor g_36325_(out[165], _26214_, _26276_);
  xor g_36326_(_18628_, _26214_, _26277_);
  xor g_36327_(out[181], _26224_, _26278_);
  xor g_36328_(_18749_, _26224_, _26279_);
  and g_36329_(_26276_, _26279_, _26280_);
  or g_36330_(_26277_, _26278_, _26281_);
  and g_36331_(_26275_, _26281_, _26282_);
  or g_36332_(_26274_, _26280_, _26283_);
  and g_36333_(_26272_, _26282_, _26285_);
  or g_36334_(_26271_, _26283_, _26286_);
  and g_36335_(_26266_, _26285_, _26287_);
  or g_36336_(_26265_, _26286_, _26288_);
  and g_36337_(_26277_, _26278_, _26289_);
  or g_36338_(_26276_, _26279_, _26290_);
  and g_36339_(_26272_, _26289_, _26291_);
  or g_36340_(_26271_, _26290_, _26292_);
  xor g_36341_(out[167], _26216_, _26293_);
  not g_36342_(_26293_, _26294_);
  xor g_36343_(out[183], _26226_, _26296_);
  not g_36344_(_26296_, _26297_);
  and g_36345_(_26294_, _26296_, _26298_);
  or g_36346_(_26293_, _26297_, _26299_);
  and g_36347_(_26268_, _26269_, _26300_);
  or g_36348_(_26267_, _26270_, _26301_);
  and g_36349_(_26292_, _26301_, _26302_);
  or g_36350_(_26291_, _26300_, _26303_);
  and g_36351_(_26299_, _26302_, _26304_);
  or g_36352_(_26298_, _26303_, _26305_);
  and g_36353_(_26288_, _26304_, _26307_);
  or g_36354_(_26287_, _26305_, _26308_);
  and g_36355_(_26293_, _26297_, _26309_);
  or g_36356_(_26294_, _26296_, _26310_);
  xor g_36357_(out[168], _26217_, _26311_);
  xor g_36358_(_18683_, _26217_, _26312_);
  xor g_36359_(out[184], _26227_, _26313_);
  xor g_36360_(_18815_, _26227_, _26314_);
  and g_36361_(_26311_, _26314_, _26315_);
  or g_36362_(_26312_, _26313_, _26316_);
  and g_36363_(_26310_, _26316_, _26318_);
  or g_36364_(_26309_, _26315_, _26319_);
  and g_36365_(_26308_, _26318_, _26320_);
  or g_36366_(_26307_, _26319_, _26321_);
  and g_36367_(_26312_, _26313_, _26322_);
  or g_36368_(_26311_, _26314_, _26323_);
  xor g_36369_(out[185], _26228_, _26324_);
  xor g_36370_(_18826_, _26228_, _26325_);
  xor g_36371_(out[169], _26219_, _26326_);
  xor g_36372_(_18694_, _26219_, _26327_);
  and g_36373_(_26325_, _26326_, _26329_);
  or g_36374_(_26324_, _26327_, _26330_);
  and g_36375_(_26323_, _26330_, _26331_);
  or g_36376_(_26322_, _26329_, _26332_);
  and g_36377_(_26321_, _26331_, _26333_);
  or g_36378_(_26320_, _26332_, _26334_);
  xor g_36379_(out[170], _26220_, _26335_);
  xor g_36380_(_18705_, _26220_, _26336_);
  xor g_36381_(out[186], _26230_, _26337_);
  xor g_36382_(_18837_, _26230_, _26338_);
  and g_36383_(_26335_, _26338_, _26340_);
  or g_36384_(_26336_, _26337_, _26341_);
  and g_36385_(_26324_, _26327_, _26342_);
  or g_36386_(_26325_, _26326_, _26343_);
  and g_36387_(_26341_, _26343_, _26344_);
  or g_36388_(_26340_, _26342_, _26345_);
  and g_36389_(_26334_, _26344_, _26346_);
  or g_36390_(_26333_, _26345_, _26347_);
  and g_36391_(_26222_, _26233_, _26348_);
  or g_36392_(_26223_, _26232_, _26349_);
  and g_36393_(_26336_, _26337_, _26351_);
  or g_36394_(_26335_, _26338_, _26352_);
  and g_36395_(_26349_, _26352_, _26353_);
  or g_36396_(_26348_, _26351_, _26354_);
  and g_36397_(_26347_, _26353_, _26355_);
  or g_36398_(_26346_, _26354_, _26356_);
  and g_36399_(_26235_, _26356_, _26357_);
  or g_36400_(_26234_, _26355_, _26358_);
  and g_36401_(_18782_, _26357_, _26359_);
  or g_36402_(out[176], _26358_, _26360_);
  and g_36403_(_18584_, _26358_, _26362_);
  or g_36404_(out[160], _26357_, _26363_);
  and g_36405_(_26360_, _26363_, _26364_);
  or g_36406_(_26359_, _26362_, _26365_);
  and g_36407_(_18914_, _26364_, _26366_);
  not g_36408_(_26366_, _26367_);
  and g_36409_(_26337_, _26357_, _26368_);
  or g_36410_(_26338_, _26358_, _26369_);
  and g_36411_(_26335_, _26358_, _26370_);
  or g_36412_(_26336_, _26357_, _26371_);
  and g_36413_(_26369_, _26371_, _26373_);
  or g_36414_(_26368_, _26370_, _26374_);
  and g_36415_(out[196], out[195], _26375_);
  or g_36416_(out[197], _26375_, _26376_);
  or g_36417_(out[198], _26376_, _26377_);
  or g_36418_(out[199], _26377_, _26378_);
  or g_36419_(out[200], _26378_, _26379_);
  and g_36420_(out[201], _26379_, _26380_);
  or g_36421_(out[202], _26380_, _26381_);
  xor g_36422_(out[202], _26380_, _26382_);
  not g_36423_(_26382_, _26384_);
  and g_36424_(_26374_, _26384_, _26385_);
  or g_36425_(_26373_, _26382_, _26386_);
  and g_36426_(_26222_, _26232_, _26387_);
  or g_36427_(_26223_, _26233_, _26388_);
  xor g_36428_(out[203], _26381_, _26389_);
  xor g_36429_(_18848_, _26381_, _26390_);
  and g_36430_(_26387_, _26390_, _26391_);
  or g_36431_(_26388_, _26389_, _26392_);
  and g_36432_(_26388_, _26389_, _26393_);
  or g_36433_(_26387_, _26390_, _26395_);
  and g_36434_(_26392_, _26395_, _26396_);
  and g_36435_(_26386_, _26396_, _26397_);
  and g_36436_(_26373_, _26382_, _26398_);
  or g_36437_(_26374_, _26384_, _26399_);
  and g_36438_(_26324_, _26357_, _26400_);
  or g_36439_(_26325_, _26358_, _26401_);
  and g_36440_(_26326_, _26358_, _26402_);
  or g_36441_(_26327_, _26357_, _26403_);
  and g_36442_(_26401_, _26403_, _26404_);
  or g_36443_(_26400_, _26402_, _26406_);
  xor g_36444_(out[201], _26379_, _26407_);
  not g_36445_(_26407_, _26408_);
  and g_36446_(_26404_, _26407_, _26409_);
  or g_36447_(_26406_, _26408_, _26410_);
  and g_36448_(_26399_, _26410_, _26411_);
  or g_36449_(_26385_, _26391_, _26412_);
  or g_36450_(_26393_, _26398_, _26413_);
  or g_36451_(_26412_, _26413_, _26414_);
  and g_36452_(_26397_, _26411_, _26415_);
  or g_36453_(_26409_, _26414_, _26417_);
  xor g_36454_(out[200], _26378_, _26418_);
  xor g_36455_(_18947_, _26378_, _26419_);
  and g_36456_(_26314_, _26357_, _26420_);
  or g_36457_(_26313_, _26358_, _26421_);
  and g_36458_(_26312_, _26358_, _26422_);
  or g_36459_(_26311_, _26357_, _26423_);
  and g_36460_(_26421_, _26423_, _26424_);
  or g_36461_(_26420_, _26422_, _26425_);
  and g_36462_(_26419_, _26424_, _26426_);
  not g_36463_(_26426_, _26428_);
  and g_36464_(_26406_, _26408_, _26429_);
  or g_36465_(_26404_, _26407_, _26430_);
  and g_36466_(_26418_, _26425_, _26431_);
  or g_36467_(_26419_, _26424_, _26432_);
  and g_36468_(_26430_, _26432_, _26433_);
  or g_36469_(_26429_, _26431_, _26434_);
  and g_36470_(_26428_, _26433_, _26435_);
  or g_36471_(_26426_, _26434_, _26436_);
  and g_36472_(_26415_, _26435_, _26437_);
  or g_36473_(_26417_, _26436_, _26439_);
  xor g_36474_(out[198], _26376_, _26440_);
  not g_36475_(_26440_, _26441_);
  or g_36476_(_26270_, _26358_, _26442_);
  or g_36477_(_26268_, _26357_, _26443_);
  and g_36478_(_26442_, _26443_, _26444_);
  xor g_36479_(out[199], _26377_, _26445_);
  xor g_36480_(_18859_, _26377_, _26446_);
  or g_36481_(_26296_, _26358_, _26447_);
  or g_36482_(_26293_, _26357_, _26448_);
  and g_36483_(_26447_, _26448_, _26450_);
  not g_36484_(_26450_, _26451_);
  and g_36485_(_26446_, _26450_, _26452_);
  or g_36486_(_26445_, _26451_, _26453_);
  and g_36487_(_26440_, _26444_, _26454_);
  not g_36488_(_26454_, _26455_);
  and g_36489_(_26445_, _26451_, _26456_);
  or g_36490_(_26446_, _26450_, _26457_);
  xor g_36491_(_26440_, _26444_, _26458_);
  xor g_36492_(_26441_, _26444_, _26459_);
  xor g_36493_(_26446_, _26450_, _26461_);
  or g_36494_(_26452_, _26456_, _26462_);
  and g_36495_(_26458_, _26461_, _26463_);
  or g_36496_(_26459_, _26462_, _26464_);
  xor g_36497_(out[196], out[195], _26465_);
  not g_36498_(_26465_, _26466_);
  and g_36499_(_26238_, _26357_, _26467_);
  or g_36500_(_26239_, _26358_, _26468_);
  and g_36501_(_26236_, _26358_, _26469_);
  or g_36502_(_26237_, _26357_, _26470_);
  and g_36503_(_26468_, _26470_, _26472_);
  or g_36504_(_26467_, _26469_, _26473_);
  and g_36505_(_26466_, _26473_, _26474_);
  or g_36506_(_26465_, _26472_, _26475_);
  xor g_36507_(out[197], _26375_, _26476_);
  xor g_36508_(_18881_, _26375_, _26477_);
  and g_36509_(_26279_, _26357_, _26478_);
  or g_36510_(_26278_, _26358_, _26479_);
  and g_36511_(_26277_, _26358_, _26480_);
  or g_36512_(_26276_, _26357_, _26481_);
  and g_36513_(_26479_, _26481_, _26483_);
  or g_36514_(_26478_, _26480_, _26484_);
  and g_36515_(_26476_, _26484_, _26485_);
  or g_36516_(_26477_, _26483_, _26486_);
  and g_36517_(_26475_, _26486_, _26487_);
  or g_36518_(_26474_, _26485_, _26488_);
  and g_36519_(_26465_, _26472_, _26489_);
  or g_36520_(_26466_, _26473_, _26490_);
  and g_36521_(_26477_, _26483_, _26491_);
  or g_36522_(_26476_, _26484_, _26492_);
  and g_36523_(_26490_, _26492_, _26494_);
  or g_36524_(_26489_, _26491_, _26495_);
  and g_36525_(_26487_, _26494_, _26496_);
  or g_36526_(_26488_, _26495_, _26497_);
  and g_36527_(_26463_, _26496_, _26498_);
  or g_36528_(_26464_, _26497_, _26499_);
  and g_36529_(_18793_, _26357_, _26500_);
  or g_36530_(out[178], _26358_, _26501_);
  and g_36531_(_18661_, _26358_, _26502_);
  or g_36532_(out[162], _26357_, _26503_);
  and g_36533_(_26501_, _26503_, _26505_);
  or g_36534_(_26500_, _26502_, _26506_);
  and g_36535_(out[163], _26358_, _26507_);
  or g_36536_(_18672_, _26357_, _26508_);
  and g_36537_(out[179], _26357_, _26509_);
  or g_36538_(_18804_, _26358_, _26510_);
  and g_36539_(_26508_, _26510_, _26511_);
  or g_36540_(_26507_, _26509_, _26512_);
  or g_36541_(_18936_, _26512_, _26513_);
  not g_36542_(_26513_, _26514_);
  and g_36543_(_18925_, _26505_, _26516_);
  or g_36544_(out[194], _26506_, _26517_);
  and g_36545_(out[192], _26365_, _26518_);
  or g_36546_(_18914_, _26364_, _26519_);
  and g_36547_(_18771_, _26357_, _26520_);
  or g_36548_(out[177], _26358_, _26521_);
  and g_36549_(_18650_, _26358_, _26522_);
  or g_36550_(out[161], _26357_, _26523_);
  and g_36551_(_26521_, _26523_, _26524_);
  or g_36552_(_26520_, _26522_, _26525_);
  and g_36553_(_18903_, _26524_, _26527_);
  or g_36554_(out[193], _26525_, _26528_);
  and g_36555_(_18936_, _26512_, _26529_);
  or g_36556_(out[195], _26511_, _26530_);
  and g_36557_(_26513_, _26530_, _26531_);
  or g_36558_(_26514_, _26529_, _26532_);
  xor g_36559_(_18925_, _26505_, _26533_);
  xor g_36560_(out[194], _26505_, _26534_);
  and g_36561_(_26531_, _26533_, _26535_);
  or g_36562_(_26532_, _26534_, _26536_);
  xor g_36563_(_18903_, _26524_, _26538_);
  xor g_36564_(out[193], _26524_, _26539_);
  and g_36565_(_26519_, _26538_, _26540_);
  or g_36566_(_26518_, _26539_, _26541_);
  and g_36567_(_26535_, _26540_, _26542_);
  or g_36568_(_26536_, _26541_, _26543_);
  and g_36569_(_26498_, _26542_, _26544_);
  or g_36570_(_26499_, _26543_, _26545_);
  and g_36571_(_26437_, _26544_, _26546_);
  or g_36572_(_26439_, _26545_, _26547_);
  and g_36573_(_26367_, _26546_, _26549_);
  or g_36574_(_26366_, _26547_, _26550_);
  and g_36575_(_26527_, _26535_, _26551_);
  or g_36576_(_26528_, _26536_, _26552_);
  and g_36577_(_26516_, _26530_, _26553_);
  or g_36578_(_26517_, _26529_, _26554_);
  and g_36579_(_26513_, _26554_, _26555_);
  or g_36580_(_26514_, _26553_, _26556_);
  and g_36581_(_26552_, _26555_, _26557_);
  or g_36582_(_26551_, _26556_, _26558_);
  and g_36583_(_26498_, _26558_, _26560_);
  or g_36584_(_26499_, _26557_, _26561_);
  and g_36585_(_26463_, _26488_, _26562_);
  or g_36586_(_26464_, _26487_, _26563_);
  and g_36587_(_26492_, _26562_, _26564_);
  or g_36588_(_26491_, _26563_, _26565_);
  and g_36589_(_26453_, _26454_, _26566_);
  or g_36590_(_26452_, _26455_, _26567_);
  and g_36591_(_26457_, _26567_, _26568_);
  or g_36592_(_26456_, _26566_, _26569_);
  and g_36593_(_26565_, _26568_, _26571_);
  or g_36594_(_26564_, _26569_, _26572_);
  and g_36595_(_26561_, _26571_, _26573_);
  or g_36596_(_26439_, _26573_, _26574_);
  and g_36597_(_26415_, _26434_, _26575_);
  or g_36598_(_26417_, _26433_, _26576_);
  and g_36599_(_26392_, _26399_, _26577_);
  or g_36600_(_26391_, _26398_, _26578_);
  and g_36601_(_26395_, _26578_, _26579_);
  or g_36602_(_26393_, _26577_, _26580_);
  and g_36603_(_26576_, _26580_, _26582_);
  or g_36604_(_26575_, _26579_, _26583_);
  and g_36605_(_26547_, _26582_, _26584_);
  or g_36606_(_26544_, _26572_, _26585_);
  or g_36607_(_26560_, _26585_, _26586_);
  and g_36608_(_26437_, _26586_, _26587_);
  and g_36609_(_26574_, _26584_, _26588_);
  or g_36610_(_26583_, _26587_, _26589_);
  and g_36611_(_26550_, _26589_, _26590_);
  or g_36612_(_26549_, _26588_, _26591_);
  or g_36613_(_26364_, _26590_, _26593_);
  not g_36614_(_26593_, _26594_);
  and g_36615_(_18914_, _26590_, _26595_);
  not g_36616_(_26595_, _26596_);
  and g_36617_(_26593_, _26596_, _26597_);
  or g_36618_(_26594_, _26595_, _26598_);
  and g_36619_(_26387_, _26389_, _26599_);
  or g_36620_(_26388_, _26390_, _26600_);
  and g_36621_(out[212], out[211], _26601_);
  or g_36622_(out[213], _26601_, _26602_);
  or g_36623_(out[214], _26602_, _26604_);
  or g_36624_(out[215], _26604_, _26605_);
  or g_36625_(out[216], _26605_, _26606_);
  and g_36626_(out[217], _26606_, _26607_);
  or g_36627_(out[218], _26607_, _26608_);
  xor g_36628_(out[219], _26608_, _26609_);
  xor g_36629_(_18958_, _26608_, _26610_);
  and g_36630_(_26599_, _26610_, _26611_);
  or g_36631_(_26600_, _26609_, _26612_);
  xor g_36632_(out[218], _26607_, _26613_);
  xor g_36633_(_19079_, _26607_, _26615_);
  or g_36634_(_26373_, _26590_, _26616_);
  not g_36635_(_26616_, _26617_);
  and g_36636_(_26382_, _26590_, _26618_);
  not g_36637_(_26618_, _26619_);
  and g_36638_(_26616_, _26619_, _26620_);
  or g_36639_(_26617_, _26618_, _26621_);
  and g_36640_(_26613_, _26620_, _26622_);
  or g_36641_(_26615_, _26621_, _26623_);
  and g_36642_(_26612_, _26623_, _26624_);
  or g_36643_(_26611_, _26622_, _26626_);
  and g_36644_(_26615_, _26621_, _26627_);
  or g_36645_(_26613_, _26620_, _26628_);
  and g_36646_(_26600_, _26609_, _26629_);
  or g_36647_(_26599_, _26610_, _26630_);
  xor g_36648_(out[217], _26606_, _26631_);
  xor g_36649_(_19068_, _26606_, _26632_);
  or g_36650_(_26404_, _26590_, _26633_);
  not g_36651_(_26633_, _26634_);
  and g_36652_(_26407_, _26590_, _26635_);
  not g_36653_(_26635_, _26637_);
  and g_36654_(_26633_, _26637_, _26638_);
  or g_36655_(_26634_, _26635_, _26639_);
  and g_36656_(_26631_, _26638_, _26640_);
  or g_36657_(_26632_, _26639_, _26641_);
  and g_36658_(_26630_, _26641_, _26642_);
  or g_36659_(_26629_, _26640_, _26643_);
  and g_36660_(_26628_, _26642_, _26644_);
  or g_36661_(_26627_, _26643_, _26645_);
  and g_36662_(_26624_, _26644_, _26646_);
  or g_36663_(_26626_, _26645_, _26648_);
  and g_36664_(_26632_, _26639_, _26649_);
  or g_36665_(_26631_, _26638_, _26650_);
  xor g_36666_(out[216], _26605_, _26651_);
  xor g_36667_(_19057_, _26605_, _26652_);
  or g_36668_(_26424_, _26590_, _26653_);
  not g_36669_(_26653_, _26654_);
  and g_36670_(_26419_, _26590_, _26655_);
  not g_36671_(_26655_, _26656_);
  and g_36672_(_26653_, _26656_, _26657_);
  or g_36673_(_26654_, _26655_, _26659_);
  and g_36674_(_26651_, _26659_, _26660_);
  or g_36675_(_26652_, _26657_, _26661_);
  and g_36676_(_26650_, _26661_, _26662_);
  or g_36677_(_26649_, _26660_, _26663_);
  and g_36678_(_26652_, _26657_, _26664_);
  or g_36679_(_26651_, _26659_, _26665_);
  and g_36680_(_26662_, _26665_, _26666_);
  or g_36681_(_26663_, _26664_, _26667_);
  and g_36682_(_26646_, _26666_, _26668_);
  or g_36683_(_26648_, _26667_, _26670_);
  xor g_36684_(out[215], _26604_, _26671_);
  xor g_36685_(_18969_, _26604_, _26672_);
  and g_36686_(_26451_, _26591_, _26673_);
  or g_36687_(_26450_, _26590_, _26674_);
  and g_36688_(_26446_, _26590_, _26675_);
  or g_36689_(_26445_, _26591_, _26676_);
  and g_36690_(_26674_, _26676_, _26677_);
  or g_36691_(_26673_, _26675_, _26678_);
  and g_36692_(_26671_, _26678_, _26679_);
  or g_36693_(_26672_, _26677_, _26681_);
  xor g_36694_(out[214], _26602_, _26682_);
  not g_36695_(_26682_, _26683_);
  or g_36696_(_26444_, _26590_, _26684_);
  not g_36697_(_26684_, _26685_);
  and g_36698_(_26440_, _26590_, _26686_);
  not g_36699_(_26686_, _26687_);
  and g_36700_(_26684_, _26687_, _26688_);
  or g_36701_(_26685_, _26686_, _26689_);
  and g_36702_(_26682_, _26688_, _26690_);
  or g_36703_(_26683_, _26689_, _26692_);
  and g_36704_(_26681_, _26692_, _26693_);
  or g_36705_(_26679_, _26690_, _26694_);
  xor g_36706_(out[213], _26601_, _26695_);
  xor g_36707_(_18991_, _26601_, _26696_);
  or g_36708_(_26483_, _26590_, _26697_);
  not g_36709_(_26697_, _26698_);
  and g_36710_(_26477_, _26590_, _26699_);
  not g_36711_(_26699_, _26700_);
  and g_36712_(_26697_, _26700_, _26701_);
  or g_36713_(_26698_, _26699_, _26703_);
  and g_36714_(_26696_, _26701_, _26704_);
  or g_36715_(_26695_, _26703_, _26705_);
  and g_36716_(_26672_, _26677_, _26706_);
  or g_36717_(_26671_, _26678_, _26707_);
  and g_36718_(_26683_, _26689_, _26708_);
  or g_36719_(_26682_, _26688_, _26709_);
  and g_36720_(_26707_, _26709_, _26710_);
  or g_36721_(_26706_, _26708_, _26711_);
  and g_36722_(_26705_, _26710_, _26712_);
  or g_36723_(_26704_, _26711_, _26714_);
  and g_36724_(_26693_, _26712_, _26715_);
  or g_36725_(_26694_, _26714_, _26716_);
  xor g_36726_(out[212], out[211], _26717_);
  xor g_36727_(_19002_, out[211], _26718_);
  and g_36728_(_26465_, _26590_, _26719_);
  not g_36729_(_26719_, _26720_);
  or g_36730_(_26472_, _26590_, _26721_);
  not g_36731_(_26721_, _26722_);
  and g_36732_(_26720_, _26721_, _26723_);
  or g_36733_(_26719_, _26722_, _26725_);
  and g_36734_(_26718_, _26725_, _26726_);
  or g_36735_(_26717_, _26723_, _26727_);
  and g_36736_(_26695_, _26703_, _26728_);
  or g_36737_(_26696_, _26701_, _26729_);
  and g_36738_(_26727_, _26729_, _26730_);
  or g_36739_(_26726_, _26728_, _26731_);
  and g_36740_(_26717_, _26723_, _26732_);
  or g_36741_(_26718_, _26725_, _26733_);
  and g_36742_(_26730_, _26733_, _26734_);
  or g_36743_(_26731_, _26732_, _26736_);
  and g_36744_(_26715_, _26734_, _26737_);
  or g_36745_(_26716_, _26736_, _26738_);
  and g_36746_(out[195], _26590_, _26739_);
  and g_36747_(_26512_, _26591_, _26740_);
  or g_36748_(_26739_, _26740_, _26741_);
  not g_36749_(_26741_, _26742_);
  or g_36750_(_19046_, _26741_, _26743_);
  not g_36751_(_26743_, _26744_);
  or g_36752_(_26505_, _26590_, _26745_);
  or g_36753_(out[194], _26591_, _26747_);
  and g_36754_(_26745_, _26747_, _26748_);
  not g_36755_(_26748_, _26749_);
  or g_36756_(out[211], _26742_, _26750_);
  not g_36757_(_26750_, _26751_);
  or g_36758_(out[210], _26749_, _26752_);
  not g_36759_(_26752_, _26753_);
  xor g_36760_(out[211], _26741_, _26754_);
  xor g_36761_(out[210], _26748_, _26755_);
  or g_36762_(_26754_, _26755_, _26756_);
  not g_36763_(_26756_, _26758_);
  or g_36764_(_26524_, _26590_, _26759_);
  not g_36765_(_26759_, _26760_);
  and g_36766_(_18903_, _26590_, _26761_);
  not g_36767_(_26761_, _26762_);
  and g_36768_(_26759_, _26762_, _26763_);
  or g_36769_(_26760_, _26761_, _26764_);
  and g_36770_(_19013_, _26763_, _26765_);
  or g_36771_(out[209], _26764_, _26766_);
  and g_36772_(out[208], _26598_, _26767_);
  or g_36773_(_19024_, _26597_, _26769_);
  xor g_36774_(_19013_, _26763_, _26770_);
  xor g_36775_(out[209], _26763_, _26771_);
  and g_36776_(_26769_, _26770_, _26772_);
  or g_36777_(_26767_, _26771_, _26773_);
  and g_36778_(_26766_, _26773_, _26774_);
  or g_36779_(_26765_, _26772_, _26775_);
  and g_36780_(_26758_, _26775_, _26776_);
  or g_36781_(_26756_, _26774_, _26777_);
  and g_36782_(_26750_, _26753_, _26778_);
  or g_36783_(_26751_, _26752_, _26780_);
  and g_36784_(_26743_, _26780_, _26781_);
  or g_36785_(_26744_, _26778_, _26782_);
  and g_36786_(_26777_, _26781_, _26783_);
  or g_36787_(_26776_, _26782_, _26784_);
  and g_36788_(_26737_, _26784_, _26785_);
  or g_36789_(_26738_, _26783_, _26786_);
  and g_36790_(_26715_, _26731_, _26787_);
  or g_36791_(_26716_, _26730_, _26788_);
  and g_36792_(_26694_, _26707_, _26789_);
  or g_36793_(_26693_, _26706_, _26791_);
  and g_36794_(_26788_, _26791_, _26792_);
  or g_36795_(_26787_, _26789_, _26793_);
  and g_36796_(_26786_, _26792_, _26794_);
  or g_36797_(_26785_, _26793_, _26795_);
  and g_36798_(_26668_, _26795_, _26796_);
  or g_36799_(_26670_, _26794_, _26797_);
  and g_36800_(_26626_, _26630_, _26798_);
  or g_36801_(_26624_, _26629_, _26799_);
  and g_36802_(_26646_, _26663_, _26800_);
  or g_36803_(_26648_, _26662_, _26802_);
  and g_36804_(_26799_, _26802_, _26803_);
  or g_36805_(_26798_, _26800_, _26804_);
  and g_36806_(_26797_, _26803_, _26805_);
  or g_36807_(_26796_, _26804_, _26806_);
  or g_36808_(out[208], _26598_, _26807_);
  or g_36809_(_26756_, _26773_, _26808_);
  not g_36810_(_26808_, _26809_);
  and g_36811_(_26668_, _26807_, _26810_);
  not g_36812_(_26810_, _26811_);
  and g_36813_(_26809_, _26810_, _26813_);
  or g_36814_(_26808_, _26811_, _26814_);
  and g_36815_(_26737_, _26813_, _26815_);
  or g_36816_(_26738_, _26814_, _26816_);
  and g_36817_(_26806_, _26816_, _26817_);
  or g_36818_(_26805_, _26815_, _26818_);
  and g_36819_(_26598_, _26818_, _26819_);
  not g_36820_(_26819_, _26820_);
  or g_36821_(out[208], _26818_, _26821_);
  not g_36822_(_26821_, _26822_);
  and g_36823_(_26820_, _26821_, _26824_);
  or g_36824_(_26819_, _26822_, _26825_);
  and g_36825_(out[211], _26817_, _26826_);
  and g_36826_(_26741_, _26818_, _26827_);
  or g_36827_(_26826_, _26827_, _26828_);
  not g_36828_(_26828_, _26829_);
  or g_36829_(_19178_, _26828_, _26830_);
  and g_36830_(_26749_, _26818_, _26831_);
  not g_36831_(_26831_, _26832_);
  or g_36832_(out[210], _26818_, _26833_);
  not g_36833_(_26833_, _09274_);
  and g_36834_(_26832_, _26833_, _09275_);
  or g_36835_(_26831_, _09274_, _09276_);
  or g_36836_(out[227], _26829_, _09277_);
  not g_36837_(_09277_, _09278_);
  or g_36838_(out[226], _09276_, _09279_);
  xor g_36839_(out[227], _26828_, _09280_);
  xor g_36840_(out[226], _09275_, _09281_);
  or g_36841_(_09280_, _09281_, _09282_);
  and g_36842_(_26764_, _26818_, _09283_);
  not g_36843_(_09283_, _09285_);
  or g_36844_(out[209], _26818_, _09286_);
  not g_36845_(_09286_, _09287_);
  and g_36846_(_09285_, _09286_, _09288_);
  or g_36847_(_09283_, _09287_, _09289_);
  or g_36848_(out[225], _09289_, _09290_);
  and g_36849_(out[224], _26825_, _09291_);
  xor g_36850_(out[225], _09288_, _09292_);
  or g_36851_(_09291_, _09292_, _09293_);
  and g_36852_(_09290_, _09293_, _09294_);
  or g_36853_(_09282_, _09294_, _09296_);
  and g_36854_(_26830_, _09279_, _09297_);
  or g_36855_(_09278_, _09297_, _09298_);
  and g_36856_(_09296_, _09298_, _09299_);
  and g_36857_(out[228], out[227], _09300_);
  or g_36858_(out[229], _09300_, _09301_);
  or g_36859_(out[230], _09301_, _09302_);
  or g_36860_(out[231], _09302_, _09303_);
  or g_36861_(out[232], _09303_, _09304_);
  and g_36862_(out[233], _09304_, _09305_);
  or g_36863_(out[234], _09305_, _09307_);
  xor g_36864_(out[234], _09305_, _09308_);
  xor g_36865_(_19211_, _09305_, _09309_);
  and g_36866_(_26613_, _26817_, _09310_);
  or g_36867_(_26615_, _26818_, _09311_);
  and g_36868_(_26621_, _26818_, _09312_);
  or g_36869_(_26620_, _26817_, _09313_);
  and g_36870_(_09311_, _09313_, _09314_);
  or g_36871_(_09310_, _09312_, _09315_);
  and g_36872_(_09308_, _09314_, _09316_);
  or g_36873_(_09309_, _09315_, _09318_);
  and g_36874_(_26599_, _26609_, _09319_);
  or g_36875_(_26600_, _26610_, _09320_);
  xor g_36876_(out[235], _09307_, _09321_);
  xor g_36877_(_19090_, _09307_, _09322_);
  and g_36878_(_09319_, _09322_, _09323_);
  or g_36879_(_09320_, _09321_, _09324_);
  and g_36880_(_09318_, _09324_, _09325_);
  or g_36881_(_09316_, _09323_, _09326_);
  and g_36882_(_09320_, _09321_, _09327_);
  or g_36883_(_09319_, _09322_, _09329_);
  and g_36884_(_09309_, _09315_, _09330_);
  or g_36885_(_09308_, _09314_, _09331_);
  and g_36886_(_09329_, _09331_, _09332_);
  or g_36887_(_09327_, _09330_, _09333_);
  and g_36888_(_26631_, _26817_, _09334_);
  or g_36889_(_26632_, _26818_, _09335_);
  and g_36890_(_26639_, _26818_, _09336_);
  or g_36891_(_26638_, _26817_, _09337_);
  and g_36892_(_09335_, _09337_, _09338_);
  or g_36893_(_09334_, _09336_, _09340_);
  xor g_36894_(out[233], _09304_, _09341_);
  xor g_36895_(_19200_, _09304_, _09342_);
  and g_36896_(_09338_, _09341_, _09343_);
  or g_36897_(_09340_, _09342_, _09344_);
  xor g_36898_(out[232], _09303_, _09345_);
  xor g_36899_(_19189_, _09303_, _09346_);
  and g_36900_(_26652_, _26817_, _09347_);
  or g_36901_(_26651_, _26818_, _09348_);
  and g_36902_(_26659_, _26818_, _09349_);
  or g_36903_(_26657_, _26817_, _09351_);
  and g_36904_(_09348_, _09351_, _09352_);
  or g_36905_(_09347_, _09349_, _09353_);
  and g_36906_(_09345_, _09353_, _09354_);
  or g_36907_(_09346_, _09352_, _09355_);
  and g_36908_(_09340_, _09342_, _09356_);
  or g_36909_(_09338_, _09341_, _09357_);
  and g_36910_(_09355_, _09357_, _09358_);
  or g_36911_(_09354_, _09356_, _09359_);
  and g_36912_(_09346_, _09352_, _09360_);
  or g_36913_(_09345_, _09353_, _09362_);
  and g_36914_(_09325_, _09332_, _09363_);
  or g_36915_(_09326_, _09333_, _09364_);
  and g_36916_(_09344_, _09362_, _09365_);
  or g_36917_(_09343_, _09360_, _09366_);
  and g_36918_(_09358_, _09365_, _09367_);
  or g_36919_(_09359_, _09366_, _09368_);
  and g_36920_(_09363_, _09367_, _09369_);
  or g_36921_(_09364_, _09368_, _09370_);
  xor g_36922_(out[231], _09302_, _09371_);
  xor g_36923_(_19101_, _09302_, _09373_);
  or g_36924_(_26671_, _26818_, _09374_);
  not g_36925_(_09374_, _09375_);
  and g_36926_(_26678_, _26818_, _09376_);
  not g_36927_(_09376_, _09377_);
  and g_36928_(_09374_, _09377_, _09378_);
  or g_36929_(_09375_, _09376_, _09379_);
  and g_36930_(_09371_, _09379_, _09380_);
  or g_36931_(_09373_, _09378_, _09381_);
  xor g_36932_(out[230], _09301_, _09382_);
  xor g_36933_(_19112_, _09301_, _09384_);
  or g_36934_(_26683_, _26818_, _09385_);
  not g_36935_(_09385_, _09386_);
  and g_36936_(_26689_, _26818_, _09387_);
  not g_36937_(_09387_, _09388_);
  and g_36938_(_09385_, _09388_, _09389_);
  or g_36939_(_09386_, _09387_, _09390_);
  and g_36940_(_09382_, _09389_, _09391_);
  or g_36941_(_09384_, _09390_, _09392_);
  and g_36942_(_09381_, _09392_, _09393_);
  or g_36943_(_09380_, _09391_, _09395_);
  and g_36944_(_09384_, _09390_, _09396_);
  or g_36945_(_09382_, _09389_, _09397_);
  and g_36946_(_09373_, _09378_, _09398_);
  or g_36947_(_09371_, _09379_, _09399_);
  and g_36948_(_09397_, _09399_, _09400_);
  or g_36949_(_09396_, _09398_, _09401_);
  and g_36950_(_09393_, _09400_, _09402_);
  or g_36951_(_09395_, _09401_, _09403_);
  xor g_36952_(out[228], out[227], _09404_);
  xor g_36953_(_19134_, out[227], _09406_);
  or g_36954_(_26718_, _26818_, _09407_);
  not g_36955_(_09407_, _09408_);
  and g_36956_(_26725_, _26818_, _09409_);
  not g_36957_(_09409_, _09410_);
  and g_36958_(_09407_, _09410_, _09411_);
  or g_36959_(_09408_, _09409_, _09412_);
  and g_36960_(_09406_, _09412_, _09413_);
  or g_36961_(_09404_, _09411_, _09414_);
  xor g_36962_(out[229], _09300_, _09415_);
  xor g_36963_(_19123_, _09300_, _09417_);
  or g_36964_(_26695_, _26818_, _09418_);
  not g_36965_(_09418_, _09419_);
  and g_36966_(_26703_, _26818_, _09420_);
  not g_36967_(_09420_, _09421_);
  and g_36968_(_09418_, _09421_, _09422_);
  or g_36969_(_09419_, _09420_, _09423_);
  and g_36970_(_09415_, _09423_, _09424_);
  or g_36971_(_09417_, _09422_, _09425_);
  and g_36972_(_09414_, _09425_, _09426_);
  or g_36973_(_09413_, _09424_, _09428_);
  and g_36974_(_09417_, _09422_, _09429_);
  or g_36975_(_09415_, _09423_, _09430_);
  and g_36976_(_09404_, _09411_, _09431_);
  or g_36977_(_09406_, _09412_, _09432_);
  and g_36978_(_09430_, _09432_, _09433_);
  or g_36979_(_09429_, _09431_, _09434_);
  and g_36980_(_09426_, _09433_, _09435_);
  or g_36981_(_09428_, _09434_, _09436_);
  and g_36982_(_09369_, _09435_, _09437_);
  or g_36983_(_09370_, _09436_, _09439_);
  and g_36984_(_09402_, _09437_, _09440_);
  or g_36985_(_09403_, _09439_, _09441_);
  or g_36986_(_09299_, _09441_, _09442_);
  or g_36987_(_09426_, _09429_, _09443_);
  or g_36988_(_09403_, _09443_, _09444_);
  or g_36989_(_09393_, _09398_, _09445_);
  and g_36990_(_09444_, _09445_, _09446_);
  or g_36991_(_09370_, _09446_, _09447_);
  or g_36992_(_09343_, _09358_, _09448_);
  or g_36993_(_09364_, _09448_, _09450_);
  or g_36994_(_09325_, _09327_, _09451_);
  and g_36995_(_09450_, _09451_, _09452_);
  and g_36996_(_09442_, _09452_, _09453_);
  and g_36997_(_09447_, _09453_, _09454_);
  and g_36998_(_19156_, _26824_, _09455_);
  or g_36999_(_09282_, _09455_, _09456_);
  or g_37000_(_09293_, _09456_, _09457_);
  not g_37001_(_09457_, _09458_);
  and g_37002_(_09440_, _09458_, _09459_);
  or g_37003_(_09454_, _09459_, _09461_);
  not g_37004_(_09461_, _09462_);
  and g_37005_(_26825_, _09461_, _09463_);
  or g_37006_(_26824_, _09462_, _09464_);
  or g_37007_(out[224], _09461_, _09465_);
  not g_37008_(_09465_, _09466_);
  and g_37009_(_09464_, _09465_, _09467_);
  or g_37010_(_09463_, _09466_, _09468_);
  and g_37011_(_09319_, _09321_, _09469_);
  or g_37012_(_09320_, _09322_, _09470_);
  and g_37013_(out[244], out[243], _09472_);
  or g_37014_(out[245], _09472_, _09473_);
  or g_37015_(out[246], _09473_, _09474_);
  or g_37016_(out[247], _09474_, _09475_);
  or g_37017_(out[248], _09475_, _09476_);
  and g_37018_(out[249], _09476_, _09477_);
  or g_37019_(out[250], _09477_, _09478_);
  xor g_37020_(out[251], _09478_, _09479_);
  xor g_37021_(_19222_, _09478_, _09480_);
  and g_37022_(_09469_, _09480_, _09481_);
  or g_37023_(_09470_, _09479_, _09483_);
  xor g_37024_(out[250], _09477_, _09484_);
  not g_37025_(_09484_, _09485_);
  and g_37026_(_09308_, _09462_, _09486_);
  or g_37027_(_09309_, _09461_, _09487_);
  and g_37028_(_09315_, _09461_, _09488_);
  or g_37029_(_09314_, _09462_, _09489_);
  and g_37030_(_09487_, _09489_, _09490_);
  or g_37031_(_09486_, _09488_, _09491_);
  and g_37032_(_09484_, _09490_, _09492_);
  or g_37033_(_09485_, _09491_, _09494_);
  and g_37034_(_09483_, _09494_, _09495_);
  or g_37035_(_09481_, _09492_, _09496_);
  and g_37036_(_09485_, _09491_, _09497_);
  or g_37037_(_09484_, _09490_, _09498_);
  and g_37038_(_09470_, _09479_, _09499_);
  or g_37039_(_09469_, _09480_, _09500_);
  and g_37040_(_09341_, _09462_, _09501_);
  or g_37041_(_09342_, _09461_, _09502_);
  and g_37042_(_09340_, _09461_, _09503_);
  or g_37043_(_09338_, _09462_, _09505_);
  and g_37044_(_09502_, _09505_, _09506_);
  or g_37045_(_09501_, _09503_, _09507_);
  xor g_37046_(out[249], _09476_, _09508_);
  not g_37047_(_09508_, _09509_);
  and g_37048_(_09506_, _09508_, _09510_);
  or g_37049_(_09507_, _09509_, _09511_);
  and g_37050_(_09500_, _09511_, _09512_);
  or g_37051_(_09499_, _09510_, _09513_);
  and g_37052_(_09498_, _09512_, _09514_);
  or g_37053_(_09497_, _09513_, _09516_);
  and g_37054_(_09495_, _09514_, _09517_);
  or g_37055_(_09496_, _09516_, _09518_);
  and g_37056_(_09507_, _09509_, _09519_);
  or g_37057_(_09506_, _09508_, _09520_);
  xor g_37058_(out[248], _09475_, _09521_);
  xor g_37059_(_19321_, _09475_, _09522_);
  or g_37060_(_09345_, _09461_, _09523_);
  not g_37061_(_09523_, _09524_);
  and g_37062_(_09353_, _09461_, _09525_);
  or g_37063_(_09352_, _09462_, _09527_);
  and g_37064_(_09523_, _09527_, _09528_);
  or g_37065_(_09524_, _09525_, _09529_);
  and g_37066_(_09521_, _09529_, _09530_);
  or g_37067_(_09522_, _09528_, _09531_);
  and g_37068_(_09520_, _09531_, _09532_);
  or g_37069_(_09519_, _09530_, _09533_);
  and g_37070_(_09522_, _09528_, _09534_);
  or g_37071_(_09521_, _09529_, _09535_);
  and g_37072_(_09532_, _09535_, _09536_);
  or g_37073_(_09533_, _09534_, _09538_);
  and g_37074_(_09517_, _09536_, _09539_);
  or g_37075_(_09518_, _09538_, _09540_);
  xor g_37076_(out[247], _09474_, _09541_);
  not g_37077_(_09541_, _09542_);
  or g_37078_(_09371_, _09461_, _09543_);
  not g_37079_(_09543_, _09544_);
  and g_37080_(_09379_, _09461_, _09545_);
  or g_37081_(_09378_, _09462_, _09546_);
  and g_37082_(_09543_, _09546_, _09547_);
  or g_37083_(_09544_, _09545_, _09549_);
  and g_37084_(_09541_, _09549_, _09550_);
  xor g_37085_(out[246], _09473_, _09551_);
  not g_37086_(_09551_, _09552_);
  and g_37087_(_09382_, _09462_, _09553_);
  or g_37088_(_09384_, _09461_, _09554_);
  and g_37089_(_09390_, _09461_, _09555_);
  or g_37090_(_09389_, _09462_, _09556_);
  and g_37091_(_09554_, _09556_, _09557_);
  or g_37092_(_09553_, _09555_, _09558_);
  and g_37093_(_09551_, _09557_, _09560_);
  or g_37094_(_09550_, _09560_, _09561_);
  and g_37095_(_09542_, _09547_, _09562_);
  or g_37096_(_09541_, _09549_, _09563_);
  and g_37097_(_09552_, _09558_, _09564_);
  or g_37098_(_09562_, _09564_, _09565_);
  xor g_37099_(_09542_, _09547_, _09566_);
  xor g_37100_(_09551_, _09557_, _09567_);
  and g_37101_(_09566_, _09567_, _09568_);
  or g_37102_(_09561_, _09565_, _09569_);
  xor g_37103_(out[245], _09472_, _09571_);
  xor g_37104_(_19255_, _09472_, _09572_);
  or g_37105_(_09415_, _09461_, _09573_);
  not g_37106_(_09573_, _09574_);
  and g_37107_(_09423_, _09461_, _09575_);
  or g_37108_(_09422_, _09462_, _09576_);
  and g_37109_(_09573_, _09576_, _09577_);
  or g_37110_(_09574_, _09575_, _09578_);
  and g_37111_(_09571_, _09578_, _09579_);
  or g_37112_(_09572_, _09577_, _09580_);
  xor g_37113_(out[244], out[243], _09582_);
  not g_37114_(_09582_, _09583_);
  and g_37115_(_09404_, _09462_, _09584_);
  or g_37116_(_09406_, _09461_, _09585_);
  and g_37117_(_09412_, _09461_, _09586_);
  or g_37118_(_09411_, _09462_, _09587_);
  and g_37119_(_09585_, _09587_, _09588_);
  or g_37120_(_09584_, _09586_, _09589_);
  and g_37121_(_09583_, _09589_, _09590_);
  or g_37122_(_09582_, _09588_, _09591_);
  and g_37123_(_09580_, _09591_, _09593_);
  or g_37124_(_09579_, _09590_, _09594_);
  and g_37125_(_09572_, _09577_, _09595_);
  or g_37126_(_09571_, _09578_, _09596_);
  and g_37127_(_09582_, _09588_, _09597_);
  or g_37128_(_09583_, _09589_, _09598_);
  and g_37129_(_09596_, _09598_, _09599_);
  or g_37130_(_09595_, _09597_, _09600_);
  and g_37131_(_09593_, _09599_, _09601_);
  or g_37132_(_09594_, _09600_, _09602_);
  and g_37133_(_09568_, _09601_, _09604_);
  or g_37134_(_09569_, _09602_, _09605_);
  and g_37135_(_09539_, _09604_, _09606_);
  or g_37136_(_09540_, _09605_, _09607_);
  and g_37137_(out[227], _09462_, _09608_);
  or g_37138_(_19178_, _09461_, _09609_);
  and g_37139_(_26828_, _09461_, _09610_);
  not g_37140_(_09610_, _09611_);
  and g_37141_(_09609_, _09611_, _09612_);
  or g_37142_(_09608_, _09610_, _09613_);
  and g_37143_(out[243], _09612_, _09615_);
  or g_37144_(_19310_, _09613_, _09616_);
  or g_37145_(_09275_, _09462_, _09617_);
  or g_37146_(out[226], _09461_, _09618_);
  and g_37147_(_09617_, _09618_, _09619_);
  not g_37148_(_09619_, _09620_);
  and g_37149_(out[242], _09620_, _09621_);
  or g_37150_(_19299_, _09619_, _09622_);
  and g_37151_(_09616_, _09622_, _09623_);
  or g_37152_(_09615_, _09621_, _09624_);
  and g_37153_(_19310_, _09613_, _09626_);
  or g_37154_(out[243], _09612_, _09627_);
  and g_37155_(_19299_, _09619_, _09628_);
  or g_37156_(out[242], _09620_, _09629_);
  and g_37157_(_09627_, _09629_, _09630_);
  or g_37158_(_09626_, _09628_, _09631_);
  and g_37159_(_09623_, _09630_, _09632_);
  or g_37160_(_09624_, _09631_, _09633_);
  and g_37161_(_09289_, _09461_, _09634_);
  or g_37162_(_09288_, _09462_, _09635_);
  or g_37163_(out[225], _09461_, _09637_);
  not g_37164_(_09637_, _09638_);
  and g_37165_(_09635_, _09637_, _09639_);
  or g_37166_(_09634_, _09638_, _09640_);
  and g_37167_(_19277_, _09639_, _09641_);
  or g_37168_(out[241], _09640_, _09642_);
  and g_37169_(out[240], _09468_, _09643_);
  or g_37170_(_19288_, _09467_, _09644_);
  xor g_37171_(_19277_, _09639_, _09645_);
  xor g_37172_(out[241], _09639_, _09646_);
  and g_37173_(_09644_, _09645_, _09648_);
  or g_37174_(_09643_, _09646_, _09649_);
  and g_37175_(_09642_, _09649_, _09650_);
  or g_37176_(_09641_, _09648_, _09651_);
  and g_37177_(_09632_, _09651_, _09652_);
  or g_37178_(_09633_, _09650_, _09653_);
  and g_37179_(_09627_, _09628_, _09654_);
  or g_37180_(_09626_, _09629_, _09655_);
  and g_37181_(_09616_, _09655_, _09656_);
  or g_37182_(_09615_, _09654_, _09657_);
  and g_37183_(_09653_, _09656_, _09659_);
  or g_37184_(_09652_, _09657_, _09660_);
  and g_37185_(_09606_, _09660_, _09661_);
  or g_37186_(_09607_, _09659_, _09662_);
  and g_37187_(_09517_, _09533_, _09663_);
  or g_37188_(_09518_, _09532_, _09664_);
  and g_37189_(_09496_, _09500_, _09665_);
  or g_37190_(_09495_, _09499_, _09666_);
  and g_37191_(_09664_, _09666_, _09667_);
  or g_37192_(_09663_, _09665_, _09668_);
  and g_37193_(_09561_, _09563_, _09670_);
  not g_37194_(_09670_, _09671_);
  or g_37195_(_09593_, _09595_, _09672_);
  and g_37196_(_09568_, _09594_, _09673_);
  and g_37197_(_09596_, _09673_, _09674_);
  or g_37198_(_09569_, _09672_, _09675_);
  and g_37199_(_09671_, _09675_, _09676_);
  or g_37200_(_09670_, _09674_, _09677_);
  and g_37201_(_09539_, _09677_, _09678_);
  or g_37202_(_09540_, _09676_, _09679_);
  or g_37203_(_09668_, _09678_, _09681_);
  and g_37204_(_09662_, _09679_, _09682_);
  and g_37205_(_09667_, _09682_, _09683_);
  or g_37206_(_09661_, _09681_, _09684_);
  and g_37207_(_19288_, _09467_, _09685_);
  or g_37208_(out[240], _09468_, _09686_);
  and g_37209_(_09632_, _09686_, _09687_);
  or g_37210_(_09633_, _09685_, _09688_);
  and g_37211_(_09648_, _09687_, _09689_);
  or g_37212_(_09649_, _09688_, _09690_);
  and g_37213_(_09606_, _09689_, _09692_);
  or g_37214_(_09607_, _09690_, _09693_);
  and g_37215_(_09684_, _09693_, _09694_);
  or g_37216_(_09683_, _09692_, _09695_);
  and g_37217_(_09468_, _09695_, _09696_);
  or g_37218_(_09467_, _09694_, _09697_);
  and g_37219_(_19288_, _09694_, _09698_);
  not g_37220_(_09698_, _09699_);
  and g_37221_(_09697_, _09699_, _09700_);
  or g_37222_(_09696_, _09698_, _09701_);
  and g_37223_(out[243], _09694_, _09703_);
  and g_37224_(_09613_, _09695_, _09704_);
  or g_37225_(_09703_, _09704_, _09705_);
  or g_37226_(_19442_, _09705_, _09706_);
  and g_37227_(_09620_, _09695_, _09707_);
  and g_37228_(_19299_, _09694_, _09708_);
  or g_37229_(_09707_, _09708_, _09709_);
  and g_37230_(_19442_, _09705_, _09710_);
  or g_37231_(out[258], _09709_, _09711_);
  xor g_37232_(out[259], _09705_, _09712_);
  xor g_37233_(_19431_, _09709_, _09714_);
  or g_37234_(_09712_, _09714_, _09715_);
  and g_37235_(_09640_, _09695_, _09716_);
  and g_37236_(_19277_, _09694_, _09717_);
  or g_37237_(_09716_, _09717_, _09718_);
  or g_37238_(out[257], _09718_, _09719_);
  and g_37239_(out[256], _09701_, _09720_);
  xor g_37240_(_19409_, _09718_, _09721_);
  or g_37241_(_09720_, _09721_, _09722_);
  and g_37242_(_09719_, _09722_, _09723_);
  or g_37243_(_09715_, _09723_, _09725_);
  or g_37244_(_09710_, _09711_, _09726_);
  and g_37245_(_09706_, _09726_, _09727_);
  and g_37246_(_09725_, _09727_, _09728_);
  not g_37247_(_09728_, _09729_);
  and g_37248_(_09469_, _09479_, _09730_);
  or g_37249_(_09470_, _09480_, _09731_);
  and g_37250_(out[260], out[259], _09732_);
  or g_37251_(out[261], _09732_, _09733_);
  or g_37252_(out[262], _09733_, _09734_);
  or g_37253_(out[263], _09734_, _09736_);
  or g_37254_(out[264], _09736_, _09737_);
  and g_37255_(out[265], _09737_, _09738_);
  or g_37256_(out[266], _09738_, _09739_);
  xor g_37257_(out[267], _09739_, _09740_);
  xor g_37258_(_19354_, _09739_, _09741_);
  and g_37259_(_09730_, _09741_, _09742_);
  or g_37260_(_09731_, _09740_, _09743_);
  xor g_37261_(out[266], _09738_, _09744_);
  xor g_37262_(_19475_, _09738_, _09745_);
  and g_37263_(_09484_, _09694_, _09747_);
  or g_37264_(_09485_, _09695_, _09748_);
  and g_37265_(_09491_, _09695_, _09749_);
  or g_37266_(_09490_, _09694_, _09750_);
  and g_37267_(_09748_, _09750_, _09751_);
  or g_37268_(_09747_, _09749_, _09752_);
  and g_37269_(_09744_, _09751_, _09753_);
  or g_37270_(_09745_, _09752_, _09754_);
  and g_37271_(_09743_, _09754_, _09755_);
  or g_37272_(_09742_, _09753_, _09756_);
  and g_37273_(_09731_, _09740_, _09758_);
  or g_37274_(_09730_, _09741_, _09759_);
  and g_37275_(_09745_, _09752_, _09760_);
  or g_37276_(_09744_, _09751_, _09761_);
  and g_37277_(_09759_, _09761_, _09762_);
  or g_37278_(_09758_, _09760_, _09763_);
  and g_37279_(_09755_, _09762_, _09764_);
  or g_37280_(_09756_, _09763_, _09765_);
  xor g_37281_(out[264], _09736_, _09766_);
  xor g_37282_(_19453_, _09736_, _09767_);
  and g_37283_(_09522_, _09694_, _09769_);
  not g_37284_(_09769_, _09770_);
  or g_37285_(_09528_, _09694_, _09771_);
  not g_37286_(_09771_, _09772_);
  and g_37287_(_09770_, _09771_, _09773_);
  or g_37288_(_09769_, _09772_, _09774_);
  and g_37289_(_09766_, _09774_, _09775_);
  or g_37290_(_09767_, _09773_, _09776_);
  and g_37291_(_09508_, _09694_, _09777_);
  not g_37292_(_09777_, _09778_);
  or g_37293_(_09506_, _09694_, _09780_);
  not g_37294_(_09780_, _09781_);
  and g_37295_(_09778_, _09780_, _09782_);
  or g_37296_(_09777_, _09781_, _09783_);
  xor g_37297_(out[265], _09737_, _09784_);
  xor g_37298_(_19464_, _09737_, _09785_);
  and g_37299_(_09783_, _09785_, _09786_);
  or g_37300_(_09782_, _09784_, _09787_);
  and g_37301_(_09776_, _09787_, _09788_);
  or g_37302_(_09775_, _09786_, _09789_);
  and g_37303_(_09782_, _09784_, _09791_);
  or g_37304_(_09783_, _09785_, _09792_);
  and g_37305_(_09767_, _09773_, _09793_);
  or g_37306_(_09766_, _09774_, _09794_);
  and g_37307_(_09792_, _09794_, _09795_);
  or g_37308_(_09791_, _09793_, _09796_);
  and g_37309_(_09788_, _09795_, _09797_);
  or g_37310_(_09789_, _09796_, _09798_);
  and g_37311_(_09764_, _09797_, _09799_);
  or g_37312_(_09765_, _09798_, _09800_);
  xor g_37313_(out[262], _09733_, _09802_);
  xor g_37314_(_19376_, _09733_, _09803_);
  and g_37315_(_09551_, _09694_, _09804_);
  or g_37316_(_09552_, _09695_, _09805_);
  and g_37317_(_09558_, _09695_, _09806_);
  or g_37318_(_09557_, _09694_, _09807_);
  and g_37319_(_09805_, _09807_, _09808_);
  or g_37320_(_09804_, _09806_, _09809_);
  and g_37321_(_09802_, _09808_, _09810_);
  or g_37322_(_09803_, _09809_, _09811_);
  xor g_37323_(out[263], _09734_, _09813_);
  not g_37324_(_09813_, _09814_);
  and g_37325_(_09542_, _09694_, _09815_);
  or g_37326_(_09541_, _09695_, _09816_);
  and g_37327_(_09549_, _09695_, _09817_);
  or g_37328_(_09547_, _09694_, _09818_);
  and g_37329_(_09816_, _09818_, _09819_);
  or g_37330_(_09815_, _09817_, _09820_);
  and g_37331_(_09813_, _09820_, _09821_);
  or g_37332_(_09814_, _09819_, _09822_);
  and g_37333_(_09811_, _09822_, _09824_);
  or g_37334_(_09810_, _09821_, _09825_);
  and g_37335_(_09814_, _09819_, _09826_);
  or g_37336_(_09813_, _09820_, _09827_);
  and g_37337_(_09803_, _09809_, _09828_);
  or g_37338_(_09802_, _09808_, _09829_);
  and g_37339_(_09827_, _09829_, _09830_);
  or g_37340_(_09826_, _09828_, _09831_);
  and g_37341_(_09824_, _09830_, _09832_);
  or g_37342_(_09825_, _09831_, _09833_);
  xor g_37343_(out[260], out[259], _09835_);
  xor g_37344_(_19398_, out[259], _09836_);
  and g_37345_(_09582_, _09694_, _09837_);
  not g_37346_(_09837_, _09838_);
  or g_37347_(_09588_, _09694_, _09839_);
  not g_37348_(_09839_, _09840_);
  and g_37349_(_09838_, _09839_, _09841_);
  or g_37350_(_09837_, _09840_, _09842_);
  and g_37351_(_09836_, _09842_, _09843_);
  or g_37352_(_09835_, _09841_, _09844_);
  xor g_37353_(out[261], _09732_, _09846_);
  xor g_37354_(_19387_, _09732_, _09847_);
  and g_37355_(_09572_, _09694_, _09848_);
  not g_37356_(_09848_, _09849_);
  or g_37357_(_09577_, _09694_, _09850_);
  not g_37358_(_09850_, _09851_);
  and g_37359_(_09849_, _09850_, _09852_);
  or g_37360_(_09848_, _09851_, _09853_);
  and g_37361_(_09846_, _09853_, _09854_);
  or g_37362_(_09847_, _09852_, _09855_);
  and g_37363_(_09844_, _09855_, _09857_);
  or g_37364_(_09843_, _09854_, _09858_);
  and g_37365_(_09847_, _09852_, _09859_);
  or g_37366_(_09846_, _09853_, _09860_);
  and g_37367_(_09835_, _09841_, _09861_);
  or g_37368_(_09836_, _09842_, _09862_);
  and g_37369_(_09860_, _09862_, _09863_);
  or g_37370_(_09859_, _09861_, _09864_);
  and g_37371_(_09857_, _09863_, _09865_);
  or g_37372_(_09858_, _09864_, _09866_);
  and g_37373_(_09832_, _09865_, _09868_);
  or g_37374_(_09833_, _09866_, _09869_);
  and g_37375_(_09799_, _09868_, _09870_);
  or g_37376_(_09800_, _09869_, _09871_);
  and g_37377_(_09729_, _09870_, _09872_);
  or g_37378_(_09728_, _09871_, _09873_);
  and g_37379_(_09756_, _09759_, _09874_);
  or g_37380_(_09755_, _09758_, _09875_);
  and g_37381_(_09789_, _09792_, _09876_);
  or g_37382_(_09788_, _09791_, _09877_);
  and g_37383_(_09764_, _09876_, _09879_);
  or g_37384_(_09765_, _09877_, _09880_);
  and g_37385_(_09875_, _09880_, _09881_);
  or g_37386_(_09874_, _09879_, _09882_);
  and g_37387_(_09825_, _09827_, _09883_);
  or g_37388_(_09824_, _09826_, _09884_);
  and g_37389_(_09858_, _09860_, _09885_);
  or g_37390_(_09857_, _09859_, _09886_);
  and g_37391_(_09832_, _09885_, _09887_);
  or g_37392_(_09833_, _09886_, _09888_);
  and g_37393_(_09884_, _09888_, _09890_);
  or g_37394_(_09883_, _09887_, _09891_);
  and g_37395_(_09799_, _09891_, _09892_);
  or g_37396_(_09800_, _09890_, _09893_);
  or g_37397_(_09882_, _09892_, _09894_);
  and g_37398_(_09873_, _09881_, _09895_);
  and g_37399_(_09893_, _09895_, _09896_);
  or g_37400_(_09872_, _09894_, _09897_);
  and g_37401_(_19420_, _09700_, _09898_);
  or g_37402_(_09715_, _09722_, _09899_);
  or g_37403_(_09898_, _09899_, _09901_);
  or g_37404_(_09871_, _09901_, _09902_);
  not g_37405_(_09902_, _09903_);
  and g_37406_(_09897_, _09902_, _09904_);
  or g_37407_(_09896_, _09903_, _09905_);
  and g_37408_(_09701_, _09905_, _09906_);
  not g_37409_(_09906_, _09907_);
  or g_37410_(out[256], _09905_, _09908_);
  not g_37411_(_09908_, _09909_);
  and g_37412_(_09907_, _09908_, _09910_);
  or g_37413_(_09906_, _09909_, _09912_);
  and g_37414_(out[276], out[275], _09913_);
  or g_37415_(out[277], _09913_, _09914_);
  or g_37416_(out[278], _09914_, _09915_);
  or g_37417_(out[279], _09915_, _09916_);
  or g_37418_(out[280], _09916_, _09917_);
  and g_37419_(out[281], _09917_, _09918_);
  or g_37420_(out[282], _09918_, _09919_);
  xor g_37421_(out[282], _09918_, _09920_);
  xor g_37422_(_19607_, _09918_, _09921_);
  and g_37423_(_09744_, _09904_, _09923_);
  or g_37424_(_09745_, _09905_, _09924_);
  and g_37425_(_09752_, _09905_, _09925_);
  or g_37426_(_09751_, _09904_, _09926_);
  and g_37427_(_09924_, _09926_, _09927_);
  or g_37428_(_09923_, _09925_, _09928_);
  and g_37429_(_09920_, _09927_, _09929_);
  or g_37430_(_09921_, _09928_, _09930_);
  and g_37431_(_09730_, _09740_, _09931_);
  or g_37432_(_09731_, _09741_, _09932_);
  xor g_37433_(out[283], _09919_, _09934_);
  xor g_37434_(_19486_, _09919_, _09935_);
  and g_37435_(_09931_, _09935_, _09936_);
  or g_37436_(_09932_, _09934_, _09937_);
  and g_37437_(_09930_, _09937_, _09938_);
  or g_37438_(_09929_, _09936_, _09939_);
  and g_37439_(_09921_, _09928_, _09940_);
  or g_37440_(_09920_, _09927_, _09941_);
  and g_37441_(_09932_, _09934_, _09942_);
  or g_37442_(_09931_, _09935_, _09943_);
  and g_37443_(_09941_, _09943_, _09945_);
  or g_37444_(_09940_, _09942_, _09946_);
  and g_37445_(_09938_, _09945_, _09947_);
  or g_37446_(_09939_, _09946_, _09948_);
  and g_37447_(_09784_, _09904_, _09949_);
  or g_37448_(_09785_, _09905_, _09950_);
  and g_37449_(_09783_, _09905_, _09951_);
  or g_37450_(_09782_, _09904_, _09952_);
  and g_37451_(_09950_, _09952_, _09953_);
  or g_37452_(_09949_, _09951_, _09954_);
  xor g_37453_(out[281], _09917_, _09956_);
  xor g_37454_(_19596_, _09917_, _09957_);
  and g_37455_(_09954_, _09957_, _09958_);
  or g_37456_(_09953_, _09956_, _09959_);
  xor g_37457_(out[280], _09916_, _09960_);
  xor g_37458_(_19585_, _09916_, _09961_);
  and g_37459_(_09767_, _09904_, _09962_);
  or g_37460_(_09766_, _09905_, _09963_);
  and g_37461_(_09774_, _09905_, _09964_);
  or g_37462_(_09773_, _09904_, _09965_);
  and g_37463_(_09963_, _09965_, _09967_);
  or g_37464_(_09962_, _09964_, _09968_);
  and g_37465_(_09960_, _09968_, _09969_);
  or g_37466_(_09961_, _09967_, _09970_);
  and g_37467_(_09959_, _09970_, _09971_);
  or g_37468_(_09958_, _09969_, _09972_);
  and g_37469_(_09953_, _09956_, _09973_);
  or g_37470_(_09954_, _09957_, _09974_);
  and g_37471_(_09961_, _09967_, _09975_);
  or g_37472_(_09960_, _09968_, _09976_);
  and g_37473_(_09974_, _09976_, _09978_);
  or g_37474_(_09973_, _09975_, _09979_);
  and g_37475_(_09971_, _09978_, _09980_);
  or g_37476_(_09972_, _09979_, _09981_);
  and g_37477_(_09947_, _09980_, _09982_);
  or g_37478_(_09948_, _09981_, _09983_);
  xor g_37479_(out[279], _09915_, _09984_);
  not g_37480_(_09984_, _09985_);
  or g_37481_(_09813_, _09905_, _09986_);
  not g_37482_(_09986_, _09987_);
  and g_37483_(_09820_, _09905_, _09989_);
  not g_37484_(_09989_, _09990_);
  and g_37485_(_09986_, _09990_, _09991_);
  or g_37486_(_09987_, _09989_, _09992_);
  and g_37487_(_09984_, _09992_, _09993_);
  or g_37488_(_09985_, _09991_, _09994_);
  xor g_37489_(out[278], _09914_, _09995_);
  xor g_37490_(_19508_, _09914_, _09996_);
  or g_37491_(_09803_, _09905_, _09997_);
  not g_37492_(_09997_, _09998_);
  and g_37493_(_09809_, _09905_, _10000_);
  not g_37494_(_10000_, _10001_);
  and g_37495_(_09997_, _10001_, _10002_);
  or g_37496_(_09998_, _10000_, _10003_);
  and g_37497_(_09995_, _10002_, _10004_);
  or g_37498_(_09996_, _10003_, _10005_);
  and g_37499_(_09994_, _10005_, _10006_);
  or g_37500_(_09993_, _10004_, _10007_);
  xor g_37501_(out[277], _09913_, _10008_);
  xor g_37502_(_19519_, _09913_, _10009_);
  and g_37503_(_09847_, _09904_, _10011_);
  or g_37504_(_09846_, _09905_, _10012_);
  and g_37505_(_09853_, _09905_, _10013_);
  or g_37506_(_09852_, _09904_, _10014_);
  and g_37507_(_10012_, _10014_, _10015_);
  or g_37508_(_10011_, _10013_, _10016_);
  and g_37509_(_10008_, _10016_, _10017_);
  or g_37510_(_10009_, _10015_, _10018_);
  xor g_37511_(out[276], out[275], _10019_);
  xor g_37512_(_19530_, out[275], _10020_);
  and g_37513_(_09835_, _09904_, _10022_);
  or g_37514_(_09836_, _09905_, _10023_);
  and g_37515_(_09842_, _09905_, _10024_);
  or g_37516_(_09841_, _09904_, _10025_);
  and g_37517_(_10023_, _10025_, _10026_);
  or g_37518_(_10022_, _10024_, _10027_);
  and g_37519_(_10020_, _10027_, _10028_);
  or g_37520_(_10019_, _10026_, _10029_);
  and g_37521_(_10018_, _10029_, _10030_);
  or g_37522_(_10017_, _10028_, _10031_);
  and g_37523_(_09996_, _10003_, _10033_);
  not g_37524_(_10033_, _10034_);
  or g_37525_(_10008_, _10016_, _10035_);
  not g_37526_(_10035_, _10036_);
  or g_37527_(_09984_, _09992_, _10037_);
  not g_37528_(_10037_, _10038_);
  or g_37529_(_10020_, _10027_, _10039_);
  not g_37530_(_10039_, _10040_);
  and g_37531_(_10006_, _10034_, _10041_);
  or g_37532_(_10007_, _10033_, _10042_);
  and g_37533_(_10037_, _10041_, _10044_);
  or g_37534_(_10038_, _10042_, _10045_);
  and g_37535_(_10030_, _10035_, _10046_);
  or g_37536_(_10031_, _10036_, _10047_);
  and g_37537_(_10039_, _10046_, _10048_);
  or g_37538_(_10040_, _10047_, _10049_);
  and g_37539_(_09982_, _10048_, _10050_);
  or g_37540_(_09983_, _10049_, _10051_);
  and g_37541_(_10044_, _10050_, _10052_);
  or g_37542_(_10045_, _10051_, _10053_);
  or g_37543_(_19442_, _09905_, _10055_);
  not g_37544_(_10055_, _10056_);
  and g_37545_(_09705_, _09905_, _10057_);
  not g_37546_(_10057_, _10058_);
  and g_37547_(_10055_, _10058_, _10059_);
  or g_37548_(_10056_, _10057_, _10060_);
  and g_37549_(out[275], _10059_, _10061_);
  or g_37550_(_19574_, _10060_, _10062_);
  and g_37551_(_09709_, _09905_, _10063_);
  and g_37552_(_19431_, _09904_, _10064_);
  or g_37553_(_10063_, _10064_, _10066_);
  not g_37554_(_10066_, _10067_);
  or g_37555_(_19563_, _10067_, _10068_);
  and g_37556_(_10062_, _10068_, _10069_);
  and g_37557_(_19574_, _10060_, _10070_);
  or g_37558_(out[275], _10059_, _10071_);
  or g_37559_(out[274], _10066_, _10072_);
  not g_37560_(_10072_, _10073_);
  and g_37561_(_10071_, _10072_, _10074_);
  or g_37562_(_10061_, _10070_, _10075_);
  xor g_37563_(_19563_, _10066_, _10077_);
  and g_37564_(_10069_, _10074_, _10078_);
  or g_37565_(_10075_, _10077_, _10079_);
  and g_37566_(_09718_, _09905_, _10080_);
  and g_37567_(_19409_, _09904_, _10081_);
  or g_37568_(_10080_, _10081_, _10082_);
  or g_37569_(out[273], _10082_, _10083_);
  not g_37570_(_10083_, _10084_);
  and g_37571_(out[272], _09912_, _10085_);
  or g_37572_(_19552_, _09910_, _10086_);
  xor g_37573_(out[273], _10082_, _10088_);
  xor g_37574_(_19541_, _10082_, _10089_);
  and g_37575_(_10086_, _10088_, _10090_);
  or g_37576_(_10085_, _10089_, _10091_);
  and g_37577_(_10083_, _10091_, _10092_);
  or g_37578_(_10084_, _10090_, _10093_);
  and g_37579_(_10078_, _10093_, _10094_);
  or g_37580_(_10079_, _10092_, _10095_);
  and g_37581_(_10071_, _10073_, _10096_);
  or g_37582_(_10070_, _10072_, _10097_);
  and g_37583_(_10062_, _10097_, _10099_);
  or g_37584_(_10061_, _10096_, _10100_);
  and g_37585_(_10095_, _10099_, _10101_);
  or g_37586_(_10094_, _10100_, _10102_);
  and g_37587_(_10052_, _10102_, _10103_);
  or g_37588_(_10053_, _10101_, _10104_);
  and g_37589_(_10031_, _10035_, _10105_);
  not g_37590_(_10105_, _10106_);
  or g_37591_(_10033_, _10106_, _10107_);
  and g_37592_(_10006_, _10107_, _10108_);
  or g_37593_(_09983_, _10038_, _10110_);
  or g_37594_(_10108_, _10110_, _10111_);
  not g_37595_(_10111_, _10112_);
  or g_37596_(_09938_, _09942_, _10113_);
  and g_37597_(_09972_, _09974_, _10114_);
  not g_37598_(_10114_, _10115_);
  or g_37599_(_09948_, _10115_, _10116_);
  and g_37600_(_10113_, _10116_, _10117_);
  not g_37601_(_10117_, _10118_);
  and g_37602_(_10104_, _10117_, _10119_);
  or g_37603_(_10103_, _10118_, _10121_);
  and g_37604_(_10111_, _10119_, _10122_);
  or g_37605_(_10112_, _10121_, _10123_);
  or g_37606_(out[272], _09912_, _10124_);
  not g_37607_(_10124_, _10125_);
  or g_37608_(_10079_, _10091_, _10126_);
  or g_37609_(_10125_, _10126_, _10127_);
  or g_37610_(_10053_, _10127_, _10128_);
  not g_37611_(_10128_, _10129_);
  and g_37612_(_10123_, _10128_, _10130_);
  or g_37613_(_10122_, _10129_, _10132_);
  or g_37614_(_09910_, _10130_, _10133_);
  or g_37615_(out[272], _10132_, _10134_);
  and g_37616_(_10133_, _10134_, _10135_);
  not g_37617_(_10135_, _10136_);
  and g_37618_(_09931_, _09934_, _10137_);
  not g_37619_(_10137_, _10138_);
  and g_37620_(out[292], out[291], _10139_);
  or g_37621_(out[293], _10139_, _10140_);
  or g_37622_(out[294], _10140_, _10141_);
  or g_37623_(out[295], _10141_, _10143_);
  or g_37624_(out[296], _10143_, _10144_);
  and g_37625_(out[297], _10144_, _10145_);
  or g_37626_(out[298], _10145_, _10146_);
  xor g_37627_(out[299], _10146_, _10147_);
  and g_37628_(_10138_, _10147_, _10148_);
  or g_37629_(_10138_, _10147_, _10149_);
  xor g_37630_(out[298], _10145_, _10150_);
  not g_37631_(_10150_, _10151_);
  and g_37632_(_09920_, _10130_, _10152_);
  and g_37633_(_09928_, _10132_, _10154_);
  or g_37634_(_10152_, _10154_, _10155_);
  not g_37635_(_10155_, _10156_);
  and g_37636_(_10150_, _10156_, _10157_);
  or g_37637_(_10151_, _10155_, _10158_);
  and g_37638_(_10149_, _10158_, _10159_);
  or g_37639_(_10148_, _10159_, _10160_);
  xor g_37640_(out[296], _10143_, _10161_);
  not g_37641_(_10161_, _10162_);
  and g_37642_(_09960_, _10130_, _10163_);
  and g_37643_(_09967_, _10132_, _10165_);
  or g_37644_(_10163_, _10165_, _10166_);
  not g_37645_(_10166_, _10167_);
  and g_37646_(_10161_, _10167_, _10168_);
  or g_37647_(_10162_, _10166_, _10169_);
  or g_37648_(_09957_, _10132_, _10170_);
  not g_37649_(_10170_, _10171_);
  and g_37650_(_09954_, _10132_, _10172_);
  not g_37651_(_10172_, _10173_);
  and g_37652_(_10170_, _10173_, _10174_);
  or g_37653_(_10171_, _10172_, _10176_);
  xor g_37654_(out[297], _10144_, _10177_);
  xor g_37655_(_19717_, _10144_, _10178_);
  and g_37656_(_10176_, _10178_, _10179_);
  or g_37657_(_10174_, _10177_, _10180_);
  and g_37658_(_10169_, _10180_, _10181_);
  or g_37659_(_10168_, _10179_, _10182_);
  xor g_37660_(out[294], _10140_, _10183_);
  or g_37661_(_09996_, _10132_, _10184_);
  or g_37662_(_10002_, _10130_, _10185_);
  and g_37663_(_10184_, _10185_, _10187_);
  and g_37664_(_10183_, _10187_, _10188_);
  xor g_37665_(out[295], _10141_, _10189_);
  or g_37666_(_09984_, _10132_, _10190_);
  not g_37667_(_10190_, _10191_);
  and g_37668_(_09992_, _10132_, _10192_);
  not g_37669_(_10192_, _10193_);
  and g_37670_(_10190_, _10193_, _10194_);
  or g_37671_(_10191_, _10192_, _10195_);
  and g_37672_(_10189_, _10195_, _10196_);
  or g_37673_(_10188_, _10196_, _10198_);
  or g_37674_(_10189_, _10195_, _10199_);
  or g_37675_(_10008_, _10132_, _10200_);
  not g_37676_(_10200_, _10201_);
  and g_37677_(_10016_, _10132_, _10202_);
  not g_37678_(_10202_, _10203_);
  and g_37679_(_10200_, _10203_, _10204_);
  or g_37680_(_10201_, _10202_, _10205_);
  xor g_37681_(out[293], _10139_, _10206_);
  or g_37682_(_10205_, _10206_, _10207_);
  xor g_37683_(_10183_, _10187_, _10209_);
  xor g_37684_(_10189_, _10195_, _10210_);
  and g_37685_(_10209_, _10210_, _10211_);
  and g_37686_(_10207_, _10211_, _10212_);
  not g_37687_(_10212_, _10213_);
  xor g_37688_(out[292], out[291], _10214_);
  not g_37689_(_10214_, _10215_);
  or g_37690_(_10020_, _10132_, _10216_);
  not g_37691_(_10216_, _10217_);
  and g_37692_(_10027_, _10132_, _10218_);
  not g_37693_(_10218_, _10220_);
  and g_37694_(_10216_, _10220_, _10221_);
  or g_37695_(_10217_, _10218_, _10222_);
  and g_37696_(_10215_, _10222_, _10223_);
  and g_37697_(_10205_, _10206_, _10224_);
  or g_37698_(_10223_, _10224_, _10225_);
  and g_37699_(_10214_, _10221_, _10226_);
  or g_37700_(_10225_, _10226_, _10227_);
  or g_37701_(_10213_, _10227_, _10228_);
  and g_37702_(out[275], _10130_, _10229_);
  and g_37703_(_10060_, _10132_, _10231_);
  or g_37704_(_10229_, _10231_, _10232_);
  or g_37705_(_19695_, _10232_, _10233_);
  and g_37706_(_10066_, _10132_, _10234_);
  and g_37707_(_19563_, _10130_, _10235_);
  or g_37708_(_10234_, _10235_, _10236_);
  or g_37709_(out[290], _10236_, _10237_);
  and g_37710_(_19695_, _10232_, _10238_);
  xor g_37711_(out[291], _10232_, _10239_);
  xor g_37712_(_19684_, _10236_, _10240_);
  or g_37713_(_10239_, _10240_, _10242_);
  and g_37714_(_10082_, _10132_, _10243_);
  and g_37715_(_19541_, _10130_, _10244_);
  or g_37716_(_10243_, _10244_, _10245_);
  or g_37717_(out[289], _10245_, _10246_);
  and g_37718_(out[288], _10136_, _10247_);
  xor g_37719_(_19673_, _10245_, _10248_);
  or g_37720_(_10247_, _10248_, _10249_);
  or g_37721_(_10242_, _10249_, _10250_);
  or g_37722_(_10237_, _10238_, _10251_);
  and g_37723_(_10233_, _10251_, _10253_);
  or g_37724_(_10242_, _10246_, _10254_);
  and g_37725_(_10253_, _10254_, _10255_);
  and g_37726_(_10250_, _10255_, _10256_);
  or g_37727_(_10228_, _10256_, _10257_);
  and g_37728_(_10212_, _10225_, _10258_);
  and g_37729_(_10198_, _10199_, _10259_);
  or g_37730_(_10258_, _10259_, _10260_);
  not g_37731_(_10260_, _10261_);
  and g_37732_(_10257_, _10261_, _10262_);
  and g_37733_(_10162_, _10166_, _10264_);
  or g_37734_(_10262_, _10264_, _10265_);
  or g_37735_(_10182_, _10264_, _10266_);
  and g_37736_(_10181_, _10265_, _10267_);
  and g_37737_(_10174_, _10177_, _10268_);
  and g_37738_(_10151_, _10155_, _10269_);
  or g_37739_(_10268_, _10269_, _10270_);
  xor g_37740_(_10137_, _10147_, _10271_);
  or g_37741_(_10157_, _10271_, _10272_);
  or g_37742_(_10270_, _10272_, _10273_);
  or g_37743_(_10267_, _10273_, _10275_);
  and g_37744_(_10160_, _10275_, _10276_);
  and g_37745_(_18573_, _10135_, _10277_);
  or g_37746_(_10228_, _10266_, _10278_);
  or g_37747_(_10273_, _10277_, _10279_);
  or g_37748_(_10250_, _10279_, _10280_);
  or g_37749_(_10278_, _10280_, _10281_);
  not g_37750_(_10281_, _10282_);
  or g_37751_(_10276_, _10282_, _10283_);
  not g_37752_(_10283_, _10284_);
  or g_37753_(_10135_, _10284_, _10286_);
  or g_37754_(out[288], _10283_, _10287_);
  and g_37755_(_10286_, _10287_, _10288_);
  not g_37756_(_10288_, _10289_);
  and g_37757_(_10245_, _10283_, _10290_);
  not g_37758_(_10290_, _10291_);
  or g_37759_(out[289], _10283_, _10292_);
  not g_37760_(_10292_, _10293_);
  and g_37761_(_10291_, _10292_, _10294_);
  or g_37762_(_10290_, _10293_, _10295_);
  and g_37763_(out[304], _10289_, _10297_);
  or g_37764_(_18562_, _10288_, _10298_);
  and g_37765_(_19794_, _10294_, _10299_);
  or g_37766_(out[305], _10295_, _10300_);
  xor g_37767_(_19794_, _10294_, _10301_);
  xor g_37768_(out[305], _10294_, _10302_);
  and g_37769_(_10298_, _10301_, _10303_);
  or g_37770_(_10297_, _10302_, _10304_);
  and g_37771_(_10232_, _10283_, _10305_);
  and g_37772_(out[291], _10284_, _10306_);
  or g_37773_(_10305_, _10306_, _10308_);
  or g_37774_(_19816_, _10308_, _10309_);
  and g_37775_(_10236_, _10283_, _10310_);
  and g_37776_(_19684_, _10284_, _10311_);
  or g_37777_(_10310_, _10311_, _10312_);
  or g_37778_(out[306], _10312_, _10313_);
  and g_37779_(_19816_, _10308_, _10314_);
  xor g_37780_(_19816_, _10308_, _10315_);
  xor g_37781_(out[307], _10308_, _10316_);
  xor g_37782_(out[306], _10312_, _10317_);
  xor g_37783_(_19805_, _10312_, _10319_);
  and g_37784_(_10315_, _10317_, _10320_);
  or g_37785_(_10316_, _10319_, _10321_);
  and g_37786_(_18562_, _10288_, _10322_);
  or g_37787_(out[304], _10289_, _10323_);
  or g_37788_(_10321_, _10322_, _10324_);
  and g_37789_(_10303_, _10323_, _10325_);
  and g_37790_(_10320_, _10325_, _10326_);
  or g_37791_(_10304_, _10324_, _10327_);
  and g_37792_(out[308], out[307], _10328_);
  or g_37793_(out[309], _10328_, _10330_);
  or g_37794_(out[310], _10330_, _10331_);
  or g_37795_(out[311], _10331_, _10332_);
  xor g_37796_(out[311], _10331_, _10333_);
  not g_37797_(_10333_, _10334_);
  and g_37798_(_10195_, _10283_, _10335_);
  or g_37799_(_10194_, _10284_, _10336_);
  or g_37800_(_10189_, _10283_, _10337_);
  not g_37801_(_10337_, _10338_);
  and g_37802_(_10336_, _10337_, _10339_);
  or g_37803_(_10335_, _10338_, _10341_);
  and g_37804_(_10333_, _10341_, _10342_);
  or g_37805_(_10334_, _10339_, _10343_);
  xor g_37806_(out[310], _10330_, _10344_);
  xor g_37807_(_19761_, _10330_, _10345_);
  and g_37808_(_10187_, _10283_, _10346_);
  not g_37809_(_10346_, _10347_);
  or g_37810_(_10183_, _10283_, _10348_);
  not g_37811_(_10348_, _10349_);
  or g_37812_(_10346_, _10349_, _10350_);
  and g_37813_(_10347_, _10348_, _10352_);
  and g_37814_(_10344_, _10350_, _10353_);
  or g_37815_(_10345_, _10352_, _10354_);
  and g_37816_(_10343_, _10354_, _10355_);
  or g_37817_(_10342_, _10353_, _10356_);
  and g_37818_(_10345_, _10352_, _10357_);
  and g_37819_(_10334_, _10339_, _10358_);
  or g_37820_(_10357_, _10358_, _10359_);
  not g_37821_(_10359_, _10360_);
  and g_37822_(_10355_, _10360_, _10361_);
  or g_37823_(_10356_, _10359_, _10363_);
  xor g_37824_(out[308], out[307], _10364_);
  xor g_37825_(_19772_, out[307], _10365_);
  or g_37826_(_10214_, _10283_, _10366_);
  or g_37827_(_10222_, _10284_, _10367_);
  and g_37828_(_10366_, _10367_, _10368_);
  not g_37829_(_10368_, _10369_);
  and g_37830_(_10365_, _10368_, _10370_);
  not g_37831_(_10370_, _10371_);
  or g_37832_(_10204_, _10284_, _10372_);
  or g_37833_(_10206_, _10283_, _10374_);
  and g_37834_(_10372_, _10374_, _10375_);
  not g_37835_(_10375_, _10376_);
  xor g_37836_(out[309], _10328_, _10377_);
  xor g_37837_(_19783_, _10328_, _10378_);
  or g_37838_(_10375_, _10378_, _10379_);
  and g_37839_(_10371_, _10379_, _10380_);
  not g_37840_(_10380_, _10381_);
  or g_37841_(_10376_, _10377_, _10382_);
  not g_37842_(_10382_, _10383_);
  or g_37843_(_10365_, _10368_, _10385_);
  and g_37844_(_10382_, _10385_, _10386_);
  and g_37845_(_10380_, _10386_, _10387_);
  and g_37846_(_10361_, _10387_, _10388_);
  not g_37847_(_10388_, _10389_);
  and g_37848_(_10137_, _10147_, _10390_);
  not g_37849_(_10390_, _10391_);
  or g_37850_(out[312], _10332_, _10392_);
  and g_37851_(out[313], _10392_, _10393_);
  or g_37852_(out[314], _10393_, _10394_);
  xor g_37853_(out[315], _10394_, _10396_);
  not g_37854_(_10396_, _10397_);
  and g_37855_(_10391_, _10396_, _10398_);
  or g_37856_(_10390_, _10397_, _10399_);
  xor g_37857_(out[314], _10393_, _10400_);
  not g_37858_(_10400_, _10401_);
  and g_37859_(_10155_, _10283_, _10402_);
  and g_37860_(_10150_, _10284_, _10403_);
  or g_37861_(_10402_, _10403_, _10404_);
  not g_37862_(_10404_, _10405_);
  and g_37863_(_10401_, _10404_, _10407_);
  or g_37864_(_10400_, _10405_, _10408_);
  and g_37865_(_10399_, _10408_, _10409_);
  or g_37866_(_10398_, _10407_, _10410_);
  and g_37867_(_10176_, _10283_, _10411_);
  or g_37868_(_10174_, _10284_, _10412_);
  and g_37869_(_10177_, _10284_, _10413_);
  or g_37870_(_10178_, _10283_, _10414_);
  and g_37871_(_10412_, _10414_, _10415_);
  or g_37872_(_10411_, _10413_, _10416_);
  xor g_37873_(out[313], _10392_, _10418_);
  xor g_37874_(_19838_, _10392_, _10419_);
  and g_37875_(_10415_, _10418_, _10420_);
  or g_37876_(_10416_, _10419_, _10421_);
  and g_37877_(_10409_, _10421_, _10422_);
  or g_37878_(_10410_, _10420_, _10423_);
  and g_37879_(_10400_, _10405_, _10424_);
  or g_37880_(_10401_, _10404_, _10425_);
  and g_37881_(_10390_, _10397_, _10426_);
  or g_37882_(_10391_, _10396_, _10427_);
  and g_37883_(_10425_, _10427_, _10429_);
  or g_37884_(_10424_, _10426_, _10430_);
  and g_37885_(_10416_, _10419_, _10431_);
  or g_37886_(_10415_, _10418_, _10432_);
  xor g_37887_(out[312], _10332_, _10433_);
  not g_37888_(_10433_, _10434_);
  and g_37889_(_10166_, _10283_, _10435_);
  and g_37890_(_10161_, _10284_, _10436_);
  or g_37891_(_10435_, _10436_, _10437_);
  not g_37892_(_10437_, _10438_);
  and g_37893_(_10434_, _10437_, _10440_);
  or g_37894_(_10433_, _10438_, _10441_);
  and g_37895_(_10432_, _10441_, _10442_);
  or g_37896_(_10431_, _10440_, _10443_);
  and g_37897_(_10433_, _10438_, _10444_);
  or g_37898_(_10434_, _10437_, _10445_);
  and g_37899_(_10442_, _10445_, _10446_);
  or g_37900_(_10443_, _10444_, _10447_);
  and g_37901_(_10429_, _10446_, _10448_);
  or g_37902_(_10430_, _10447_, _10449_);
  and g_37903_(_10422_, _10448_, _10451_);
  or g_37904_(_10423_, _10449_, _10452_);
  or g_37905_(_10389_, _10452_, _10453_);
  and g_37906_(_10326_, _10388_, _10454_);
  and g_37907_(_10451_, _10454_, _10455_);
  or g_37908_(_10327_, _10453_, _10456_);
  and g_37909_(_10300_, _10304_, _10457_);
  or g_37910_(_10299_, _10303_, _10458_);
  and g_37911_(_10320_, _10458_, _10459_);
  or g_37912_(_10321_, _10457_, _10460_);
  or g_37913_(_10313_, _10314_, _10462_);
  and g_37914_(_10309_, _10462_, _10463_);
  not g_37915_(_10463_, _10464_);
  and g_37916_(_10460_, _10463_, _10465_);
  or g_37917_(_10459_, _10464_, _10466_);
  or g_37918_(_10453_, _10465_, _10467_);
  and g_37919_(_10399_, _10430_, _10468_);
  or g_37920_(_10398_, _10429_, _10469_);
  and g_37921_(_10432_, _10445_, _10470_);
  or g_37922_(_10431_, _10444_, _10471_);
  and g_37923_(_10422_, _10471_, _10473_);
  or g_37924_(_10423_, _10470_, _10474_);
  and g_37925_(_10469_, _10474_, _10475_);
  or g_37926_(_10468_, _10473_, _10476_);
  or g_37927_(_10355_, _10358_, _10477_);
  not g_37928_(_10477_, _10478_);
  and g_37929_(_10361_, _10381_, _10479_);
  or g_37930_(_10363_, _10380_, _10480_);
  and g_37931_(_10382_, _10479_, _10481_);
  or g_37932_(_10383_, _10480_, _10482_);
  and g_37933_(_10477_, _10482_, _10484_);
  or g_37934_(_10478_, _10481_, _10485_);
  or g_37935_(_10452_, _10484_, _10486_);
  and g_37936_(_10475_, _10486_, _10487_);
  and g_37937_(_10388_, _10466_, _10488_);
  or g_37938_(_10485_, _10488_, _10489_);
  and g_37939_(_10451_, _10489_, _10490_);
  and g_37940_(_10467_, _10487_, _10491_);
  or g_37941_(_10476_, _10490_, _10492_);
  and g_37942_(_10456_, _10492_, _10493_);
  or g_37943_(_10455_, _10491_, _10495_);
  or g_37944_(_10288_, _10493_, _10496_);
  or g_37945_(out[304], _10495_, _10497_);
  and g_37946_(_10496_, _10497_, _10498_);
  xor g_37947_(_26213_, _10498_, _10499_);
  and g_37948_(_26051_, _26061_, _10500_);
  and g_37949_(_10390_, _10396_, _10501_);
  xor g_37950_(_10500_, _10501_, _10502_);
  or g_37951_(_26143_, _26210_, _10503_);
  or g_37952_(_26147_, _26209_, _10504_);
  and g_37953_(_10503_, _10504_, _10506_);
  or g_37954_(_10375_, _10493_, _10507_);
  or g_37955_(_10377_, _10495_, _10508_);
  and g_37956_(_10507_, _10508_, _10509_);
  and g_37957_(_26095_, _26209_, _10510_);
  and g_37958_(_26100_, _26210_, _10511_);
  or g_37959_(_10510_, _10511_, _10512_);
  or g_37960_(_10437_, _10493_, _10513_);
  or g_37961_(_10433_, _10495_, _10514_);
  and g_37962_(_10513_, _10514_, _10515_);
  xor g_37963_(_10512_, _10515_, _10517_);
  and g_37964_(_26124_, _26209_, _10518_);
  and g_37965_(_26128_, _26210_, _10519_);
  or g_37966_(_10518_, _10519_, _10520_);
  or g_37967_(_10334_, _10495_, _10521_);
  or g_37968_(_10341_, _10493_, _10522_);
  and g_37969_(_10521_, _10522_, _10523_);
  xor g_37970_(_10520_, _10523_, _10524_);
  and g_37971_(_26066_, _26209_, _10525_);
  and g_37972_(_26070_, _26210_, _10526_);
  or g_37973_(_10525_, _10526_, _10528_);
  and g_37974_(_10400_, _10493_, _10529_);
  and g_37975_(_10404_, _10495_, _10530_);
  or g_37976_(_10529_, _10530_, _10531_);
  or g_37977_(_26115_, _26210_, _10532_);
  or g_37978_(_26120_, _26209_, _10533_);
  and g_37979_(_10532_, _10533_, _10534_);
  or g_37980_(_10345_, _10495_, _10535_);
  or g_37981_(_10350_, _10493_, _10536_);
  and g_37982_(_10535_, _10536_, _10537_);
  and g_37983_(_26091_, _26209_, _10539_);
  or g_37984_(_26092_, _26210_, _10540_);
  and g_37985_(_26090_, _26210_, _10541_);
  or g_37986_(_26089_, _26209_, _10542_);
  and g_37987_(_10540_, _10542_, _10543_);
  or g_37988_(_10539_, _10541_, _10544_);
  and g_37989_(_10416_, _10495_, _10545_);
  or g_37990_(_10415_, _10493_, _10546_);
  and g_37991_(_10418_, _10493_, _10547_);
  or g_37992_(_10419_, _10495_, _10548_);
  and g_37993_(_10546_, _10548_, _10550_);
  or g_37994_(_10545_, _10547_, _10551_);
  and g_37995_(_10544_, _10550_, _10552_);
  or g_37996_(_26028_, _26209_, _10553_);
  or g_37997_(out[146], _26210_, _10554_);
  and g_37998_(_10553_, _10554_, _10555_);
  and g_37999_(_10312_, _10495_, _10556_);
  and g_38000_(_19805_, _10493_, _10557_);
  or g_38001_(_10556_, _10557_, _10558_);
  or g_38002_(_10555_, _10558_, _10559_);
  not g_38003_(_10559_, _10561_);
  and g_38004_(_26038_, _26210_, _10562_);
  or g_38005_(_26039_, _26209_, _10563_);
  and g_38006_(_21103_, _26209_, _10564_);
  or g_38007_(out[145], _26210_, _10565_);
  and g_38008_(_10563_, _10565_, _10566_);
  or g_38009_(_10562_, _10564_, _10567_);
  and g_38010_(_10295_, _10495_, _10568_);
  or g_38011_(_10294_, _10493_, _10569_);
  and g_38012_(_19794_, _10493_, _10570_);
  or g_38013_(out[305], _10495_, _10572_);
  and g_38014_(_10569_, _10572_, _10573_);
  or g_38015_(_10568_, _10570_, _10574_);
  and g_38016_(_10567_, _10573_, _10575_);
  and g_38017_(_10566_, _10574_, _10576_);
  and g_38018_(_10543_, _10551_, _10577_);
  and g_38019_(out[147], _26209_, _10578_);
  and g_38020_(_26022_, _26210_, _10579_);
  or g_38021_(_10578_, _10579_, _10580_);
  and g_38022_(out[307], _10493_, _10581_);
  and g_38023_(_10308_, _10495_, _10583_);
  or g_38024_(_10581_, _10583_, _10584_);
  or g_38025_(_26151_, _26210_, _10585_);
  or g_38026_(_26156_, _26209_, _10586_);
  and g_38027_(_10585_, _10586_, _10587_);
  and g_38028_(_10364_, _10493_, _10588_);
  not g_38029_(_10588_, _10589_);
  or g_38030_(_10369_, _10493_, _10590_);
  not g_38031_(_10590_, _10591_);
  and g_38032_(_10589_, _10590_, _10592_);
  or g_38033_(_10588_, _10591_, _10594_);
  and g_38034_(_10555_, _10558_, _10595_);
  xor g_38035_(_10506_, _10509_, _10596_);
  or g_38036_(_10517_, _10596_, _10597_);
  not g_38037_(_10597_, _10598_);
  xor g_38038_(_10587_, _10594_, _10599_);
  xor g_38039_(_10587_, _10592_, _10600_);
  and g_38040_(_10559_, _10600_, _10601_);
  or g_38041_(_10561_, _10599_, _10602_);
  and g_38042_(_10598_, _10601_, _10603_);
  or g_38043_(_10597_, _10602_, _10605_);
  xor g_38044_(_10534_, _10537_, _10606_);
  or g_38045_(_10524_, _10606_, _10607_);
  or g_38046_(_10502_, _10577_, _10608_);
  or g_38047_(_10499_, _10608_, _10609_);
  or g_38048_(_10607_, _10609_, _10610_);
  xor g_38049_(_10528_, _10531_, _10611_);
  xor g_38050_(_10580_, _10584_, _10612_);
  or g_38051_(_10611_, _10612_, _10613_);
  or g_38052_(_10552_, _10576_, _10614_);
  or g_38053_(_10575_, _10595_, _10616_);
  or g_38054_(_10614_, _10616_, _10617_);
  or g_38055_(_10613_, _10617_, _10618_);
  or g_38056_(_10610_, _10618_, _10619_);
  not g_38057_(_10619_, _10620_);
  and g_38058_(_10603_, _10620_, _10621_);
  or g_38059_(_10605_, _10619_, _10622_);
  or g_38060_(out[138], _22141_, _10623_);
  xor g_38061_(out[138], _22141_, _10624_);
  not g_38062_(_10624_, _10625_);
  or g_38063_(out[106], _21710_, _10627_);
  xor g_38064_(out[106], _21710_, _10628_);
  xor g_38065_(_20784_, _21710_, _10629_);
  or g_38066_(out[42], _20786_, _10630_);
  not g_38067_(_10630_, _10631_);
  xor g_38068_(out[43], _10630_, _10632_);
  xor g_38069_(_20135_, _10630_, _10633_);
  or g_38070_(out[26], _20583_, _10634_);
  xor g_38071_(out[27], _10634_, _10635_);
  not g_38072_(_10635_, _10636_);
  or g_38073_(out[10], _20580_, _10638_);
  xor g_38074_(out[10], _20580_, _10639_);
  xor g_38075_(_19992_, _20580_, _10640_);
  xor g_38076_(out[26], _20583_, _10641_);
  xor g_38077_(_20124_, _20583_, _10642_);
  and g_38078_(_10640_, _10641_, _10643_);
  or g_38079_(_10639_, _10642_, _10644_);
  and g_38080_(_10639_, _10642_, _10645_);
  or g_38081_(_10640_, _10641_, _10646_);
  and g_38082_(_20590_, _20722_, _10647_);
  or g_38083_(_20589_, _20721_, _10649_);
  and g_38084_(_10646_, _10649_, _10650_);
  or g_38085_(_10645_, _10647_, _10651_);
  and g_38086_(_10644_, _10651_, _10652_);
  or g_38087_(_10643_, _10650_, _10653_);
  xor g_38088_(out[11], _10638_, _10654_);
  not g_38089_(_10654_, _10655_);
  and g_38090_(_10635_, _10655_, _10656_);
  or g_38091_(_10636_, _10654_, _10657_);
  and g_38092_(_10653_, _10657_, _10658_);
  or g_38093_(_10652_, _10656_, _10660_);
  and g_38094_(_10636_, _10654_, _10661_);
  or g_38095_(_10635_, _10655_, _10662_);
  and g_38096_(_20720_, _10662_, _10663_);
  or g_38097_(_20719_, _10661_, _10664_);
  and g_38098_(_10660_, _10663_, _10665_);
  or g_38099_(_10658_, _10664_, _10666_);
  and g_38100_(_20689_, _10666_, _10667_);
  or g_38101_(_20688_, _10665_, _10668_);
  or g_38102_(_10635_, _10668_, _10669_);
  or g_38103_(_10654_, _10667_, _10671_);
  and g_38104_(_10669_, _10671_, _10672_);
  not g_38105_(_10672_, _10673_);
  and g_38106_(_10632_, _10672_, _10674_);
  or g_38107_(_10633_, _10673_, _10675_);
  or g_38108_(out[58], _21003_, _10676_);
  xor g_38109_(out[59], _10676_, _10677_);
  xor g_38110_(_20267_, _10676_, _10678_);
  and g_38111_(_10674_, _10677_, _10679_);
  or g_38112_(_10675_, _10678_, _10680_);
  or g_38113_(out[74], _21216_, _10682_);
  xor g_38114_(out[75], _10682_, _10683_);
  xor g_38115_(_20399_, _10682_, _10684_);
  and g_38116_(_10679_, _10683_, _10685_);
  or g_38117_(_10680_, _10684_, _10686_);
  or g_38118_(out[90], _21467_, _10687_);
  xor g_38119_(out[91], _10687_, _10688_);
  xor g_38120_(_20531_, _10687_, _10689_);
  and g_38121_(_10685_, _10689_, _10690_);
  or g_38122_(_10686_, _10688_, _10691_);
  xor g_38123_(out[90], _21467_, _10693_);
  xor g_38124_(_20652_, _21467_, _10694_);
  xor g_38125_(out[58], _21003_, _10695_);
  xor g_38126_(_20388_, _21003_, _10696_);
  and g_38127_(_10674_, _10678_, _10697_);
  or g_38128_(_10675_, _10677_, _10698_);
  and g_38129_(out[42], _20786_, _10699_);
  xor g_38130_(out[42], _20786_, _10700_);
  or g_38131_(_10631_, _10699_, _10701_);
  or g_38132_(_10640_, _10667_, _10702_);
  or g_38133_(_10642_, _10668_, _10704_);
  and g_38134_(_10702_, _10704_, _10705_);
  not g_38135_(_10705_, _10706_);
  or g_38136_(_10701_, _10706_, _10707_);
  not g_38137_(_10707_, _10708_);
  and g_38138_(_10633_, _10672_, _10709_);
  or g_38139_(_10632_, _10673_, _10710_);
  and g_38140_(_10632_, _10673_, _10711_);
  or g_38141_(_10633_, _10672_, _10712_);
  xor g_38142_(_10633_, _10672_, _10713_);
  xor g_38143_(_10632_, _10672_, _10715_);
  xor g_38144_(_10700_, _10705_, _10716_);
  xor g_38145_(_10701_, _10705_, _10717_);
  and g_38146_(_10713_, _10716_, _10718_);
  or g_38147_(_10715_, _10717_, _10719_);
  and g_38148_(_20581_, _10668_, _10720_);
  or g_38149_(_20582_, _10667_, _10721_);
  and g_38150_(_20584_, _10667_, _10722_);
  or g_38151_(_20585_, _10668_, _10723_);
  and g_38152_(_10721_, _10723_, _10724_);
  or g_38153_(_10720_, _10722_, _10726_);
  and g_38154_(_20788_, _10726_, _10727_);
  or g_38155_(_20787_, _10724_, _10728_);
  and g_38156_(_20596_, _10667_, _10729_);
  or g_38157_(_20595_, _10668_, _10730_);
  and g_38158_(_20594_, _10668_, _10731_);
  or g_38159_(_20593_, _10667_, _10732_);
  and g_38160_(_10730_, _10732_, _10733_);
  or g_38161_(_10729_, _10731_, _10734_);
  and g_38162_(_20792_, _10733_, _10735_);
  or g_38163_(_20791_, _10734_, _10737_);
  and g_38164_(_10728_, _10737_, _10738_);
  or g_38165_(_10727_, _10735_, _10739_);
  and g_38166_(_20787_, _10724_, _10740_);
  or g_38167_(_20788_, _10726_, _10741_);
  and g_38168_(_20791_, _10734_, _10742_);
  or g_38169_(_20792_, _10733_, _10743_);
  and g_38170_(_10741_, _10743_, _10744_);
  or g_38171_(_10740_, _10742_, _10745_);
  and g_38172_(_10718_, _10744_, _10746_);
  or g_38173_(_10719_, _10745_, _10748_);
  and g_38174_(_10738_, _10746_, _10749_);
  or g_38175_(_10739_, _10748_, _10750_);
  and g_38176_(_20640_, _10667_, _10751_);
  or g_38177_(_20639_, _10668_, _10752_);
  and g_38178_(_20545_, _10668_, _10753_);
  or g_38179_(_20544_, _10667_, _10754_);
  and g_38180_(_10752_, _10754_, _10755_);
  or g_38181_(_10751_, _10753_, _10756_);
  and g_38182_(_20840_, _10755_, _10757_);
  or g_38183_(_20838_, _10756_, _10759_);
  and g_38184_(_20645_, _10668_, _10760_);
  or g_38185_(_20644_, _10667_, _10761_);
  and g_38186_(_20647_, _10667_, _10762_);
  or g_38187_(_20646_, _10668_, _10763_);
  and g_38188_(_10761_, _10763_, _10764_);
  or g_38189_(_10760_, _10762_, _10765_);
  and g_38190_(_20844_, _10764_, _10766_);
  or g_38191_(_20843_, _10765_, _10767_);
  and g_38192_(_10759_, _10767_, _10768_);
  or g_38193_(_10757_, _10766_, _10770_);
  and g_38194_(_20843_, _10765_, _10771_);
  or g_38195_(_20844_, _10764_, _10772_);
  or g_38196_(_20613_, _10667_, _10773_);
  or g_38197_(_20615_, _10668_, _10774_);
  and g_38198_(_10773_, _10774_, _10775_);
  not g_38199_(_10775_, _10776_);
  and g_38200_(_20620_, _10668_, _10777_);
  and g_38201_(_20622_, _10667_, _10778_);
  or g_38202_(_10777_, _10778_, _10779_);
  or g_38203_(_20825_, _10779_, _10781_);
  and g_38204_(_20825_, _10779_, _10782_);
  or g_38205_(_20815_, _10776_, _10783_);
  xor g_38206_(_20825_, _10779_, _10784_);
  xor g_38207_(_20824_, _10779_, _10785_);
  xor g_38208_(_20816_, _10775_, _10786_);
  xor g_38209_(_20815_, _10775_, _10787_);
  and g_38210_(_10784_, _10786_, _10788_);
  or g_38211_(_10785_, _10787_, _10789_);
  or g_38212_(_10771_, _10789_, _10790_);
  or g_38213_(_10768_, _10790_, _10792_);
  or g_38214_(_10782_, _10783_, _10793_);
  and g_38215_(_10781_, _10793_, _10794_);
  and g_38216_(_10792_, _10794_, _10795_);
  or g_38217_(_10750_, _10795_, _10796_);
  not g_38218_(_10796_, _10797_);
  and g_38219_(_10718_, _10739_, _10798_);
  or g_38220_(_10719_, _10738_, _10799_);
  and g_38221_(_10741_, _10798_, _10800_);
  or g_38222_(_10740_, _10799_, _10801_);
  and g_38223_(_10708_, _10712_, _10803_);
  or g_38224_(_10707_, _10711_, _10804_);
  and g_38225_(_10710_, _10804_, _10805_);
  or g_38226_(_10709_, _10800_, _10806_);
  and g_38227_(_10801_, _10805_, _10807_);
  or g_38228_(_10803_, _10806_, _10808_);
  and g_38229_(_22401_, _10667_, _10809_);
  and g_38230_(_22434_, _10668_, _10810_);
  or g_38231_(_10809_, _10810_, _10811_);
  not g_38232_(_10811_, _10812_);
  and g_38233_(_24183_, _10812_, _10814_);
  or g_38234_(_24194_, _10811_, _10815_);
  and g_38235_(_20692_, _10667_, _10816_);
  or g_38236_(_20693_, _10668_, _10817_);
  and g_38237_(_20690_, _10668_, _10818_);
  or g_38238_(_20691_, _10667_, _10819_);
  and g_38239_(_10817_, _10819_, _10820_);
  or g_38240_(_10816_, _10818_, _10821_);
  and g_38241_(_20876_, _10820_, _10822_);
  or g_38242_(_20877_, _10821_, _10823_);
  and g_38243_(_10815_, _10823_, _10825_);
  or g_38244_(_10814_, _10822_, _10826_);
  and g_38245_(out[17], _10667_, _10827_);
  or g_38246_(_20058_, _10668_, _10828_);
  and g_38247_(out[1], _10668_, _10829_);
  or g_38248_(_19926_, _10667_, _10830_);
  and g_38249_(_10828_, _10830_, _10831_);
  or g_38250_(_10827_, _10829_, _10832_);
  and g_38251_(out[33], _10831_, _10833_);
  or g_38252_(_20190_, _10832_, _10834_);
  and g_38253_(_19937_, _10668_, _10836_);
  or g_38254_(out[0], _10667_, _10837_);
  and g_38255_(_20069_, _10667_, _10838_);
  or g_38256_(out[16], _10668_, _10839_);
  and g_38257_(_10837_, _10839_, _10840_);
  or g_38258_(_10836_, _10838_, _10841_);
  and g_38259_(out[32], _10841_, _10842_);
  or g_38260_(_20201_, _10840_, _10843_);
  xor g_38261_(out[33], _10831_, _10844_);
  xor g_38262_(_20190_, _10831_, _10845_);
  and g_38263_(_10843_, _10844_, _10847_);
  or g_38264_(_10842_, _10845_, _10848_);
  and g_38265_(_10834_, _10848_, _10849_);
  or g_38266_(_10833_, _10847_, _10850_);
  xor g_38267_(_24194_, _10811_, _10851_);
  xor g_38268_(_24183_, _10811_, _10852_);
  and g_38269_(_20838_, _10756_, _10853_);
  or g_38270_(_20840_, _10755_, _10854_);
  and g_38271_(_20877_, _10821_, _10855_);
  or g_38272_(_20876_, _10820_, _10856_);
  and g_38273_(_10823_, _10856_, _10858_);
  or g_38274_(_10822_, _10855_, _10859_);
  and g_38275_(_10851_, _10858_, _10860_);
  or g_38276_(_10852_, _10859_, _10861_);
  and g_38277_(_10850_, _10860_, _10862_);
  or g_38278_(_10849_, _10861_, _10863_);
  and g_38279_(_10826_, _10856_, _10864_);
  or g_38280_(_10825_, _10855_, _10865_);
  and g_38281_(_10863_, _10865_, _10866_);
  or g_38282_(_10862_, _10864_, _10867_);
  and g_38283_(_10772_, _10854_, _10869_);
  or g_38284_(_10771_, _10853_, _10870_);
  and g_38285_(_10768_, _10869_, _10871_);
  or g_38286_(_10770_, _10870_, _10872_);
  and g_38287_(_10788_, _10871_, _10873_);
  or g_38288_(_10789_, _10872_, _10874_);
  and g_38289_(_10749_, _10873_, _10875_);
  or g_38290_(_10750_, _10874_, _10876_);
  and g_38291_(_10867_, _10875_, _10877_);
  or g_38292_(_10866_, _10876_, _10878_);
  and g_38293_(_10807_, _10878_, _10880_);
  or g_38294_(_10808_, _10877_, _10881_);
  and g_38295_(_10796_, _10880_, _10882_);
  or g_38296_(_10797_, _10881_, _10883_);
  and g_38297_(_20201_, _10840_, _10884_);
  or g_38298_(out[32], _10841_, _10885_);
  and g_38299_(_10847_, _10860_, _10886_);
  or g_38300_(_10848_, _10861_, _10887_);
  and g_38301_(_10873_, _10886_, _10888_);
  or g_38302_(_10874_, _10887_, _10889_);
  and g_38303_(_10749_, _10888_, _10891_);
  or g_38304_(_10750_, _10889_, _10892_);
  and g_38305_(_10885_, _10891_, _10893_);
  or g_38306_(_10884_, _10892_, _10894_);
  and g_38307_(_10883_, _10894_, _10895_);
  or g_38308_(_10882_, _10893_, _10896_);
  and g_38309_(_10700_, _10895_, _10897_);
  or g_38310_(_10701_, _10896_, _10898_);
  or g_38311_(_10705_, _10895_, _10899_);
  not g_38312_(_10899_, _10900_);
  and g_38313_(_10898_, _10899_, _10902_);
  or g_38314_(_10897_, _10900_, _10903_);
  and g_38315_(_10695_, _10902_, _10904_);
  or g_38316_(_10696_, _10903_, _10905_);
  and g_38317_(_10698_, _10905_, _10906_);
  or g_38318_(_10697_, _10904_, _10907_);
  and g_38319_(_10696_, _10903_, _10908_);
  or g_38320_(_10695_, _10902_, _10909_);
  and g_38321_(_10675_, _10677_, _10910_);
  or g_38322_(_10674_, _10678_, _10911_);
  and g_38323_(_10909_, _10911_, _10913_);
  or g_38324_(_10908_, _10910_, _10914_);
  and g_38325_(_10906_, _10913_, _10915_);
  or g_38326_(_10907_, _10914_, _10916_);
  and g_38327_(_20791_, _10895_, _10917_);
  not g_38328_(_10917_, _10918_);
  or g_38329_(_10734_, _10895_, _10919_);
  not g_38330_(_10919_, _10920_);
  and g_38331_(_10918_, _10919_, _10921_);
  or g_38332_(_10917_, _10920_, _10922_);
  and g_38333_(_21010_, _10922_, _10924_);
  or g_38334_(_21009_, _10921_, _10925_);
  and g_38335_(_20787_, _10895_, _10926_);
  not g_38336_(_10926_, _10927_);
  or g_38337_(_10724_, _10895_, _10928_);
  not g_38338_(_10928_, _10929_);
  and g_38339_(_10927_, _10928_, _10930_);
  or g_38340_(_10926_, _10929_, _10931_);
  and g_38341_(_21006_, _10931_, _10932_);
  or g_38342_(_21005_, _10930_, _10933_);
  and g_38343_(_10925_, _10933_, _10935_);
  or g_38344_(_10924_, _10932_, _10936_);
  and g_38345_(_21005_, _10930_, _10937_);
  or g_38346_(_21006_, _10931_, _10938_);
  and g_38347_(_21009_, _10921_, _10939_);
  or g_38348_(_21010_, _10922_, _10940_);
  and g_38349_(_10938_, _10940_, _10941_);
  or g_38350_(_10937_, _10939_, _10942_);
  and g_38351_(_10935_, _10941_, _10943_);
  or g_38352_(_10936_, _10942_, _10944_);
  and g_38353_(_10915_, _10943_, _10946_);
  or g_38354_(_10916_, _10944_, _10947_);
  or g_38355_(_20815_, _10896_, _10948_);
  or g_38356_(_10775_, _10895_, _10949_);
  and g_38357_(_10948_, _10949_, _10950_);
  not g_38358_(_10950_, _10951_);
  and g_38359_(_21032_, _10950_, _10952_);
  or g_38360_(_21031_, _10951_, _10953_);
  or g_38361_(_20824_, _10896_, _10954_);
  or g_38362_(_10779_, _10895_, _10955_);
  and g_38363_(_10954_, _10955_, _10957_);
  not g_38364_(_10957_, _10958_);
  and g_38365_(_21038_, _10957_, _10959_);
  or g_38366_(_21036_, _10958_, _10960_);
  xor g_38367_(_21032_, _10950_, _10961_);
  xor g_38368_(_21031_, _10950_, _10962_);
  and g_38369_(_10960_, _10961_, _10963_);
  or g_38370_(_10959_, _10962_, _10964_);
  and g_38371_(_20838_, _10895_, _10965_);
  not g_38372_(_10965_, _10966_);
  or g_38373_(_10756_, _10895_, _10968_);
  not g_38374_(_10968_, _10969_);
  and g_38375_(_10966_, _10968_, _10970_);
  or g_38376_(_10965_, _10969_, _10971_);
  and g_38377_(_21066_, _10971_, _10972_);
  or g_38378_(_21065_, _10970_, _10973_);
  and g_38379_(_20843_, _10895_, _10974_);
  not g_38380_(_10974_, _10975_);
  or g_38381_(_10765_, _10895_, _10976_);
  not g_38382_(_10976_, _10977_);
  and g_38383_(_10975_, _10976_, _10979_);
  or g_38384_(_10974_, _10977_, _10980_);
  and g_38385_(_21047_, _10980_, _10981_);
  or g_38386_(_21046_, _10979_, _10982_);
  and g_38387_(_10973_, _10982_, _10983_);
  or g_38388_(_10972_, _10981_, _10984_);
  and g_38389_(_21065_, _10970_, _10985_);
  or g_38390_(_21066_, _10971_, _10986_);
  and g_38391_(_21036_, _10958_, _10987_);
  or g_38392_(_21038_, _10957_, _10988_);
  and g_38393_(_21046_, _10979_, _10990_);
  or g_38394_(_21047_, _10980_, _10991_);
  and g_38395_(_10988_, _10991_, _10992_);
  or g_38396_(_10987_, _10990_, _10993_);
  and g_38397_(_10986_, _10992_, _10994_);
  or g_38398_(_10985_, _10993_, _10995_);
  and g_38399_(_10983_, _10994_, _10996_);
  or g_38400_(_10984_, _10995_, _10997_);
  and g_38401_(_10963_, _10996_, _10998_);
  or g_38402_(_10964_, _10997_, _10999_);
  and g_38403_(_24183_, _10895_, _11001_);
  or g_38404_(_24194_, _10896_, _11002_);
  and g_38405_(_10811_, _10896_, _11003_);
  or g_38406_(_10812_, _10895_, _11004_);
  and g_38407_(_11002_, _11004_, _11005_);
  or g_38408_(_11001_, _11003_, _11006_);
  and g_38409_(_10230_, _11005_, _11007_);
  or g_38410_(_10241_, _11006_, _11008_);
  xor g_38411_(_10230_, _11005_, _11009_);
  xor g_38412_(_10241_, _11005_, _11010_);
  and g_38413_(_20877_, _10895_, _11012_);
  or g_38414_(_20876_, _10896_, _11013_);
  and g_38415_(_10820_, _10896_, _11014_);
  or g_38416_(_10821_, _10895_, _11015_);
  and g_38417_(_11013_, _11015_, _11016_);
  or g_38418_(_11012_, _11014_, _11017_);
  and g_38419_(_21082_, _11016_, _11018_);
  or g_38420_(_21080_, _11017_, _11019_);
  or g_38421_(_21082_, _11016_, _11020_);
  not g_38422_(_11020_, _11021_);
  and g_38423_(_11009_, _11020_, _11023_);
  or g_38424_(_11010_, _11021_, _11024_);
  and g_38425_(_11019_, _11023_, _11025_);
  or g_38426_(_11018_, _11024_, _11026_);
  and g_38427_(out[33], _10895_, _11027_);
  not g_38428_(_11027_, _11028_);
  and g_38429_(_10832_, _10896_, _11029_);
  or g_38430_(_10831_, _10895_, _11030_);
  and g_38431_(_11028_, _11030_, _11031_);
  or g_38432_(_11027_, _11029_, _11032_);
  or g_38433_(_10840_, _10895_, _11034_);
  not g_38434_(_11034_, _11035_);
  and g_38435_(_20201_, _10895_, _11036_);
  or g_38436_(out[32], _10896_, _11037_);
  and g_38437_(_11034_, _11037_, _11038_);
  or g_38438_(_11035_, _11036_, _11039_);
  and g_38439_(out[48], _11039_, _11040_);
  or g_38440_(_20333_, _11038_, _11041_);
  and g_38441_(out[49], _11031_, _11042_);
  or g_38442_(_20322_, _11032_, _11043_);
  xor g_38443_(_20322_, _11032_, _11045_);
  xor g_38444_(out[49], _11032_, _11046_);
  and g_38445_(_11041_, _11045_, _11047_);
  or g_38446_(_11040_, _11046_, _11048_);
  and g_38447_(_11025_, _11047_, _11049_);
  or g_38448_(_11026_, _11048_, _11050_);
  and g_38449_(_11025_, _11042_, _11051_);
  or g_38450_(_11026_, _11043_, _11052_);
  and g_38451_(_11007_, _11019_, _11053_);
  or g_38452_(_11008_, _11018_, _11054_);
  and g_38453_(_11020_, _11054_, _11056_);
  or g_38454_(_11021_, _11053_, _11057_);
  and g_38455_(_11052_, _11056_, _11058_);
  or g_38456_(_11051_, _11057_, _11059_);
  and g_38457_(_11050_, _11058_, _11060_);
  or g_38458_(_11049_, _11059_, _11061_);
  and g_38459_(_10998_, _11061_, _11062_);
  or g_38460_(_10999_, _11060_, _11063_);
  and g_38461_(_10952_, _10960_, _11064_);
  or g_38462_(_10953_, _10959_, _11065_);
  and g_38463_(_10988_, _11065_, _11067_);
  or g_38464_(_10987_, _11064_, _11068_);
  and g_38465_(_10984_, _10991_, _11069_);
  or g_38466_(_10983_, _10990_, _11070_);
  and g_38467_(_10963_, _11069_, _11071_);
  or g_38468_(_10964_, _11070_, _11072_);
  and g_38469_(_11067_, _11072_, _11073_);
  or g_38470_(_11068_, _11071_, _11074_);
  and g_38471_(_11063_, _11073_, _11075_);
  or g_38472_(_11062_, _11074_, _11076_);
  and g_38473_(_10946_, _11076_, _11078_);
  or g_38474_(_10947_, _11075_, _11079_);
  and g_38475_(_10907_, _10911_, _11080_);
  or g_38476_(_10906_, _10910_, _11081_);
  and g_38477_(_10936_, _10938_, _11082_);
  or g_38478_(_10935_, _10937_, _11083_);
  and g_38479_(_10915_, _11082_, _11084_);
  or g_38480_(_10916_, _11083_, _11085_);
  and g_38481_(_11081_, _11085_, _11086_);
  or g_38482_(_11080_, _11084_, _11087_);
  and g_38483_(_11079_, _11086_, _11089_);
  or g_38484_(_11078_, _11087_, _11090_);
  and g_38485_(_20333_, _11038_, _11091_);
  or g_38486_(out[48], _11039_, _11092_);
  and g_38487_(_10946_, _11092_, _11093_);
  or g_38488_(_10947_, _11091_, _11094_);
  and g_38489_(_11049_, _11093_, _11095_);
  or g_38490_(_11050_, _11094_, _11096_);
  and g_38491_(_10998_, _11095_, _11097_);
  or g_38492_(_10999_, _11096_, _11098_);
  and g_38493_(_11090_, _11098_, _11100_);
  or g_38494_(_11089_, _11097_, _11101_);
  and g_38495_(_10695_, _11100_, _11102_);
  or g_38496_(_10696_, _11101_, _11103_);
  and g_38497_(_10903_, _11101_, _11104_);
  not g_38498_(_11104_, _11105_);
  and g_38499_(_11103_, _11105_, _11106_);
  or g_38500_(_11102_, _11104_, _11107_);
  xor g_38501_(out[74], _21216_, _11108_);
  xor g_38502_(_20520_, _21216_, _11109_);
  and g_38503_(_11106_, _11108_, _11111_);
  or g_38504_(_11107_, _11109_, _11112_);
  and g_38505_(_10679_, _10684_, _11113_);
  or g_38506_(_10680_, _10683_, _11114_);
  and g_38507_(_11112_, _11114_, _11115_);
  or g_38508_(_11111_, _11113_, _11116_);
  and g_38509_(_11107_, _11109_, _11117_);
  or g_38510_(_11106_, _11108_, _11118_);
  and g_38511_(_10680_, _10683_, _11119_);
  or g_38512_(_10679_, _10684_, _11120_);
  or g_38513_(_11117_, _11119_, _11122_);
  and g_38514_(_11115_, _11120_, _11123_);
  and g_38515_(_11118_, _11123_, _11124_);
  or g_38516_(_11116_, _11122_, _11125_);
  or g_38517_(_21036_, _11101_, _11126_);
  or g_38518_(_10957_, _11100_, _11127_);
  and g_38519_(_11126_, _11127_, _11128_);
  not g_38520_(_11128_, _11129_);
  or g_38521_(_21269_, _11128_, _11130_);
  and g_38522_(_21269_, _11128_, _11131_);
  xor g_38523_(_21269_, _11128_, _11133_);
  xor g_38524_(_21267_, _11128_, _11134_);
  or g_38525_(_21031_, _11101_, _11135_);
  or g_38526_(_10950_, _11100_, _11136_);
  and g_38527_(_11135_, _11136_, _11137_);
  not g_38528_(_11137_, _11138_);
  or g_38529_(_21256_, _11138_, _11139_);
  or g_38530_(_21047_, _11101_, _11140_);
  not g_38531_(_11140_, _11141_);
  and g_38532_(_10980_, _11101_, _11142_);
  not g_38533_(_11142_, _11144_);
  and g_38534_(_11140_, _11144_, _11145_);
  or g_38535_(_11141_, _11142_, _11146_);
  and g_38536_(_21292_, _11145_, _11147_);
  or g_38537_(_21293_, _11146_, _11148_);
  xor g_38538_(_21258_, _11137_, _11149_);
  xor g_38539_(_21256_, _11137_, _11150_);
  and g_38540_(_11133_, _11149_, _11151_);
  or g_38541_(_11134_, _11150_, _11152_);
  and g_38542_(_11148_, _11151_, _11153_);
  or g_38543_(_11147_, _11152_, _11155_);
  and g_38544_(_21065_, _11100_, _11156_);
  or g_38545_(_21066_, _11101_, _11157_);
  and g_38546_(_10971_, _11101_, _11158_);
  not g_38547_(_11158_, _11159_);
  and g_38548_(_11157_, _11159_, _11160_);
  or g_38549_(_11156_, _11158_, _11161_);
  and g_38550_(_21288_, _11161_, _11162_);
  or g_38551_(_21287_, _11160_, _11163_);
  and g_38552_(_21293_, _11146_, _11164_);
  or g_38553_(_21292_, _11145_, _11166_);
  and g_38554_(_11163_, _11166_, _11167_);
  or g_38555_(_11162_, _11164_, _11168_);
  and g_38556_(_21287_, _11160_, _11169_);
  or g_38557_(_21288_, _11161_, _11170_);
  and g_38558_(_11167_, _11170_, _11171_);
  or g_38559_(_11168_, _11169_, _11172_);
  and g_38560_(_11153_, _11171_, _11173_);
  or g_38561_(_11155_, _11172_, _11174_);
  or g_38562_(_11016_, _11100_, _11175_);
  or g_38563_(_21080_, _11101_, _11177_);
  and g_38564_(_11175_, _11177_, _11178_);
  not g_38565_(_11178_, _11179_);
  or g_38566_(_21319_, _11178_, _11180_);
  and g_38567_(_11006_, _11101_, _11181_);
  and g_38568_(_10230_, _11100_, _11182_);
  or g_38569_(_11181_, _11182_, _11183_);
  not g_38570_(_11183_, _11184_);
  and g_38571_(_21319_, _11178_, _11185_);
  or g_38572_(_12540_, _11183_, _11186_);
  xor g_38573_(_21319_, _11178_, _11188_);
  xor g_38574_(_21318_, _11178_, _11189_);
  xor g_38575_(_12540_, _11183_, _11190_);
  xor g_38576_(_12529_, _11183_, _11191_);
  and g_38577_(_11188_, _11190_, _11192_);
  or g_38578_(_11189_, _11191_, _11193_);
  or g_38579_(_20322_, _11101_, _11194_);
  or g_38580_(_11031_, _11100_, _11195_);
  and g_38581_(_11194_, _11195_, _11196_);
  and g_38582_(out[65], _11196_, _11197_);
  not g_38583_(_11197_, _11199_);
  and g_38584_(_11039_, _11101_, _11200_);
  or g_38585_(_11038_, _11100_, _11201_);
  and g_38586_(_20333_, _11100_, _11202_);
  or g_38587_(out[48], _11101_, _11203_);
  and g_38588_(_11201_, _11203_, _11204_);
  or g_38589_(_11200_, _11202_, _11205_);
  and g_38590_(out[64], _11205_, _11206_);
  or g_38591_(_20465_, _11204_, _11207_);
  xor g_38592_(out[65], _11196_, _11208_);
  xor g_38593_(_20454_, _11196_, _11210_);
  and g_38594_(_11207_, _11208_, _11211_);
  or g_38595_(_11206_, _11210_, _11212_);
  and g_38596_(_11199_, _11212_, _11213_);
  or g_38597_(_11197_, _11211_, _11214_);
  and g_38598_(_11192_, _11214_, _11215_);
  or g_38599_(_11193_, _11213_, _11216_);
  or g_38600_(_11185_, _11186_, _11217_);
  and g_38601_(_11180_, _11217_, _11218_);
  not g_38602_(_11218_, _11219_);
  and g_38603_(_11216_, _11218_, _11221_);
  or g_38604_(_11215_, _11219_, _11222_);
  and g_38605_(_11173_, _11222_, _11223_);
  or g_38606_(_11174_, _11221_, _11224_);
  and g_38607_(_11153_, _11168_, _11225_);
  or g_38608_(_11155_, _11167_, _11226_);
  or g_38609_(_11131_, _11139_, _11227_);
  and g_38610_(_11130_, _11227_, _11228_);
  not g_38611_(_11228_, _11229_);
  and g_38612_(_11226_, _11228_, _11230_);
  or g_38613_(_11225_, _11229_, _11232_);
  and g_38614_(_11224_, _11230_, _11233_);
  or g_38615_(_11223_, _11232_, _11234_);
  or g_38616_(_21006_, _11101_, _11235_);
  not g_38617_(_11235_, _11236_);
  and g_38618_(_10931_, _11101_, _11237_);
  not g_38619_(_11237_, _11238_);
  and g_38620_(_11235_, _11238_, _11239_);
  or g_38621_(_11236_, _11237_, _11240_);
  and g_38622_(_21218_, _11240_, _11241_);
  or g_38623_(_21217_, _11239_, _11243_);
  or g_38624_(_21010_, _11101_, _11244_);
  not g_38625_(_11244_, _11245_);
  and g_38626_(_10922_, _11101_, _11246_);
  not g_38627_(_11246_, _11247_);
  and g_38628_(_11244_, _11247_, _11248_);
  or g_38629_(_11245_, _11246_, _11249_);
  and g_38630_(_21229_, _11249_, _11250_);
  or g_38631_(_21228_, _11248_, _11251_);
  and g_38632_(_11243_, _11251_, _11252_);
  or g_38633_(_11241_, _11250_, _11254_);
  and g_38634_(_21228_, _11248_, _11255_);
  or g_38635_(_21229_, _11249_, _11256_);
  and g_38636_(_21217_, _11239_, _11257_);
  or g_38637_(_21218_, _11240_, _11258_);
  and g_38638_(_11256_, _11258_, _11259_);
  or g_38639_(_11255_, _11257_, _11260_);
  and g_38640_(_11252_, _11259_, _11261_);
  or g_38641_(_11254_, _11260_, _11262_);
  and g_38642_(_11234_, _11261_, _11263_);
  or g_38643_(_11233_, _11262_, _11265_);
  and g_38644_(_11254_, _11258_, _11266_);
  or g_38645_(_11252_, _11257_, _11267_);
  and g_38646_(_11265_, _11267_, _11268_);
  or g_38647_(_11263_, _11266_, _11269_);
  and g_38648_(_11124_, _11269_, _11270_);
  or g_38649_(_11125_, _11268_, _11271_);
  and g_38650_(_11116_, _11120_, _11272_);
  or g_38651_(_11115_, _11119_, _11273_);
  and g_38652_(_11271_, _11273_, _11274_);
  or g_38653_(_11270_, _11272_, _11276_);
  and g_38654_(_11192_, _11211_, _11277_);
  or g_38655_(_11193_, _11212_, _11278_);
  and g_38656_(_11261_, _11277_, _11279_);
  or g_38657_(_11262_, _11278_, _11280_);
  and g_38658_(_20465_, _11204_, _11281_);
  or g_38659_(out[64], _11205_, _11282_);
  and g_38660_(_11124_, _11282_, _11283_);
  or g_38661_(_11125_, _11281_, _11284_);
  and g_38662_(_11279_, _11283_, _11285_);
  or g_38663_(_11280_, _11284_, _11287_);
  and g_38664_(_11173_, _11285_, _11288_);
  or g_38665_(_11174_, _11287_, _11289_);
  and g_38666_(_11276_, _11289_, _11290_);
  or g_38667_(_11274_, _11288_, _11291_);
  and g_38668_(_11107_, _11291_, _11292_);
  not g_38669_(_11292_, _11293_);
  and g_38670_(_11108_, _11290_, _11294_);
  or g_38671_(_11109_, _11291_, _11295_);
  and g_38672_(_11293_, _11295_, _11296_);
  or g_38673_(_11292_, _11294_, _11298_);
  and g_38674_(_10693_, _11296_, _11299_);
  or g_38675_(_10694_, _11298_, _11300_);
  and g_38676_(_10691_, _11300_, _11301_);
  or g_38677_(_10690_, _11299_, _11302_);
  and g_38678_(_10686_, _10688_, _11303_);
  or g_38679_(_10685_, _10689_, _11304_);
  and g_38680_(_10694_, _11298_, _11305_);
  or g_38681_(_10693_, _11296_, _11306_);
  or g_38682_(_11303_, _11305_, _11307_);
  and g_38683_(_11301_, _11306_, _11309_);
  and g_38684_(_11304_, _11309_, _11310_);
  or g_38685_(_11302_, _11307_, _11311_);
  and g_38686_(_11249_, _11291_, _11312_);
  not g_38687_(_11312_, _11313_);
  or g_38688_(_21229_, _11291_, _11314_);
  not g_38689_(_11314_, _11315_);
  and g_38690_(_11313_, _11314_, _11316_);
  or g_38691_(_11312_, _11315_, _11317_);
  and g_38692_(_21475_, _11317_, _11318_);
  or g_38693_(_21474_, _11316_, _11320_);
  or g_38694_(_21218_, _11291_, _11321_);
  not g_38695_(_11321_, _11322_);
  and g_38696_(_11240_, _11291_, _11323_);
  not g_38697_(_11323_, _11324_);
  and g_38698_(_11321_, _11324_, _11325_);
  or g_38699_(_11322_, _11323_, _11326_);
  and g_38700_(_21469_, _11326_, _11327_);
  or g_38701_(_21468_, _11325_, _11328_);
  and g_38702_(_11320_, _11328_, _11329_);
  or g_38703_(_11318_, _11327_, _11331_);
  and g_38704_(_21468_, _11325_, _11332_);
  or g_38705_(_21469_, _11326_, _11333_);
  and g_38706_(_21474_, _11316_, _11334_);
  or g_38707_(_21475_, _11317_, _11335_);
  and g_38708_(_11333_, _11335_, _11336_);
  or g_38709_(_11332_, _11334_, _11337_);
  and g_38710_(_11329_, _11336_, _11338_);
  or g_38711_(_11331_, _11337_, _11339_);
  and g_38712_(_11310_, _11338_, _11340_);
  or g_38713_(_11311_, _11339_, _11342_);
  or g_38714_(_11137_, _11290_, _11343_);
  or g_38715_(_21256_, _11291_, _11344_);
  and g_38716_(_11343_, _11344_, _11345_);
  not g_38717_(_11345_, _11346_);
  and g_38718_(_21526_, _11345_, _11347_);
  or g_38719_(_21525_, _11346_, _11348_);
  and g_38720_(_11129_, _11291_, _11349_);
  or g_38721_(_11128_, _11290_, _11350_);
  and g_38722_(_21269_, _11290_, _11351_);
  or g_38723_(_21267_, _11291_, _11353_);
  and g_38724_(_11350_, _11353_, _11354_);
  or g_38725_(_11349_, _11351_, _11355_);
  and g_38726_(_21512_, _11355_, _11356_);
  or g_38727_(_21513_, _11354_, _11357_);
  and g_38728_(_21513_, _11354_, _11358_);
  or g_38729_(_21512_, _11355_, _11359_);
  and g_38730_(_11146_, _11291_, _11360_);
  not g_38731_(_11360_, _11361_);
  or g_38732_(_21293_, _11291_, _11362_);
  not g_38733_(_11362_, _11364_);
  and g_38734_(_11361_, _11362_, _11365_);
  or g_38735_(_11360_, _11364_, _11366_);
  or g_38736_(_21548_, _11366_, _11367_);
  not g_38737_(_11367_, _11368_);
  xor g_38738_(_21526_, _11345_, _11369_);
  xor g_38739_(_21525_, _11345_, _11370_);
  and g_38740_(_11359_, _11369_, _11371_);
  or g_38741_(_11358_, _11370_, _11372_);
  and g_38742_(_11357_, _11371_, _11373_);
  or g_38743_(_11356_, _11372_, _11375_);
  and g_38744_(_11367_, _11373_, _11376_);
  or g_38745_(_11368_, _11375_, _11377_);
  or g_38746_(_21288_, _11291_, _11378_);
  not g_38747_(_11378_, _11379_);
  and g_38748_(_11161_, _11291_, _11380_);
  not g_38749_(_11380_, _11381_);
  and g_38750_(_11378_, _11381_, _11382_);
  or g_38751_(_11379_, _11380_, _11383_);
  and g_38752_(_21561_, _11383_, _11384_);
  or g_38753_(_21560_, _11382_, _11386_);
  and g_38754_(_21548_, _11366_, _11387_);
  or g_38755_(_21547_, _11365_, _11388_);
  and g_38756_(_11386_, _11388_, _11389_);
  or g_38757_(_11384_, _11387_, _11390_);
  or g_38758_(_21561_, _11383_, _11391_);
  not g_38759_(_11391_, _11392_);
  and g_38760_(_11389_, _11391_, _11393_);
  or g_38761_(_11390_, _11392_, _11394_);
  and g_38762_(_11376_, _11393_, _11395_);
  or g_38763_(_11377_, _11394_, _11397_);
  and g_38764_(_21319_, _11290_, _11398_);
  or g_38765_(_21318_, _11291_, _11399_);
  and g_38766_(_11179_, _11291_, _11400_);
  or g_38767_(_11178_, _11290_, _11401_);
  and g_38768_(_11399_, _11401_, _11402_);
  or g_38769_(_11398_, _11400_, _11403_);
  or g_38770_(_21572_, _11402_, _11404_);
  not g_38771_(_11404_, _11405_);
  and g_38772_(_21572_, _11402_, _11406_);
  or g_38773_(_21571_, _11403_, _11408_);
  and g_38774_(_11404_, _11408_, _11409_);
  xor g_38775_(_21571_, _11402_, _11410_);
  and g_38776_(_11183_, _11291_, _11411_);
  or g_38777_(_11184_, _11290_, _11412_);
  and g_38778_(_12529_, _11290_, _11413_);
  or g_38779_(_12540_, _11291_, _11414_);
  and g_38780_(_11412_, _11414_, _11415_);
  or g_38781_(_11411_, _11413_, _11416_);
  and g_38782_(_14575_, _11415_, _11417_);
  or g_38783_(_14586_, _11416_, _11419_);
  xor g_38784_(_14575_, _11415_, _11420_);
  xor g_38785_(_14586_, _11415_, _11421_);
  and g_38786_(_11409_, _11420_, _11422_);
  or g_38787_(_11410_, _11421_, _11423_);
  and g_38788_(_11196_, _11291_, _11424_);
  not g_38789_(_11424_, _11425_);
  and g_38790_(_20454_, _11290_, _11426_);
  or g_38791_(out[65], _11291_, _11427_);
  or g_38792_(_11424_, _11426_, _11428_);
  and g_38793_(_11425_, _11427_, _11430_);
  and g_38794_(_11205_, _11291_, _11431_);
  or g_38795_(_11204_, _11290_, _11432_);
  or g_38796_(out[64], _11291_, _11433_);
  not g_38797_(_11433_, _11434_);
  and g_38798_(_11432_, _11433_, _11435_);
  or g_38799_(_11431_, _11434_, _11436_);
  and g_38800_(out[80], _11436_, _11437_);
  or g_38801_(_20597_, _11435_, _11438_);
  and g_38802_(out[81], _11428_, _11439_);
  or g_38803_(_20586_, _11430_, _11441_);
  xor g_38804_(out[81], _11428_, _11442_);
  xor g_38805_(_20586_, _11428_, _11443_);
  and g_38806_(_11438_, _11442_, _11444_);
  or g_38807_(_11437_, _11443_, _11445_);
  and g_38808_(_11422_, _11444_, _11446_);
  or g_38809_(_11423_, _11445_, _11447_);
  and g_38810_(_11422_, _11439_, _11448_);
  or g_38811_(_11423_, _11441_, _11449_);
  and g_38812_(_11408_, _11417_, _11450_);
  or g_38813_(_11406_, _11419_, _11452_);
  and g_38814_(_11404_, _11452_, _11453_);
  or g_38815_(_11405_, _11450_, _11454_);
  and g_38816_(_11449_, _11453_, _11455_);
  or g_38817_(_11448_, _11454_, _11456_);
  and g_38818_(_11447_, _11455_, _11457_);
  or g_38819_(_11446_, _11456_, _11458_);
  and g_38820_(_11395_, _11458_, _11459_);
  or g_38821_(_11397_, _11457_, _11460_);
  and g_38822_(_11376_, _11390_, _11461_);
  or g_38823_(_11377_, _11389_, _11463_);
  and g_38824_(_11347_, _11359_, _11464_);
  or g_38825_(_11348_, _11358_, _11465_);
  and g_38826_(_11357_, _11465_, _11466_);
  or g_38827_(_11356_, _11464_, _11467_);
  and g_38828_(_11463_, _11466_, _11468_);
  or g_38829_(_11461_, _11467_, _11469_);
  and g_38830_(_11460_, _11468_, _11470_);
  or g_38831_(_11459_, _11469_, _11471_);
  and g_38832_(_11340_, _11471_, _11472_);
  or g_38833_(_11342_, _11470_, _11474_);
  and g_38834_(_11302_, _11304_, _11475_);
  or g_38835_(_11301_, _11303_, _11476_);
  and g_38836_(_11331_, _11333_, _11477_);
  or g_38837_(_11329_, _11332_, _11478_);
  and g_38838_(_11310_, _11477_, _11479_);
  or g_38839_(_11311_, _11478_, _11480_);
  and g_38840_(_11476_, _11480_, _11481_);
  or g_38841_(_11475_, _11479_, _11482_);
  and g_38842_(_11474_, _11481_, _11483_);
  or g_38843_(_11472_, _11482_, _11485_);
  and g_38844_(_20597_, _11435_, _11486_);
  or g_38845_(out[80], _11436_, _11487_);
  or g_38846_(_11342_, _11447_, _11488_);
  or g_38847_(_11397_, _11488_, _11489_);
  not g_38848_(_11489_, _11490_);
  and g_38849_(_11487_, _11490_, _11491_);
  or g_38850_(_11486_, _11489_, _11492_);
  and g_38851_(_11485_, _11492_, _11493_);
  or g_38852_(_11483_, _11491_, _11494_);
  or g_38853_(_21571_, _11494_, _11496_);
  or g_38854_(_11402_, _11493_, _11497_);
  and g_38855_(_11496_, _11497_, _11498_);
  or g_38856_(_21790_, _11498_, _11499_);
  and g_38857_(_11416_, _11494_, _11500_);
  and g_38858_(_14575_, _11493_, _11501_);
  or g_38859_(_11500_, _11501_, _11502_);
  or g_38860_(_17006_, _11502_, _11503_);
  and g_38861_(_11499_, _11503_, _11504_);
  and g_38862_(_21790_, _11498_, _11505_);
  xor g_38863_(_21789_, _11498_, _11507_);
  xor g_38864_(_16995_, _11502_, _11508_);
  or g_38865_(_11507_, _11508_, _11509_);
  and g_38866_(out[81], _11493_, _11510_);
  and g_38867_(_11430_, _11494_, _11511_);
  or g_38868_(_11510_, _11511_, _11512_);
  or g_38869_(_20718_, _11512_, _11513_);
  and g_38870_(_11436_, _11494_, _11514_);
  not g_38871_(_11514_, _11515_);
  or g_38872_(out[80], _11494_, _11516_);
  not g_38873_(_11516_, _11518_);
  and g_38874_(_11515_, _11516_, _11519_);
  or g_38875_(_11514_, _11518_, _11520_);
  and g_38876_(out[96], _11520_, _11521_);
  xor g_38877_(out[97], _11512_, _11522_);
  or g_38878_(_11521_, _11522_, _11523_);
  and g_38879_(_11513_, _11523_, _11524_);
  or g_38880_(_11509_, _11524_, _11525_);
  or g_38881_(_11504_, _11505_, _11526_);
  and g_38882_(_11525_, _11526_, _11527_);
  and g_38883_(_21474_, _11493_, _11529_);
  or g_38884_(_21475_, _11494_, _11530_);
  and g_38885_(_11317_, _11494_, _11531_);
  or g_38886_(_11316_, _11493_, _11532_);
  and g_38887_(_11530_, _11532_, _11533_);
  or g_38888_(_11529_, _11531_, _11534_);
  and g_38889_(_21720_, _11534_, _11535_);
  or g_38890_(_21718_, _11533_, _11536_);
  and g_38891_(_21468_, _11493_, _11537_);
  or g_38892_(_21469_, _11494_, _11538_);
  and g_38893_(_11326_, _11494_, _11540_);
  or g_38894_(_11325_, _11493_, _11541_);
  and g_38895_(_11538_, _11541_, _11542_);
  or g_38896_(_11537_, _11540_, _11543_);
  and g_38897_(_21712_, _11543_, _11544_);
  or g_38898_(_21711_, _11542_, _11545_);
  and g_38899_(_11536_, _11545_, _11546_);
  or g_38900_(_11535_, _11544_, _11547_);
  and g_38901_(_10685_, _10688_, _11548_);
  or g_38902_(_10686_, _10689_, _11549_);
  xor g_38903_(out[107], _10627_, _11551_);
  xor g_38904_(_20663_, _10627_, _11552_);
  and g_38905_(_11549_, _11551_, _11553_);
  or g_38906_(_11548_, _11552_, _11554_);
  and g_38907_(_21718_, _11533_, _11555_);
  or g_38908_(_21720_, _11534_, _11556_);
  and g_38909_(_11554_, _11556_, _11557_);
  or g_38910_(_11553_, _11555_, _11558_);
  and g_38911_(_11546_, _11557_, _11559_);
  or g_38912_(_11547_, _11558_, _11560_);
  and g_38913_(_10693_, _11493_, _11562_);
  or g_38914_(_10694_, _11494_, _11563_);
  and g_38915_(_11298_, _11494_, _11564_);
  or g_38916_(_11296_, _11493_, _11565_);
  and g_38917_(_11563_, _11565_, _11566_);
  or g_38918_(_11562_, _11564_, _11567_);
  and g_38919_(_10629_, _11567_, _11568_);
  or g_38920_(_10628_, _11566_, _11569_);
  and g_38921_(_21711_, _11542_, _11570_);
  or g_38922_(_21712_, _11543_, _11571_);
  and g_38923_(_11569_, _11571_, _11573_);
  or g_38924_(_11568_, _11570_, _11574_);
  and g_38925_(_10628_, _11566_, _11575_);
  or g_38926_(_10629_, _11567_, _11576_);
  and g_38927_(_11548_, _11552_, _11577_);
  or g_38928_(_11549_, _11551_, _11578_);
  and g_38929_(_11576_, _11578_, _11579_);
  or g_38930_(_11575_, _11577_, _11580_);
  and g_38931_(_11573_, _11579_, _11581_);
  or g_38932_(_11574_, _11580_, _11582_);
  and g_38933_(_11559_, _11581_, _11584_);
  or g_38934_(_11560_, _11582_, _11585_);
  or g_38935_(_21525_, _11494_, _11586_);
  or g_38936_(_11345_, _11493_, _11587_);
  and g_38937_(_11586_, _11587_, _11588_);
  and g_38938_(_21748_, _11588_, _11589_);
  xor g_38939_(_21748_, _11588_, _11590_);
  xor g_38940_(_21747_, _11588_, _11591_);
  or g_38941_(_21512_, _11494_, _11592_);
  not g_38942_(_11592_, _11593_);
  and g_38943_(_11355_, _11494_, _11595_);
  not g_38944_(_11595_, _11596_);
  and g_38945_(_11592_, _11596_, _11597_);
  or g_38946_(_11593_, _11595_, _11598_);
  or g_38947_(_21754_, _11598_, _11599_);
  and g_38948_(_21754_, _11598_, _11600_);
  xor g_38949_(_21755_, _11597_, _11601_);
  xor g_38950_(_21754_, _11597_, _11602_);
  and g_38951_(_11590_, _11601_, _11603_);
  or g_38952_(_11591_, _11602_, _11604_);
  or g_38953_(_21548_, _11494_, _11606_);
  not g_38954_(_11606_, _11607_);
  and g_38955_(_11366_, _11494_, _11608_);
  not g_38956_(_11608_, _11609_);
  and g_38957_(_11606_, _11609_, _11610_);
  or g_38958_(_11607_, _11608_, _11611_);
  and g_38959_(_21739_, _11611_, _11612_);
  or g_38960_(_21738_, _11610_, _11613_);
  or g_38961_(_21561_, _11494_, _11614_);
  not g_38962_(_11614_, _11615_);
  and g_38963_(_11383_, _11494_, _11617_);
  not g_38964_(_11617_, _11618_);
  and g_38965_(_11614_, _11618_, _11619_);
  or g_38966_(_11615_, _11617_, _11620_);
  and g_38967_(_21775_, _11620_, _11621_);
  or g_38968_(_21773_, _11619_, _11622_);
  and g_38969_(_11613_, _11622_, _11623_);
  or g_38970_(_11612_, _11621_, _11624_);
  and g_38971_(_21738_, _11610_, _11625_);
  or g_38972_(_21739_, _11611_, _11626_);
  and g_38973_(_21773_, _11619_, _11628_);
  or g_38974_(_21775_, _11620_, _11629_);
  and g_38975_(_11626_, _11629_, _11630_);
  or g_38976_(_11625_, _11628_, _11631_);
  and g_38977_(_11623_, _11630_, _11632_);
  or g_38978_(_11624_, _11631_, _11633_);
  and g_38979_(_11603_, _11632_, _11634_);
  or g_38980_(_11604_, _11633_, _11635_);
  and g_38981_(_11584_, _11634_, _11636_);
  or g_38982_(_11585_, _11635_, _11637_);
  or g_38983_(_11527_, _11637_, _11639_);
  not g_38984_(_11639_, _11640_);
  and g_38985_(_11624_, _11626_, _11641_);
  or g_38986_(_11623_, _11625_, _11642_);
  and g_38987_(_11603_, _11641_, _11643_);
  or g_38988_(_11604_, _11642_, _11644_);
  and g_38989_(_11589_, _11599_, _11645_);
  or g_38990_(_11600_, _11645_, _11646_);
  not g_38991_(_11646_, _11647_);
  and g_38992_(_11644_, _11647_, _11648_);
  or g_38993_(_11643_, _11646_, _11650_);
  and g_38994_(_11584_, _11650_, _11651_);
  or g_38995_(_11585_, _11648_, _11652_);
  and g_38996_(_11547_, _11573_, _11653_);
  or g_38997_(_11546_, _11574_, _11654_);
  and g_38998_(_11579_, _11654_, _11655_);
  or g_38999_(_11580_, _11653_, _11656_);
  and g_39000_(_11554_, _11656_, _11657_);
  or g_39001_(_11553_, _11655_, _11658_);
  and g_39002_(_11652_, _11658_, _11659_);
  or g_39003_(_11651_, _11657_, _11661_);
  and g_39004_(_11639_, _11659_, _11662_);
  or g_39005_(_11640_, _11661_, _11663_);
  and g_39006_(_20729_, _11519_, _11664_);
  or g_39007_(out[96], _11520_, _11665_);
  or g_39008_(_11509_, _11523_, _11666_);
  not g_39009_(_11666_, _11667_);
  and g_39010_(_11665_, _11667_, _11668_);
  or g_39011_(_11664_, _11666_, _11669_);
  and g_39012_(_11636_, _11668_, _11670_);
  or g_39013_(_11637_, _11669_, _11672_);
  and g_39014_(_11663_, _11672_, _11673_);
  or g_39015_(_11662_, _11670_, _11674_);
  and g_39016_(_10628_, _11673_, _11675_);
  and g_39017_(_11567_, _11674_, _11676_);
  or g_39018_(_11675_, _11676_, _11677_);
  not g_39019_(_11677_, _11678_);
  and g_39020_(_11548_, _11551_, _11679_);
  or g_39021_(_11549_, _11552_, _11680_);
  or g_39022_(out[122], _21900_, _11681_);
  xor g_39023_(out[123], _11681_, _11683_);
  xor g_39024_(_20795_, _11681_, _11684_);
  and g_39025_(_11679_, _11684_, _11685_);
  or g_39026_(_11680_, _11683_, _11686_);
  xor g_39027_(out[122], _21900_, _11687_);
  xor g_39028_(_20905_, _21900_, _11688_);
  and g_39029_(_11678_, _11687_, _11689_);
  or g_39030_(_11677_, _11688_, _11690_);
  and g_39031_(_11686_, _11690_, _11691_);
  or g_39032_(_11685_, _11689_, _11692_);
  and g_39033_(_11677_, _11688_, _11694_);
  or g_39034_(_11678_, _11687_, _11695_);
  and g_39035_(_11680_, _11683_, _11696_);
  or g_39036_(_11679_, _11684_, _11697_);
  or g_39037_(_11694_, _11696_, _11698_);
  and g_39038_(_11691_, _11697_, _11699_);
  and g_39039_(_11695_, _11699_, _11700_);
  or g_39040_(_11692_, _11698_, _11701_);
  and g_39041_(_21718_, _11673_, _11702_);
  and g_39042_(_11534_, _11674_, _11703_);
  or g_39043_(_11702_, _11703_, _11705_);
  not g_39044_(_11705_, _11706_);
  and g_39045_(_21912_, _11705_, _11707_);
  or g_39046_(_21911_, _11706_, _11708_);
  and g_39047_(_21711_, _11673_, _11709_);
  and g_39048_(_11543_, _11674_, _11710_);
  or g_39049_(_11709_, _11710_, _11711_);
  not g_39050_(_11711_, _11712_);
  and g_39051_(_21902_, _11711_, _11713_);
  or g_39052_(_21901_, _11712_, _11714_);
  and g_39053_(_11708_, _11714_, _11716_);
  or g_39054_(_11707_, _11713_, _11717_);
  and g_39055_(_21901_, _11712_, _11718_);
  or g_39056_(_21902_, _11711_, _11719_);
  and g_39057_(_21911_, _11706_, _11720_);
  or g_39058_(_21912_, _11705_, _11721_);
  and g_39059_(_11719_, _11721_, _11722_);
  or g_39060_(_11718_, _11720_, _11723_);
  and g_39061_(_11716_, _11722_, _11724_);
  or g_39062_(_11717_, _11723_, _11725_);
  and g_39063_(_11700_, _11724_, _11727_);
  or g_39064_(_11701_, _11725_, _11728_);
  and g_39065_(_21755_, _11673_, _11729_);
  or g_39066_(_21754_, _11674_, _11730_);
  and g_39067_(_11598_, _11674_, _11731_);
  or g_39068_(_11597_, _11673_, _11732_);
  and g_39069_(_11730_, _11732_, _11733_);
  or g_39070_(_11729_, _11731_, _11734_);
  and g_39071_(_21938_, _11734_, _11735_);
  or g_39072_(_21938_, _11734_, _11736_);
  xor g_39073_(_21940_, _11733_, _11738_);
  xor g_39074_(_21938_, _11733_, _11739_);
  and g_39075_(_21738_, _11673_, _11740_);
  and g_39076_(_11611_, _11674_, _11741_);
  or g_39077_(_11740_, _11741_, _11742_);
  not g_39078_(_11742_, _11743_);
  and g_39079_(_21946_, _11743_, _11744_);
  or g_39080_(_21947_, _11742_, _11745_);
  or g_39081_(_21747_, _11674_, _11746_);
  or g_39082_(_11588_, _11673_, _11747_);
  and g_39083_(_11746_, _11747_, _11749_);
  and g_39084_(_21930_, _11749_, _11750_);
  xor g_39085_(_21930_, _11749_, _11751_);
  xor g_39086_(_21929_, _11749_, _11752_);
  and g_39087_(_11738_, _11751_, _11753_);
  or g_39088_(_11739_, _11752_, _11754_);
  and g_39089_(_11745_, _11753_, _11755_);
  or g_39090_(_11744_, _11754_, _11756_);
  or g_39091_(_21775_, _11674_, _11757_);
  not g_39092_(_11757_, _11758_);
  and g_39093_(_11620_, _11674_, _11760_);
  not g_39094_(_11760_, _11761_);
  and g_39095_(_11757_, _11761_, _11762_);
  or g_39096_(_11758_, _11760_, _11763_);
  and g_39097_(_21962_, _11763_, _11764_);
  or g_39098_(_21960_, _11762_, _11765_);
  and g_39099_(_21947_, _11742_, _11766_);
  or g_39100_(_21946_, _11743_, _11767_);
  and g_39101_(_11765_, _11767_, _11768_);
  or g_39102_(_11764_, _11766_, _11769_);
  and g_39103_(_21960_, _11762_, _11771_);
  or g_39104_(_21962_, _11763_, _11772_);
  and g_39105_(_11768_, _11772_, _11773_);
  or g_39106_(_11769_, _11771_, _11774_);
  and g_39107_(_11755_, _11773_, _11775_);
  or g_39108_(_11756_, _11774_, _11776_);
  or g_39109_(_21789_, _11674_, _11777_);
  or g_39110_(_11498_, _11673_, _11778_);
  and g_39111_(_11777_, _11778_, _11779_);
  or g_39112_(_21967_, _11779_, _11780_);
  and g_39113_(_21967_, _11779_, _11782_);
  xor g_39114_(_21967_, _11779_, _11783_);
  xor g_39115_(_21966_, _11779_, _11784_);
  and g_39116_(_11502_, _11674_, _11785_);
  and g_39117_(_16995_, _11673_, _11786_);
  or g_39118_(_11785_, _11786_, _11787_);
  or g_39119_(_17989_, _11787_, _11788_);
  xor g_39120_(_17989_, _11787_, _11789_);
  xor g_39121_(_17988_, _11787_, _11790_);
  and g_39122_(_11783_, _11789_, _11791_);
  or g_39123_(_11784_, _11790_, _11793_);
  and g_39124_(out[97], _11673_, _11794_);
  and g_39125_(_11512_, _11674_, _11795_);
  or g_39126_(_11794_, _11795_, _11796_);
  or g_39127_(_20850_, _11796_, _11797_);
  or g_39128_(_11793_, _11797_, _11798_);
  and g_39129_(_11780_, _11788_, _11799_);
  or g_39130_(_11782_, _11799_, _11800_);
  or g_39131_(_11756_, _11768_, _11801_);
  and g_39132_(_11736_, _11750_, _11802_);
  or g_39133_(_11735_, _11802_, _11804_);
  not g_39134_(_11804_, _11805_);
  and g_39135_(_11801_, _11805_, _11806_);
  and g_39136_(_11520_, _11674_, _11807_);
  and g_39137_(_20729_, _11673_, _11808_);
  or g_39138_(_11807_, _11808_, _11809_);
  and g_39139_(out[112], _11809_, _11810_);
  xor g_39140_(out[113], _11796_, _11811_);
  or g_39141_(_11810_, _11811_, _11812_);
  not g_39142_(_11812_, _11813_);
  and g_39143_(_11791_, _11813_, _11815_);
  or g_39144_(_11793_, _11812_, _11816_);
  and g_39145_(_11775_, _11815_, _11817_);
  and g_39146_(_11800_, _11816_, _11818_);
  and g_39147_(_11798_, _11818_, _11819_);
  or g_39148_(_11776_, _11819_, _11820_);
  and g_39149_(_11806_, _11820_, _11821_);
  or g_39150_(_11728_, _11821_, _11822_);
  or g_39151_(_11691_, _11696_, _11823_);
  or g_39152_(_11716_, _11718_, _11824_);
  or g_39153_(_11701_, _11824_, _11826_);
  and g_39154_(_11823_, _11826_, _11827_);
  and g_39155_(_11822_, _11827_, _11828_);
  or g_39156_(out[112], _11809_, _11829_);
  and g_39157_(_11727_, _11829_, _11830_);
  and g_39158_(_11817_, _11830_, _11831_);
  or g_39159_(_11828_, _11831_, _11832_);
  not g_39160_(_11832_, _11833_);
  and g_39161_(_11677_, _11832_, _11834_);
  and g_39162_(_11687_, _11833_, _11835_);
  or g_39163_(_11834_, _11835_, _11837_);
  or g_39164_(_10625_, _11837_, _11838_);
  and g_39165_(_11679_, _11683_, _11839_);
  not g_39166_(_11839_, _11840_);
  xor g_39167_(out[139], _10623_, _11841_);
  or g_39168_(_11840_, _11841_, _11842_);
  and g_39169_(_11840_, _11841_, _11843_);
  xor g_39170_(_11839_, _11841_, _11844_);
  xor g_39171_(_10624_, _11837_, _11845_);
  or g_39172_(_11844_, _11845_, _11846_);
  not g_39173_(_11846_, _11848_);
  and g_39174_(_21911_, _11833_, _11849_);
  and g_39175_(_11705_, _11832_, _11850_);
  or g_39176_(_11849_, _11850_, _11851_);
  not g_39177_(_11851_, _11852_);
  or g_39178_(_22152_, _11852_, _11853_);
  and g_39179_(_21901_, _11833_, _11854_);
  and g_39180_(_11711_, _11832_, _11855_);
  or g_39181_(_11854_, _11855_, _11856_);
  not g_39182_(_11856_, _11857_);
  or g_39183_(_22142_, _11857_, _11859_);
  and g_39184_(_11853_, _11859_, _11860_);
  not g_39185_(_11860_, _11861_);
  and g_39186_(_22142_, _11857_, _11862_);
  not g_39187_(_11862_, _11863_);
  and g_39188_(_22152_, _11852_, _11864_);
  or g_39189_(_22153_, _11851_, _11865_);
  or g_39190_(_11862_, _11864_, _11866_);
  or g_39191_(_11861_, _11866_, _11867_);
  and g_39192_(_11860_, _11863_, _11868_);
  and g_39193_(_11848_, _11865_, _11870_);
  and g_39194_(_11868_, _11870_, _11871_);
  or g_39195_(_11846_, _11867_, _11872_);
  or g_39196_(_21929_, _11832_, _11873_);
  or g_39197_(_11749_, _11833_, _11874_);
  and g_39198_(_11873_, _11874_, _11875_);
  not g_39199_(_11875_, _11876_);
  or g_39200_(_21938_, _11832_, _11877_);
  not g_39201_(_11877_, _11878_);
  and g_39202_(_11734_, _11832_, _11879_);
  or g_39203_(_11733_, _11833_, _11881_);
  and g_39204_(_11877_, _11881_, _11882_);
  or g_39205_(_11878_, _11879_, _11883_);
  or g_39206_(_22173_, _11882_, _11884_);
  or g_39207_(_22178_, _11876_, _11885_);
  and g_39208_(_22173_, _11882_, _11886_);
  and g_39209_(_21946_, _11833_, _11887_);
  or g_39210_(_21947_, _11832_, _11888_);
  and g_39211_(_11742_, _11832_, _11889_);
  not g_39212_(_11889_, _11890_);
  and g_39213_(_11888_, _11890_, _11892_);
  or g_39214_(_11887_, _11889_, _11893_);
  and g_39215_(_22040_, _11892_, _11894_);
  xor g_39216_(_22178_, _11875_, _11895_);
  xor g_39217_(_22172_, _11882_, _11896_);
  or g_39218_(_11895_, _11896_, _11897_);
  or g_39219_(_11894_, _11897_, _11898_);
  not g_39220_(_11898_, _11899_);
  and g_39221_(_21960_, _11833_, _11900_);
  and g_39222_(_11763_, _11832_, _11901_);
  or g_39223_(_11900_, _11901_, _11903_);
  not g_39224_(_11903_, _11904_);
  or g_39225_(_20536_, _11904_, _11905_);
  or g_39226_(_22040_, _11892_, _11906_);
  and g_39227_(_11905_, _11906_, _11907_);
  or g_39228_(_20537_, _11903_, _11908_);
  and g_39229_(_11907_, _11908_, _11909_);
  not g_39230_(_11909_, _11910_);
  and g_39231_(_11899_, _11909_, _11911_);
  or g_39232_(_11898_, _11910_, _11912_);
  and g_39233_(out[113], _11833_, _11914_);
  and g_39234_(_11796_, _11832_, _11915_);
  or g_39235_(_11914_, _11915_, _11916_);
  or g_39236_(_20971_, _11916_, _11917_);
  or g_39237_(_21966_, _11832_, _11918_);
  or g_39238_(_11779_, _11833_, _11919_);
  and g_39239_(_11918_, _11919_, _11920_);
  or g_39240_(_20530_, _11920_, _11921_);
  and g_39241_(_20530_, _11920_, _11922_);
  xor g_39242_(_20529_, _11920_, _11923_);
  and g_39243_(_17988_, _11833_, _11925_);
  and g_39244_(_11787_, _11832_, _11926_);
  or g_39245_(_11925_, _11926_, _11927_);
  or g_39246_(_18128_, _11927_, _11928_);
  xor g_39247_(_18127_, _11927_, _11929_);
  or g_39248_(_11923_, _11929_, _11930_);
  or g_39249_(_11917_, _11930_, _11931_);
  and g_39250_(_11809_, _11832_, _11932_);
  and g_39251_(_19860_, _11833_, _11933_);
  or g_39252_(_11932_, _11933_, _11934_);
  and g_39253_(out[128], _11934_, _11936_);
  xor g_39254_(out[129], _11916_, _11937_);
  or g_39255_(_11936_, _11937_, _11938_);
  or g_39256_(_11930_, _11938_, _11939_);
  not g_39257_(_11939_, _11940_);
  and g_39258_(_11921_, _11928_, _11941_);
  or g_39259_(_11922_, _11941_, _11942_);
  and g_39260_(_11931_, _11942_, _11943_);
  and g_39261_(_11939_, _11943_, _11944_);
  or g_39262_(_11912_, _11944_, _11945_);
  or g_39263_(_11898_, _11907_, _11947_);
  or g_39264_(_11885_, _11886_, _11948_);
  and g_39265_(_11884_, _11948_, _11949_);
  and g_39266_(_11947_, _11949_, _11950_);
  and g_39267_(_11945_, _11950_, _11951_);
  or g_39268_(_11872_, _11951_, _11952_);
  or g_39269_(_11846_, _11862_, _11953_);
  or g_39270_(_11860_, _11953_, _11954_);
  or g_39271_(_11838_, _11843_, _11955_);
  and g_39272_(_11842_, _11955_, _11956_);
  and g_39273_(_11954_, _11956_, _11958_);
  and g_39274_(_11952_, _11958_, _11959_);
  or g_39275_(out[128], _11934_, _11960_);
  and g_39276_(_11871_, _11960_, _11961_);
  and g_39277_(_11940_, _11961_, _11962_);
  and g_39278_(_11911_, _11962_, _11963_);
  or g_39279_(_11959_, _11963_, _11964_);
  not g_39280_(_11964_, _11965_);
  or g_39281_(_22172_, _11964_, _11966_);
  not g_39282_(_11966_, _11967_);
  and g_39283_(_11883_, _11964_, _11969_);
  or g_39284_(_11882_, _11965_, _11970_);
  and g_39285_(_11966_, _11970_, _11971_);
  or g_39286_(_11967_, _11969_, _11972_);
  and g_39287_(_11839_, _11841_, _11973_);
  not g_39288_(_11973_, _11974_);
  or g_39289_(out[154], _22339_, _11975_);
  xor g_39290_(out[155], _11975_, _11976_);
  not g_39291_(_11976_, _11977_);
  and g_39292_(_11973_, _11977_, _11978_);
  or g_39293_(_11974_, _11976_, _11980_);
  xor g_39294_(out[154], _22339_, _11981_);
  xor g_39295_(_21169_, _22339_, _11982_);
  and g_39296_(_10624_, _11965_, _11983_);
  or g_39297_(_10625_, _11964_, _11984_);
  and g_39298_(_11837_, _11964_, _11985_);
  not g_39299_(_11985_, _11986_);
  and g_39300_(_11984_, _11986_, _11987_);
  or g_39301_(_11983_, _11985_, _11988_);
  and g_39302_(_11981_, _11987_, _11989_);
  or g_39303_(_11982_, _11988_, _11991_);
  and g_39304_(_11980_, _11991_, _11992_);
  or g_39305_(_11978_, _11989_, _11993_);
  and g_39306_(_11982_, _11988_, _11994_);
  or g_39307_(_11981_, _11987_, _11995_);
  and g_39308_(_11974_, _11976_, _11996_);
  or g_39309_(_11973_, _11977_, _11997_);
  and g_39310_(_11995_, _11997_, _11998_);
  or g_39311_(_11994_, _11996_, _11999_);
  and g_39312_(_11992_, _11998_, _12000_);
  or g_39313_(_11993_, _11999_, _12002_);
  and g_39314_(_22142_, _11965_, _12003_);
  and g_39315_(_11856_, _11964_, _12004_);
  or g_39316_(_12003_, _12004_, _12005_);
  not g_39317_(_12005_, _12006_);
  and g_39318_(_22341_, _12005_, _12007_);
  or g_39319_(_22340_, _12006_, _12008_);
  and g_39320_(_22152_, _11965_, _12009_);
  or g_39321_(_22153_, _11964_, _12010_);
  and g_39322_(_11851_, _11964_, _12011_);
  not g_39323_(_12011_, _12013_);
  or g_39324_(_12009_, _12011_, _12014_);
  and g_39325_(_12010_, _12013_, _12015_);
  and g_39326_(_22328_, _12014_, _12016_);
  or g_39327_(_22327_, _12015_, _12017_);
  and g_39328_(_12008_, _12017_, _12018_);
  or g_39329_(_12007_, _12016_, _12019_);
  and g_39330_(_22327_, _12015_, _12020_);
  or g_39331_(_22328_, _12014_, _12021_);
  and g_39332_(_22340_, _12006_, _12022_);
  or g_39333_(_22341_, _12005_, _12024_);
  and g_39334_(_12021_, _12024_, _12025_);
  or g_39335_(_12019_, _12020_, _12026_);
  and g_39336_(_12018_, _12025_, _12027_);
  or g_39337_(_12022_, _12026_, _12028_);
  and g_39338_(_12000_, _12027_, _12029_);
  or g_39339_(_12002_, _12028_, _12030_);
  or g_39340_(_22178_, _11964_, _12031_);
  or g_39341_(_11875_, _11965_, _12032_);
  and g_39342_(_12031_, _12032_, _12033_);
  and g_39343_(_22275_, _12033_, _12035_);
  and g_39344_(_22040_, _11965_, _12036_);
  or g_39345_(_22041_, _11964_, _12037_);
  and g_39346_(_11893_, _11964_, _12038_);
  or g_39347_(_11892_, _11965_, _12039_);
  and g_39348_(_12037_, _12039_, _12040_);
  or g_39349_(_12036_, _12038_, _12041_);
  and g_39350_(_22282_, _12040_, _12042_);
  or g_39351_(_22283_, _12041_, _12043_);
  and g_39352_(_22267_, _11972_, _12044_);
  or g_39353_(_22267_, _11972_, _12046_);
  xor g_39354_(_22275_, _12033_, _12047_);
  xor g_39355_(_22274_, _12033_, _12048_);
  xor g_39356_(_22268_, _11971_, _12049_);
  xor g_39357_(_22267_, _11971_, _12050_);
  and g_39358_(_12047_, _12049_, _12051_);
  or g_39359_(_12048_, _12050_, _12052_);
  and g_39360_(_12043_, _12051_, _12053_);
  or g_39361_(_12042_, _12052_, _12054_);
  or g_39362_(_20536_, _11964_, _12055_);
  or g_39363_(_11903_, _11965_, _12057_);
  and g_39364_(_12055_, _12057_, _12058_);
  not g_39365_(_12058_, _12059_);
  and g_39366_(_22358_, _12058_, _12060_);
  or g_39367_(_22356_, _12059_, _12061_);
  and g_39368_(_22283_, _12041_, _12062_);
  or g_39369_(_22282_, _12040_, _12063_);
  and g_39370_(_12061_, _12063_, _12064_);
  or g_39371_(_12060_, _12062_, _12065_);
  and g_39372_(_22356_, _12059_, _12066_);
  or g_39373_(_22358_, _12058_, _12068_);
  and g_39374_(_12064_, _12068_, _12069_);
  or g_39375_(_12065_, _12066_, _12070_);
  and g_39376_(_12053_, _12069_, _12071_);
  or g_39377_(_12054_, _12070_, _12072_);
  or g_39378_(_20529_, _11964_, _12073_);
  or g_39379_(_11920_, _11965_, _12074_);
  and g_39380_(_12073_, _12074_, _12075_);
  and g_39381_(_20526_, _12075_, _12076_);
  not g_39382_(_12076_, _12077_);
  and g_39383_(_11927_, _11964_, _12079_);
  and g_39384_(_18127_, _11965_, _12080_);
  or g_39385_(_12079_, _12080_, _12081_);
  not g_39386_(_12081_, _12082_);
  or g_39387_(_18338_, _12081_, _12083_);
  or g_39388_(_20526_, _12075_, _12084_);
  and g_39389_(_12083_, _12084_, _12085_);
  or g_39390_(_12076_, _12085_, _12086_);
  not g_39391_(_12086_, _12087_);
  and g_39392_(_18338_, _12081_, _12088_);
  or g_39393_(_18337_, _12082_, _12090_);
  and g_39394_(_12077_, _12090_, _12091_);
  or g_39395_(_12076_, _12088_, _12092_);
  and g_39396_(out[129], _11965_, _12093_);
  and g_39397_(_11916_, _11964_, _12094_);
  or g_39398_(_12093_, _12094_, _12095_);
  or g_39399_(_21103_, _12095_, _12096_);
  not g_39400_(_12096_, _12097_);
  and g_39401_(_11934_, _11964_, _12098_);
  not g_39402_(_12098_, _12099_);
  or g_39403_(out[128], _11964_, _12101_);
  not g_39404_(_12101_, _12102_);
  and g_39405_(_12099_, _12101_, _12103_);
  or g_39406_(_12098_, _12102_, _12104_);
  and g_39407_(out[144], _12104_, _12105_);
  or g_39408_(_21114_, _12103_, _12106_);
  xor g_39409_(_21103_, _12095_, _12107_);
  xor g_39410_(out[145], _12095_, _12108_);
  and g_39411_(_12106_, _12107_, _12109_);
  or g_39412_(_12105_, _12108_, _12110_);
  and g_39413_(_12096_, _12110_, _12112_);
  or g_39414_(_12097_, _12109_, _12113_);
  and g_39415_(_12091_, _12113_, _12114_);
  or g_39416_(_12092_, _12112_, _12115_);
  and g_39417_(_12086_, _12115_, _12116_);
  or g_39418_(_12087_, _12114_, _12117_);
  and g_39419_(_12071_, _12117_, _12118_);
  or g_39420_(_12072_, _12116_, _12119_);
  and g_39421_(_12053_, _12065_, _12120_);
  or g_39422_(_12054_, _12064_, _12121_);
  or g_39423_(_12035_, _12044_, _12123_);
  and g_39424_(_12046_, _12123_, _12124_);
  not g_39425_(_12124_, _12125_);
  and g_39426_(_12121_, _12125_, _12126_);
  or g_39427_(_12120_, _12124_, _12127_);
  and g_39428_(_12119_, _12126_, _12128_);
  or g_39429_(_12118_, _12127_, _12129_);
  and g_39430_(_12029_, _12129_, _12130_);
  or g_39431_(_12030_, _12128_, _12131_);
  and g_39432_(_11993_, _11997_, _12132_);
  or g_39433_(_11992_, _11996_, _12134_);
  and g_39434_(_12019_, _12024_, _12135_);
  or g_39435_(_12002_, _12018_, _12136_);
  and g_39436_(_12000_, _12135_, _12137_);
  or g_39437_(_12022_, _12136_, _12138_);
  and g_39438_(_12134_, _12138_, _12139_);
  or g_39439_(_12132_, _12137_, _12140_);
  and g_39440_(_12131_, _12139_, _12141_);
  or g_39441_(_12130_, _12140_, _12142_);
  and g_39442_(_21114_, _12103_, _12143_);
  not g_39443_(_12143_, _12145_);
  and g_39444_(_12085_, _12145_, _12146_);
  and g_39445_(_12091_, _12146_, _12147_);
  and g_39446_(_12109_, _12147_, _12148_);
  not g_39447_(_12148_, _12149_);
  and g_39448_(_12071_, _12148_, _12150_);
  or g_39449_(_12030_, _12072_, _12151_);
  and g_39450_(_12029_, _12150_, _12152_);
  or g_39451_(_12149_, _12151_, _12153_);
  and g_39452_(_12142_, _12153_, _12154_);
  or g_39453_(_12141_, _12152_, _12156_);
  and g_39454_(_11972_, _12156_, _12157_);
  or g_39455_(_11971_, _12154_, _12158_);
  and g_39456_(_22268_, _12154_, _12159_);
  not g_39457_(_12159_, _12160_);
  and g_39458_(_12158_, _12160_, _12161_);
  or g_39459_(_12157_, _12159_, _12162_);
  or g_39460_(out[202], _22625_, _12163_);
  xor g_39461_(out[203], _12163_, _12164_);
  xor g_39462_(_18848_, _12163_, _12165_);
  or g_39463_(out[186], _22492_, _12167_);
  xor g_39464_(out[187], _12167_, _12168_);
  not g_39465_(_12168_, _12169_);
  or g_39466_(out[170], _22488_, _12170_);
  xor g_39467_(out[171], _12170_, _12171_);
  not g_39468_(_12171_, _12172_);
  and g_39469_(_12168_, _12172_, _12173_);
  or g_39470_(_12169_, _12171_, _12174_);
  xor g_39471_(out[186], _22492_, _12175_);
  xor g_39472_(_18837_, _22492_, _12176_);
  xor g_39473_(out[170], _22488_, _12178_);
  xor g_39474_(_18705_, _22488_, _12179_);
  and g_39475_(_12175_, _12179_, _12180_);
  or g_39476_(_12176_, _12178_, _12181_);
  and g_39477_(_12176_, _12178_, _12182_);
  or g_39478_(_12175_, _12179_, _12183_);
  and g_39479_(_22498_, _22595_, _12184_);
  or g_39480_(_22497_, _22594_, _12185_);
  and g_39481_(_12183_, _12185_, _12186_);
  or g_39482_(_12182_, _12184_, _12187_);
  and g_39483_(_12181_, _12187_, _12189_);
  or g_39484_(_12180_, _12186_, _12190_);
  and g_39485_(_12169_, _12171_, _12191_);
  or g_39486_(_12168_, _12172_, _12192_);
  and g_39487_(_12189_, _12192_, _12193_);
  or g_39488_(_12190_, _12191_, _12194_);
  and g_39489_(_12174_, _12194_, _12195_);
  or g_39490_(_12173_, _12193_, _12196_);
  and g_39491_(_22593_, _12196_, _12197_);
  or g_39492_(_22592_, _12195_, _12198_);
  and g_39493_(_22573_, _12198_, _12200_);
  or g_39494_(_22572_, _12197_, _12201_);
  or g_39495_(_12168_, _12201_, _12202_);
  or g_39496_(_12171_, _12200_, _12203_);
  and g_39497_(_12202_, _12203_, _12204_);
  not g_39498_(_12204_, _12205_);
  and g_39499_(_12164_, _12204_, _12206_);
  or g_39500_(_12165_, _12205_, _12207_);
  or g_39501_(out[218], _22919_, _12208_);
  xor g_39502_(out[219], _12208_, _12209_);
  xor g_39503_(_18958_, _12208_, _12211_);
  and g_39504_(_12206_, _12209_, _12212_);
  or g_39505_(_12207_, _12211_, _12213_);
  or g_39506_(out[234], _23068_, _12214_);
  xor g_39507_(out[235], _12214_, _12215_);
  xor g_39508_(_19090_, _12214_, _12216_);
  and g_39509_(_12212_, _12215_, _12217_);
  or g_39510_(_12213_, _12216_, _12218_);
  or g_39511_(out[250], _23280_, _12219_);
  xor g_39512_(out[251], _12219_, _12220_);
  xor g_39513_(_19222_, _12219_, _12222_);
  and g_39514_(_12217_, _12220_, _12223_);
  or g_39515_(_12218_, _12222_, _12224_);
  or g_39516_(out[266], _23565_, _12225_);
  xor g_39517_(out[267], _12225_, _12226_);
  xor g_39518_(_19354_, _12225_, _12227_);
  and g_39519_(_12223_, _12226_, _12228_);
  or g_39520_(_12224_, _12227_, _12229_);
  or g_39521_(out[282], _23690_, _12230_);
  xor g_39522_(out[283], _12230_, _12231_);
  xor g_39523_(_19486_, _12230_, _12233_);
  and g_39524_(_12228_, _12231_, _12234_);
  not g_39525_(_12234_, _12235_);
  or g_39526_(out[298], _23894_, _12236_);
  xor g_39527_(out[299], _12236_, _12237_);
  not g_39528_(_12237_, _12238_);
  and g_39529_(_12235_, _12237_, _12239_);
  or g_39530_(_12234_, _12238_, _12240_);
  xor g_39531_(out[282], _23690_, _12241_);
  xor g_39532_(_19607_, _23690_, _12242_);
  xor g_39533_(out[250], _23280_, _12244_);
  xor g_39534_(_19343_, _23280_, _12245_);
  xor g_39535_(out[234], _23068_, _12246_);
  xor g_39536_(out[218], _22919_, _12247_);
  xor g_39537_(_19079_, _22919_, _12248_);
  xor g_39538_(out[202], _22625_, _12249_);
  not g_39539_(_12249_, _12250_);
  or g_39540_(_22521_, _12200_, _12251_);
  or g_39541_(_22524_, _12201_, _12252_);
  and g_39542_(_12251_, _12252_, _12253_);
  and g_39543_(_22553_, _12200_, _12255_);
  or g_39544_(_22552_, _12201_, _12256_);
  and g_39545_(_22551_, _12201_, _12257_);
  or g_39546_(_22550_, _12200_, _12258_);
  and g_39547_(_12256_, _12258_, _12259_);
  or g_39548_(_12255_, _12257_, _12260_);
  and g_39549_(_22700_, _12260_, _12261_);
  or g_39550_(_22701_, _12259_, _12262_);
  or g_39551_(_22528_, _12201_, _12263_);
  or g_39552_(_22527_, _12200_, _12264_);
  and g_39553_(_12263_, _12264_, _12266_);
  not g_39554_(_12266_, _12267_);
  and g_39555_(_22666_, _12266_, _12268_);
  or g_39556_(_22666_, _12266_, _12269_);
  and g_39557_(_22677_, _12253_, _12270_);
  xor g_39558_(_22666_, _12266_, _12271_);
  xor g_39559_(_22667_, _12266_, _12272_);
  xor g_39560_(_22677_, _12253_, _12273_);
  xor g_39561_(_22675_, _12253_, _12274_);
  and g_39562_(_12271_, _12273_, _12275_);
  or g_39563_(_12272_, _12274_, _12277_);
  and g_39564_(_12262_, _12275_, _12278_);
  or g_39565_(_12261_, _12277_, _12279_);
  and g_39566_(_22547_, _12200_, _12280_);
  or g_39567_(_22546_, _12201_, _12281_);
  and g_39568_(_22542_, _12201_, _12282_);
  or g_39569_(_22541_, _12200_, _12283_);
  and g_39570_(_12281_, _12283_, _12284_);
  or g_39571_(_12280_, _12282_, _12285_);
  and g_39572_(_22690_, _12284_, _12286_);
  or g_39573_(_22689_, _12285_, _12288_);
  and g_39574_(_22701_, _12259_, _12289_);
  or g_39575_(_22700_, _12260_, _12290_);
  and g_39576_(_12288_, _12290_, _12291_);
  or g_39577_(_12286_, _12289_, _12292_);
  and g_39578_(_22689_, _12285_, _12293_);
  or g_39579_(_22690_, _12284_, _12294_);
  and g_39580_(_12291_, _12294_, _12295_);
  or g_39581_(_12292_, _12293_, _12296_);
  and g_39582_(_12278_, _12295_, _12297_);
  or g_39583_(_12279_, _12296_, _12299_);
  or g_39584_(_12176_, _12201_, _12300_);
  or g_39585_(_12179_, _12200_, _12301_);
  and g_39586_(_12300_, _12301_, _12302_);
  or g_39587_(_12165_, _12204_, _12303_);
  and g_39588_(_12249_, _12302_, _12304_);
  and g_39589_(_12165_, _12204_, _12305_);
  and g_39590_(_22493_, _12200_, _12306_);
  or g_39591_(_22494_, _12201_, _12307_);
  and g_39592_(_22490_, _12201_, _12308_);
  or g_39593_(_22491_, _12200_, _12310_);
  and g_39594_(_12307_, _12310_, _12311_);
  or g_39595_(_12306_, _12308_, _12312_);
  or g_39596_(_22627_, _12312_, _12313_);
  or g_39597_(_22502_, _12200_, _12314_);
  or g_39598_(_22504_, _12201_, _12315_);
  and g_39599_(_12314_, _12315_, _12316_);
  not g_39600_(_12316_, _12317_);
  and g_39601_(_22627_, _12312_, _12318_);
  and g_39602_(_22647_, _12316_, _12319_);
  or g_39603_(_12318_, _12319_, _12321_);
  xor g_39604_(_22626_, _12311_, _12322_);
  xor g_39605_(_22627_, _12311_, _12323_);
  xor g_39606_(_12249_, _12302_, _12324_);
  xor g_39607_(_12250_, _12302_, _12325_);
  xor g_39608_(_12165_, _12204_, _12326_);
  xor g_39609_(_12164_, _12204_, _12327_);
  and g_39610_(_12324_, _12326_, _12328_);
  or g_39611_(_12325_, _12327_, _12329_);
  xor g_39612_(_22647_, _12316_, _12330_);
  xor g_39613_(_22646_, _12316_, _12332_);
  and g_39614_(_12328_, _12330_, _12333_);
  or g_39615_(_12329_, _12332_, _12334_);
  and g_39616_(_12322_, _12333_, _12335_);
  or g_39617_(_12323_, _12334_, _12336_);
  and g_39618_(_12297_, _12335_, _12337_);
  or g_39619_(_12299_, _12336_, _12338_);
  and g_39620_(out[177], _12200_, _12339_);
  or g_39621_(_18771_, _12201_, _12340_);
  and g_39622_(out[161], _12201_, _12341_);
  or g_39623_(_18650_, _12200_, _12343_);
  and g_39624_(_12340_, _12343_, _12344_);
  or g_39625_(_12339_, _12341_, _12345_);
  and g_39626_(_18584_, _12201_, _12346_);
  or g_39627_(out[160], _12200_, _12347_);
  and g_39628_(_18782_, _12200_, _12348_);
  or g_39629_(out[176], _12201_, _12349_);
  and g_39630_(_12347_, _12349_, _12350_);
  or g_39631_(_12346_, _12348_, _12351_);
  and g_39632_(out[192], _12351_, _12352_);
  or g_39633_(_18914_, _12350_, _12354_);
  and g_39634_(out[193], _12344_, _12355_);
  or g_39635_(_18903_, _12345_, _12356_);
  xor g_39636_(out[193], _12344_, _12357_);
  xor g_39637_(_18903_, _12344_, _12358_);
  and g_39638_(_12354_, _12357_, _12359_);
  or g_39639_(_12352_, _12358_, _12360_);
  and g_39640_(_18465_, _12200_, _12361_);
  and g_39641_(_18468_, _12201_, _12362_);
  or g_39642_(_12361_, _12362_, _12363_);
  not g_39643_(_12363_, _12365_);
  or g_39644_(_18743_, _12363_, _12366_);
  xor g_39645_(_18743_, _12363_, _12367_);
  xor g_39646_(_18742_, _12363_, _12368_);
  and g_39647_(_22576_, _12200_, _12369_);
  or g_39648_(_22578_, _12201_, _12370_);
  and g_39649_(_22574_, _12201_, _12371_);
  or g_39650_(_22575_, _12200_, _12372_);
  and g_39651_(_12370_, _12372_, _12373_);
  or g_39652_(_12369_, _12371_, _12374_);
  and g_39653_(_22727_, _12374_, _12376_);
  or g_39654_(_22727_, _12374_, _12377_);
  xor g_39655_(_22726_, _12373_, _12378_);
  xor g_39656_(_22727_, _12373_, _12379_);
  and g_39657_(_18914_, _12350_, _12380_);
  or g_39658_(_12379_, _12380_, _12381_);
  or g_39659_(_12368_, _12381_, _12382_);
  not g_39660_(_12382_, _12383_);
  and g_39661_(_12359_, _12383_, _12384_);
  or g_39662_(_12360_, _12382_, _12385_);
  and g_39663_(_12367_, _12378_, _12387_);
  or g_39664_(_12368_, _12379_, _12388_);
  and g_39665_(_12337_, _12384_, _12389_);
  or g_39666_(_12338_, _12385_, _12390_);
  and g_39667_(_12366_, _12377_, _12391_);
  and g_39668_(_12356_, _12360_, _12392_);
  or g_39669_(_12355_, _12359_, _12393_);
  and g_39670_(_12387_, _12393_, _12394_);
  or g_39671_(_12388_, _12392_, _12395_);
  or g_39672_(_12376_, _12391_, _12396_);
  not g_39673_(_12396_, _12398_);
  and g_39674_(_12395_, _12396_, _12399_);
  or g_39675_(_12394_, _12398_, _12400_);
  and g_39676_(_12337_, _12400_, _12401_);
  or g_39677_(_12338_, _12399_, _12402_);
  and g_39678_(_12321_, _12328_, _12403_);
  and g_39679_(_12313_, _12403_, _12404_);
  not g_39680_(_12404_, _12405_);
  and g_39681_(_12303_, _12304_, _12406_);
  or g_39682_(_12305_, _12406_, _12407_);
  not g_39683_(_12407_, _12409_);
  and g_39684_(_12405_, _12409_, _12410_);
  or g_39685_(_12404_, _12407_, _12411_);
  and g_39686_(_12278_, _12292_, _12412_);
  or g_39687_(_12279_, _12291_, _12413_);
  and g_39688_(_12269_, _12270_, _12414_);
  or g_39689_(_12268_, _12414_, _12415_);
  not g_39690_(_12415_, _12416_);
  and g_39691_(_12413_, _12416_, _12417_);
  or g_39692_(_12412_, _12415_, _12418_);
  and g_39693_(_12335_, _12418_, _12420_);
  or g_39694_(_12336_, _12417_, _12421_);
  and g_39695_(_12402_, _12410_, _12422_);
  or g_39696_(_12401_, _12411_, _12423_);
  and g_39697_(_12421_, _12422_, _12424_);
  or g_39698_(_12420_, _12423_, _12425_);
  and g_39699_(_12390_, _12425_, _12426_);
  or g_39700_(_12389_, _12424_, _12427_);
  and g_39701_(_12249_, _12426_, _12428_);
  not g_39702_(_12428_, _12429_);
  or g_39703_(_12302_, _12426_, _12431_);
  not g_39704_(_12431_, _12432_);
  and g_39705_(_12429_, _12431_, _12433_);
  or g_39706_(_12428_, _12432_, _12434_);
  and g_39707_(_12247_, _12433_, _12435_);
  or g_39708_(_12248_, _12434_, _12436_);
  and g_39709_(_12206_, _12211_, _12437_);
  or g_39710_(_12207_, _12209_, _12438_);
  and g_39711_(_12436_, _12438_, _12439_);
  or g_39712_(_12435_, _12437_, _12440_);
  and g_39713_(_12207_, _12209_, _12442_);
  or g_39714_(_12206_, _12211_, _12443_);
  and g_39715_(_12248_, _12434_, _12444_);
  or g_39716_(_12247_, _12433_, _12445_);
  and g_39717_(_12443_, _12445_, _12446_);
  or g_39718_(_12442_, _12444_, _12447_);
  and g_39719_(_12439_, _12446_, _12448_);
  or g_39720_(_12440_, _12447_, _12449_);
  and g_39721_(_22626_, _12426_, _12450_);
  not g_39722_(_12450_, _12451_);
  or g_39723_(_12311_, _12426_, _12453_);
  not g_39724_(_12453_, _12454_);
  and g_39725_(_12451_, _12453_, _12455_);
  or g_39726_(_12450_, _12454_, _12456_);
  and g_39727_(_22921_, _12456_, _12457_);
  or g_39728_(_22920_, _12455_, _12458_);
  and g_39729_(_22646_, _12426_, _12459_);
  not g_39730_(_12459_, _12460_);
  and g_39731_(_12316_, _12427_, _12461_);
  or g_39732_(_12317_, _12426_, _12462_);
  and g_39733_(_12460_, _12462_, _12464_);
  or g_39734_(_12459_, _12461_, _12465_);
  and g_39735_(_22906_, _12465_, _12466_);
  or g_39736_(_22905_, _12464_, _12467_);
  and g_39737_(_12458_, _12467_, _12468_);
  or g_39738_(_12457_, _12466_, _12469_);
  and g_39739_(_22920_, _12455_, _12470_);
  or g_39740_(_22921_, _12456_, _12471_);
  and g_39741_(_22905_, _12464_, _12472_);
  or g_39742_(_22906_, _12465_, _12473_);
  and g_39743_(_12471_, _12473_, _12475_);
  or g_39744_(_12470_, _12472_, _12476_);
  and g_39745_(_12468_, _12475_, _12477_);
  or g_39746_(_12469_, _12476_, _12478_);
  and g_39747_(_12448_, _12477_, _12479_);
  or g_39748_(_12449_, _12478_, _12480_);
  or g_39749_(_22666_, _12427_, _12481_);
  or g_39750_(_12267_, _12426_, _12482_);
  and g_39751_(_12481_, _12482_, _12483_);
  not g_39752_(_12483_, _12484_);
  and g_39753_(_22843_, _12483_, _12486_);
  or g_39754_(_22842_, _12484_, _12487_);
  and g_39755_(_22689_, _12426_, _12488_);
  or g_39756_(_22690_, _12427_, _12489_);
  and g_39757_(_12284_, _12427_, _12490_);
  or g_39758_(_12285_, _12426_, _12491_);
  and g_39759_(_12489_, _12491_, _12492_);
  or g_39760_(_12488_, _12490_, _12493_);
  and g_39761_(_22861_, _12493_, _12494_);
  or g_39762_(_22860_, _12492_, _12495_);
  and g_39763_(_22700_, _12426_, _12497_);
  or g_39764_(_22701_, _12427_, _12498_);
  and g_39765_(_12259_, _12427_, _12499_);
  or g_39766_(_12260_, _12426_, _12500_);
  and g_39767_(_12498_, _12500_, _12501_);
  or g_39768_(_12497_, _12499_, _12502_);
  and g_39769_(_22834_, _12502_, _12503_);
  or g_39770_(_22833_, _12501_, _12504_);
  and g_39771_(_12495_, _12504_, _12505_);
  or g_39772_(_12494_, _12503_, _12506_);
  or g_39773_(_22675_, _12427_, _12508_);
  or g_39774_(_12253_, _12426_, _12509_);
  and g_39775_(_12508_, _12509_, _12510_);
  and g_39776_(_22827_, _12510_, _12511_);
  not g_39777_(_12511_, _12512_);
  xor g_39778_(_22827_, _12510_, _12513_);
  xor g_39779_(_22826_, _12510_, _12514_);
  and g_39780_(_22842_, _12484_, _12515_);
  or g_39781_(_22843_, _12483_, _12516_);
  and g_39782_(_22833_, _12501_, _12517_);
  or g_39783_(_22834_, _12502_, _12519_);
  and g_39784_(_12487_, _12516_, _12520_);
  or g_39785_(_12486_, _12515_, _12521_);
  and g_39786_(_12513_, _12520_, _12522_);
  or g_39787_(_12514_, _12521_, _12523_);
  and g_39788_(_12519_, _12522_, _12524_);
  or g_39789_(_12517_, _12523_, _12525_);
  and g_39790_(_12506_, _12524_, _12526_);
  or g_39791_(_12505_, _12525_, _12527_);
  and g_39792_(_12487_, _12511_, _12528_);
  or g_39793_(_12486_, _12512_, _12530_);
  and g_39794_(_12516_, _12530_, _12531_);
  or g_39795_(_12515_, _12528_, _12532_);
  or g_39796_(_12526_, _12532_, _12533_);
  and g_39797_(_12527_, _12531_, _12534_);
  and g_39798_(_22860_, _12492_, _12535_);
  or g_39799_(_22861_, _12493_, _12536_);
  and g_39800_(_12505_, _12536_, _12537_);
  or g_39801_(_12506_, _12535_, _12538_);
  and g_39802_(_12524_, _12537_, _12539_);
  or g_39803_(_12525_, _12538_, _12541_);
  and g_39804_(out[193], _12426_, _12542_);
  or g_39805_(_18903_, _12427_, _12543_);
  and g_39806_(_12345_, _12427_, _12544_);
  or g_39807_(_12344_, _12426_, _12545_);
  and g_39808_(_12543_, _12545_, _12546_);
  or g_39809_(_12542_, _12544_, _12547_);
  and g_39810_(out[209], _12546_, _12548_);
  or g_39811_(_19013_, _12547_, _12549_);
  xor g_39812_(out[209], _12546_, _12550_);
  and g_39813_(_18742_, _12426_, _12552_);
  or g_39814_(_18743_, _12427_, _12553_);
  and g_39815_(_12363_, _12427_, _12554_);
  or g_39816_(_12365_, _12426_, _12555_);
  and g_39817_(_12553_, _12555_, _12556_);
  or g_39818_(_12552_, _12554_, _12557_);
  and g_39819_(_18851_, _12557_, _12558_);
  or g_39820_(_18850_, _12556_, _12559_);
  and g_39821_(_12550_, _12559_, _12560_);
  not g_39822_(_12560_, _12561_);
  and g_39823_(_18850_, _12556_, _12563_);
  or g_39824_(_18851_, _12557_, _12564_);
  and g_39825_(_22727_, _12426_, _12565_);
  or g_39826_(_22726_, _12427_, _12566_);
  and g_39827_(_12373_, _12427_, _12567_);
  or g_39828_(_12374_, _12426_, _12568_);
  and g_39829_(_12566_, _12568_, _12569_);
  or g_39830_(_12565_, _12567_, _12570_);
  and g_39831_(_22963_, _12570_, _12571_);
  or g_39832_(_22964_, _12569_, _12572_);
  and g_39833_(_12564_, _12572_, _12574_);
  or g_39834_(_12563_, _12571_, _12575_);
  or g_39835_(_12350_, _12426_, _12576_);
  not g_39836_(_12576_, _12577_);
  and g_39837_(_18914_, _12426_, _12578_);
  or g_39838_(out[192], _12427_, _12579_);
  and g_39839_(_12576_, _12579_, _12580_);
  or g_39840_(_12577_, _12578_, _12581_);
  and g_39841_(out[208], _12581_, _12582_);
  or g_39842_(_19024_, _12580_, _12583_);
  and g_39843_(_22964_, _12569_, _12585_);
  or g_39844_(_22963_, _12570_, _12586_);
  and g_39845_(_12583_, _12586_, _12587_);
  or g_39846_(_12582_, _12585_, _12588_);
  and g_39847_(_12574_, _12587_, _12589_);
  or g_39848_(_12575_, _12588_, _12590_);
  and g_39849_(_12560_, _12589_, _12591_);
  or g_39850_(_12561_, _12590_, _12592_);
  and g_39851_(_12548_, _12559_, _12593_);
  or g_39852_(_12549_, _12558_, _12594_);
  and g_39853_(_12574_, _12594_, _12596_);
  or g_39854_(_12575_, _12593_, _12597_);
  and g_39855_(_12586_, _12597_, _12598_);
  or g_39856_(_12585_, _12596_, _12599_);
  and g_39857_(_12592_, _12599_, _12600_);
  or g_39858_(_12591_, _12598_, _12601_);
  and g_39859_(_12539_, _12601_, _12602_);
  or g_39860_(_12541_, _12600_, _12603_);
  and g_39861_(_12539_, _12591_, _12604_);
  or g_39862_(_12541_, _12592_, _12605_);
  and g_39863_(_12534_, _12603_, _12607_);
  or g_39864_(_12533_, _12602_, _12608_);
  and g_39865_(_12479_, _12608_, _12609_);
  or g_39866_(_12480_, _12607_, _12610_);
  and g_39867_(_12469_, _12471_, _12611_);
  or g_39868_(_12468_, _12470_, _12612_);
  and g_39869_(_12448_, _12611_, _12613_);
  or g_39870_(_12449_, _12612_, _12614_);
  and g_39871_(_12440_, _12443_, _12615_);
  or g_39872_(_12439_, _12442_, _12616_);
  and g_39873_(_12614_, _12616_, _12618_);
  or g_39874_(_12613_, _12615_, _12619_);
  and g_39875_(_12610_, _12618_, _12620_);
  or g_39876_(_12609_, _12619_, _12621_);
  and g_39877_(_19024_, _12580_, _12622_);
  or g_39878_(out[208], _12581_, _12623_);
  and g_39879_(_12479_, _12623_, _12624_);
  or g_39880_(_12480_, _12622_, _12625_);
  and g_39881_(_12604_, _12624_, _12626_);
  or g_39882_(_12605_, _12625_, _12627_);
  and g_39883_(_12621_, _12627_, _12629_);
  or g_39884_(_12620_, _12626_, _12630_);
  or g_39885_(_12248_, _12630_, _12631_);
  not g_39886_(_12631_, _12632_);
  and g_39887_(_12434_, _12630_, _12633_);
  not g_39888_(_12633_, _12634_);
  and g_39889_(_12631_, _12634_, _12635_);
  or g_39890_(_12632_, _12633_, _12636_);
  and g_39891_(_12246_, _12635_, _12637_);
  and g_39892_(_12212_, _12216_, _12638_);
  or g_39893_(_12212_, _12216_, _12640_);
  xor g_39894_(_12212_, _12216_, _12641_);
  or g_39895_(_22921_, _12630_, _12642_);
  not g_39896_(_12642_, _12643_);
  and g_39897_(_12456_, _12630_, _12644_);
  not g_39898_(_12644_, _12645_);
  and g_39899_(_12642_, _12645_, _12646_);
  or g_39900_(_12643_, _12644_, _12647_);
  or g_39901_(_23070_, _12647_, _12648_);
  xor g_39902_(_12246_, _12635_, _12649_);
  and g_39903_(_12641_, _12649_, _12651_);
  and g_39904_(_12648_, _12651_, _12652_);
  and g_39905_(_23070_, _12647_, _12653_);
  or g_39906_(_23069_, _12646_, _12654_);
  or g_39907_(_22906_, _12630_, _12655_);
  not g_39908_(_12655_, _12656_);
  and g_39909_(_12465_, _12630_, _12657_);
  not g_39910_(_12657_, _12658_);
  and g_39911_(_12655_, _12658_, _12659_);
  or g_39912_(_12656_, _12657_, _12660_);
  and g_39913_(_23079_, _12660_, _12662_);
  or g_39914_(_23078_, _12659_, _12663_);
  and g_39915_(_12654_, _12663_, _12664_);
  or g_39916_(_12653_, _12662_, _12665_);
  or g_39917_(_23079_, _12660_, _12666_);
  and g_39918_(_12664_, _12666_, _12667_);
  and g_39919_(_12652_, _12667_, _12668_);
  or g_39920_(_22842_, _12630_, _12669_);
  or g_39921_(_12483_, _12629_, _12670_);
  and g_39922_(_12669_, _12670_, _12671_);
  or g_39923_(_23101_, _12671_, _12673_);
  and g_39924_(_23101_, _12671_, _12674_);
  xor g_39925_(_23100_, _12671_, _12675_);
  or g_39926_(_22826_, _12630_, _12676_);
  or g_39927_(_12510_, _12629_, _12677_);
  and g_39928_(_12676_, _12677_, _12678_);
  not g_39929_(_12678_, _12679_);
  or g_39930_(_23107_, _12679_, _12680_);
  or g_39931_(_22834_, _12630_, _12681_);
  not g_39932_(_12681_, _12682_);
  and g_39933_(_12502_, _12630_, _12684_);
  not g_39934_(_12684_, _12685_);
  and g_39935_(_12681_, _12685_, _12686_);
  or g_39936_(_12682_, _12684_, _12687_);
  and g_39937_(_23131_, _12686_, _12688_);
  xor g_39938_(_23107_, _12678_, _12689_);
  or g_39939_(_12675_, _12689_, _12690_);
  or g_39940_(_12688_, _12690_, _12691_);
  not g_39941_(_12691_, _12692_);
  or g_39942_(_22861_, _12630_, _12693_);
  not g_39943_(_12693_, _12695_);
  and g_39944_(_12493_, _12630_, _12696_);
  not g_39945_(_12696_, _12697_);
  and g_39946_(_12693_, _12697_, _12698_);
  or g_39947_(_12695_, _12696_, _12699_);
  or g_39948_(_23123_, _12698_, _12700_);
  or g_39949_(_23131_, _12686_, _12701_);
  and g_39950_(_12700_, _12701_, _12702_);
  or g_39951_(_23124_, _12699_, _12703_);
  and g_39952_(_12702_, _12703_, _12704_);
  and g_39953_(_12692_, _12704_, _12706_);
  or g_39954_(_19013_, _12630_, _12707_);
  or g_39955_(_12546_, _12629_, _12708_);
  and g_39956_(_12707_, _12708_, _12709_);
  and g_39957_(out[225], _12709_, _12710_);
  and g_39958_(_22964_, _12629_, _12711_);
  or g_39959_(_22963_, _12630_, _12712_);
  and g_39960_(_12570_, _12630_, _12713_);
  or g_39961_(_12569_, _12629_, _12714_);
  and g_39962_(_12712_, _12714_, _12715_);
  or g_39963_(_12711_, _12713_, _12717_);
  and g_39964_(_23154_, _12715_, _12718_);
  not g_39965_(_12718_, _12719_);
  or g_39966_(_12556_, _12629_, _12720_);
  or g_39967_(_18851_, _12630_, _12721_);
  and g_39968_(_12720_, _12721_, _12722_);
  and g_39969_(_19230_, _12722_, _12723_);
  and g_39970_(_23153_, _12717_, _12724_);
  xor g_39971_(_23154_, _12715_, _12725_);
  xor g_39972_(_19230_, _12722_, _12726_);
  and g_39973_(_12725_, _12726_, _12728_);
  and g_39974_(_12710_, _12728_, _12729_);
  xor g_39975_(out[225], _12709_, _12730_);
  and g_39976_(_12581_, _12630_, _12731_);
  not g_39977_(_12731_, _12732_);
  or g_39978_(out[208], _12630_, _12733_);
  not g_39979_(_12733_, _12734_);
  and g_39980_(_12732_, _12733_, _12735_);
  or g_39981_(_12731_, _12734_, _12736_);
  or g_39982_(_19156_, _12735_, _12737_);
  and g_39983_(_12730_, _12737_, _12739_);
  and g_39984_(_12728_, _12739_, _12740_);
  or g_39985_(_12723_, _12724_, _12741_);
  and g_39986_(_12719_, _12741_, _12742_);
  or g_39987_(_12729_, _12742_, _12743_);
  or g_39988_(_12740_, _12743_, _12744_);
  and g_39989_(_12706_, _12744_, _12745_);
  or g_39990_(_12691_, _12702_, _12746_);
  or g_39991_(_12674_, _12680_, _12747_);
  and g_39992_(_12673_, _12747_, _12748_);
  and g_39993_(_12746_, _12748_, _12750_);
  not g_39994_(_12750_, _12751_);
  or g_39995_(_12745_, _12751_, _12752_);
  and g_39996_(_12668_, _12752_, _12753_);
  and g_39997_(_12652_, _12665_, _12754_);
  and g_39998_(_12637_, _12640_, _12755_);
  or g_39999_(_12638_, _12755_, _12756_);
  or g_40000_(_12754_, _12756_, _12757_);
  or g_40001_(_12753_, _12757_, _12758_);
  or g_40002_(out[224], _12736_, _12759_);
  and g_40003_(_12668_, _12759_, _12761_);
  and g_40004_(_12706_, _12761_, _12762_);
  and g_40005_(_12740_, _12762_, _12763_);
  not g_40006_(_12763_, _12764_);
  and g_40007_(_12758_, _12764_, _12765_);
  not g_40008_(_12765_, _12766_);
  and g_40009_(_12246_, _12765_, _12767_);
  not g_40010_(_12767_, _12768_);
  and g_40011_(_12636_, _12766_, _12769_);
  or g_40012_(_12635_, _12765_, _12770_);
  and g_40013_(_12768_, _12770_, _12772_);
  or g_40014_(_12767_, _12769_, _12773_);
  and g_40015_(_12244_, _12772_, _12774_);
  or g_40016_(_12245_, _12773_, _12775_);
  and g_40017_(_12217_, _12222_, _12776_);
  or g_40018_(_12218_, _12220_, _12777_);
  and g_40019_(_12775_, _12777_, _12778_);
  or g_40020_(_12774_, _12776_, _12779_);
  and g_40021_(_12218_, _12220_, _12780_);
  or g_40022_(_12217_, _12222_, _12781_);
  and g_40023_(_12245_, _12773_, _12783_);
  or g_40024_(_12244_, _12772_, _12784_);
  and g_40025_(_12781_, _12784_, _12785_);
  or g_40026_(_12780_, _12783_, _12786_);
  and g_40027_(_12778_, _12785_, _12787_);
  or g_40028_(_12779_, _12786_, _12788_);
  and g_40029_(_23069_, _12765_, _12789_);
  not g_40030_(_12789_, _12790_);
  and g_40031_(_12647_, _12766_, _12791_);
  or g_40032_(_12646_, _12765_, _12792_);
  and g_40033_(_12790_, _12792_, _12794_);
  or g_40034_(_12789_, _12791_, _12795_);
  and g_40035_(_23283_, _12795_, _12796_);
  or g_40036_(_23282_, _12794_, _12797_);
  and g_40037_(_23078_, _12765_, _12798_);
  not g_40038_(_12798_, _12799_);
  and g_40039_(_12660_, _12766_, _12800_);
  or g_40040_(_12659_, _12765_, _12801_);
  and g_40041_(_12799_, _12801_, _12802_);
  or g_40042_(_12798_, _12800_, _12803_);
  and g_40043_(_23271_, _12803_, _12805_);
  or g_40044_(_23269_, _12802_, _12806_);
  and g_40045_(_12797_, _12806_, _12807_);
  or g_40046_(_12796_, _12805_, _12808_);
  and g_40047_(_23282_, _12794_, _12809_);
  or g_40048_(_23283_, _12795_, _12810_);
  and g_40049_(_23269_, _12802_, _12811_);
  or g_40050_(_23271_, _12803_, _12812_);
  and g_40051_(_12810_, _12812_, _12813_);
  or g_40052_(_12809_, _12811_, _12814_);
  and g_40053_(_12807_, _12813_, _12816_);
  or g_40054_(_12808_, _12814_, _12817_);
  and g_40055_(_12787_, _12816_, _12818_);
  or g_40056_(_12788_, _12817_, _12819_);
  and g_40057_(_23101_, _12765_, _12820_);
  not g_40058_(_12820_, _12821_);
  or g_40059_(_12671_, _12765_, _12822_);
  not g_40060_(_12822_, _12823_);
  and g_40061_(_12821_, _12822_, _12824_);
  or g_40062_(_12820_, _12823_, _12825_);
  and g_40063_(_23315_, _12825_, _12827_);
  or g_40064_(_23316_, _12824_, _12828_);
  and g_40065_(_23108_, _12765_, _12829_);
  or g_40066_(_23107_, _12766_, _12830_);
  or g_40067_(_12678_, _12765_, _12831_);
  not g_40068_(_12831_, _12832_);
  and g_40069_(_12830_, _12831_, _12833_);
  or g_40070_(_12829_, _12832_, _12834_);
  and g_40071_(_23307_, _12833_, _12835_);
  or g_40072_(_23306_, _12834_, _12836_);
  and g_40073_(_12828_, _12836_, _12838_);
  or g_40074_(_12827_, _12835_, _12839_);
  and g_40075_(_23316_, _12824_, _12840_);
  not g_40076_(_12840_, _12841_);
  and g_40077_(_23306_, _12834_, _12842_);
  or g_40078_(_23307_, _12833_, _12843_);
  or g_40079_(_12840_, _12842_, _12844_);
  and g_40080_(_12838_, _12843_, _12845_);
  and g_40081_(_12841_, _12845_, _12846_);
  or g_40082_(_12839_, _12844_, _12847_);
  and g_40083_(_12698_, _12766_, _12849_);
  or g_40084_(_12699_, _12765_, _12850_);
  and g_40085_(_23124_, _12765_, _12851_);
  not g_40086_(_12851_, _12852_);
  or g_40087_(_12849_, _12851_, _12853_);
  and g_40088_(_12850_, _12852_, _12854_);
  or g_40089_(_23354_, _12853_, _12855_);
  and g_40090_(_23131_, _12765_, _12856_);
  not g_40091_(_12856_, _12857_);
  and g_40092_(_12687_, _12766_, _12858_);
  or g_40093_(_12686_, _12765_, _12860_);
  and g_40094_(_12857_, _12860_, _12861_);
  or g_40095_(_12856_, _12858_, _12862_);
  and g_40096_(_23332_, _12861_, _12863_);
  or g_40097_(_23333_, _12862_, _12864_);
  or g_40098_(_23332_, _12861_, _12865_);
  xor g_40099_(_23354_, _12853_, _12866_);
  and g_40100_(_12864_, _12866_, _12867_);
  and g_40101_(_12865_, _12867_, _12868_);
  and g_40102_(_12846_, _12868_, _12869_);
  not g_40103_(_12869_, _12871_);
  and g_40104_(_12818_, _12869_, _12872_);
  or g_40105_(_12819_, _12871_, _12873_);
  and g_40106_(out[225], _12765_, _12874_);
  not g_40107_(_12874_, _12875_);
  or g_40108_(_12709_, _12765_, _12876_);
  not g_40109_(_12876_, _12877_);
  and g_40110_(_12875_, _12876_, _12878_);
  or g_40111_(_12874_, _12877_, _12879_);
  or g_40112_(_19277_, _12879_, _12880_);
  or g_40113_(_23153_, _12766_, _12882_);
  or g_40114_(_12715_, _12765_, _12883_);
  and g_40115_(_12882_, _12883_, _12884_);
  and g_40116_(_23377_, _12884_, _12885_);
  or g_40117_(_12722_, _12765_, _12886_);
  or g_40118_(_19231_, _12766_, _12887_);
  and g_40119_(_12886_, _12887_, _12888_);
  not g_40120_(_12888_, _12889_);
  or g_40121_(_19444_, _12889_, _12890_);
  or g_40122_(_23377_, _12884_, _12891_);
  xor g_40123_(_23377_, _12884_, _12893_);
  xor g_40124_(_23376_, _12884_, _12894_);
  xor g_40125_(_19443_, _12888_, _12895_);
  xor g_40126_(_19444_, _12888_, _12896_);
  and g_40127_(_12893_, _12895_, _12897_);
  or g_40128_(_12894_, _12896_, _12898_);
  or g_40129_(_12880_, _12898_, _12899_);
  or g_40130_(out[241], _12878_, _12900_);
  and g_40131_(_12736_, _12766_, _12901_);
  or g_40132_(_12735_, _12765_, _12902_);
  or g_40133_(out[224], _12766_, _12904_);
  not g_40134_(_12904_, _12905_);
  and g_40135_(_12902_, _12904_, _12906_);
  or g_40136_(_12901_, _12905_, _12907_);
  and g_40137_(out[240], _12907_, _12908_);
  or g_40138_(_19288_, _12906_, _12909_);
  and g_40139_(_12900_, _12909_, _12910_);
  and g_40140_(_12880_, _12910_, _12911_);
  xor g_40141_(_19277_, _12878_, _12912_);
  or g_40142_(_12898_, _12908_, _12913_);
  and g_40143_(_12897_, _12911_, _12915_);
  or g_40144_(_12912_, _12913_, _12916_);
  or g_40145_(_12885_, _12890_, _12917_);
  and g_40146_(_12891_, _12917_, _12918_);
  and g_40147_(_12916_, _12918_, _12919_);
  and g_40148_(_12899_, _12919_, _12920_);
  or g_40149_(_12873_, _12920_, _12921_);
  or g_40150_(_12838_, _12840_, _12922_);
  and g_40151_(_12855_, _12865_, _12923_);
  or g_40152_(_12863_, _12923_, _12924_);
  or g_40153_(_12847_, _12924_, _12926_);
  and g_40154_(_12922_, _12926_, _12927_);
  or g_40155_(_12819_, _12927_, _12928_);
  or g_40156_(_12778_, _12780_, _12929_);
  or g_40157_(_12807_, _12809_, _12930_);
  or g_40158_(_12788_, _12930_, _12931_);
  and g_40159_(_12929_, _12931_, _12932_);
  and g_40160_(_12928_, _12932_, _12933_);
  and g_40161_(_12921_, _12933_, _12934_);
  or g_40162_(out[240], _12907_, _12935_);
  and g_40163_(_12915_, _12935_, _12937_);
  and g_40164_(_12872_, _12937_, _12938_);
  or g_40165_(_12934_, _12938_, _12939_);
  not g_40166_(_12939_, _12940_);
  and g_40167_(_12244_, _12940_, _12941_);
  or g_40168_(_12245_, _12939_, _12942_);
  and g_40169_(_12773_, _12939_, _12943_);
  or g_40170_(_12772_, _12940_, _12944_);
  and g_40171_(_12942_, _12944_, _12945_);
  or g_40172_(_12941_, _12943_, _12946_);
  and g_40173_(_12224_, _12226_, _12948_);
  or g_40174_(_12223_, _12227_, _12949_);
  xor g_40175_(out[266], _23565_, _12950_);
  xor g_40176_(_19475_, _23565_, _12951_);
  and g_40177_(_12945_, _12950_, _12952_);
  or g_40178_(_12946_, _12951_, _12953_);
  and g_40179_(_12223_, _12227_, _12954_);
  or g_40180_(_12224_, _12226_, _12955_);
  and g_40181_(_12953_, _12955_, _12956_);
  or g_40182_(_12952_, _12954_, _12957_);
  and g_40183_(_12949_, _12957_, _12959_);
  or g_40184_(_12948_, _12956_, _12960_);
  and g_40185_(_23269_, _12940_, _12961_);
  or g_40186_(_23271_, _12939_, _12962_);
  and g_40187_(_12803_, _12939_, _12963_);
  or g_40188_(_12802_, _12940_, _12964_);
  and g_40189_(_12962_, _12964_, _12965_);
  or g_40190_(_12961_, _12963_, _12966_);
  and g_40191_(_23572_, _12966_, _12967_);
  or g_40192_(_23571_, _12965_, _12968_);
  and g_40193_(_23282_, _12940_, _12970_);
  or g_40194_(_23283_, _12939_, _12971_);
  and g_40195_(_12795_, _12939_, _12972_);
  or g_40196_(_12794_, _12940_, _12973_);
  and g_40197_(_12971_, _12973_, _12974_);
  or g_40198_(_12970_, _12972_, _12975_);
  and g_40199_(_23568_, _12975_, _12976_);
  or g_40200_(_23566_, _12974_, _12977_);
  and g_40201_(_12968_, _12977_, _12978_);
  or g_40202_(_12967_, _12976_, _12979_);
  and g_40203_(_12833_, _12939_, _12981_);
  not g_40204_(_12981_, _12982_);
  and g_40205_(_23306_, _12940_, _12983_);
  or g_40206_(_23307_, _12939_, _12984_);
  or g_40207_(_12981_, _12983_, _12985_);
  and g_40208_(_12982_, _12984_, _12986_);
  and g_40209_(_23594_, _12985_, _12987_);
  or g_40210_(_23593_, _12986_, _12988_);
  and g_40211_(_12824_, _12939_, _12989_);
  not g_40212_(_12989_, _12990_);
  and g_40213_(_23315_, _12940_, _12992_);
  or g_40214_(_23316_, _12939_, _12993_);
  or g_40215_(_12989_, _12992_, _12994_);
  and g_40216_(_12990_, _12993_, _12995_);
  and g_40217_(_23599_, _12994_, _12996_);
  or g_40218_(_23598_, _12995_, _12997_);
  and g_40219_(_23598_, _12995_, _12998_);
  or g_40220_(_23599_, _12994_, _12999_);
  and g_40221_(_23332_, _12940_, _13000_);
  or g_40222_(_23333_, _12939_, _13001_);
  and g_40223_(_12862_, _12939_, _13003_);
  or g_40224_(_12861_, _12940_, _13004_);
  and g_40225_(_13001_, _13004_, _13005_);
  or g_40226_(_13000_, _13003_, _13006_);
  and g_40227_(_23476_, _13005_, _13007_);
  or g_40228_(_23477_, _13006_, _13008_);
  xor g_40229_(_23594_, _12985_, _13009_);
  xor g_40230_(_23593_, _12985_, _13010_);
  and g_40231_(_12997_, _13009_, _13011_);
  or g_40232_(_12996_, _13010_, _13012_);
  and g_40233_(_12999_, _13011_, _13014_);
  or g_40234_(_12998_, _13012_, _13015_);
  and g_40235_(_13008_, _13014_, _13016_);
  or g_40236_(_13007_, _13015_, _13017_);
  and g_40237_(_23354_, _12940_, _13018_);
  or g_40238_(_23355_, _12939_, _13019_);
  and g_40239_(_12854_, _12939_, _13020_);
  or g_40240_(_12853_, _12940_, _13021_);
  and g_40241_(_13019_, _13021_, _13022_);
  or g_40242_(_13018_, _13020_, _13023_);
  and g_40243_(_23467_, _13023_, _13025_);
  or g_40244_(_23466_, _13022_, _13026_);
  and g_40245_(_23477_, _13006_, _13027_);
  or g_40246_(_23476_, _13005_, _13028_);
  and g_40247_(_13026_, _13028_, _13029_);
  or g_40248_(_13025_, _13027_, _13030_);
  and g_40249_(_23466_, _13022_, _13031_);
  or g_40250_(_23467_, _13023_, _13032_);
  and g_40251_(_13029_, _13032_, _13033_);
  or g_40252_(_13030_, _13031_, _13034_);
  and g_40253_(_13016_, _13033_, _13036_);
  or g_40254_(_13017_, _13034_, _13037_);
  and g_40255_(_12884_, _12939_, _13038_);
  not g_40256_(_13038_, _13039_);
  and g_40257_(_23376_, _12940_, _13040_);
  or g_40258_(_23377_, _12939_, _13041_);
  or g_40259_(_13038_, _13040_, _13042_);
  and g_40260_(_13039_, _13041_, _13043_);
  and g_40261_(_23492_, _13043_, _13044_);
  or g_40262_(_23492_, _13043_, _13045_);
  or g_40263_(_19444_, _12939_, _13047_);
  or g_40264_(_12888_, _12940_, _13048_);
  and g_40265_(_13047_, _13048_, _13049_);
  and g_40266_(_19674_, _13049_, _13050_);
  and g_40267_(_13045_, _13050_, _13051_);
  or g_40268_(_13044_, _13051_, _13052_);
  not g_40269_(_13052_, _13053_);
  and g_40270_(out[241], _12940_, _13054_);
  or g_40271_(_19277_, _12939_, _13055_);
  and g_40272_(_12879_, _12939_, _13056_);
  or g_40273_(_12878_, _12940_, _13058_);
  and g_40274_(_13055_, _13058_, _13059_);
  or g_40275_(_13054_, _13056_, _13060_);
  or g_40276_(_19409_, _13060_, _13061_);
  not g_40277_(_13061_, _13062_);
  and g_40278_(_12907_, _12939_, _13063_);
  or g_40279_(_12906_, _12940_, _13064_);
  or g_40280_(out[240], _12939_, _13065_);
  not g_40281_(_13065_, _13066_);
  and g_40282_(_13064_, _13065_, _13067_);
  or g_40283_(_13063_, _13066_, _13069_);
  and g_40284_(out[256], _13069_, _13070_);
  or g_40285_(_19420_, _13067_, _13071_);
  or g_40286_(out[257], _13059_, _13072_);
  and g_40287_(_13071_, _13072_, _13073_);
  xor g_40288_(_19409_, _13059_, _13074_);
  or g_40289_(_13070_, _13074_, _13075_);
  and g_40290_(_13061_, _13075_, _13076_);
  or g_40291_(_13062_, _13073_, _13077_);
  xor g_40292_(_19674_, _13049_, _13078_);
  xor g_40293_(_19675_, _13049_, _13080_);
  xor g_40294_(_23493_, _13042_, _13081_);
  xor g_40295_(_23492_, _13042_, _13082_);
  and g_40296_(_13078_, _13081_, _13083_);
  or g_40297_(_13080_, _13082_, _13084_);
  and g_40298_(_13077_, _13083_, _13085_);
  or g_40299_(_13076_, _13084_, _13086_);
  and g_40300_(_13053_, _13086_, _13087_);
  or g_40301_(_13052_, _13085_, _13088_);
  and g_40302_(_13036_, _13088_, _13089_);
  or g_40303_(_13037_, _13087_, _13091_);
  and g_40304_(_13016_, _13030_, _13092_);
  or g_40305_(_13017_, _13029_, _13093_);
  and g_40306_(_12987_, _12997_, _13094_);
  or g_40307_(_12988_, _12996_, _13095_);
  and g_40308_(_12999_, _13095_, _13096_);
  or g_40309_(_12998_, _13094_, _13097_);
  and g_40310_(_13093_, _13096_, _13098_);
  or g_40311_(_13092_, _13097_, _13099_);
  and g_40312_(_13091_, _13098_, _13100_);
  or g_40313_(_13089_, _13099_, _13102_);
  and g_40314_(_23571_, _12965_, _13103_);
  or g_40315_(_23572_, _12966_, _13104_);
  and g_40316_(_13102_, _13104_, _13105_);
  or g_40317_(_13100_, _13103_, _13106_);
  and g_40318_(_12978_, _13106_, _13107_);
  or g_40319_(_12979_, _13105_, _13108_);
  and g_40320_(_23566_, _12974_, _13109_);
  or g_40321_(_23568_, _12975_, _13110_);
  and g_40322_(_12946_, _12951_, _13111_);
  or g_40323_(_12945_, _12950_, _13113_);
  and g_40324_(_13110_, _13113_, _13114_);
  or g_40325_(_13109_, _13111_, _13115_);
  and g_40326_(_12949_, _13114_, _13116_);
  or g_40327_(_12948_, _13115_, _13117_);
  and g_40328_(_13108_, _13116_, _13118_);
  or g_40329_(_13107_, _13117_, _13119_);
  and g_40330_(_12960_, _13119_, _13120_);
  or g_40331_(_12959_, _13118_, _13121_);
  and g_40332_(_19420_, _13067_, _13122_);
  or g_40333_(out[256], _13069_, _13124_);
  and g_40334_(_13116_, _13124_, _13125_);
  or g_40335_(_13117_, _13122_, _13126_);
  or g_40336_(_12979_, _13084_, _13127_);
  or g_40337_(_13075_, _13103_, _13128_);
  or g_40338_(_13127_, _13128_, _13129_);
  not g_40339_(_13129_, _13130_);
  and g_40340_(_13036_, _13130_, _13131_);
  or g_40341_(_13037_, _13129_, _13132_);
  and g_40342_(_13125_, _13131_, _13133_);
  or g_40343_(_13126_, _13132_, _13135_);
  and g_40344_(_12956_, _13133_, _13136_);
  or g_40345_(_12957_, _13135_, _13137_);
  and g_40346_(_13121_, _13137_, _13138_);
  or g_40347_(_13120_, _13136_, _13139_);
  and g_40348_(_12946_, _13139_, _13140_);
  not g_40349_(_13140_, _13141_);
  or g_40350_(_12951_, _13139_, _13142_);
  not g_40351_(_13142_, _13143_);
  and g_40352_(_13141_, _13142_, _13144_);
  or g_40353_(_13140_, _13143_, _13146_);
  and g_40354_(_12242_, _13146_, _13147_);
  or g_40355_(_12241_, _13144_, _13148_);
  and g_40356_(_12241_, _13144_, _13149_);
  or g_40357_(_12242_, _13146_, _13150_);
  and g_40358_(_12228_, _12233_, _13151_);
  or g_40359_(_12229_, _12231_, _13152_);
  and g_40360_(_12229_, _12231_, _13153_);
  or g_40361_(_12228_, _12233_, _13154_);
  and g_40362_(_13148_, _13152_, _13155_);
  or g_40363_(_13147_, _13151_, _13157_);
  and g_40364_(_13150_, _13154_, _13158_);
  or g_40365_(_13149_, _13153_, _13159_);
  and g_40366_(_13155_, _13158_, _13160_);
  or g_40367_(_13157_, _13159_, _13161_);
  and g_40368_(_12966_, _13139_, _13162_);
  not g_40369_(_13162_, _13163_);
  or g_40370_(_23572_, _13139_, _13164_);
  not g_40371_(_13164_, _13165_);
  and g_40372_(_13163_, _13164_, _13166_);
  or g_40373_(_13162_, _13165_, _13168_);
  and g_40374_(_23703_, _13168_, _13169_);
  or g_40375_(_23702_, _13166_, _13170_);
  and g_40376_(_23566_, _13138_, _13171_);
  and g_40377_(_12975_, _13139_, _13172_);
  or g_40378_(_13171_, _13172_, _13173_);
  not g_40379_(_13173_, _13174_);
  and g_40380_(_23692_, _13173_, _13175_);
  or g_40381_(_23691_, _13174_, _13176_);
  and g_40382_(_13170_, _13176_, _13177_);
  or g_40383_(_13169_, _13175_, _13179_);
  and g_40384_(_23691_, _13174_, _13180_);
  or g_40385_(_23692_, _13173_, _13181_);
  and g_40386_(_23702_, _13166_, _13182_);
  or g_40387_(_23703_, _13168_, _13183_);
  and g_40388_(_13181_, _13183_, _13184_);
  or g_40389_(_13180_, _13182_, _13185_);
  and g_40390_(_13177_, _13184_, _13186_);
  or g_40391_(_13179_, _13185_, _13187_);
  and g_40392_(_13160_, _13186_, _13188_);
  or g_40393_(_13161_, _13187_, _13190_);
  or g_40394_(_12985_, _13138_, _13191_);
  or g_40395_(_23593_, _13139_, _13192_);
  and g_40396_(_13191_, _13192_, _13193_);
  not g_40397_(_13193_, _13194_);
  and g_40398_(_23729_, _13193_, _13195_);
  or g_40399_(_23728_, _13194_, _13196_);
  or g_40400_(_23598_, _13139_, _13197_);
  not g_40401_(_13197_, _13198_);
  and g_40402_(_12995_, _13139_, _13199_);
  not g_40403_(_13199_, _13201_);
  and g_40404_(_13197_, _13201_, _13202_);
  or g_40405_(_13198_, _13199_, _13203_);
  and g_40406_(_23731_, _13203_, _13204_);
  or g_40407_(_23733_, _13202_, _13205_);
  and g_40408_(_23733_, _13202_, _13206_);
  or g_40409_(_23731_, _13203_, _13207_);
  xor g_40410_(_23729_, _13193_, _13208_);
  xor g_40411_(_23728_, _13193_, _13209_);
  and g_40412_(_13205_, _13207_, _13210_);
  or g_40413_(_13204_, _13206_, _13212_);
  and g_40414_(_13208_, _13210_, _13213_);
  or g_40415_(_13209_, _13212_, _13214_);
  or g_40416_(_23467_, _13139_, _13215_);
  not g_40417_(_13215_, _13216_);
  and g_40418_(_13023_, _13139_, _13217_);
  not g_40419_(_13217_, _13218_);
  and g_40420_(_13215_, _13218_, _13219_);
  or g_40421_(_13216_, _13217_, _13220_);
  and g_40422_(_23749_, _13220_, _13221_);
  or g_40423_(_23748_, _13219_, _13223_);
  xor g_40424_(_23748_, _13219_, _13224_);
  xor g_40425_(_23749_, _13219_, _13225_);
  and g_40426_(_13006_, _13139_, _13226_);
  not g_40427_(_13226_, _13227_);
  or g_40428_(_23477_, _13139_, _13228_);
  not g_40429_(_13228_, _13229_);
  and g_40430_(_13227_, _13228_, _13230_);
  or g_40431_(_13226_, _13229_, _13231_);
  and g_40432_(_23759_, _13230_, _13232_);
  or g_40433_(_23760_, _13231_, _13234_);
  and g_40434_(_23760_, _13231_, _13235_);
  or g_40435_(_23759_, _13230_, _13236_);
  and g_40436_(_13234_, _13236_, _13237_);
  or g_40437_(_13232_, _13235_, _13238_);
  and g_40438_(_13224_, _13237_, _13239_);
  or g_40439_(_13225_, _13238_, _13240_);
  and g_40440_(_13213_, _13239_, _13241_);
  or g_40441_(_13214_, _13240_, _13242_);
  and g_40442_(out[257], _13138_, _13243_);
  and g_40443_(_13060_, _13139_, _13245_);
  or g_40444_(_13243_, _13245_, _13246_);
  not g_40445_(_13246_, _13247_);
  and g_40446_(out[273], _13247_, _13248_);
  or g_40447_(_19541_, _13246_, _13249_);
  and g_40448_(_23493_, _13138_, _13250_);
  or g_40449_(_23492_, _13139_, _13251_);
  and g_40450_(_13043_, _13139_, _13252_);
  or g_40451_(_13042_, _13138_, _13253_);
  and g_40452_(_13251_, _13253_, _13254_);
  or g_40453_(_13250_, _13252_, _13256_);
  and g_40454_(_23785_, _13256_, _13257_);
  or g_40455_(_23786_, _13254_, _13258_);
  and g_40456_(_23786_, _13254_, _13259_);
  or g_40457_(_23785_, _13256_, _13260_);
  and g_40458_(_13258_, _13260_, _13261_);
  or g_40459_(_13257_, _13259_, _13262_);
  or g_40460_(_19675_, _13139_, _13263_);
  or g_40461_(_13049_, _13138_, _13264_);
  and g_40462_(_13263_, _13264_, _13265_);
  not g_40463_(_13265_, _13267_);
  and g_40464_(_19886_, _13265_, _13268_);
  or g_40465_(_19887_, _13267_, _13269_);
  xor g_40466_(_19886_, _13265_, _13270_);
  xor g_40467_(_19887_, _13265_, _13271_);
  and g_40468_(_13261_, _13270_, _13272_);
  or g_40469_(_13262_, _13271_, _13273_);
  and g_40470_(_13248_, _13272_, _13274_);
  or g_40471_(_13249_, _13273_, _13275_);
  and g_40472_(_13260_, _13268_, _13276_);
  or g_40473_(_13259_, _13269_, _13278_);
  and g_40474_(_13258_, _13278_, _13279_);
  or g_40475_(_13257_, _13276_, _13280_);
  and g_40476_(_13275_, _13279_, _13281_);
  or g_40477_(_13274_, _13280_, _13282_);
  and g_40478_(_13241_, _13282_, _13283_);
  or g_40479_(_13242_, _13281_, _13284_);
  and g_40480_(_13223_, _13236_, _13285_);
  or g_40481_(_13221_, _13235_, _13286_);
  and g_40482_(_13234_, _13286_, _13287_);
  or g_40483_(_13232_, _13285_, _13289_);
  and g_40484_(_13213_, _13287_, _13290_);
  or g_40485_(_13214_, _13289_, _13291_);
  and g_40486_(_13195_, _13207_, _13292_);
  or g_40487_(_13196_, _13206_, _13293_);
  and g_40488_(_13205_, _13293_, _13294_);
  or g_40489_(_13204_, _13292_, _13295_);
  and g_40490_(_13291_, _13294_, _13296_);
  or g_40491_(_13290_, _13295_, _13297_);
  and g_40492_(_13069_, _13139_, _13298_);
  not g_40493_(_13298_, _13300_);
  or g_40494_(out[256], _13139_, _13301_);
  not g_40495_(_13301_, _13302_);
  and g_40496_(_13300_, _13301_, _13303_);
  or g_40497_(_13298_, _13302_, _13304_);
  and g_40498_(out[272], _13304_, _13305_);
  xor g_40499_(out[273], _13246_, _13306_);
  or g_40500_(_13305_, _13306_, _13307_);
  or g_40501_(_13273_, _13307_, _13308_);
  not g_40502_(_13308_, _13309_);
  and g_40503_(_13241_, _13309_, _13311_);
  or g_40504_(_13242_, _13308_, _13312_);
  and g_40505_(_13284_, _13296_, _13313_);
  or g_40506_(_13283_, _13297_, _13314_);
  and g_40507_(_13312_, _13313_, _13315_);
  or g_40508_(_13311_, _13314_, _13316_);
  and g_40509_(_13188_, _13316_, _13317_);
  or g_40510_(_13190_, _13315_, _13318_);
  and g_40511_(_13179_, _13181_, _13319_);
  or g_40512_(_13177_, _13180_, _13320_);
  and g_40513_(_13160_, _13319_, _13322_);
  or g_40514_(_13161_, _13320_, _13323_);
  and g_40515_(_13149_, _13154_, _13324_);
  or g_40516_(_13150_, _13153_, _13325_);
  and g_40517_(_13152_, _13325_, _13326_);
  or g_40518_(_13151_, _13324_, _13327_);
  and g_40519_(_13323_, _13326_, _13328_);
  or g_40520_(_13322_, _13327_, _13329_);
  and g_40521_(_13318_, _13328_, _13330_);
  or g_40522_(_13317_, _13329_, _13331_);
  and g_40523_(_19552_, _13303_, _13333_);
  or g_40524_(out[272], _13304_, _13334_);
  and g_40525_(_13188_, _13334_, _13335_);
  or g_40526_(_13190_, _13333_, _13336_);
  and g_40527_(_13311_, _13335_, _13337_);
  or g_40528_(_13312_, _13336_, _13338_);
  and g_40529_(_13331_, _13338_, _13339_);
  or g_40530_(_13330_, _13337_, _13340_);
  and g_40531_(_23691_, _13339_, _13341_);
  and g_40532_(_13173_, _13340_, _13342_);
  or g_40533_(_13341_, _13342_, _13344_);
  not g_40534_(_13344_, _13345_);
  and g_40535_(_23895_, _13345_, _13346_);
  or g_40536_(_23896_, _13344_, _13347_);
  xor g_40537_(out[298], _23894_, _13348_);
  xor g_40538_(_19728_, _23894_, _13349_);
  or g_40539_(_12242_, _13340_, _13350_);
  not g_40540_(_13350_, _13351_);
  and g_40541_(_13146_, _13340_, _13352_);
  not g_40542_(_13352_, _13353_);
  and g_40543_(_13350_, _13353_, _13355_);
  or g_40544_(_13351_, _13352_, _13356_);
  and g_40545_(_13349_, _13356_, _13357_);
  or g_40546_(_13348_, _13355_, _13358_);
  or g_40547_(_23703_, _13340_, _13359_);
  not g_40548_(_13359_, _13360_);
  and g_40549_(_13168_, _13340_, _13361_);
  not g_40550_(_13361_, _13362_);
  and g_40551_(_13359_, _13362_, _13363_);
  or g_40552_(_13360_, _13361_, _13364_);
  and g_40553_(_23906_, _13363_, _13366_);
  or g_40554_(_23907_, _13364_, _13367_);
  and g_40555_(_12234_, _12238_, _13368_);
  or g_40556_(_12235_, _12237_, _13369_);
  and g_40557_(_13348_, _13355_, _13370_);
  or g_40558_(_13349_, _13356_, _13371_);
  and g_40559_(_13369_, _13371_, _13372_);
  or g_40560_(_13368_, _13370_, _13373_);
  and g_40561_(_23907_, _13364_, _13374_);
  or g_40562_(_23906_, _13363_, _13375_);
  and g_40563_(_23896_, _13344_, _13377_);
  or g_40564_(_23895_, _13345_, _13378_);
  and g_40565_(_13375_, _13378_, _13379_);
  or g_40566_(_13374_, _13377_, _13380_);
  and g_40567_(_12240_, _13358_, _13381_);
  or g_40568_(_12239_, _13357_, _13382_);
  and g_40569_(_13372_, _13381_, _13383_);
  or g_40570_(_13373_, _13382_, _13384_);
  and g_40571_(_13347_, _13367_, _13385_);
  or g_40572_(_13346_, _13366_, _13386_);
  and g_40573_(_13379_, _13385_, _13388_);
  or g_40574_(_13380_, _13386_, _13389_);
  and g_40575_(_13383_, _13388_, _13390_);
  or g_40576_(_13384_, _13389_, _13391_);
  and g_40577_(_13203_, _13340_, _13392_);
  or g_40578_(_13202_, _13339_, _13393_);
  and g_40579_(_23733_, _13339_, _13394_);
  or g_40580_(_23731_, _13340_, _13395_);
  and g_40581_(_13393_, _13395_, _13396_);
  or g_40582_(_13392_, _13394_, _13397_);
  and g_40583_(_23936_, _13397_, _13399_);
  or g_40584_(_23937_, _13396_, _13400_);
  and g_40585_(_23937_, _13396_, _13401_);
  or g_40586_(_23936_, _13397_, _13402_);
  and g_40587_(_13400_, _13402_, _13403_);
  or g_40588_(_13399_, _13401_, _13404_);
  or g_40589_(_13193_, _13339_, _13405_);
  or g_40590_(_23728_, _13340_, _13406_);
  and g_40591_(_13405_, _13406_, _13407_);
  not g_40592_(_13407_, _13408_);
  and g_40593_(_22421_, _13407_, _13410_);
  or g_40594_(_22420_, _13408_, _13411_);
  xor g_40595_(_22421_, _13407_, _13412_);
  xor g_40596_(_22420_, _13407_, _13413_);
  and g_40597_(_13403_, _13412_, _13414_);
  or g_40598_(_13404_, _13413_, _13415_);
  and g_40599_(_23748_, _13339_, _13416_);
  and g_40600_(_13220_, _13340_, _13417_);
  or g_40601_(_13416_, _13417_, _13418_);
  not g_40602_(_13418_, _13419_);
  and g_40603_(_23954_, _13418_, _13421_);
  or g_40604_(_23953_, _13419_, _13422_);
  or g_40605_(_23760_, _13340_, _13423_);
  not g_40606_(_13423_, _13424_);
  and g_40607_(_13231_, _13340_, _13425_);
  not g_40608_(_13425_, _13426_);
  and g_40609_(_13423_, _13426_, _13427_);
  or g_40610_(_13424_, _13425_, _13428_);
  and g_40611_(_23960_, _13428_, _13429_);
  or g_40612_(_23959_, _13427_, _13430_);
  and g_40613_(_13422_, _13430_, _13432_);
  or g_40614_(_13421_, _13429_, _13433_);
  and g_40615_(_23959_, _13427_, _13434_);
  or g_40616_(_23960_, _13428_, _13435_);
  and g_40617_(_23953_, _13419_, _13436_);
  or g_40618_(_23954_, _13418_, _13437_);
  and g_40619_(_13435_, _13437_, _13438_);
  or g_40620_(_13434_, _13436_, _13439_);
  and g_40621_(_13432_, _13438_, _13440_);
  or g_40622_(_13433_, _13439_, _13441_);
  and g_40623_(_13414_, _13440_, _13443_);
  or g_40624_(_13415_, _13441_, _13444_);
  and g_40625_(_13390_, _13443_, _13445_);
  or g_40626_(_13391_, _13444_, _13446_);
  or g_40627_(_23785_, _13340_, _13447_);
  or g_40628_(_13254_, _13339_, _13448_);
  and g_40629_(_13447_, _13448_, _13449_);
  or g_40630_(_23979_, _13449_, _13450_);
  not g_40631_(_13450_, _13451_);
  and g_40632_(_13267_, _13340_, _13452_);
  and g_40633_(_19886_, _13339_, _13454_);
  or g_40634_(_13452_, _13454_, _13455_);
  and g_40635_(_23979_, _13449_, _13456_);
  not g_40636_(_13456_, _13457_);
  or g_40637_(_20108_, _13455_, _13458_);
  and g_40638_(_13450_, _13457_, _13459_);
  or g_40639_(_13451_, _13456_, _13460_);
  xor g_40640_(_20108_, _13455_, _13461_);
  xor g_40641_(_20107_, _13455_, _13462_);
  and g_40642_(_13459_, _13461_, _13463_);
  or g_40643_(_13460_, _13462_, _13465_);
  and g_40644_(out[273], _13339_, _13466_);
  and g_40645_(_13246_, _13340_, _13467_);
  or g_40646_(_13466_, _13467_, _13468_);
  not g_40647_(_13468_, _13469_);
  and g_40648_(out[289], _13469_, _13470_);
  or g_40649_(_19673_, _13468_, _13471_);
  or g_40650_(_13303_, _13339_, _13472_);
  or g_40651_(out[272], _13340_, _13473_);
  and g_40652_(_13472_, _13473_, _13474_);
  not g_40653_(_13474_, _13476_);
  and g_40654_(out[288], _13476_, _13477_);
  or g_40655_(_18573_, _13474_, _13478_);
  xor g_40656_(_19673_, _13468_, _13479_);
  xor g_40657_(out[289], _13468_, _13480_);
  and g_40658_(_13478_, _13479_, _13481_);
  or g_40659_(_13477_, _13480_, _13482_);
  and g_40660_(_13471_, _13482_, _13483_);
  or g_40661_(_13470_, _13481_, _13484_);
  and g_40662_(_13463_, _13484_, _13485_);
  or g_40663_(_13465_, _13483_, _13487_);
  or g_40664_(_13456_, _13458_, _13488_);
  and g_40665_(_13450_, _13488_, _13489_);
  not g_40666_(_13489_, _13490_);
  and g_40667_(_13487_, _13489_, _13491_);
  or g_40668_(_13485_, _13490_, _13492_);
  and g_40669_(_13445_, _13492_, _13493_);
  or g_40670_(_13446_, _13491_, _13494_);
  and g_40671_(_13414_, _13433_, _13495_);
  or g_40672_(_13415_, _13432_, _13496_);
  and g_40673_(_13435_, _13495_, _13498_);
  or g_40674_(_13434_, _13496_, _13499_);
  and g_40675_(_13402_, _13410_, _13500_);
  or g_40676_(_13401_, _13411_, _13501_);
  and g_40677_(_13400_, _13501_, _13502_);
  or g_40678_(_13399_, _13500_, _13503_);
  and g_40679_(_13499_, _13502_, _13504_);
  or g_40680_(_13498_, _13503_, _13505_);
  and g_40681_(_13390_, _13505_, _13506_);
  or g_40682_(_13391_, _13504_, _13507_);
  and g_40683_(_13347_, _13358_, _13509_);
  or g_40684_(_13346_, _13357_, _13510_);
  and g_40685_(_13380_, _13509_, _13511_);
  or g_40686_(_13379_, _13510_, _13512_);
  and g_40687_(_13372_, _13512_, _13513_);
  or g_40688_(_13373_, _13511_, _13514_);
  and g_40689_(_12240_, _13514_, _13515_);
  or g_40690_(_12239_, _13513_, _13516_);
  and g_40691_(_13507_, _13516_, _13517_);
  or g_40692_(_13506_, _13515_, _13518_);
  and g_40693_(_13494_, _13517_, _13520_);
  or g_40694_(_13493_, _13518_, _13521_);
  and g_40695_(_18573_, _13474_, _13522_);
  or g_40696_(out[288], _13476_, _13523_);
  and g_40697_(_13463_, _13523_, _13524_);
  or g_40698_(_13465_, _13522_, _13525_);
  and g_40699_(_13481_, _13524_, _13526_);
  or g_40700_(_13482_, _13525_, _13527_);
  and g_40701_(_13445_, _13526_, _13528_);
  or g_40702_(_13446_, _13527_, _13529_);
  and g_40703_(_13521_, _13529_, _13531_);
  or g_40704_(_13520_, _13528_, _13532_);
  or g_40705_(_23978_, _13532_, _13533_);
  or g_40706_(_13449_, _13531_, _13534_);
  and g_40707_(_13533_, _13534_, _13535_);
  or g_40708_(_24164_, _13535_, _13536_);
  and g_40709_(_24164_, _13535_, _13537_);
  xor g_40710_(_24163_, _13535_, _13538_);
  and g_40711_(_20107_, _13531_, _13539_);
  and g_40712_(_13455_, _13532_, _13540_);
  or g_40713_(_13539_, _13540_, _13542_);
  or g_40714_(_20294_, _13542_, _13543_);
  xor g_40715_(_20293_, _13542_, _13544_);
  or g_40716_(_13538_, _13544_, _13545_);
  and g_40717_(out[289], _13531_, _13546_);
  and g_40718_(_13468_, _13532_, _13547_);
  or g_40719_(_13546_, _13547_, _13548_);
  or g_40720_(_19794_, _13548_, _13549_);
  or g_40721_(_13474_, _13531_, _13550_);
  or g_40722_(out[288], _13532_, _13551_);
  and g_40723_(_13550_, _13551_, _13553_);
  not g_40724_(_13553_, _13554_);
  and g_40725_(out[304], _13554_, _13555_);
  xor g_40726_(out[305], _13548_, _13556_);
  or g_40727_(_13555_, _13556_, _13557_);
  and g_40728_(_13549_, _13557_, _13558_);
  or g_40729_(_13545_, _13558_, _13559_);
  and g_40730_(_13536_, _13543_, _13560_);
  or g_40731_(_13537_, _13560_, _13561_);
  and g_40732_(_13559_, _13561_, _13562_);
  not g_40733_(_13562_, _13564_);
  or g_40734_(out[314], _24121_, _13565_);
  xor g_40735_(out[314], _24121_, _13566_);
  xor g_40736_(_19849_, _24121_, _13567_);
  and g_40737_(_13348_, _13531_, _13568_);
  or g_40738_(_13349_, _13532_, _13569_);
  and g_40739_(_13356_, _13532_, _13570_);
  or g_40740_(_13355_, _13531_, _13571_);
  and g_40741_(_13569_, _13571_, _13572_);
  or g_40742_(_13568_, _13570_, _13573_);
  and g_40743_(_13567_, _13573_, _13575_);
  or g_40744_(_13566_, _13572_, _13576_);
  and g_40745_(_12234_, _12237_, _13577_);
  not g_40746_(_13577_, _13578_);
  xor g_40747_(out[315], _13565_, _13579_);
  not g_40748_(_13579_, _13580_);
  and g_40749_(_13578_, _13579_, _13581_);
  or g_40750_(_13577_, _13580_, _13582_);
  and g_40751_(_13576_, _13582_, _13583_);
  or g_40752_(_13575_, _13581_, _13584_);
  and g_40753_(_23907_, _13531_, _13586_);
  or g_40754_(_23906_, _13532_, _13587_);
  and g_40755_(_13363_, _13532_, _13588_);
  or g_40756_(_13364_, _13531_, _13589_);
  and g_40757_(_13587_, _13589_, _13590_);
  or g_40758_(_13586_, _13588_, _13591_);
  and g_40759_(_24116_, _13591_, _13592_);
  or g_40760_(_24118_, _13590_, _13593_);
  and g_40761_(_23895_, _13531_, _13594_);
  and g_40762_(_13344_, _13532_, _13595_);
  or g_40763_(_13594_, _13595_, _13597_);
  not g_40764_(_13597_, _13598_);
  and g_40765_(_24122_, _13598_, _13599_);
  or g_40766_(_24123_, _13597_, _13600_);
  and g_40767_(_13593_, _13600_, _13601_);
  or g_40768_(_13592_, _13599_, _13602_);
  and g_40769_(_13566_, _13572_, _13603_);
  or g_40770_(_13567_, _13573_, _13604_);
  and g_40771_(_13577_, _13580_, _13605_);
  or g_40772_(_13578_, _13579_, _13606_);
  and g_40773_(_13604_, _13606_, _13608_);
  or g_40774_(_13603_, _13605_, _13609_);
  and g_40775_(_24123_, _13597_, _13610_);
  or g_40776_(_24122_, _13598_, _13611_);
  and g_40777_(_24118_, _13590_, _13612_);
  or g_40778_(_24116_, _13591_, _13613_);
  and g_40779_(_13611_, _13613_, _13614_);
  or g_40780_(_13610_, _13612_, _13615_);
  and g_40781_(_13583_, _13608_, _13616_);
  or g_40782_(_13584_, _13609_, _13617_);
  and g_40783_(_13601_, _13614_, _13619_);
  or g_40784_(_13602_, _13615_, _13620_);
  and g_40785_(_13616_, _13619_, _13621_);
  or g_40786_(_13617_, _13620_, _13622_);
  or g_40787_(_22420_, _13532_, _13623_);
  or g_40788_(_13407_, _13531_, _13624_);
  and g_40789_(_13623_, _13624_, _13625_);
  and g_40790_(_22413_, _13625_, _13626_);
  xor g_40791_(_22413_, _13625_, _13627_);
  xor g_40792_(_22411_, _13625_, _13628_);
  and g_40793_(_23937_, _13531_, _13630_);
  or g_40794_(_23936_, _13532_, _13631_);
  and g_40795_(_13397_, _13532_, _13632_);
  or g_40796_(_13396_, _13531_, _13633_);
  and g_40797_(_13631_, _13633_, _13634_);
  or g_40798_(_13630_, _13632_, _13635_);
  and g_40799_(_24056_, _13635_, _13636_);
  or g_40800_(_24056_, _13635_, _13637_);
  xor g_40801_(_24057_, _13634_, _13638_);
  xor g_40802_(_24056_, _13634_, _13639_);
  and g_40803_(_13627_, _13638_, _13641_);
  or g_40804_(_13628_, _13639_, _13642_);
  and g_40805_(_23959_, _13531_, _13643_);
  or g_40806_(_23960_, _13532_, _13644_);
  and g_40807_(_13428_, _13532_, _13645_);
  or g_40808_(_13427_, _13531_, _13646_);
  and g_40809_(_13644_, _13646_, _13647_);
  or g_40810_(_13643_, _13645_, _13648_);
  and g_40811_(_24068_, _13648_, _13649_);
  or g_40812_(_24067_, _13647_, _13650_);
  or g_40813_(_23953_, _13532_, _13652_);
  or g_40814_(_13418_, _13531_, _13653_);
  and g_40815_(_13652_, _13653_, _13654_);
  not g_40816_(_13654_, _13655_);
  and g_40817_(_24142_, _13654_, _13656_);
  or g_40818_(_24141_, _13655_, _13657_);
  and g_40819_(_13650_, _13657_, _13658_);
  or g_40820_(_13649_, _13656_, _13659_);
  and g_40821_(_24067_, _13647_, _13660_);
  or g_40822_(_24068_, _13648_, _13661_);
  and g_40823_(_24141_, _13655_, _13663_);
  or g_40824_(_13660_, _13663_, _13664_);
  or g_40825_(_13659_, _13664_, _13665_);
  or g_40826_(_13642_, _13665_, _13666_);
  not g_40827_(_13666_, _13667_);
  and g_40828_(_13621_, _13667_, _13668_);
  or g_40829_(_13622_, _13666_, _13669_);
  and g_40830_(_13564_, _13668_, _13670_);
  or g_40831_(_13562_, _13669_, _13671_);
  and g_40832_(_13641_, _13661_, _13672_);
  or g_40833_(_13642_, _13660_, _13674_);
  and g_40834_(_13659_, _13672_, _13675_);
  or g_40835_(_13658_, _13674_, _13676_);
  and g_40836_(_13626_, _13637_, _13677_);
  or g_40837_(_13636_, _13677_, _13678_);
  not g_40838_(_13678_, _13679_);
  and g_40839_(_13676_, _13679_, _13680_);
  or g_40840_(_13675_, _13678_, _13681_);
  and g_40841_(_13621_, _13681_, _13682_);
  or g_40842_(_13622_, _13680_, _13683_);
  and g_40843_(_13576_, _13600_, _13685_);
  or g_40844_(_13575_, _13599_, _13686_);
  and g_40845_(_13615_, _13685_, _13687_);
  or g_40846_(_13614_, _13686_, _13688_);
  and g_40847_(_13608_, _13688_, _13689_);
  or g_40848_(_13609_, _13687_, _13690_);
  and g_40849_(_13582_, _13690_, _13691_);
  or g_40850_(_13581_, _13689_, _13692_);
  and g_40851_(_13683_, _13692_, _13693_);
  or g_40852_(_13682_, _13691_, _13694_);
  and g_40853_(_13671_, _13693_, _13696_);
  or g_40854_(_13670_, _13694_, _13697_);
  and g_40855_(_18562_, _13553_, _13698_);
  or g_40856_(out[304], _13554_, _13699_);
  or g_40857_(_13545_, _13557_, _13700_);
  not g_40858_(_13700_, _13701_);
  and g_40859_(_13668_, _13701_, _13702_);
  or g_40860_(_13669_, _13700_, _13703_);
  and g_40861_(_13699_, _13702_, _13704_);
  or g_40862_(_13698_, _13703_, _13705_);
  and g_40863_(_13697_, _13705_, _13707_);
  or g_40864_(_13696_, _13704_, _13708_);
  and g_40865_(_24057_, _13707_, _13709_);
  or g_40866_(_24056_, _13708_, _13710_);
  and g_40867_(_13635_, _13708_, _13711_);
  or g_40868_(_13634_, _13707_, _13712_);
  and g_40869_(_13710_, _13712_, _13713_);
  or g_40870_(_13709_, _13711_, _13714_);
  and g_40871_(_12162_, _13713_, _13715_);
  and g_40872_(_12161_, _13714_, _13716_);
  or g_40873_(_12040_, _12154_, _13718_);
  not g_40874_(_13718_, _13719_);
  and g_40875_(_22282_, _12154_, _13720_);
  or g_40876_(_22283_, _12156_, _13721_);
  and g_40877_(_13718_, _13721_, _13722_);
  or g_40878_(_13719_, _13720_, _13723_);
  and g_40879_(_24067_, _13707_, _13724_);
  or g_40880_(_24068_, _13708_, _13725_);
  and g_40881_(_13648_, _13708_, _13726_);
  or g_40882_(_13647_, _13707_, _13727_);
  and g_40883_(_13725_, _13727_, _13729_);
  or g_40884_(_13724_, _13726_, _13730_);
  and g_40885_(_13722_, _13730_, _13731_);
  and g_40886_(_12095_, _12156_, _13732_);
  and g_40887_(out[145], _12154_, _13733_);
  or g_40888_(_13732_, _13733_, _13734_);
  and g_40889_(out[305], _13707_, _13735_);
  and g_40890_(_13548_, _13708_, _13736_);
  or g_40891_(_13735_, _13736_, _13737_);
  or g_40892_(_12103_, _12154_, _13738_);
  or g_40893_(out[144], _12156_, _13740_);
  and g_40894_(_13738_, _13740_, _13741_);
  or g_40895_(_13553_, _13707_, _13742_);
  or g_40896_(out[304], _13708_, _13743_);
  and g_40897_(_13742_, _13743_, _13744_);
  xor g_40898_(_13741_, _13744_, _13745_);
  and g_40899_(_11973_, _11976_, _13746_);
  and g_40900_(_13577_, _13579_, _13747_);
  xor g_40901_(_13746_, _13747_, _13748_);
  and g_40902_(_18337_, _12154_, _13749_);
  and g_40903_(_12081_, _12156_, _13751_);
  or g_40904_(_13749_, _13751_, _13752_);
  and g_40905_(_20293_, _13707_, _13753_);
  and g_40906_(_13542_, _13708_, _13754_);
  or g_40907_(_13753_, _13754_, _13755_);
  xor g_40908_(_13752_, _13755_, _13756_);
  and g_40909_(_22328_, _12154_, _13757_);
  or g_40910_(_22327_, _12156_, _13758_);
  or g_40911_(_12014_, _12154_, _13759_);
  not g_40912_(_13759_, _13760_);
  and g_40913_(_13758_, _13759_, _13762_);
  or g_40914_(_13757_, _13760_, _13763_);
  and g_40915_(_24118_, _13707_, _13764_);
  or g_40916_(_24116_, _13708_, _13765_);
  and g_40917_(_13591_, _13708_, _13766_);
  or g_40918_(_13590_, _13707_, _13767_);
  and g_40919_(_13765_, _13767_, _13768_);
  or g_40920_(_13764_, _13766_, _13769_);
  and g_40921_(_13763_, _13768_, _13770_);
  and g_40922_(_13723_, _13729_, _13771_);
  or g_40923_(_22341_, _12156_, _13773_);
  or g_40924_(_12006_, _12154_, _13774_);
  and g_40925_(_13773_, _13774_, _13775_);
  or g_40926_(_24123_, _13708_, _13776_);
  or g_40927_(_13598_, _13707_, _13777_);
  and g_40928_(_13776_, _13777_, _13778_);
  xor g_40929_(_13775_, _13778_, _13779_);
  or g_40930_(_12075_, _12154_, _13780_);
  or g_40931_(_20525_, _12156_, _13781_);
  and g_40932_(_13780_, _13781_, _13782_);
  or g_40933_(_24163_, _13708_, _13784_);
  or g_40934_(_13535_, _13707_, _13785_);
  and g_40935_(_13784_, _13785_, _13786_);
  xor g_40936_(_13782_, _13786_, _13787_);
  or g_40937_(_22356_, _12156_, _13788_);
  or g_40938_(_12058_, _12154_, _13789_);
  and g_40939_(_13788_, _13789_, _13790_);
  or g_40940_(_24141_, _13708_, _13791_);
  or g_40941_(_13654_, _13707_, _13792_);
  and g_40942_(_13791_, _13792_, _13793_);
  and g_40943_(_13762_, _13769_, _13795_);
  and g_40944_(_11981_, _12154_, _13796_);
  or g_40945_(_11982_, _12156_, _13797_);
  or g_40946_(_11987_, _12154_, _13798_);
  not g_40947_(_13798_, _13799_);
  and g_40948_(_13797_, _13798_, _13800_);
  or g_40949_(_13796_, _13799_, _13801_);
  and g_40950_(_13566_, _13707_, _13802_);
  or g_40951_(_13567_, _13708_, _13803_);
  and g_40952_(_13573_, _13708_, _13804_);
  or g_40953_(_13572_, _13707_, _13806_);
  and g_40954_(_13803_, _13806_, _13807_);
  or g_40955_(_13802_, _13804_, _13808_);
  and g_40956_(_13800_, _13808_, _13809_);
  or g_40957_(_22274_, _12156_, _13810_);
  or g_40958_(_12033_, _12154_, _13811_);
  and g_40959_(_13810_, _13811_, _13812_);
  or g_40960_(_22411_, _13708_, _13813_);
  or g_40961_(_13625_, _13707_, _13814_);
  and g_40962_(_13813_, _13814_, _13815_);
  and g_40963_(_13801_, _13807_, _13817_);
  or g_40964_(_13748_, _13770_, _13818_);
  or g_40965_(_13779_, _13818_, _13819_);
  or g_40966_(_13716_, _13817_, _13820_);
  or g_40967_(_13771_, _13820_, _13821_);
  or g_40968_(_13819_, _13821_, _13822_);
  xor g_40969_(_13812_, _13815_, _13823_);
  or g_40970_(_13756_, _13823_, _13824_);
  xor g_40971_(_13734_, _13737_, _13825_);
  or g_40972_(_13745_, _13825_, _13826_);
  or g_40973_(_13824_, _13826_, _13828_);
  or g_40974_(_13715_, _13795_, _13829_);
  or g_40975_(_13787_, _13829_, _13830_);
  xor g_40976_(_13790_, _13793_, _13831_);
  or g_40977_(_13731_, _13809_, _13832_);
  or g_40978_(_13831_, _13832_, _13833_);
  or g_40979_(_13830_, _13833_, _13834_);
  or g_40980_(_13828_, _13834_, _13835_);
  or g_40981_(_13822_, _13835_, _13836_);
  not g_40982_(_13836_, _13837_);
  or g_40983_(out[145], out[144], _13839_);
  or g_40984_(out[144], _18336_, _13840_);
  and g_40985_(out[147], _13840_, _13841_);
  and g_40986_(_26054_, _13840_, _13842_);
  and g_40987_(out[149], _13842_, _13843_);
  or g_40988_(out[150], _13843_, _13844_);
  and g_40989_(out[151], _13844_, _13845_);
  and g_40990_(out[152], _13845_, _13846_);
  xor g_40991_(out[152], _13845_, _13847_);
  xor g_40992_(out[151], _13844_, _13848_);
  or g_40993_(out[97], out[96], _13850_);
  or g_40994_(out[96], _16984_, _13851_);
  and g_40995_(out[99], _13851_, _13852_);
  and g_40996_(_25530_, _13851_, _13853_);
  and g_40997_(out[101], _13853_, _13854_);
  or g_40998_(out[102], _13854_, _13855_);
  and g_40999_(out[103], _13855_, _13856_);
  xor g_41000_(out[103], _13855_, _13857_);
  xor g_41001_(_20674_, _13855_, _13858_);
  and g_41002_(out[104], _13856_, _13859_);
  xor g_41003_(out[104], _13856_, _13861_);
  xor g_41004_(_20762_, _13856_, _13862_);
  or g_41005_(out[81], out[80], _13863_);
  or g_41006_(out[80], _14564_, _13864_);
  and g_41007_(out[83], _13864_, _13865_);
  and g_41008_(_25273_, _13864_, _13866_);
  and g_41009_(out[85], _13866_, _13867_);
  or g_41010_(out[86], _13867_, _13868_);
  and g_41011_(out[87], _13868_, _13869_);
  and g_41012_(out[88], _13869_, _13870_);
  xor g_41013_(out[88], _13869_, _13872_);
  xor g_41014_(_20630_, _13869_, _13873_);
  or g_41015_(out[89], _13870_, _13874_);
  xor g_41016_(out[89], _13870_, _13875_);
  xor g_41017_(_20641_, _13870_, _13876_);
  or g_41018_(out[65], out[64], _13877_);
  or g_41019_(out[64], _12518_, _13878_);
  and g_41020_(out[67], _13878_, _13879_);
  and g_41021_(_25039_, _13878_, _13880_);
  and g_41022_(out[69], _13880_, _13881_);
  or g_41023_(out[70], _13881_, _13883_);
  and g_41024_(out[71], _13883_, _13884_);
  and g_41025_(out[72], _13884_, _13885_);
  or g_41026_(out[73], _13885_, _13886_);
  xor g_41027_(out[73], _13885_, _13887_);
  xor g_41028_(_20509_, _13885_, _13888_);
  or g_41029_(out[49], out[48], _13889_);
  or g_41030_(out[48], _10219_, _13890_);
  and g_41031_(out[51], _13890_, _13891_);
  and g_41032_(_24803_, _13890_, _13892_);
  and g_41033_(out[53], _13892_, _13894_);
  or g_41034_(out[54], _13894_, _13895_);
  and g_41035_(out[55], _13895_, _13896_);
  and g_41036_(out[56], _13896_, _13897_);
  or g_41037_(out[57], _13897_, _13898_);
  and g_41038_(out[58], _13898_, _13899_);
  xor g_41039_(out[59], _13899_, _13900_);
  xor g_41040_(_20267_, _13899_, _13901_);
  xor g_41041_(out[51], _13890_, _13902_);
  xor g_41042_(_20355_, _13890_, _13903_);
  or g_41043_(out[33], out[32], _13905_);
  or g_41044_(out[32], _24172_, _13906_);
  and g_41045_(out[35], _13906_, _13907_);
  xor g_41046_(out[35], _13906_, _13908_);
  xor g_41047_(_20223_, _13906_, _13909_);
  and g_41048_(_24571_, _13906_, _13910_);
  and g_41049_(out[37], _13910_, _13911_);
  or g_41050_(out[38], _13911_, _13912_);
  and g_41051_(out[39], _13912_, _13913_);
  xor g_41052_(out[39], _13912_, _13914_);
  xor g_41053_(_20146_, _13912_, _13916_);
  and g_41054_(out[8], _20665_, _13917_);
  or g_41055_(out[9], _13917_, _13918_);
  xor g_41056_(out[9], _13917_, _13919_);
  xor g_41057_(_19981_, _13917_, _13920_);
  and g_41058_(out[24], _20669_, _13921_);
  or g_41059_(out[25], _13921_, _13922_);
  xor g_41060_(out[25], _13921_, _13923_);
  xor g_41061_(_20113_, _13921_, _13924_);
  and g_41062_(_13919_, _13924_, _13925_);
  or g_41063_(_13920_, _13923_, _13927_);
  and g_41064_(out[26], _13922_, _13928_);
  xor g_41065_(out[26], _13922_, _13929_);
  xor g_41066_(_20124_, _13922_, _13930_);
  and g_41067_(out[10], _13918_, _13931_);
  xor g_41068_(out[10], _13918_, _13932_);
  xor g_41069_(_19992_, _13918_, _13933_);
  and g_41070_(_13929_, _13933_, _13934_);
  or g_41071_(_13930_, _13932_, _13935_);
  and g_41072_(_13927_, _13935_, _13936_);
  or g_41073_(_13925_, _13934_, _13938_);
  xor g_41074_(out[8], _20665_, _13939_);
  xor g_41075_(_19970_, _20665_, _13940_);
  xor g_41076_(out[24], _20669_, _13941_);
  xor g_41077_(_20102_, _20669_, _13942_);
  and g_41078_(_13939_, _13942_, _13943_);
  or g_41079_(_13940_, _13941_, _13944_);
  and g_41080_(_13920_, _13923_, _13945_);
  or g_41081_(_13919_, _13924_, _13946_);
  and g_41082_(_13944_, _13946_, _13947_);
  or g_41083_(_13943_, _13945_, _13949_);
  and g_41084_(_20673_, _20682_, _13950_);
  or g_41085_(_20672_, _20681_, _13951_);
  xor g_41086_(out[19], _23127_, _13952_);
  xor g_41087_(_20091_, _23127_, _13953_);
  xor g_41088_(out[3], _23039_, _13954_);
  xor g_41089_(_19959_, _23039_, _13955_);
  and g_41090_(_13953_, _13954_, _13956_);
  or g_41091_(_13952_, _13955_, _13957_);
  xor g_41092_(out[2], _23017_, _13958_);
  xor g_41093_(_19948_, _23017_, _13960_);
  xor g_41094_(out[18], _23105_, _13961_);
  xor g_41095_(_20080_, _23105_, _13962_);
  and g_41096_(_13958_, _13962_, _13963_);
  or g_41097_(_13960_, _13961_, _13964_);
  and g_41098_(out[1], _22621_, _13965_);
  or g_41099_(_19926_, _22610_, _13966_);
  and g_41100_(out[17], _13966_, _13967_);
  or g_41101_(_20058_, _13965_, _13968_);
  and g_41102_(_23105_, _13968_, _13969_);
  or g_41103_(_23116_, _13967_, _13971_);
  and g_41104_(_13960_, _13961_, _13972_);
  or g_41105_(_13958_, _13962_, _13973_);
  and g_41106_(_23017_, _13973_, _13974_);
  or g_41107_(_23028_, _13972_, _13975_);
  and g_41108_(_13971_, _13974_, _13976_);
  or g_41109_(_13969_, _13975_, _13977_);
  and g_41110_(_13964_, _13977_, _13978_);
  or g_41111_(_13963_, _13976_, _13979_);
  and g_41112_(_13957_, _13979_, _13980_);
  or g_41113_(_13956_, _13978_, _13982_);
  and g_41114_(_13952_, _13955_, _13983_);
  or g_41115_(_13953_, _13954_, _13984_);
  and g_41116_(_23204_, _13984_, _13985_);
  or g_41117_(_23193_, _13983_, _13986_);
  and g_41118_(_13982_, _13985_, _13987_);
  or g_41119_(_13980_, _13986_, _13988_);
  and g_41120_(_23347_, _13988_, _13989_);
  or g_41121_(_23358_, _13987_, _13990_);
  and g_41122_(_23292_, _20684_, _13991_);
  or g_41123_(_23281_, _20683_, _13993_);
  and g_41124_(_22819_, _23204_, _13994_);
  or g_41125_(_22830_, _23193_, _13995_);
  and g_41126_(_23347_, _13994_, _13996_);
  or g_41127_(_23358_, _13995_, _13997_);
  and g_41128_(_13991_, _13997_, _13998_);
  or g_41129_(_13993_, _13996_, _13999_);
  and g_41130_(_13990_, _13998_, _14000_);
  or g_41131_(_13989_, _13999_, _14001_);
  and g_41132_(_13950_, _14001_, _14002_);
  or g_41133_(_13951_, _14000_, _14004_);
  and g_41134_(_13940_, _13941_, _14005_);
  or g_41135_(_13939_, _13942_, _14006_);
  and g_41136_(_20676_, _14006_, _14007_);
  or g_41137_(_20675_, _14005_, _14008_);
  and g_41138_(_14004_, _14007_, _14009_);
  or g_41139_(_14002_, _14008_, _14010_);
  and g_41140_(_13947_, _14010_, _14011_);
  or g_41141_(_13949_, _14009_, _14012_);
  and g_41142_(_13936_, _14012_, _14013_);
  or g_41143_(_13938_, _14011_, _14015_);
  xor g_41144_(out[27], _13928_, _14016_);
  xor g_41145_(_20003_, _13928_, _14017_);
  xor g_41146_(out[11], _13931_, _14018_);
  xor g_41147_(_19871_, _13931_, _14019_);
  and g_41148_(_14017_, _14018_, _14020_);
  or g_41149_(_14016_, _14019_, _14021_);
  and g_41150_(_13930_, _13932_, _14022_);
  or g_41151_(_13929_, _13933_, _14023_);
  and g_41152_(_14021_, _14023_, _14024_);
  or g_41153_(_14020_, _14022_, _14026_);
  and g_41154_(_14015_, _14024_, _14027_);
  or g_41155_(_14013_, _14026_, _14028_);
  and g_41156_(_14016_, _14019_, _14029_);
  or g_41157_(_14017_, _14018_, _14030_);
  and g_41158_(_14028_, _14030_, _14031_);
  or g_41159_(_14027_, _14029_, _14032_);
  and g_41160_(_20667_, _14032_, _14033_);
  or g_41161_(_20666_, _14031_, _14034_);
  and g_41162_(_20671_, _14031_, _14035_);
  or g_41163_(_20670_, _14032_, _14037_);
  and g_41164_(_14034_, _14037_, _14038_);
  or g_41165_(_14033_, _14035_, _14039_);
  and g_41166_(_13914_, _14039_, _14040_);
  or g_41167_(_13916_, _14038_, _14041_);
  xor g_41168_(out[38], _13911_, _14042_);
  xor g_41169_(_20157_, _13911_, _14043_);
  and g_41170_(_20677_, _14032_, _14044_);
  or g_41171_(_20678_, _14031_, _14045_);
  and g_41172_(_20679_, _14031_, _14046_);
  or g_41173_(_20680_, _14032_, _14048_);
  and g_41174_(_14045_, _14048_, _14049_);
  or g_41175_(_14044_, _14046_, _14050_);
  and g_41176_(_14042_, _14049_, _14051_);
  or g_41177_(_14043_, _14050_, _14052_);
  xor g_41178_(_20190_, out[32], _14053_);
  not g_41179_(_14053_, _14054_);
  xor g_41180_(out[17], out[16], _14055_);
  xor g_41181_(_20058_, out[16], _14056_);
  and g_41182_(_14031_, _14055_, _14057_);
  or g_41183_(_14032_, _14056_, _14059_);
  xor g_41184_(out[1], out[0], _14060_);
  xor g_41185_(_19926_, out[0], _14061_);
  and g_41186_(_14032_, _14060_, _14062_);
  or g_41187_(_14031_, _14061_, _14063_);
  and g_41188_(_14059_, _14063_, _14064_);
  or g_41189_(_14057_, _14062_, _14065_);
  and g_41190_(_14054_, _14064_, _14066_);
  or g_41191_(_14053_, _14065_, _14067_);
  and g_41192_(out[16], _14031_, _14068_);
  or g_41193_(_20069_, _14032_, _14070_);
  and g_41194_(out[0], _14032_, _14071_);
  or g_41195_(_19937_, _14031_, _14072_);
  and g_41196_(_14070_, _14072_, _14073_);
  or g_41197_(_14068_, _14071_, _14074_);
  and g_41198_(out[32], _14073_, _14075_);
  or g_41199_(_20201_, _14074_, _14076_);
  and g_41200_(_14067_, _14076_, _14077_);
  or g_41201_(_14066_, _14075_, _14078_);
  xor g_41202_(out[34], _13905_, _14079_);
  xor g_41203_(_20212_, _13905_, _14081_);
  and g_41204_(_13961_, _14031_, _14082_);
  or g_41205_(_13962_, _14032_, _14083_);
  and g_41206_(_13958_, _14032_, _14084_);
  or g_41207_(_13960_, _14031_, _14085_);
  and g_41208_(_14083_, _14085_, _14086_);
  or g_41209_(_14082_, _14084_, _14087_);
  and g_41210_(_14081_, _14087_, _14088_);
  or g_41211_(_14079_, _14086_, _14089_);
  and g_41212_(out[33], _14065_, _14090_);
  or g_41213_(_20190_, _14064_, _14092_);
  and g_41214_(_14089_, _14092_, _14093_);
  or g_41215_(_14088_, _14090_, _14094_);
  and g_41216_(_14078_, _14093_, _14095_);
  or g_41217_(_14077_, _14094_, _14096_);
  and g_41218_(_13955_, _14032_, _14097_);
  or g_41219_(_13954_, _14031_, _14098_);
  and g_41220_(_13953_, _14031_, _14099_);
  or g_41221_(_13952_, _14032_, _14100_);
  and g_41222_(_14098_, _14100_, _14101_);
  or g_41223_(_14097_, _14099_, _14103_);
  and g_41224_(_13909_, _14101_, _14104_);
  or g_41225_(_13908_, _14103_, _14105_);
  and g_41226_(_14079_, _14086_, _14106_);
  or g_41227_(_14081_, _14087_, _14107_);
  and g_41228_(_14105_, _14107_, _14108_);
  or g_41229_(_14104_, _14106_, _14109_);
  and g_41230_(_14096_, _14108_, _14110_);
  or g_41231_(_14095_, _14109_, _14111_);
  xor g_41232_(out[36], _13907_, _14112_);
  xor g_41233_(_20179_, _13907_, _14114_);
  and g_41234_(_23182_, _14031_, _14115_);
  or g_41235_(_23171_, _14032_, _14116_);
  and g_41236_(_23094_, _14032_, _14117_);
  or g_41237_(_23083_, _14031_, _14118_);
  and g_41238_(_14116_, _14118_, _14119_);
  or g_41239_(_14115_, _14117_, _14120_);
  and g_41240_(_14112_, _14120_, _14121_);
  or g_41241_(_14114_, _14119_, _14122_);
  and g_41242_(_13908_, _14103_, _14123_);
  or g_41243_(_13909_, _14101_, _14125_);
  and g_41244_(_14122_, _14125_, _14126_);
  or g_41245_(_14121_, _14123_, _14127_);
  and g_41246_(_14111_, _14126_, _14128_);
  or g_41247_(_14110_, _14127_, _14129_);
  xor g_41248_(out[37], _13910_, _14130_);
  xor g_41249_(_20168_, _13910_, _14131_);
  and g_41250_(_23270_, _14031_, _14132_);
  or g_41251_(_23259_, _14032_, _14133_);
  and g_41252_(_23237_, _14032_, _14134_);
  or g_41253_(_23226_, _14031_, _14136_);
  and g_41254_(_14133_, _14136_, _14137_);
  or g_41255_(_14132_, _14134_, _14138_);
  and g_41256_(_14131_, _14137_, _14139_);
  or g_41257_(_14130_, _14138_, _14140_);
  and g_41258_(_14114_, _14119_, _14141_);
  or g_41259_(_14112_, _14120_, _14142_);
  and g_41260_(_14140_, _14142_, _14143_);
  or g_41261_(_14139_, _14141_, _14144_);
  and g_41262_(_14129_, _14143_, _14145_);
  or g_41263_(_14128_, _14144_, _14147_);
  and g_41264_(_14043_, _14050_, _14148_);
  or g_41265_(_14042_, _14049_, _14149_);
  and g_41266_(_14130_, _14138_, _14150_);
  or g_41267_(_14131_, _14137_, _14151_);
  and g_41268_(_14149_, _14151_, _14152_);
  or g_41269_(_14148_, _14150_, _14153_);
  and g_41270_(_14147_, _14152_, _14154_);
  or g_41271_(_14145_, _14153_, _14155_);
  and g_41272_(_14052_, _14155_, _14156_);
  or g_41273_(_14051_, _14154_, _14158_);
  and g_41274_(_14041_, _14158_, _14159_);
  or g_41275_(_14040_, _14156_, _14160_);
  and g_41276_(out[40], _13913_, _14161_);
  or g_41277_(out[41], _14161_, _14162_);
  and g_41278_(out[42], _14162_, _14163_);
  xor g_41279_(out[42], _14162_, _14164_);
  not g_41280_(_14164_, _14165_);
  and g_41281_(_13932_, _14032_, _14166_);
  or g_41282_(_13933_, _14031_, _14167_);
  and g_41283_(_13929_, _14031_, _14169_);
  or g_41284_(_13930_, _14032_, _14170_);
  and g_41285_(_14167_, _14170_, _14171_);
  or g_41286_(_14166_, _14169_, _14172_);
  and g_41287_(_14164_, _14171_, _14173_);
  and g_41288_(_14016_, _14018_, _14174_);
  or g_41289_(_14017_, _14019_, _14175_);
  xor g_41290_(out[43], _14163_, _14176_);
  not g_41291_(_14176_, _14177_);
  and g_41292_(_14175_, _14176_, _14178_);
  or g_41293_(_14173_, _14178_, _14180_);
  and g_41294_(_14165_, _14172_, _14181_);
  and g_41295_(_14174_, _14177_, _14182_);
  or g_41296_(_14175_, _14176_, _14183_);
  or g_41297_(_14181_, _14182_, _14184_);
  xor g_41298_(_14164_, _14171_, _14185_);
  xor g_41299_(_14175_, _14176_, _14186_);
  and g_41300_(_14185_, _14186_, _14187_);
  or g_41301_(_14180_, _14184_, _14188_);
  xor g_41302_(out[40], _13913_, _14189_);
  not g_41303_(_14189_, _14191_);
  and g_41304_(_13939_, _14032_, _14192_);
  or g_41305_(_13940_, _14031_, _14193_);
  and g_41306_(_13941_, _14031_, _14194_);
  or g_41307_(_13942_, _14032_, _14195_);
  and g_41308_(_14193_, _14195_, _14196_);
  or g_41309_(_14192_, _14194_, _14197_);
  and g_41310_(_14189_, _14196_, _14198_);
  and g_41311_(_14191_, _14197_, _14199_);
  xor g_41312_(_14189_, _14196_, _14200_);
  and g_41313_(_13916_, _14038_, _14202_);
  or g_41314_(_13914_, _14039_, _14203_);
  xor g_41315_(out[41], _14161_, _14204_);
  xor g_41316_(_20245_, _14161_, _14205_);
  and g_41317_(_13919_, _14032_, _14206_);
  or g_41318_(_13920_, _14031_, _14207_);
  and g_41319_(_13923_, _14031_, _14208_);
  or g_41320_(_13924_, _14032_, _14209_);
  and g_41321_(_14207_, _14209_, _14210_);
  or g_41322_(_14206_, _14208_, _14211_);
  and g_41323_(_14205_, _14211_, _14213_);
  or g_41324_(_14204_, _14210_, _14214_);
  and g_41325_(_14203_, _14214_, _14215_);
  or g_41326_(_14202_, _14213_, _14216_);
  and g_41327_(_14204_, _14210_, _14217_);
  or g_41328_(_14205_, _14211_, _14218_);
  and g_41329_(_14215_, _14218_, _14219_);
  and g_41330_(_14200_, _14219_, _14220_);
  or g_41331_(_14199_, _14217_, _14221_);
  or g_41332_(_14216_, _14221_, _14222_);
  or g_41333_(_14188_, _14222_, _14224_);
  and g_41334_(_14187_, _14220_, _14225_);
  or g_41335_(_14198_, _14224_, _14226_);
  and g_41336_(_14160_, _14225_, _14227_);
  or g_41337_(_14159_, _14226_, _14228_);
  or g_41338_(_14198_, _14213_, _14229_);
  and g_41339_(_14187_, _14229_, _14230_);
  and g_41340_(_14218_, _14230_, _14231_);
  and g_41341_(_14180_, _14183_, _14232_);
  or g_41342_(_14231_, _14232_, _14233_);
  not g_41343_(_14233_, _14235_);
  and g_41344_(_14228_, _14235_, _14236_);
  or g_41345_(_14227_, _14233_, _14237_);
  or g_41346_(_13908_, _14237_, _14238_);
  not g_41347_(_14238_, _14239_);
  and g_41348_(_14103_, _14237_, _14240_);
  or g_41349_(_14101_, _14236_, _14241_);
  and g_41350_(_14238_, _14241_, _14242_);
  or g_41351_(_14239_, _14240_, _14243_);
  and g_41352_(_13903_, _14242_, _14244_);
  or g_41353_(_13902_, _14243_, _14246_);
  xor g_41354_(out[50], _13889_, _14247_);
  not g_41355_(_14247_, _14248_);
  and g_41356_(_14079_, _14236_, _14249_);
  or g_41357_(_14081_, _14237_, _14250_);
  and g_41358_(_14087_, _14237_, _14251_);
  not g_41359_(_14251_, _14252_);
  and g_41360_(_14250_, _14252_, _14253_);
  or g_41361_(_14249_, _14251_, _14254_);
  and g_41362_(_14247_, _14253_, _14255_);
  or g_41363_(_14248_, _14254_, _14257_);
  and g_41364_(_14246_, _14257_, _14258_);
  or g_41365_(_14244_, _14255_, _14259_);
  and g_41366_(_13902_, _14243_, _14260_);
  or g_41367_(_13903_, _14242_, _14261_);
  and g_41368_(_14248_, _14254_, _14262_);
  or g_41369_(_14247_, _14253_, _14263_);
  and g_41370_(_14261_, _14263_, _14264_);
  or g_41371_(_14260_, _14262_, _14265_);
  and g_41372_(_14258_, _14264_, _14266_);
  or g_41373_(_14259_, _14265_, _14268_);
  xor g_41374_(out[49], out[48], _14269_);
  xor g_41375_(_20322_, out[48], _14270_);
  or g_41376_(_14053_, _14237_, _14271_);
  or g_41377_(_14064_, _14236_, _14272_);
  and g_41378_(_14271_, _14272_, _14273_);
  and g_41379_(_14269_, _14273_, _14274_);
  not g_41380_(_14274_, _14275_);
  and g_41381_(out[32], _14236_, _14276_);
  or g_41382_(_20201_, _14237_, _14277_);
  and g_41383_(_14074_, _14237_, _14279_);
  not g_41384_(_14279_, _14280_);
  and g_41385_(_14277_, _14280_, _14281_);
  or g_41386_(_14276_, _14279_, _14282_);
  and g_41387_(_20333_, _14282_, _14283_);
  or g_41388_(out[48], _14281_, _14284_);
  xor g_41389_(_14269_, _14273_, _14285_);
  xor g_41390_(_14270_, _14273_, _14286_);
  and g_41391_(_14284_, _14285_, _14287_);
  or g_41392_(_14283_, _14286_, _14288_);
  and g_41393_(_14275_, _14288_, _14290_);
  or g_41394_(_14274_, _14287_, _14291_);
  and g_41395_(_14266_, _14291_, _14292_);
  or g_41396_(_14268_, _14290_, _14293_);
  and g_41397_(_14259_, _14261_, _14294_);
  or g_41398_(_14258_, _14260_, _14295_);
  and g_41399_(_14293_, _14295_, _14296_);
  or g_41400_(_14292_, _14294_, _14297_);
  xor g_41401_(out[58], _13898_, _14298_);
  xor g_41402_(_20388_, _13898_, _14299_);
  and g_41403_(_14171_, _14237_, _14301_);
  or g_41404_(_14172_, _14236_, _14302_);
  and g_41405_(_14165_, _14236_, _14303_);
  or g_41406_(_14164_, _14237_, _14304_);
  and g_41407_(_14302_, _14304_, _14305_);
  or g_41408_(_14301_, _14303_, _14306_);
  and g_41409_(_14298_, _14306_, _14307_);
  or g_41410_(_14299_, _14305_, _14308_);
  and g_41411_(_14174_, _14176_, _14309_);
  or g_41412_(_14175_, _14177_, _14310_);
  and g_41413_(_13900_, _14310_, _14312_);
  or g_41414_(_13901_, _14309_, _14313_);
  and g_41415_(_14308_, _14313_, _14314_);
  or g_41416_(_14307_, _14312_, _14315_);
  xor g_41417_(out[56], _13896_, _14316_);
  xor g_41418_(_20366_, _13896_, _14317_);
  and g_41419_(_14196_, _14237_, _14318_);
  or g_41420_(_14197_, _14236_, _14319_);
  and g_41421_(_14191_, _14236_, _14320_);
  or g_41422_(_14189_, _14237_, _14321_);
  and g_41423_(_14319_, _14321_, _14323_);
  or g_41424_(_14318_, _14320_, _14324_);
  and g_41425_(_14316_, _14324_, _14325_);
  or g_41426_(_14317_, _14323_, _14326_);
  xor g_41427_(out[57], _13897_, _14327_);
  xor g_41428_(_20377_, _13897_, _14328_);
  and g_41429_(_14211_, _14237_, _14329_);
  or g_41430_(_14210_, _14236_, _14330_);
  and g_41431_(_14204_, _14236_, _14331_);
  or g_41432_(_14205_, _14237_, _14332_);
  and g_41433_(_14330_, _14332_, _14334_);
  or g_41434_(_14329_, _14331_, _14335_);
  and g_41435_(_14328_, _14335_, _14336_);
  or g_41436_(_14327_, _14334_, _14337_);
  and g_41437_(_14326_, _14337_, _14338_);
  or g_41438_(_14325_, _14336_, _14339_);
  and g_41439_(_14314_, _14338_, _14340_);
  or g_41440_(_14315_, _14339_, _14341_);
  and g_41441_(_13901_, _14309_, _14342_);
  or g_41442_(_13900_, _14310_, _14343_);
  and g_41443_(_14299_, _14305_, _14345_);
  or g_41444_(_14298_, _14306_, _14346_);
  and g_41445_(_14343_, _14346_, _14347_);
  or g_41446_(_14342_, _14345_, _14348_);
  and g_41447_(_14327_, _14334_, _14349_);
  or g_41448_(_14328_, _14335_, _14350_);
  and g_41449_(_14317_, _14323_, _14351_);
  or g_41450_(_14316_, _14324_, _14352_);
  and g_41451_(_14350_, _14352_, _14353_);
  or g_41452_(_14349_, _14351_, _14354_);
  and g_41453_(_14347_, _14353_, _14356_);
  or g_41454_(_14348_, _14354_, _14357_);
  and g_41455_(_14340_, _14356_, _14358_);
  or g_41456_(_14341_, _14357_, _14359_);
  xor g_41457_(out[55], _13895_, _14360_);
  xor g_41458_(_20278_, _13895_, _14361_);
  and g_41459_(_14039_, _14237_, _14362_);
  or g_41460_(_14038_, _14236_, _14363_);
  and g_41461_(_13916_, _14236_, _14364_);
  or g_41462_(_13914_, _14237_, _14365_);
  and g_41463_(_14363_, _14365_, _14367_);
  or g_41464_(_14362_, _14364_, _14368_);
  and g_41465_(_14361_, _14367_, _14369_);
  or g_41466_(_14360_, _14368_, _14370_);
  xor g_41467_(out[54], _13894_, _14371_);
  xor g_41468_(_20289_, _13894_, _14372_);
  and g_41469_(_14050_, _14237_, _14373_);
  or g_41470_(_14049_, _14236_, _14374_);
  and g_41471_(_14042_, _14236_, _14375_);
  or g_41472_(_14043_, _14237_, _14376_);
  and g_41473_(_14374_, _14376_, _14378_);
  or g_41474_(_14373_, _14375_, _14379_);
  and g_41475_(_14371_, _14378_, _14380_);
  or g_41476_(_14372_, _14379_, _14381_);
  and g_41477_(_14370_, _14381_, _14382_);
  or g_41478_(_14369_, _14380_, _14383_);
  and g_41479_(_14372_, _14379_, _14384_);
  or g_41480_(_14371_, _14378_, _14385_);
  and g_41481_(_14360_, _14368_, _14386_);
  or g_41482_(_14361_, _14367_, _14387_);
  and g_41483_(_14385_, _14387_, _14389_);
  or g_41484_(_14384_, _14386_, _14390_);
  and g_41485_(_14382_, _14389_, _14391_);
  or g_41486_(_14383_, _14390_, _14392_);
  xor g_41487_(out[52], _13891_, _14393_);
  xor g_41488_(_20311_, _13891_, _14394_);
  and g_41489_(_14114_, _14236_, _14395_);
  or g_41490_(_14112_, _14237_, _14396_);
  and g_41491_(_14120_, _14237_, _14397_);
  or g_41492_(_14119_, _14236_, _14398_);
  and g_41493_(_14396_, _14398_, _14400_);
  or g_41494_(_14395_, _14397_, _14401_);
  and g_41495_(_14394_, _14400_, _14402_);
  or g_41496_(_14393_, _14401_, _14403_);
  xor g_41497_(out[53], _13892_, _14404_);
  xor g_41498_(_20300_, _13892_, _14405_);
  and g_41499_(_14131_, _14236_, _14406_);
  or g_41500_(_14130_, _14237_, _14407_);
  and g_41501_(_14138_, _14237_, _14408_);
  or g_41502_(_14137_, _14236_, _14409_);
  and g_41503_(_14407_, _14409_, _14411_);
  or g_41504_(_14406_, _14408_, _14412_);
  and g_41505_(_14405_, _14411_, _14413_);
  or g_41506_(_14404_, _14412_, _14414_);
  and g_41507_(_14403_, _14414_, _14415_);
  or g_41508_(_14402_, _14413_, _14416_);
  and g_41509_(_14404_, _14412_, _14417_);
  or g_41510_(_14405_, _14411_, _14418_);
  and g_41511_(_14393_, _14401_, _14419_);
  or g_41512_(_14394_, _14400_, _14420_);
  and g_41513_(_14418_, _14420_, _14422_);
  or g_41514_(_14417_, _14419_, _14423_);
  and g_41515_(_14415_, _14422_, _14424_);
  or g_41516_(_14416_, _14423_, _14425_);
  and g_41517_(_14391_, _14424_, _14426_);
  or g_41518_(_14392_, _14425_, _14427_);
  and g_41519_(_14358_, _14426_, _14428_);
  or g_41520_(_14359_, _14427_, _14429_);
  and g_41521_(_14297_, _14428_, _14430_);
  or g_41522_(_14296_, _14429_, _14431_);
  and g_41523_(_14383_, _14387_, _14433_);
  or g_41524_(_14382_, _14386_, _14434_);
  and g_41525_(_14416_, _14418_, _14435_);
  or g_41526_(_14415_, _14417_, _14436_);
  and g_41527_(_14391_, _14435_, _14437_);
  or g_41528_(_14392_, _14436_, _14438_);
  and g_41529_(_14434_, _14438_, _14439_);
  or g_41530_(_14433_, _14437_, _14440_);
  and g_41531_(_14358_, _14440_, _14441_);
  or g_41532_(_14359_, _14439_, _14442_);
  and g_41533_(_14308_, _14337_, _14444_);
  or g_41534_(_14307_, _14336_, _14445_);
  and g_41535_(_14354_, _14444_, _14446_);
  or g_41536_(_14353_, _14445_, _14447_);
  and g_41537_(_14347_, _14447_, _14448_);
  or g_41538_(_14348_, _14446_, _14449_);
  and g_41539_(_14313_, _14449_, _14450_);
  or g_41540_(_14312_, _14448_, _14451_);
  and g_41541_(_14442_, _14451_, _14452_);
  or g_41542_(_14441_, _14450_, _14453_);
  and g_41543_(_14431_, _14452_, _14455_);
  or g_41544_(_14430_, _14453_, _14456_);
  and g_41545_(out[48], _14281_, _14457_);
  or g_41546_(_20333_, _14282_, _14458_);
  and g_41547_(_14266_, _14287_, _14459_);
  or g_41548_(_14268_, _14288_, _14460_);
  and g_41549_(_14428_, _14459_, _14461_);
  or g_41550_(_14429_, _14460_, _14462_);
  and g_41551_(_14458_, _14461_, _14463_);
  or g_41552_(_14457_, _14462_, _14464_);
  and g_41553_(_14456_, _14464_, _14466_);
  or g_41554_(_14455_, _14463_, _14467_);
  and g_41555_(_13901_, _14466_, _14468_);
  or g_41556_(_13900_, _14467_, _14469_);
  and g_41557_(_14310_, _14467_, _14470_);
  or g_41558_(_14309_, _14466_, _14471_);
  and g_41559_(_14469_, _14471_, _14472_);
  or g_41560_(_14468_, _14470_, _14473_);
  and g_41561_(out[74], _13886_, _14474_);
  xor g_41562_(out[75], _14474_, _14475_);
  xor g_41563_(_20399_, _14474_, _14477_);
  and g_41564_(_14472_, _14477_, _14478_);
  or g_41565_(_14473_, _14475_, _14479_);
  xor g_41566_(out[74], _13886_, _14480_);
  xor g_41567_(_20520_, _13886_, _14481_);
  and g_41568_(_14299_, _14466_, _14482_);
  or g_41569_(_14298_, _14467_, _14483_);
  and g_41570_(_14306_, _14467_, _14484_);
  or g_41571_(_14305_, _14466_, _14485_);
  and g_41572_(_14483_, _14485_, _14486_);
  or g_41573_(_14482_, _14484_, _14488_);
  and g_41574_(_14481_, _14486_, _14489_);
  or g_41575_(_14480_, _14488_, _14490_);
  and g_41576_(_14479_, _14490_, _14491_);
  or g_41577_(_14478_, _14489_, _14492_);
  and g_41578_(_14473_, _14475_, _14493_);
  or g_41579_(_14472_, _14477_, _14494_);
  and g_41580_(_14480_, _14488_, _14495_);
  or g_41581_(_14481_, _14486_, _14496_);
  and g_41582_(_14494_, _14496_, _14497_);
  or g_41583_(_14493_, _14495_, _14499_);
  and g_41584_(_14327_, _14466_, _14500_);
  or g_41585_(_14328_, _14467_, _14501_);
  and g_41586_(_14335_, _14467_, _14502_);
  or g_41587_(_14334_, _14466_, _14503_);
  and g_41588_(_14501_, _14503_, _14504_);
  or g_41589_(_14500_, _14502_, _14505_);
  and g_41590_(_13888_, _14505_, _14506_);
  or g_41591_(_13887_, _14504_, _14507_);
  and g_41592_(_14491_, _14497_, _14508_);
  or g_41593_(_14492_, _14499_, _14510_);
  and g_41594_(_14507_, _14508_, _14511_);
  or g_41595_(_14506_, _14510_, _14512_);
  xor g_41596_(out[72], _13884_, _14513_);
  xor g_41597_(_20498_, _13884_, _14514_);
  and g_41598_(_14317_, _14466_, _14515_);
  or g_41599_(_14316_, _14467_, _14516_);
  and g_41600_(_14324_, _14467_, _14517_);
  or g_41601_(_14323_, _14466_, _14518_);
  and g_41602_(_14516_, _14518_, _14519_);
  or g_41603_(_14515_, _14517_, _14521_);
  and g_41604_(_14513_, _14521_, _14522_);
  or g_41605_(_14514_, _14519_, _14523_);
  and g_41606_(_13887_, _14504_, _14524_);
  or g_41607_(_13888_, _14505_, _14525_);
  and g_41608_(_14514_, _14519_, _14526_);
  or g_41609_(_14513_, _14521_, _14527_);
  and g_41610_(_14525_, _14527_, _14528_);
  or g_41611_(_14524_, _14526_, _14529_);
  and g_41612_(_14523_, _14528_, _14530_);
  or g_41613_(_14522_, _14529_, _14532_);
  and g_41614_(_14511_, _14530_, _14533_);
  or g_41615_(_14512_, _14532_, _14534_);
  xor g_41616_(out[66], _13877_, _14535_);
  xor g_41617_(_20476_, _13877_, _14536_);
  and g_41618_(_14247_, _14466_, _14537_);
  not g_41619_(_14537_, _14538_);
  and g_41620_(_14254_, _14467_, _14539_);
  or g_41621_(_14253_, _14466_, _14540_);
  and g_41622_(_14538_, _14540_, _14541_);
  or g_41623_(_14537_, _14539_, _14543_);
  and g_41624_(_14535_, _14541_, _14544_);
  or g_41625_(_14536_, _14543_, _14545_);
  xor g_41626_(out[67], _13878_, _14546_);
  xor g_41627_(_20487_, _13878_, _14547_);
  and g_41628_(_13903_, _14466_, _14548_);
  or g_41629_(_13902_, _14467_, _14549_);
  and g_41630_(_14243_, _14467_, _14550_);
  or g_41631_(_14242_, _14466_, _14551_);
  and g_41632_(_14549_, _14551_, _14552_);
  or g_41633_(_14548_, _14550_, _14554_);
  and g_41634_(_14547_, _14552_, _14555_);
  or g_41635_(_14546_, _14554_, _14556_);
  and g_41636_(_14545_, _14556_, _14557_);
  or g_41637_(_14544_, _14555_, _14558_);
  xor g_41638_(out[65], out[64], _14559_);
  not g_41639_(_14559_, _14560_);
  or g_41640_(_14270_, _14467_, _14561_);
  or g_41641_(_14273_, _14466_, _14562_);
  and g_41642_(_14561_, _14562_, _14563_);
  not g_41643_(_14563_, _14565_);
  and g_41644_(_14559_, _14563_, _14566_);
  not g_41645_(_14566_, _14567_);
  and g_41646_(out[48], _14466_, _14568_);
  or g_41647_(_20333_, _14467_, _14569_);
  and g_41648_(_14282_, _14467_, _14570_);
  or g_41649_(_14281_, _14466_, _14571_);
  and g_41650_(_14569_, _14571_, _14572_);
  or g_41651_(_14568_, _14570_, _14573_);
  and g_41652_(_20465_, _14573_, _14574_);
  or g_41653_(out[64], _14572_, _14576_);
  xor g_41654_(_14559_, _14563_, _14577_);
  xor g_41655_(_14560_, _14563_, _14578_);
  and g_41656_(_14576_, _14577_, _14579_);
  or g_41657_(_14574_, _14578_, _14580_);
  and g_41658_(_14567_, _14580_, _14581_);
  or g_41659_(_14566_, _14579_, _14582_);
  and g_41660_(_14536_, _14543_, _14583_);
  or g_41661_(_14535_, _14541_, _14584_);
  and g_41662_(_14582_, _14584_, _14585_);
  or g_41663_(_14581_, _14583_, _14587_);
  and g_41664_(_14557_, _14587_, _14588_);
  or g_41665_(_14558_, _14585_, _14589_);
  xor g_41666_(out[71], _13883_, _14590_);
  not g_41667_(_14590_, _14591_);
  and g_41668_(_14361_, _14466_, _14592_);
  or g_41669_(_14360_, _14467_, _14593_);
  and g_41670_(_14368_, _14467_, _14594_);
  or g_41671_(_14367_, _14466_, _14595_);
  and g_41672_(_14593_, _14595_, _14596_);
  or g_41673_(_14592_, _14594_, _14598_);
  or g_41674_(_14590_, _14598_, _14599_);
  xor g_41675_(out[70], _13881_, _14600_);
  not g_41676_(_14600_, _14601_);
  and g_41677_(_14371_, _14466_, _14602_);
  or g_41678_(_14372_, _14467_, _14603_);
  and g_41679_(_14379_, _14467_, _14604_);
  or g_41680_(_14378_, _14466_, _14605_);
  and g_41681_(_14603_, _14605_, _14606_);
  or g_41682_(_14602_, _14604_, _14607_);
  or g_41683_(_14601_, _14607_, _14609_);
  and g_41684_(_14599_, _14609_, _14610_);
  and g_41685_(_14590_, _14598_, _14611_);
  or g_41686_(_14591_, _14596_, _14612_);
  or g_41687_(_14600_, _14606_, _14613_);
  and g_41688_(_14612_, _14613_, _14614_);
  xor g_41689_(_14590_, _14596_, _14615_);
  xor g_41690_(_14601_, _14606_, _14616_);
  and g_41691_(_14610_, _14614_, _14617_);
  or g_41692_(_14615_, _14616_, _14618_);
  xor g_41693_(out[69], _13880_, _14620_);
  xor g_41694_(_20432_, _13880_, _14621_);
  and g_41695_(_14405_, _14466_, _14622_);
  or g_41696_(_14404_, _14467_, _14623_);
  and g_41697_(_14412_, _14467_, _14624_);
  or g_41698_(_14411_, _14466_, _14625_);
  and g_41699_(_14623_, _14625_, _14626_);
  or g_41700_(_14622_, _14624_, _14627_);
  and g_41701_(_14621_, _14626_, _14628_);
  or g_41702_(_14620_, _14627_, _14629_);
  xor g_41703_(out[68], _13879_, _14631_);
  xor g_41704_(_20443_, _13879_, _14632_);
  and g_41705_(_14394_, _14466_, _14633_);
  or g_41706_(_14393_, _14467_, _14634_);
  and g_41707_(_14401_, _14467_, _14635_);
  or g_41708_(_14400_, _14466_, _14636_);
  and g_41709_(_14634_, _14636_, _14637_);
  or g_41710_(_14633_, _14635_, _14638_);
  and g_41711_(_14632_, _14637_, _14639_);
  or g_41712_(_14631_, _14638_, _14640_);
  and g_41713_(_14629_, _14640_, _14642_);
  or g_41714_(_14628_, _14639_, _14643_);
  and g_41715_(_14631_, _14638_, _14644_);
  or g_41716_(_14632_, _14637_, _14645_);
  and g_41717_(_14546_, _14554_, _14646_);
  or g_41718_(_14547_, _14552_, _14647_);
  and g_41719_(_14620_, _14627_, _14648_);
  or g_41720_(_14621_, _14626_, _14649_);
  and g_41721_(_14645_, _14649_, _14650_);
  or g_41722_(_14644_, _14648_, _14651_);
  and g_41723_(_14642_, _14650_, _14653_);
  or g_41724_(_14643_, _14651_, _14654_);
  and g_41725_(_14617_, _14653_, _14655_);
  or g_41726_(_14618_, _14654_, _14656_);
  and g_41727_(_14647_, _14655_, _14657_);
  or g_41728_(_14646_, _14656_, _14658_);
  and g_41729_(_14589_, _14657_, _14659_);
  or g_41730_(_14588_, _14658_, _14660_);
  or g_41731_(_14610_, _14611_, _14661_);
  or g_41732_(_14642_, _14648_, _14662_);
  or g_41733_(_14618_, _14662_, _14664_);
  and g_41734_(_14661_, _14664_, _14665_);
  not g_41735_(_14665_, _14666_);
  and g_41736_(_14660_, _14665_, _14667_);
  or g_41737_(_14659_, _14666_, _14668_);
  and g_41738_(_14533_, _14668_, _14669_);
  or g_41739_(_14534_, _14667_, _14670_);
  and g_41740_(_14492_, _14494_, _14671_);
  or g_41741_(_14491_, _14493_, _14672_);
  and g_41742_(_14511_, _14529_, _14673_);
  or g_41743_(_14512_, _14528_, _14675_);
  and g_41744_(_14672_, _14675_, _14676_);
  or g_41745_(_14671_, _14673_, _14677_);
  and g_41746_(_14670_, _14676_, _14678_);
  or g_41747_(_14669_, _14677_, _14679_);
  and g_41748_(out[64], _14572_, _14680_);
  or g_41749_(_20465_, _14573_, _14681_);
  and g_41750_(_14584_, _14681_, _14682_);
  or g_41751_(_14583_, _14680_, _14683_);
  and g_41752_(_14557_, _14682_, _14684_);
  or g_41753_(_14558_, _14683_, _14686_);
  and g_41754_(_14579_, _14684_, _14687_);
  or g_41755_(_14580_, _14686_, _14688_);
  and g_41756_(_14533_, _14687_, _14689_);
  or g_41757_(_14534_, _14688_, _14690_);
  and g_41758_(_14657_, _14689_, _14691_);
  or g_41759_(_14658_, _14690_, _14692_);
  and g_41760_(_14679_, _14692_, _14693_);
  or g_41761_(_14678_, _14691_, _14694_);
  and g_41762_(_13887_, _14693_, _14695_);
  or g_41763_(_13888_, _14694_, _14697_);
  and g_41764_(_14505_, _14694_, _14698_);
  or g_41765_(_14504_, _14693_, _14699_);
  and g_41766_(_14697_, _14699_, _14700_);
  or g_41767_(_14695_, _14698_, _14701_);
  and g_41768_(_13876_, _14701_, _14702_);
  or g_41769_(_13875_, _14700_, _14703_);
  and g_41770_(_14513_, _14693_, _14704_);
  or g_41771_(_14514_, _14694_, _14705_);
  and g_41772_(_14519_, _14694_, _14706_);
  or g_41773_(_14521_, _14693_, _14708_);
  and g_41774_(_14705_, _14708_, _14709_);
  or g_41775_(_14704_, _14706_, _14710_);
  and g_41776_(_13872_, _14709_, _14711_);
  or g_41777_(_13873_, _14710_, _14712_);
  and g_41778_(_14703_, _14712_, _14713_);
  or g_41779_(_14702_, _14711_, _14714_);
  and g_41780_(out[64], _14693_, _14715_);
  or g_41781_(_20465_, _14694_, _14716_);
  and g_41782_(_14573_, _14694_, _14717_);
  or g_41783_(_14572_, _14693_, _14719_);
  and g_41784_(_14716_, _14719_, _14720_);
  or g_41785_(_14715_, _14717_, _14721_);
  and g_41786_(out[80], _14720_, _14722_);
  or g_41787_(_20597_, _14721_, _14723_);
  and g_41788_(_14560_, _14693_, _14724_);
  or g_41789_(_14559_, _14694_, _14725_);
  and g_41790_(_14563_, _14694_, _14726_);
  or g_41791_(_14565_, _14693_, _14727_);
  and g_41792_(_14725_, _14727_, _14728_);
  or g_41793_(_14724_, _14726_, _14730_);
  and g_41794_(out[81], _14728_, _14731_);
  or g_41795_(_20586_, _14730_, _14732_);
  xor g_41796_(out[81], out[80], _14733_);
  xor g_41797_(_20586_, out[80], _14734_);
  and g_41798_(_14722_, _14732_, _14735_);
  or g_41799_(_14723_, _14731_, _14736_);
  xor g_41800_(out[82], _13863_, _14737_);
  xor g_41801_(_20608_, _13863_, _14738_);
  and g_41802_(_14536_, _14693_, _14739_);
  or g_41803_(_14535_, _14694_, _14741_);
  and g_41804_(_14541_, _14694_, _14742_);
  or g_41805_(_14543_, _14693_, _14743_);
  and g_41806_(_14741_, _14743_, _14744_);
  or g_41807_(_14739_, _14742_, _14745_);
  and g_41808_(_14737_, _14745_, _14746_);
  or g_41809_(_14738_, _14744_, _14747_);
  and g_41810_(_14730_, _14733_, _14748_);
  or g_41811_(_14728_, _14734_, _14749_);
  and g_41812_(_14747_, _14749_, _14750_);
  or g_41813_(_14746_, _14748_, _14752_);
  and g_41814_(_14736_, _14750_, _14753_);
  or g_41815_(_14735_, _14752_, _14754_);
  xor g_41816_(out[83], _13864_, _14755_);
  xor g_41817_(_20619_, _13864_, _14756_);
  and g_41818_(_14546_, _14693_, _14757_);
  or g_41819_(_14547_, _14694_, _14758_);
  and g_41820_(_14552_, _14694_, _14759_);
  or g_41821_(_14554_, _14693_, _14760_);
  and g_41822_(_14758_, _14760_, _14761_);
  or g_41823_(_14757_, _14759_, _14763_);
  and g_41824_(_14755_, _14761_, _14764_);
  or g_41825_(_14756_, _14763_, _14765_);
  and g_41826_(_14738_, _14744_, _14766_);
  or g_41827_(_14737_, _14745_, _14767_);
  and g_41828_(_14765_, _14767_, _14768_);
  or g_41829_(_14764_, _14766_, _14769_);
  and g_41830_(_14754_, _14768_, _14770_);
  or g_41831_(_14753_, _14769_, _14771_);
  xor g_41832_(out[84], _13865_, _14772_);
  xor g_41833_(_20575_, _13865_, _14774_);
  and g_41834_(_14631_, _14693_, _14775_);
  or g_41835_(_14632_, _14694_, _14776_);
  and g_41836_(_14637_, _14694_, _14777_);
  or g_41837_(_14638_, _14693_, _14778_);
  and g_41838_(_14776_, _14778_, _14779_);
  or g_41839_(_14775_, _14777_, _14780_);
  and g_41840_(_14774_, _14780_, _14781_);
  or g_41841_(_14772_, _14779_, _14782_);
  and g_41842_(_14756_, _14763_, _14783_);
  or g_41843_(_14755_, _14761_, _14785_);
  and g_41844_(_14782_, _14785_, _14786_);
  or g_41845_(_14781_, _14783_, _14787_);
  and g_41846_(_14771_, _14786_, _14788_);
  or g_41847_(_14770_, _14787_, _14789_);
  xor g_41848_(out[85], _13866_, _14790_);
  xor g_41849_(_20564_, _13866_, _14791_);
  and g_41850_(_14620_, _14693_, _14792_);
  or g_41851_(_14621_, _14694_, _14793_);
  and g_41852_(_14626_, _14694_, _14794_);
  or g_41853_(_14627_, _14693_, _14796_);
  and g_41854_(_14793_, _14796_, _14797_);
  or g_41855_(_14792_, _14794_, _14798_);
  and g_41856_(_14790_, _14797_, _14799_);
  or g_41857_(_14791_, _14798_, _14800_);
  and g_41858_(_14772_, _14779_, _14801_);
  or g_41859_(_14774_, _14780_, _14802_);
  and g_41860_(_14800_, _14802_, _14803_);
  or g_41861_(_14799_, _14801_, _14804_);
  and g_41862_(_14789_, _14803_, _14805_);
  or g_41863_(_14788_, _14804_, _14807_);
  xor g_41864_(out[86], _13867_, _14808_);
  xor g_41865_(_20553_, _13867_, _14809_);
  and g_41866_(_14601_, _14693_, _14810_);
  or g_41867_(_14600_, _14694_, _14811_);
  and g_41868_(_14606_, _14694_, _14812_);
  or g_41869_(_14607_, _14693_, _14813_);
  and g_41870_(_14811_, _14813_, _14814_);
  or g_41871_(_14810_, _14812_, _14815_);
  and g_41872_(_14808_, _14815_, _14816_);
  or g_41873_(_14809_, _14814_, _14818_);
  and g_41874_(_14791_, _14798_, _14819_);
  or g_41875_(_14790_, _14797_, _14820_);
  and g_41876_(_14818_, _14820_, _14821_);
  or g_41877_(_14816_, _14819_, _14822_);
  and g_41878_(_14807_, _14821_, _14823_);
  or g_41879_(_14805_, _14822_, _14824_);
  xor g_41880_(out[87], _13868_, _14825_);
  xor g_41881_(_20542_, _13868_, _14826_);
  and g_41882_(_14591_, _14693_, _14827_);
  or g_41883_(_14590_, _14694_, _14829_);
  and g_41884_(_14598_, _14694_, _14830_);
  or g_41885_(_14596_, _14693_, _14831_);
  and g_41886_(_14829_, _14831_, _14832_);
  or g_41887_(_14827_, _14830_, _14833_);
  and g_41888_(_14825_, _14833_, _14834_);
  or g_41889_(_14826_, _14832_, _14835_);
  and g_41890_(_14809_, _14814_, _14836_);
  or g_41891_(_14808_, _14815_, _14837_);
  and g_41892_(_14835_, _14837_, _14838_);
  or g_41893_(_14834_, _14836_, _14840_);
  and g_41894_(_14824_, _14838_, _14841_);
  or g_41895_(_14823_, _14840_, _14842_);
  and g_41896_(_14826_, _14832_, _14843_);
  or g_41897_(_14825_, _14833_, _14844_);
  and g_41898_(_13873_, _14710_, _14845_);
  or g_41899_(_13872_, _14709_, _14846_);
  and g_41900_(_14844_, _14846_, _14847_);
  or g_41901_(_14843_, _14845_, _14848_);
  and g_41902_(out[90], _13874_, _14849_);
  xor g_41903_(out[90], _13874_, _14851_);
  not g_41904_(_14851_, _14852_);
  and g_41905_(_14480_, _14693_, _14853_);
  or g_41906_(_14481_, _14694_, _14854_);
  and g_41907_(_14486_, _14694_, _14855_);
  or g_41908_(_14488_, _14693_, _14856_);
  and g_41909_(_14854_, _14856_, _14857_);
  or g_41910_(_14853_, _14855_, _14858_);
  and g_41911_(_14851_, _14857_, _14859_);
  or g_41912_(_14852_, _14858_, _14860_);
  and g_41913_(_14477_, _14693_, _14862_);
  or g_41914_(_14475_, _14694_, _14863_);
  and g_41915_(_14473_, _14694_, _14864_);
  or g_41916_(_14472_, _14693_, _14865_);
  and g_41917_(_14863_, _14865_, _14866_);
  or g_41918_(_14862_, _14864_, _14867_);
  xor g_41919_(out[91], _14849_, _14868_);
  xor g_41920_(_20531_, _14849_, _14869_);
  and g_41921_(_14867_, _14868_, _14870_);
  or g_41922_(_14866_, _14869_, _14871_);
  and g_41923_(_14866_, _14869_, _14873_);
  or g_41924_(_14867_, _14868_, _14874_);
  and g_41925_(_13875_, _14700_, _14875_);
  or g_41926_(_13876_, _14701_, _14876_);
  xor g_41927_(_14851_, _14857_, _14877_);
  xor g_41928_(_14852_, _14857_, _14878_);
  and g_41929_(_14871_, _14874_, _14879_);
  or g_41930_(_14870_, _14873_, _14880_);
  and g_41931_(_14877_, _14879_, _14881_);
  or g_41932_(_14878_, _14880_, _14882_);
  and g_41933_(_14714_, _14876_, _14884_);
  or g_41934_(_14713_, _14875_, _14885_);
  and g_41935_(_14713_, _14876_, _14886_);
  or g_41936_(_14714_, _14875_, _14887_);
  and g_41937_(_14847_, _14886_, _14888_);
  or g_41938_(_14848_, _14887_, _14889_);
  and g_41939_(_14881_, _14888_, _14890_);
  or g_41940_(_14882_, _14889_, _14891_);
  and g_41941_(_14842_, _14890_, _14892_);
  or g_41942_(_14841_, _14891_, _14893_);
  and g_41943_(_14859_, _14874_, _14895_);
  or g_41944_(_14860_, _14873_, _14896_);
  and g_41945_(_14881_, _14884_, _14897_);
  or g_41946_(_14882_, _14885_, _14898_);
  and g_41947_(_14871_, _14898_, _14899_);
  or g_41948_(_14870_, _14897_, _14900_);
  and g_41949_(_14896_, _14899_, _14901_);
  or g_41950_(_14895_, _14900_, _14902_);
  and g_41951_(_14893_, _14901_, _14903_);
  or g_41952_(_14892_, _14902_, _14904_);
  and g_41953_(_13872_, _14903_, _14906_);
  or g_41954_(_13873_, _14904_, _14907_);
  and g_41955_(_14710_, _14904_, _14908_);
  or g_41956_(_14709_, _14903_, _14909_);
  and g_41957_(_14907_, _14909_, _14910_);
  or g_41958_(_14906_, _14908_, _14911_);
  and g_41959_(_13862_, _14911_, _14912_);
  or g_41960_(_13861_, _14910_, _14913_);
  or g_41961_(out[105], _13859_, _14914_);
  xor g_41962_(out[105], _13859_, _14915_);
  xor g_41963_(_20773_, _13859_, _14917_);
  and g_41964_(_13876_, _14903_, _14918_);
  or g_41965_(_13875_, _14904_, _14919_);
  and g_41966_(_14700_, _14904_, _14920_);
  or g_41967_(_14701_, _14903_, _14921_);
  and g_41968_(_14919_, _14921_, _14922_);
  or g_41969_(_14918_, _14920_, _14923_);
  and g_41970_(_14915_, _14923_, _14924_);
  or g_41971_(_14917_, _14922_, _14925_);
  and g_41972_(_14913_, _14925_, _14926_);
  or g_41973_(_14912_, _14924_, _14928_);
  and g_41974_(_14866_, _14868_, _14929_);
  or g_41975_(_14867_, _14869_, _14930_);
  and g_41976_(out[106], _14914_, _14931_);
  xor g_41977_(out[107], _14931_, _14932_);
  xor g_41978_(_20663_, _14931_, _14933_);
  and g_41979_(_14930_, _14932_, _14934_);
  or g_41980_(_14929_, _14933_, _14935_);
  and g_41981_(_13861_, _14910_, _14936_);
  or g_41982_(_13862_, _14911_, _14937_);
  and g_41983_(_14935_, _14937_, _14939_);
  or g_41984_(_14934_, _14936_, _14940_);
  and g_41985_(_14926_, _14939_, _14941_);
  or g_41986_(_14928_, _14940_, _14942_);
  xor g_41987_(out[106], _14914_, _14943_);
  xor g_41988_(_20784_, _14914_, _14944_);
  and g_41989_(_14852_, _14903_, _14945_);
  or g_41990_(_14851_, _14904_, _14946_);
  and g_41991_(_14857_, _14904_, _14947_);
  or g_41992_(_14858_, _14903_, _14948_);
  and g_41993_(_14946_, _14948_, _14950_);
  or g_41994_(_14945_, _14947_, _14951_);
  and g_41995_(_14944_, _14950_, _14952_);
  or g_41996_(_14943_, _14951_, _14953_);
  and g_41997_(_14929_, _14933_, _14954_);
  or g_41998_(_14930_, _14932_, _14955_);
  and g_41999_(_14953_, _14955_, _14956_);
  or g_42000_(_14952_, _14954_, _14957_);
  and g_42001_(_14943_, _14951_, _14958_);
  or g_42002_(_14944_, _14950_, _14959_);
  and g_42003_(_14917_, _14922_, _14961_);
  or g_42004_(_14915_, _14923_, _14962_);
  and g_42005_(_14959_, _14962_, _14963_);
  or g_42006_(_14958_, _14961_, _14964_);
  and g_42007_(_14956_, _14963_, _14965_);
  or g_42008_(_14957_, _14964_, _14966_);
  and g_42009_(_14941_, _14965_, _14967_);
  or g_42010_(_14942_, _14966_, _14968_);
  and g_42011_(_14825_, _14903_, _14969_);
  or g_42012_(_14826_, _14904_, _14970_);
  and g_42013_(_14832_, _14904_, _14972_);
  or g_42014_(_14833_, _14903_, _14973_);
  and g_42015_(_14970_, _14973_, _14974_);
  or g_42016_(_14969_, _14972_, _14975_);
  and g_42017_(_13857_, _14974_, _14976_);
  or g_42018_(_13858_, _14975_, _14977_);
  xor g_42019_(out[102], _13854_, _14978_);
  xor g_42020_(_20685_, _13854_, _14979_);
  and g_42021_(_14808_, _14903_, _14980_);
  or g_42022_(_14809_, _14904_, _14981_);
  and g_42023_(_14814_, _14904_, _14983_);
  or g_42024_(_14815_, _14903_, _14984_);
  and g_42025_(_14981_, _14984_, _14985_);
  or g_42026_(_14980_, _14983_, _14986_);
  and g_42027_(_14979_, _14986_, _14987_);
  or g_42028_(_14978_, _14985_, _14988_);
  and g_42029_(_14977_, _14988_, _14989_);
  or g_42030_(_14976_, _14987_, _14990_);
  xor g_42031_(out[101], _13853_, _14991_);
  xor g_42032_(_20696_, _13853_, _14992_);
  and g_42033_(_14798_, _14904_, _14994_);
  or g_42034_(_14797_, _14903_, _14995_);
  and g_42035_(_14790_, _14903_, _14996_);
  or g_42036_(_14791_, _14904_, _14997_);
  and g_42037_(_14995_, _14997_, _14998_);
  or g_42038_(_14994_, _14996_, _14999_);
  and g_42039_(_14991_, _14998_, _15000_);
  or g_42040_(_14992_, _14999_, _15001_);
  and g_42041_(_14989_, _15001_, _15002_);
  or g_42042_(_14990_, _15000_, _15003_);
  and g_42043_(_14978_, _14985_, _15005_);
  or g_42044_(_14979_, _14986_, _15006_);
  and g_42045_(_13858_, _14975_, _15007_);
  or g_42046_(_13857_, _14974_, _15008_);
  and g_42047_(_15006_, _15008_, _15009_);
  or g_42048_(_15005_, _15007_, _15010_);
  xor g_42049_(out[100], _13852_, _15011_);
  xor g_42050_(_20707_, _13852_, _15012_);
  and g_42051_(_14772_, _14903_, _15013_);
  or g_42052_(_14774_, _14904_, _15014_);
  and g_42053_(_14780_, _14904_, _15016_);
  or g_42054_(_14779_, _14903_, _15017_);
  and g_42055_(_15014_, _15017_, _15018_);
  or g_42056_(_15013_, _15016_, _15019_);
  and g_42057_(_15011_, _15018_, _15020_);
  or g_42058_(_15012_, _15019_, _15021_);
  and g_42059_(_14992_, _14999_, _15022_);
  or g_42060_(_14991_, _14998_, _15023_);
  and g_42061_(_15012_, _15019_, _15024_);
  or g_42062_(_15011_, _15018_, _15025_);
  and g_42063_(_15023_, _15025_, _15027_);
  or g_42064_(_15022_, _15024_, _15028_);
  and g_42065_(_15021_, _15027_, _15029_);
  or g_42066_(_15020_, _15028_, _15030_);
  and g_42067_(_14989_, _15009_, _15031_);
  or g_42068_(_14990_, _15010_, _15032_);
  and g_42069_(_15001_, _15029_, _15033_);
  or g_42070_(_15000_, _15030_, _15034_);
  and g_42071_(_14967_, _15033_, _15035_);
  or g_42072_(_14968_, _15034_, _15036_);
  and g_42073_(_15031_, _15035_, _15038_);
  or g_42074_(_15032_, _15036_, _15039_);
  xor g_42075_(out[98], _13850_, _15040_);
  not g_42076_(_15040_, _15041_);
  and g_42077_(_14737_, _14903_, _15042_);
  or g_42078_(_14738_, _14904_, _15043_);
  and g_42079_(_14744_, _14904_, _15044_);
  or g_42080_(_14745_, _14903_, _15045_);
  and g_42081_(_15043_, _15045_, _15046_);
  or g_42082_(_15042_, _15044_, _15047_);
  and g_42083_(_15040_, _15046_, _15049_);
  or g_42084_(_15041_, _15047_, _15050_);
  xor g_42085_(out[99], _13851_, _15051_);
  xor g_42086_(_20751_, _13851_, _15052_);
  and g_42087_(_14763_, _14904_, _15053_);
  or g_42088_(_14761_, _14903_, _15054_);
  and g_42089_(_14755_, _14903_, _15055_);
  or g_42090_(_14756_, _14904_, _15056_);
  and g_42091_(_15054_, _15056_, _15057_);
  or g_42092_(_15053_, _15055_, _15058_);
  and g_42093_(_15052_, _15058_, _15060_);
  or g_42094_(_15051_, _15057_, _15061_);
  and g_42095_(_15050_, _15061_, _15062_);
  or g_42096_(_15049_, _15060_, _15063_);
  and g_42097_(_15051_, _15057_, _15064_);
  or g_42098_(_15052_, _15058_, _15065_);
  and g_42099_(_15041_, _15047_, _15066_);
  or g_42100_(_15040_, _15046_, _15067_);
  and g_42101_(_15065_, _15067_, _15068_);
  or g_42102_(_15064_, _15066_, _15069_);
  and g_42103_(_15062_, _15068_, _15071_);
  or g_42104_(_15063_, _15069_, _15072_);
  xor g_42105_(out[97], out[96], _15073_);
  not g_42106_(_15073_, _15074_);
  and g_42107_(_14733_, _14903_, _15075_);
  or g_42108_(_14734_, _14904_, _15076_);
  and g_42109_(_14728_, _14904_, _15077_);
  or g_42110_(_14730_, _14903_, _15078_);
  and g_42111_(_15076_, _15078_, _15079_);
  or g_42112_(_15075_, _15077_, _15080_);
  and g_42113_(_15073_, _15079_, _15082_);
  or g_42114_(_15074_, _15080_, _15083_);
  and g_42115_(_14721_, _14904_, _15084_);
  or g_42116_(_14720_, _14903_, _15085_);
  and g_42117_(out[80], _14903_, _15086_);
  or g_42118_(_20597_, _14904_, _15087_);
  and g_42119_(_15085_, _15087_, _15088_);
  or g_42120_(_15084_, _15086_, _15089_);
  and g_42121_(_20729_, _15089_, _15090_);
  or g_42122_(out[96], _15088_, _15091_);
  xor g_42123_(_15073_, _15079_, _15093_);
  xor g_42124_(_15074_, _15079_, _15094_);
  and g_42125_(_15091_, _15093_, _15095_);
  or g_42126_(_15090_, _15094_, _15096_);
  and g_42127_(_15083_, _15096_, _15097_);
  or g_42128_(_15082_, _15095_, _15098_);
  and g_42129_(_15071_, _15098_, _15099_);
  or g_42130_(_15072_, _15097_, _15100_);
  and g_42131_(_15063_, _15065_, _15101_);
  or g_42132_(_15062_, _15064_, _15102_);
  and g_42133_(_15100_, _15102_, _15104_);
  or g_42134_(_15099_, _15101_, _15105_);
  and g_42135_(_15038_, _15105_, _15106_);
  or g_42136_(_15039_, _15104_, _15107_);
  and g_42137_(_14977_, _15010_, _15108_);
  or g_42138_(_14976_, _15009_, _15109_);
  and g_42139_(_15002_, _15028_, _15110_);
  or g_42140_(_15003_, _15027_, _15111_);
  and g_42141_(_15109_, _15111_, _15112_);
  or g_42142_(_15108_, _15110_, _15113_);
  and g_42143_(_14967_, _15113_, _15115_);
  or g_42144_(_14968_, _15112_, _15116_);
  and g_42145_(_14928_, _14963_, _15117_);
  or g_42146_(_14926_, _14964_, _15118_);
  and g_42147_(_14956_, _15118_, _15119_);
  or g_42148_(_14957_, _15117_, _15120_);
  and g_42149_(_14935_, _15120_, _15121_);
  or g_42150_(_14934_, _15119_, _15122_);
  and g_42151_(_15116_, _15122_, _15123_);
  or g_42152_(_15115_, _15121_, _15124_);
  and g_42153_(_15107_, _15123_, _15126_);
  or g_42154_(_15106_, _15124_, _15127_);
  and g_42155_(out[96], _15088_, _15128_);
  or g_42156_(_20729_, _15089_, _15129_);
  and g_42157_(_15071_, _15129_, _15130_);
  or g_42158_(_15072_, _15128_, _15131_);
  and g_42159_(_15095_, _15130_, _15132_);
  or g_42160_(_15096_, _15131_, _15133_);
  and g_42161_(_15038_, _15132_, _15134_);
  or g_42162_(_15039_, _15133_, _15135_);
  and g_42163_(_15127_, _15135_, _15137_);
  or g_42164_(_15126_, _15134_, _15138_);
  and g_42165_(_13857_, _15137_, _15139_);
  or g_42166_(_13858_, _15138_, _15140_);
  and g_42167_(_14975_, _15138_, _15141_);
  or g_42168_(_14974_, _15137_, _15142_);
  and g_42169_(_15140_, _15142_, _15143_);
  or g_42170_(_15139_, _15141_, _15144_);
  and g_42171_(_14929_, _14932_, _15145_);
  or g_42172_(_14930_, _14933_, _15146_);
  or g_42173_(out[112], out[113], _15148_);
  or g_42174_(out[112], _17987_, _15149_);
  and g_42175_(out[115], _15149_, _15150_);
  and g_42176_(_25705_, _15149_, _15151_);
  and g_42177_(out[117], _15151_, _15152_);
  or g_42178_(out[118], _15152_, _15153_);
  and g_42179_(out[119], _15153_, _15154_);
  and g_42180_(out[120], _15154_, _15155_);
  or g_42181_(out[121], _15155_, _15156_);
  and g_42182_(out[122], _15156_, _15157_);
  xor g_42183_(out[123], _15157_, _15159_);
  xor g_42184_(_20795_, _15157_, _15160_);
  and g_42185_(_15145_, _15160_, _15161_);
  or g_42186_(_15146_, _15159_, _15162_);
  and g_42187_(_15146_, _15159_, _15163_);
  or g_42188_(_15145_, _15160_, _15164_);
  xor g_42189_(out[122], _15156_, _15165_);
  not g_42190_(_15165_, _15166_);
  and g_42191_(_14944_, _15137_, _15167_);
  or g_42192_(_14943_, _15138_, _15168_);
  and g_42193_(_14951_, _15138_, _15170_);
  or g_42194_(_14950_, _15137_, _15171_);
  and g_42195_(_15168_, _15171_, _15172_);
  or g_42196_(_15167_, _15170_, _15173_);
  and g_42197_(_15165_, _15173_, _15174_);
  or g_42198_(_15166_, _15172_, _15175_);
  and g_42199_(_15164_, _15175_, _15176_);
  or g_42200_(_15163_, _15174_, _15177_);
  and g_42201_(_15166_, _15172_, _15178_);
  or g_42202_(_15165_, _15173_, _15179_);
  xor g_42203_(out[121], _15155_, _15181_);
  not g_42204_(_15181_, _15182_);
  and g_42205_(_14915_, _15137_, _15183_);
  or g_42206_(_14917_, _15138_, _15184_);
  and g_42207_(_14922_, _15138_, _15185_);
  or g_42208_(_14923_, _15137_, _15186_);
  and g_42209_(_15184_, _15186_, _15187_);
  or g_42210_(_15183_, _15185_, _15188_);
  and g_42211_(_15182_, _15188_, _15189_);
  or g_42212_(_15181_, _15187_, _15190_);
  and g_42213_(_15181_, _15187_, _15192_);
  or g_42214_(_15182_, _15188_, _15193_);
  xor g_42215_(out[120], _15154_, _15194_);
  not g_42216_(_15194_, _15195_);
  and g_42217_(_13861_, _15137_, _15196_);
  or g_42218_(_13862_, _15138_, _15197_);
  and g_42219_(_14911_, _15138_, _15198_);
  or g_42220_(_14910_, _15137_, _15199_);
  and g_42221_(_15197_, _15199_, _15200_);
  or g_42222_(_15196_, _15198_, _15201_);
  and g_42223_(_15194_, _15200_, _15203_);
  or g_42224_(_15195_, _15201_, _15204_);
  and g_42225_(_15193_, _15203_, _15205_);
  or g_42226_(_15192_, _15204_, _15206_);
  and g_42227_(_15190_, _15206_, _15207_);
  or g_42228_(_15189_, _15205_, _15208_);
  and g_42229_(out[96], _15137_, _15209_);
  or g_42230_(_20729_, _15138_, _15210_);
  and g_42231_(_15089_, _15138_, _15211_);
  or g_42232_(_15088_, _15137_, _15212_);
  and g_42233_(_15210_, _15212_, _15214_);
  or g_42234_(_15209_, _15211_, _15215_);
  and g_42235_(out[112], _15214_, _15216_);
  or g_42236_(_19860_, _15215_, _15217_);
  and g_42237_(_15073_, _15137_, _15218_);
  or g_42238_(_15074_, _15138_, _15219_);
  and g_42239_(_15080_, _15138_, _15220_);
  or g_42240_(_15079_, _15137_, _15221_);
  and g_42241_(_15219_, _15221_, _15222_);
  or g_42242_(_15218_, _15220_, _15223_);
  and g_42243_(out[113], _15223_, _15225_);
  or g_42244_(_20850_, _15222_, _15226_);
  xor g_42245_(out[112], out[113], _15227_);
  xor g_42246_(_19860_, out[113], _15228_);
  and g_42247_(_15216_, _15226_, _15229_);
  or g_42248_(_15217_, _15225_, _15230_);
  xor g_42249_(out[114], _15148_, _15231_);
  xor g_42250_(_20861_, _15148_, _15232_);
  and g_42251_(_15040_, _15137_, _15233_);
  or g_42252_(_15041_, _15138_, _15234_);
  and g_42253_(_15047_, _15138_, _15236_);
  or g_42254_(_15046_, _15137_, _15237_);
  and g_42255_(_15234_, _15237_, _15238_);
  or g_42256_(_15233_, _15236_, _15239_);
  and g_42257_(_15231_, _15238_, _15240_);
  or g_42258_(_15232_, _15239_, _15241_);
  and g_42259_(_15222_, _15227_, _15242_);
  or g_42260_(_15223_, _15228_, _15243_);
  and g_42261_(_15241_, _15243_, _15244_);
  or g_42262_(_15240_, _15242_, _15245_);
  and g_42263_(_15230_, _15244_, _15247_);
  or g_42264_(_15229_, _15245_, _15248_);
  xor g_42265_(out[115], _15149_, _15249_);
  xor g_42266_(_20872_, _15149_, _15250_);
  and g_42267_(_15051_, _15137_, _15251_);
  or g_42268_(_15052_, _15138_, _15252_);
  and g_42269_(_15058_, _15138_, _15253_);
  or g_42270_(_15057_, _15137_, _15254_);
  and g_42271_(_15252_, _15254_, _15255_);
  or g_42272_(_15251_, _15253_, _15256_);
  and g_42273_(_15249_, _15255_, _15258_);
  or g_42274_(_15250_, _15256_, _15259_);
  and g_42275_(_15232_, _15239_, _15260_);
  or g_42276_(_15231_, _15238_, _15261_);
  and g_42277_(_15259_, _15261_, _15262_);
  or g_42278_(_15258_, _15260_, _15263_);
  and g_42279_(_15248_, _15262_, _15264_);
  or g_42280_(_15247_, _15263_, _15265_);
  xor g_42281_(out[116], _15150_, _15266_);
  xor g_42282_(_20839_, _15150_, _15267_);
  and g_42283_(_15011_, _15137_, _15269_);
  and g_42284_(_15019_, _15138_, _15270_);
  or g_42285_(_15269_, _15270_, _15271_);
  not g_42286_(_15271_, _15272_);
  and g_42287_(_15267_, _15271_, _15273_);
  or g_42288_(_15266_, _15272_, _15274_);
  and g_42289_(_15250_, _15256_, _15275_);
  or g_42290_(_15249_, _15255_, _15276_);
  and g_42291_(_15274_, _15276_, _15277_);
  or g_42292_(_15273_, _15275_, _15278_);
  and g_42293_(_15265_, _15277_, _15280_);
  or g_42294_(_15264_, _15278_, _15281_);
  xor g_42295_(out[117], _15151_, _15282_);
  xor g_42296_(_20828_, _15151_, _15283_);
  and g_42297_(_14999_, _15138_, _15284_);
  and g_42298_(_14991_, _15137_, _15285_);
  or g_42299_(_15284_, _15285_, _15286_);
  not g_42300_(_15286_, _15287_);
  or g_42301_(_15283_, _15286_, _15288_);
  or g_42302_(_15267_, _15271_, _15289_);
  and g_42303_(_15288_, _15289_, _15291_);
  not g_42304_(_15291_, _15292_);
  and g_42305_(_15281_, _15291_, _15293_);
  or g_42306_(_15280_, _15292_, _15294_);
  xor g_42307_(out[118], _15152_, _15295_);
  xor g_42308_(_20817_, _15152_, _15296_);
  and g_42309_(_14978_, _15137_, _15297_);
  or g_42310_(_14979_, _15138_, _15298_);
  and g_42311_(_14986_, _15138_, _15299_);
  or g_42312_(_14985_, _15137_, _15300_);
  and g_42313_(_15298_, _15300_, _15302_);
  or g_42314_(_15297_, _15299_, _15303_);
  and g_42315_(_15295_, _15302_, _15304_);
  or g_42316_(_15296_, _15303_, _15305_);
  and g_42317_(_15283_, _15286_, _15306_);
  or g_42318_(_15282_, _15287_, _15307_);
  and g_42319_(_15305_, _15307_, _15308_);
  or g_42320_(_15304_, _15306_, _15309_);
  and g_42321_(_15294_, _15308_, _15310_);
  or g_42322_(_15293_, _15309_, _15311_);
  xor g_42323_(out[119], _15153_, _15313_);
  xor g_42324_(_20806_, _15153_, _15314_);
  and g_42325_(_15143_, _15313_, _15315_);
  or g_42326_(_15144_, _15314_, _15316_);
  and g_42327_(_15296_, _15303_, _15317_);
  or g_42328_(_15295_, _15302_, _15318_);
  and g_42329_(_15316_, _15318_, _15319_);
  or g_42330_(_15315_, _15317_, _15320_);
  and g_42331_(_15311_, _15319_, _15321_);
  or g_42332_(_15310_, _15320_, _15322_);
  and g_42333_(_15195_, _15201_, _15324_);
  or g_42334_(_15194_, _15200_, _15325_);
  and g_42335_(_15144_, _15314_, _15326_);
  or g_42336_(_15143_, _15313_, _15327_);
  and g_42337_(_15193_, _15325_, _15328_);
  or g_42338_(_15192_, _15324_, _15329_);
  and g_42339_(_15204_, _15327_, _15330_);
  or g_42340_(_15203_, _15326_, _15331_);
  and g_42341_(_15190_, _15330_, _15332_);
  or g_42342_(_15189_, _15331_, _15333_);
  and g_42343_(_15328_, _15332_, _15335_);
  or g_42344_(_15329_, _15333_, _15336_);
  and g_42345_(_15162_, _15179_, _15337_);
  or g_42346_(_15161_, _15178_, _15338_);
  and g_42347_(_15176_, _15337_, _15339_);
  or g_42348_(_15177_, _15338_, _15340_);
  and g_42349_(_15335_, _15339_, _15341_);
  or g_42350_(_15336_, _15340_, _15342_);
  and g_42351_(_15322_, _15341_, _15343_);
  or g_42352_(_15321_, _15342_, _15344_);
  and g_42353_(_15162_, _15174_, _15346_);
  or g_42354_(_15161_, _15175_, _15347_);
  and g_42355_(_15208_, _15339_, _15348_);
  or g_42356_(_15207_, _15340_, _15349_);
  and g_42357_(_15347_, _15349_, _15350_);
  or g_42358_(_15346_, _15348_, _15351_);
  and g_42359_(_15164_, _15350_, _15352_);
  or g_42360_(_15163_, _15351_, _15353_);
  or g_42361_(_15343_, _15353_, _15354_);
  and g_42362_(_15344_, _15352_, _15355_);
  and g_42363_(_15144_, _15354_, _15357_);
  or g_42364_(_15143_, _15355_, _15358_);
  and g_42365_(_15313_, _15355_, _15359_);
  or g_42366_(_15314_, _15354_, _15360_);
  and g_42367_(_15358_, _15360_, _15361_);
  or g_42368_(_15357_, _15359_, _15362_);
  or g_42369_(out[129], out[128], _15363_);
  or g_42370_(out[128], _18126_, _15364_);
  and g_42371_(out[131], _15364_, _15365_);
  and g_42372_(_25856_, _15364_, _15366_);
  and g_42373_(out[133], _15366_, _15368_);
  or g_42374_(out[134], _15368_, _15369_);
  and g_42375_(out[135], _15369_, _15370_);
  and g_42376_(out[136], _15370_, _15371_);
  or g_42377_(out[137], _15371_, _15372_);
  and g_42378_(out[138], _15372_, _15373_);
  xor g_42379_(out[138], _15372_, _15374_);
  xor g_42380_(_21037_, _15372_, _15375_);
  and g_42381_(_15173_, _15354_, _15376_);
  and g_42382_(_15166_, _15355_, _15377_);
  or g_42383_(_15376_, _15377_, _15379_);
  not g_42384_(_15379_, _15380_);
  and g_42385_(_15375_, _15380_, _15381_);
  or g_42386_(_15374_, _15379_, _15382_);
  and g_42387_(_15145_, _15159_, _15383_);
  or g_42388_(_15146_, _15160_, _15384_);
  xor g_42389_(out[139], _15373_, _15385_);
  xor g_42390_(_20916_, _15373_, _15386_);
  and g_42391_(_15383_, _15386_, _15387_);
  or g_42392_(_15384_, _15385_, _15388_);
  and g_42393_(_15382_, _15388_, _15390_);
  or g_42394_(_15381_, _15387_, _15391_);
  and g_42395_(_15374_, _15379_, _15392_);
  or g_42396_(_15375_, _15380_, _15393_);
  and g_42397_(_15384_, _15385_, _15394_);
  or g_42398_(_15383_, _15386_, _15395_);
  and g_42399_(_15393_, _15395_, _15396_);
  or g_42400_(_15392_, _15394_, _15397_);
  and g_42401_(_15390_, _15396_, _15398_);
  or g_42402_(_15391_, _15397_, _15399_);
  xor g_42403_(out[137], _15371_, _15401_);
  xor g_42404_(_21026_, _15371_, _15402_);
  and g_42405_(_15187_, _15354_, _15403_);
  not g_42406_(_15403_, _15404_);
  or g_42407_(_15181_, _15354_, _15405_);
  not g_42408_(_15405_, _15406_);
  and g_42409_(_15404_, _15405_, _15407_);
  or g_42410_(_15403_, _15406_, _15408_);
  and g_42411_(_15401_, _15408_, _15409_);
  or g_42412_(_15402_, _15407_, _15410_);
  xor g_42413_(out[136], _15370_, _15412_);
  xor g_42414_(_21015_, _15370_, _15413_);
  and g_42415_(_15200_, _15354_, _15414_);
  and g_42416_(_15195_, _15355_, _15415_);
  or g_42417_(_15414_, _15415_, _15416_);
  not g_42418_(_15416_, _15417_);
  and g_42419_(_15413_, _15417_, _15418_);
  or g_42420_(_15412_, _15416_, _15419_);
  and g_42421_(_15410_, _15419_, _15420_);
  or g_42422_(_15409_, _15418_, _15421_);
  and g_42423_(_15412_, _15416_, _15423_);
  or g_42424_(_15413_, _15417_, _15424_);
  and g_42425_(_15402_, _15407_, _15425_);
  or g_42426_(_15401_, _15408_, _15426_);
  and g_42427_(_15424_, _15426_, _15427_);
  or g_42428_(_15423_, _15425_, _15428_);
  and g_42429_(_15420_, _15427_, _15429_);
  or g_42430_(_15421_, _15428_, _15430_);
  xor g_42431_(out[135], _15369_, _15431_);
  xor g_42432_(_20927_, _15369_, _15432_);
  and g_42433_(_15361_, _15431_, _15434_);
  or g_42434_(_15362_, _15432_, _15435_);
  xor g_42435_(out[134], _15368_, _15436_);
  xor g_42436_(_20938_, _15368_, _15437_);
  and g_42437_(_15303_, _15354_, _15438_);
  or g_42438_(_15302_, _15355_, _15439_);
  and g_42439_(_15295_, _15355_, _15440_);
  or g_42440_(_15296_, _15354_, _15441_);
  and g_42441_(_15439_, _15441_, _15442_);
  or g_42442_(_15438_, _15440_, _15443_);
  and g_42443_(_15436_, _15442_, _15445_);
  or g_42444_(_15437_, _15443_, _15446_);
  and g_42445_(_15362_, _15432_, _15447_);
  or g_42446_(_15361_, _15431_, _15448_);
  and g_42447_(_15446_, _15448_, _15449_);
  or g_42448_(_15445_, _15447_, _15450_);
  xor g_42449_(out[133], _15366_, _15451_);
  xor g_42450_(_20949_, _15366_, _15452_);
  and g_42451_(_15286_, _15354_, _15453_);
  not g_42452_(_15453_, _15454_);
  or g_42453_(_15283_, _15354_, _15456_);
  not g_42454_(_15456_, _15457_);
  and g_42455_(_15454_, _15456_, _15458_);
  or g_42456_(_15453_, _15457_, _15459_);
  and g_42457_(_15452_, _15459_, _15460_);
  or g_42458_(_15451_, _15458_, _15461_);
  xor g_42459_(out[132], _15365_, _15462_);
  xor g_42460_(_20960_, _15365_, _15463_);
  or g_42461_(_15267_, _15354_, _15464_);
  not g_42462_(_15464_, _15465_);
  and g_42463_(_15271_, _15354_, _15467_);
  not g_42464_(_15467_, _15468_);
  and g_42465_(_15464_, _15468_, _15469_);
  or g_42466_(_15465_, _15467_, _15470_);
  and g_42467_(_15463_, _15470_, _15471_);
  or g_42468_(_15462_, _15469_, _15472_);
  and g_42469_(_15461_, _15472_, _15473_);
  or g_42470_(_15460_, _15471_, _15474_);
  and g_42471_(_15451_, _15458_, _15475_);
  or g_42472_(_15452_, _15459_, _15476_);
  and g_42473_(_15437_, _15443_, _15478_);
  or g_42474_(_15436_, _15442_, _15479_);
  and g_42475_(_15476_, _15479_, _15480_);
  or g_42476_(_15475_, _15478_, _15481_);
  or g_42477_(_15473_, _15481_, _15482_);
  and g_42478_(_15449_, _15482_, _15483_);
  or g_42479_(_15434_, _15483_, _15484_);
  not g_42480_(_15484_, _15485_);
  and g_42481_(_15462_, _15469_, _15486_);
  or g_42482_(_15463_, _15470_, _15487_);
  and g_42483_(_15435_, _15487_, _15489_);
  or g_42484_(_15434_, _15486_, _15490_);
  and g_42485_(_15449_, _15489_, _15491_);
  or g_42486_(_15450_, _15490_, _15492_);
  and g_42487_(_15473_, _15480_, _15493_);
  or g_42488_(_15474_, _15481_, _15494_);
  and g_42489_(_15491_, _15493_, _15495_);
  or g_42490_(_15492_, _15494_, _15496_);
  xor g_42491_(out[130], _15363_, _15497_);
  not g_42492_(_15497_, _15498_);
  or g_42493_(_15232_, _15354_, _15500_);
  not g_42494_(_15500_, _15501_);
  and g_42495_(_15239_, _15354_, _15502_);
  not g_42496_(_15502_, _15503_);
  and g_42497_(_15500_, _15503_, _15504_);
  or g_42498_(_15501_, _15502_, _15505_);
  and g_42499_(_15497_, _15504_, _15506_);
  or g_42500_(_15498_, _15505_, _15507_);
  xor g_42501_(out[131], _15364_, _15508_);
  xor g_42502_(_21004_, _15364_, _15509_);
  or g_42503_(_15250_, _15354_, _15511_);
  not g_42504_(_15511_, _15512_);
  and g_42505_(_15256_, _15354_, _15513_);
  not g_42506_(_15513_, _15514_);
  and g_42507_(_15511_, _15514_, _15515_);
  or g_42508_(_15512_, _15513_, _15516_);
  and g_42509_(_15509_, _15516_, _15517_);
  or g_42510_(_15508_, _15515_, _15518_);
  and g_42511_(_15507_, _15518_, _15519_);
  or g_42512_(_15506_, _15517_, _15520_);
  and g_42513_(_15508_, _15515_, _15522_);
  not g_42514_(_15522_, _15523_);
  and g_42515_(_15498_, _15505_, _15524_);
  or g_42516_(_15522_, _15524_, _15525_);
  xor g_42517_(_15497_, _15504_, _15526_);
  xor g_42518_(_15508_, _15515_, _15527_);
  and g_42519_(_15526_, _15527_, _15528_);
  or g_42520_(_15520_, _15525_, _15529_);
  or g_42521_(out[112], _15354_, _15530_);
  not g_42522_(_15530_, _15531_);
  and g_42523_(_15214_, _15354_, _15533_);
  not g_42524_(_15533_, _15534_);
  and g_42525_(_15530_, _15534_, _15535_);
  or g_42526_(_15531_, _15533_, _15536_);
  and g_42527_(_20982_, _15535_, _15537_);
  or g_42528_(out[128], _15536_, _15538_);
  xor g_42529_(out[129], out[128], _15539_);
  not g_42530_(_15539_, _15540_);
  or g_42531_(_15228_, _15354_, _15541_);
  not g_42532_(_15541_, _15542_);
  and g_42533_(_15223_, _15354_, _15544_);
  not g_42534_(_15544_, _15545_);
  and g_42535_(_15541_, _15545_, _15546_);
  or g_42536_(_15542_, _15544_, _15547_);
  and g_42537_(_15539_, _15546_, _15548_);
  or g_42538_(_15540_, _15547_, _15549_);
  xor g_42539_(_15539_, _15546_, _15550_);
  xor g_42540_(_15540_, _15546_, _15551_);
  and g_42541_(_15538_, _15550_, _15552_);
  or g_42542_(_15537_, _15551_, _15553_);
  and g_42543_(_15528_, _15552_, _15555_);
  or g_42544_(_15529_, _15553_, _15556_);
  and g_42545_(_15520_, _15523_, _15557_);
  or g_42546_(_15519_, _15522_, _15558_);
  and g_42547_(_15528_, _15548_, _15559_);
  or g_42548_(_15557_, _15559_, _15560_);
  and g_42549_(_15549_, _15553_, _15561_);
  or g_42550_(_15529_, _15561_, _15562_);
  and g_42551_(_15558_, _15562_, _15563_);
  or g_42552_(_15555_, _15560_, _15564_);
  and g_42553_(_15495_, _15564_, _15566_);
  or g_42554_(_15496_, _15563_, _15567_);
  and g_42555_(_15484_, _15567_, _15568_);
  or g_42556_(_15485_, _15566_, _15569_);
  and g_42557_(_15429_, _15569_, _15570_);
  or g_42558_(_15430_, _15568_, _15571_);
  and g_42559_(_15421_, _15426_, _15572_);
  or g_42560_(_15420_, _15425_, _15573_);
  and g_42561_(_15571_, _15573_, _15574_);
  or g_42562_(_15570_, _15572_, _15575_);
  and g_42563_(_15398_, _15575_, _15577_);
  or g_42564_(_15399_, _15574_, _15578_);
  and g_42565_(_15391_, _15395_, _15579_);
  or g_42566_(_15390_, _15394_, _15580_);
  and g_42567_(_15578_, _15580_, _15581_);
  or g_42568_(_15577_, _15579_, _15582_);
  and g_42569_(out[128], _15536_, _15583_);
  or g_42570_(_20982_, _15535_, _15584_);
  and g_42571_(_15398_, _15584_, _15585_);
  or g_42572_(_15399_, _15583_, _15586_);
  and g_42573_(_15429_, _15585_, _15588_);
  or g_42574_(_15430_, _15586_, _15589_);
  and g_42575_(_15495_, _15555_, _15590_);
  or g_42576_(_15496_, _15556_, _15591_);
  and g_42577_(_15588_, _15590_, _15592_);
  or g_42578_(_15589_, _15591_, _15593_);
  and g_42579_(_15582_, _15593_, _15594_);
  or g_42580_(_15581_, _15592_, _15595_);
  and g_42581_(_15361_, _15595_, _15596_);
  and g_42582_(_15432_, _15594_, _15597_);
  or g_42583_(_15596_, _15597_, _15599_);
  and g_42584_(_13848_, _15599_, _15600_);
  not g_42585_(_15600_, _15601_);
  xor g_42586_(out[150], _13843_, _15602_);
  xor g_42587_(_21070_, _13843_, _15603_);
  and g_42588_(_15443_, _15595_, _15604_);
  or g_42589_(_15442_, _15594_, _15605_);
  and g_42590_(_15436_, _15594_, _15606_);
  or g_42591_(_15437_, _15595_, _15607_);
  and g_42592_(_15605_, _15607_, _15608_);
  or g_42593_(_15604_, _15606_, _15610_);
  and g_42594_(_15602_, _15608_, _15611_);
  or g_42595_(_15603_, _15610_, _15612_);
  xor g_42596_(out[149], _13842_, _15613_);
  xor g_42597_(_21092_, _13842_, _15614_);
  and g_42598_(_15458_, _15595_, _15615_);
  or g_42599_(_15459_, _15594_, _15616_);
  and g_42600_(_15452_, _15594_, _15617_);
  or g_42601_(_15451_, _15595_, _15618_);
  and g_42602_(_15616_, _15618_, _15619_);
  or g_42603_(_15615_, _15617_, _15621_);
  and g_42604_(_15614_, _15619_, _15622_);
  or g_42605_(_15613_, _15621_, _15623_);
  xor g_42606_(out[148], _13841_, _15624_);
  and g_42607_(_15463_, _15594_, _15625_);
  and g_42608_(_15469_, _15595_, _15626_);
  or g_42609_(_15625_, _15626_, _15627_);
  and g_42610_(_15624_, _15627_, _15628_);
  not g_42611_(_15628_, _15629_);
  and g_42612_(_15535_, _15595_, _15630_);
  or g_42613_(_15536_, _15594_, _15632_);
  and g_42614_(out[128], _15594_, _15633_);
  or g_42615_(_20982_, _15595_, _15634_);
  and g_42616_(_15632_, _15634_, _15635_);
  or g_42617_(_15630_, _15633_, _15636_);
  and g_42618_(out[144], _15635_, _15637_);
  or g_42619_(_21114_, _15636_, _15638_);
  and g_42620_(_15539_, _15594_, _15639_);
  or g_42621_(_15540_, _15595_, _15640_);
  and g_42622_(_15547_, _15595_, _15641_);
  or g_42623_(_15546_, _15594_, _15643_);
  and g_42624_(_15640_, _15643_, _15644_);
  or g_42625_(_15639_, _15641_, _15645_);
  and g_42626_(out[145], _15645_, _15646_);
  or g_42627_(_21103_, _15644_, _15647_);
  xor g_42628_(_21103_, out[144], _15648_);
  and g_42629_(_15637_, _15647_, _15649_);
  or g_42630_(_15638_, _15646_, _15650_);
  xor g_42631_(out[146], _13839_, _15651_);
  xor g_42632_(_21125_, _13839_, _15652_);
  and g_42633_(_15505_, _15595_, _15654_);
  or g_42634_(_15504_, _15594_, _15655_);
  and g_42635_(_15497_, _15594_, _15656_);
  or g_42636_(_15498_, _15595_, _15657_);
  and g_42637_(_15655_, _15657_, _15658_);
  or g_42638_(_15654_, _15656_, _15659_);
  and g_42639_(_15651_, _15658_, _15660_);
  or g_42640_(_15652_, _15659_, _15661_);
  or g_42641_(_15645_, _15648_, _15662_);
  not g_42642_(_15662_, _15663_);
  and g_42643_(_15661_, _15662_, _15665_);
  or g_42644_(_15649_, _15663_, _15666_);
  and g_42645_(_15650_, _15665_, _15667_);
  or g_42646_(_15660_, _15666_, _15668_);
  xor g_42647_(out[147], _13840_, _15669_);
  and g_42648_(_15509_, _15594_, _15670_);
  and g_42649_(_15515_, _15595_, _15671_);
  or g_42650_(_15670_, _15671_, _15672_);
  and g_42651_(_15669_, _15672_, _15673_);
  not g_42652_(_15673_, _15674_);
  and g_42653_(_15652_, _15659_, _15676_);
  or g_42654_(_15651_, _15658_, _15677_);
  and g_42655_(_15674_, _15677_, _15678_);
  or g_42656_(_15673_, _15676_, _15679_);
  and g_42657_(_15668_, _15678_, _15680_);
  or g_42658_(_15667_, _15679_, _15681_);
  or g_42659_(_15624_, _15627_, _15682_);
  or g_42660_(_15669_, _15672_, _15683_);
  and g_42661_(_15682_, _15683_, _15684_);
  not g_42662_(_15684_, _15685_);
  and g_42663_(_15681_, _15684_, _15687_);
  or g_42664_(_15680_, _15685_, _15688_);
  and g_42665_(_15629_, _15688_, _15689_);
  or g_42666_(_15628_, _15687_, _15690_);
  and g_42667_(_15623_, _15690_, _15691_);
  or g_42668_(_15622_, _15689_, _15692_);
  and g_42669_(_15603_, _15610_, _15693_);
  or g_42670_(_15602_, _15608_, _15694_);
  and g_42671_(_15613_, _15621_, _15695_);
  or g_42672_(_15614_, _15619_, _15696_);
  and g_42673_(_15694_, _15696_, _15698_);
  or g_42674_(_15693_, _15695_, _15699_);
  and g_42675_(_15692_, _15698_, _15700_);
  or g_42676_(_15691_, _15699_, _15701_);
  and g_42677_(_15612_, _15701_, _15702_);
  or g_42678_(_15611_, _15700_, _15703_);
  and g_42679_(_15601_, _15703_, _15704_);
  or g_42680_(_15600_, _15702_, _15705_);
  or g_42681_(out[153], _13846_, _15706_);
  and g_42682_(out[154], _15706_, _15707_);
  xor g_42683_(out[154], _15706_, _15709_);
  and g_42684_(_15379_, _15595_, _15710_);
  and g_42685_(_15375_, _15594_, _15711_);
  or g_42686_(_15710_, _15711_, _15712_);
  and g_42687_(_15709_, _15712_, _15713_);
  not g_42688_(_15713_, _15714_);
  and g_42689_(_15383_, _15385_, _15715_);
  or g_42690_(_15384_, _15386_, _15716_);
  xor g_42691_(out[155], _15707_, _15717_);
  xor g_42692_(_21048_, _15707_, _15718_);
  and g_42693_(_15716_, _15717_, _15720_);
  or g_42694_(_15715_, _15718_, _15721_);
  and g_42695_(_15714_, _15721_, _15722_);
  or g_42696_(_15713_, _15720_, _15723_);
  or g_42697_(_15716_, _15717_, _15724_);
  or g_42698_(_15709_, _15712_, _15725_);
  and g_42699_(_15724_, _15725_, _15726_);
  and g_42700_(_15722_, _15726_, _15727_);
  and g_42701_(_15416_, _15595_, _15728_);
  and g_42702_(_15413_, _15594_, _15729_);
  or g_42703_(_15728_, _15729_, _15731_);
  or g_42704_(_13848_, _15599_, _15732_);
  xor g_42705_(out[153], _13846_, _15733_);
  xor g_42706_(_21158_, _13846_, _15734_);
  and g_42707_(_15407_, _15595_, _15735_);
  and g_42708_(_15401_, _15594_, _15736_);
  or g_42709_(_15735_, _15736_, _15737_);
  or g_42710_(_15734_, _15737_, _15738_);
  and g_42711_(_15734_, _15737_, _15739_);
  and g_42712_(_13847_, _15731_, _15740_);
  or g_42713_(_15739_, _15740_, _15742_);
  xor g_42714_(_15734_, _15737_, _15743_);
  xor g_42715_(_13847_, _15731_, _15744_);
  and g_42716_(_15743_, _15744_, _15745_);
  and g_42717_(_15727_, _15745_, _15746_);
  and g_42718_(_15732_, _15746_, _15747_);
  not g_42719_(_15747_, _15748_);
  and g_42720_(_15705_, _15747_, _15749_);
  or g_42721_(_15704_, _15748_, _15750_);
  and g_42722_(_15738_, _15742_, _15751_);
  and g_42723_(_15727_, _15751_, _15753_);
  and g_42724_(_15723_, _15724_, _15754_);
  or g_42725_(_15753_, _15754_, _15755_);
  not g_42726_(_15755_, _15756_);
  and g_42727_(_15750_, _15756_, _15757_);
  or g_42728_(_15749_, _15755_, _15758_);
  or g_42729_(_13847_, _15758_, _15759_);
  not g_42730_(_15759_, _15760_);
  and g_42731_(_15731_, _15758_, _15761_);
  or g_42732_(_15760_, _15761_, _15762_);
  or g_42733_(out[304], out[305], _15764_);
  or g_42734_(out[304], _20292_, _15765_);
  and g_42735_(out[307], _15765_, _15766_);
  and g_42736_(_10328_, _15765_, _15767_);
  and g_42737_(out[309], _15767_, _15768_);
  or g_42738_(out[310], _15768_, _15769_);
  and g_42739_(out[311], _15769_, _15770_);
  and g_42740_(out[312], _15770_, _15771_);
  xor g_42741_(_19827_, _15770_, _15772_);
  xor g_42742_(out[306], _15764_, _15773_);
  not g_42743_(_15773_, _15775_);
  or g_42744_(out[288], out[289], _15776_);
  or g_42745_(out[288], _20106_, _15777_);
  xor g_42746_(out[290], _15776_, _15778_);
  xor g_42747_(_19684_, _15776_, _15779_);
  and g_42748_(out[291], _15777_, _15780_);
  and g_42749_(_10139_, _15777_, _15781_);
  and g_42750_(out[293], _15781_, _15782_);
  or g_42751_(out[294], _15782_, _15783_);
  and g_42752_(out[295], _15783_, _15784_);
  xor g_42753_(out[295], _15783_, _15786_);
  xor g_42754_(_19629_, _15783_, _15787_);
  or g_42755_(out[273], out[272], _15788_);
  or g_42756_(out[272], _19885_, _15789_);
  and g_42757_(out[275], _15789_, _15790_);
  and g_42758_(_09913_, _15789_, _15791_);
  and g_42759_(out[277], _15791_, _15792_);
  or g_42760_(out[278], _15792_, _15793_);
  and g_42761_(out[279], _15793_, _15794_);
  xor g_42762_(out[279], _15793_, _15795_);
  xor g_42763_(_19497_, _15793_, _15797_);
  xor g_42764_(out[275], _15789_, _15798_);
  xor g_42765_(_19574_, _15789_, _15799_);
  or g_42766_(out[257], out[256], _15800_);
  or g_42767_(out[256], _19672_, _15801_);
  and g_42768_(out[259], _15801_, _15802_);
  xor g_42769_(out[259], _15801_, _15803_);
  xor g_42770_(_19442_, _15801_, _15804_);
  and g_42771_(_09732_, _15801_, _15805_);
  and g_42772_(out[261], _15805_, _15806_);
  or g_42773_(out[262], _15806_, _15808_);
  and g_42774_(out[263], _15808_, _15809_);
  xor g_42775_(out[263], _15808_, _15810_);
  xor g_42776_(_19365_, _15808_, _15811_);
  or g_42777_(out[160], _18467_, _15812_);
  and g_42778_(out[163], _15812_, _15813_);
  not g_42779_(_15813_, _15814_);
  and g_42780_(_26214_, _15812_, _15815_);
  and g_42781_(out[165], _15815_, _15816_);
  or g_42782_(out[166], _15816_, _15817_);
  and g_42783_(out[167], _15817_, _15819_);
  xor g_42784_(out[167], _15817_, _15820_);
  xor g_42785_(_18606_, _15817_, _15821_);
  and g_42786_(out[168], _15819_, _15822_);
  or g_42787_(out[169], _15822_, _15823_);
  and g_42788_(out[170], _15823_, _15824_);
  xor g_42789_(out[171], _15824_, _15825_);
  xor g_42790_(_18595_, _15824_, _15826_);
  and g_42791_(_18771_, _18782_, _15827_);
  or g_42792_(out[177], out[176], _15828_);
  or g_42793_(out[176], _18463_, _15830_);
  and g_42794_(out[179], _15830_, _15831_);
  and g_42795_(_26224_, _15830_, _15832_);
  and g_42796_(out[181], _15832_, _15833_);
  or g_42797_(out[182], _15833_, _15834_);
  and g_42798_(out[183], _15834_, _15835_);
  and g_42799_(out[184], _15835_, _15836_);
  or g_42800_(out[185], _15836_, _15837_);
  and g_42801_(out[186], _15837_, _15838_);
  xor g_42802_(out[187], _15838_, _15839_);
  xor g_42803_(_18716_, _15838_, _15841_);
  and g_42804_(_15826_, _15839_, _15842_);
  or g_42805_(_15825_, _15841_, _15843_);
  xor g_42806_(out[166], _15816_, _15844_);
  xor g_42807_(_18617_, _15816_, _15845_);
  xor g_42808_(out[182], _15833_, _15846_);
  xor g_42809_(_18738_, _15833_, _15847_);
  and g_42810_(_15844_, _15847_, _15848_);
  or g_42811_(_15845_, _15846_, _15849_);
  xor g_42812_(out[165], _15815_, _15850_);
  xor g_42813_(_18628_, _15815_, _15852_);
  xor g_42814_(out[181], _15832_, _15853_);
  xor g_42815_(_18749_, _15832_, _15854_);
  and g_42816_(_15850_, _15854_, _15855_);
  or g_42817_(_15852_, _15853_, _15856_);
  and g_42818_(out[161], out[177], _15857_);
  not g_42819_(_15857_, _15858_);
  and g_42820_(_18507_, _15857_, _15859_);
  or g_42821_(_18506_, _15858_, _15860_);
  and g_42822_(out[160], _18650_, _15861_);
  or g_42823_(_18584_, out[161], _15863_);
  and g_42824_(_15828_, _15863_, _15864_);
  or g_42825_(_15827_, _15861_, _15865_);
  and g_42826_(_15860_, _15864_, _15866_);
  or g_42827_(_15859_, _15865_, _15867_);
  xor g_42828_(out[178], _15828_, _15868_);
  xor g_42829_(_18793_, _15828_, _15869_);
  or g_42830_(out[160], _18468_, _15870_);
  not g_42831_(_15870_, _15871_);
  and g_42832_(out[160], out[162], _15872_);
  not g_42833_(_15872_, _15874_);
  or g_42834_(_15871_, _15872_, _15875_);
  and g_42835_(_15870_, _15874_, _15876_);
  or g_42836_(out[160], _22444_, _15877_);
  not g_42837_(_15877_, _15878_);
  and g_42838_(_15814_, _15877_, _15879_);
  or g_42839_(_15813_, _15878_, _15880_);
  xor g_42840_(out[179], _15830_, _15881_);
  xor g_42841_(_18804_, _15830_, _15882_);
  and g_42842_(_15880_, _15881_, _15883_);
  or g_42843_(_15879_, _15882_, _15885_);
  and g_42844_(_15867_, _15869_, _15886_);
  or g_42845_(_15866_, _15868_, _15887_);
  and g_42846_(_15866_, _15868_, _15888_);
  or g_42847_(_15867_, _15869_, _15889_);
  and g_42848_(_15876_, _15889_, _15890_);
  or g_42849_(_15875_, _15888_, _15891_);
  and g_42850_(_15887_, _15891_, _15892_);
  or g_42851_(_15886_, _15890_, _15893_);
  and g_42852_(_15885_, _15892_, _15894_);
  or g_42853_(_15883_, _15893_, _15896_);
  and g_42854_(_15879_, _15882_, _15897_);
  or g_42855_(_15880_, _15881_, _15898_);
  xor g_42856_(out[164], _15813_, _15899_);
  xor g_42857_(_18639_, _15813_, _15900_);
  xor g_42858_(out[180], _15831_, _15901_);
  xor g_42859_(_18760_, _15831_, _15902_);
  and g_42860_(_15899_, _15902_, _15903_);
  or g_42861_(_15900_, _15901_, _15904_);
  and g_42862_(_15898_, _15904_, _15905_);
  or g_42863_(_15897_, _15903_, _15907_);
  and g_42864_(_15896_, _15905_, _15908_);
  or g_42865_(_15894_, _15907_, _15909_);
  and g_42866_(_15900_, _15901_, _15910_);
  or g_42867_(_15899_, _15902_, _15911_);
  and g_42868_(_15852_, _15853_, _15912_);
  or g_42869_(_15850_, _15854_, _15913_);
  and g_42870_(_15911_, _15913_, _15914_);
  or g_42871_(_15910_, _15912_, _15915_);
  and g_42872_(_15909_, _15914_, _15916_);
  or g_42873_(_15908_, _15915_, _15918_);
  and g_42874_(_15856_, _15918_, _15919_);
  or g_42875_(_15855_, _15916_, _15920_);
  and g_42876_(_15849_, _15920_, _15921_);
  or g_42877_(_15848_, _15919_, _15922_);
  xor g_42878_(out[183], _15834_, _15923_);
  xor g_42879_(_18727_, _15834_, _15924_);
  and g_42880_(_15820_, _15924_, _15925_);
  or g_42881_(_15821_, _15923_, _15926_);
  and g_42882_(_15845_, _15846_, _15927_);
  or g_42883_(_15844_, _15847_, _15929_);
  and g_42884_(_15926_, _15929_, _15930_);
  or g_42885_(_15925_, _15927_, _15931_);
  and g_42886_(_15922_, _15930_, _15932_);
  or g_42887_(_15921_, _15931_, _15933_);
  xor g_42888_(out[168], _15819_, _15934_);
  xor g_42889_(_18683_, _15819_, _15935_);
  xor g_42890_(out[184], _15835_, _15936_);
  xor g_42891_(_18815_, _15835_, _15937_);
  and g_42892_(_15935_, _15936_, _15938_);
  or g_42893_(_15934_, _15937_, _15940_);
  and g_42894_(_15821_, _15923_, _15941_);
  or g_42895_(_15820_, _15924_, _15942_);
  and g_42896_(_15940_, _15942_, _15943_);
  or g_42897_(_15938_, _15941_, _15944_);
  and g_42898_(_15933_, _15943_, _15945_);
  or g_42899_(_15932_, _15944_, _15946_);
  xor g_42900_(out[169], _15822_, _15947_);
  xor g_42901_(_18694_, _15822_, _15948_);
  xor g_42902_(out[185], _15836_, _15949_);
  xor g_42903_(_18826_, _15836_, _15951_);
  and g_42904_(_15948_, _15949_, _15952_);
  or g_42905_(_15947_, _15951_, _15953_);
  and g_42906_(_15934_, _15937_, _15954_);
  or g_42907_(_15935_, _15936_, _15955_);
  and g_42908_(_15953_, _15955_, _15956_);
  or g_42909_(_15952_, _15954_, _15957_);
  and g_42910_(_15946_, _15956_, _15958_);
  or g_42911_(_15945_, _15957_, _15959_);
  and g_42912_(_15947_, _15951_, _15960_);
  or g_42913_(_15948_, _15949_, _15962_);
  xor g_42914_(out[186], _15837_, _15963_);
  xor g_42915_(_18837_, _15837_, _15964_);
  xor g_42916_(out[170], _15823_, _15965_);
  xor g_42917_(_18705_, _15823_, _15966_);
  and g_42918_(_15963_, _15966_, _15967_);
  or g_42919_(_15964_, _15965_, _15968_);
  and g_42920_(_15962_, _15968_, _15969_);
  or g_42921_(_15960_, _15967_, _15970_);
  and g_42922_(_15959_, _15969_, _15971_);
  or g_42923_(_15958_, _15970_, _15973_);
  and g_42924_(_15964_, _15965_, _15974_);
  or g_42925_(_15963_, _15966_, _15975_);
  and g_42926_(_15825_, _15841_, _15976_);
  or g_42927_(_15826_, _15839_, _15977_);
  and g_42928_(_15975_, _15977_, _15978_);
  or g_42929_(_15974_, _15976_, _15979_);
  and g_42930_(_15973_, _15978_, _15980_);
  or g_42931_(_15971_, _15979_, _15981_);
  and g_42932_(_15843_, _15981_, _15982_);
  or g_42933_(_15842_, _15980_, _15984_);
  and g_42934_(_15821_, _15984_, _15985_);
  or g_42935_(_15820_, _15982_, _15986_);
  and g_42936_(_15924_, _15982_, _15987_);
  or g_42937_(_15923_, _15984_, _15988_);
  and g_42938_(_15986_, _15988_, _15989_);
  or g_42939_(_15985_, _15987_, _15990_);
  or g_42940_(out[193], out[192], _15991_);
  or g_42941_(out[192], _18741_, _15992_);
  and g_42942_(out[195], _15992_, _15993_);
  and g_42943_(_26375_, _15992_, _15995_);
  and g_42944_(out[197], _15995_, _15996_);
  or g_42945_(out[198], _15996_, _15997_);
  and g_42946_(out[199], _15997_, _15998_);
  xor g_42947_(out[199], _15997_, _15999_);
  xor g_42948_(_18859_, _15997_, _16000_);
  and g_42949_(_15990_, _15999_, _16001_);
  or g_42950_(_15989_, _16000_, _16002_);
  xor g_42951_(out[198], _15996_, _16003_);
  xor g_42952_(_18870_, _15996_, _16004_);
  and g_42953_(_15844_, _15984_, _16006_);
  or g_42954_(_15845_, _15982_, _16007_);
  and g_42955_(_15846_, _15982_, _16008_);
  or g_42956_(_15847_, _15984_, _16009_);
  and g_42957_(_16007_, _16009_, _16010_);
  or g_42958_(_16006_, _16008_, _16011_);
  and g_42959_(_16004_, _16011_, _16012_);
  or g_42960_(_16003_, _16010_, _16013_);
  xor g_42961_(out[197], _15995_, _16014_);
  xor g_42962_(_18881_, _15995_, _16015_);
  and g_42963_(_15852_, _15984_, _16017_);
  or g_42964_(_15850_, _15982_, _16018_);
  and g_42965_(_15854_, _15982_, _16019_);
  or g_42966_(_15853_, _15984_, _16020_);
  and g_42967_(_16018_, _16020_, _16021_);
  or g_42968_(_16017_, _16019_, _16022_);
  and g_42969_(_16015_, _16021_, _16023_);
  or g_42970_(_16014_, _16022_, _16024_);
  xor g_42971_(out[196], _15993_, _16025_);
  xor g_42972_(_18892_, _15993_, _16026_);
  and g_42973_(_15900_, _15984_, _16028_);
  or g_42974_(_15899_, _15982_, _16029_);
  and g_42975_(_15902_, _15982_, _16030_);
  or g_42976_(_15901_, _15984_, _16031_);
  and g_42977_(_16029_, _16031_, _16032_);
  or g_42978_(_16028_, _16030_, _16033_);
  and g_42979_(_16026_, _16032_, _16034_);
  or g_42980_(_16025_, _16033_, _16035_);
  xor g_42981_(out[195], _15992_, _16036_);
  xor g_42982_(_18936_, _15992_, _16037_);
  and g_42983_(_15880_, _15984_, _16039_);
  or g_42984_(_15879_, _15982_, _16040_);
  and g_42985_(_15882_, _15982_, _16041_);
  or g_42986_(_15881_, _15984_, _16042_);
  and g_42987_(_16040_, _16042_, _16043_);
  or g_42988_(_16039_, _16041_, _16044_);
  and g_42989_(_16036_, _16044_, _16045_);
  or g_42990_(_16037_, _16043_, _16046_);
  and g_42991_(_16037_, _16043_, _16047_);
  or g_42992_(_16036_, _16044_, _16048_);
  xor g_42993_(out[194], _15991_, _16050_);
  xor g_42994_(_18925_, _15991_, _16051_);
  and g_42995_(_15868_, _15982_, _16052_);
  or g_42996_(_15869_, _15984_, _16053_);
  and g_42997_(_15876_, _15984_, _16054_);
  or g_42998_(_15875_, _15982_, _16055_);
  and g_42999_(_16053_, _16055_, _16056_);
  or g_43000_(_16052_, _16054_, _16057_);
  and g_43001_(_16050_, _16056_, _16058_);
  or g_43002_(_16051_, _16057_, _16059_);
  xor g_43003_(_18584_, out[161], _16061_);
  xor g_43004_(out[160], out[161], _16062_);
  and g_43005_(_15984_, _16062_, _16063_);
  or g_43006_(_15982_, _16061_, _16064_);
  xor g_43007_(out[177], out[176], _16065_);
  xor g_43008_(_18771_, out[176], _16066_);
  and g_43009_(_15982_, _16065_, _16067_);
  or g_43010_(_15984_, _16066_, _16068_);
  and g_43011_(_16064_, _16068_, _16069_);
  or g_43012_(_16063_, _16067_, _16070_);
  and g_43013_(out[193], _16070_, _16072_);
  not g_43014_(_16072_, _16073_);
  xor g_43015_(out[193], out[192], _16074_);
  xor g_43016_(_18903_, out[192], _16075_);
  and g_43017_(_16069_, _16074_, _16076_);
  or g_43018_(_16070_, _16075_, _16077_);
  and g_43019_(out[176], _15982_, _16078_);
  or g_43020_(_18782_, _15984_, _16079_);
  and g_43021_(out[160], _15984_, _16080_);
  or g_43022_(_18584_, _15982_, _16081_);
  and g_43023_(_16079_, _16081_, _16083_);
  or g_43024_(_16078_, _16080_, _16084_);
  and g_43025_(out[192], _16083_, _16085_);
  or g_43026_(_18914_, _16084_, _16086_);
  and g_43027_(_16077_, _16086_, _16087_);
  or g_43028_(_16076_, _16085_, _16088_);
  and g_43029_(_16073_, _16088_, _16089_);
  or g_43030_(_16072_, _16087_, _16090_);
  and g_43031_(_16059_, _16090_, _16091_);
  or g_43032_(_16058_, _16089_, _16092_);
  and g_43033_(_16051_, _16057_, _16094_);
  or g_43034_(_16050_, _16056_, _16095_);
  and g_43035_(_16046_, _16095_, _16096_);
  or g_43036_(_16045_, _16094_, _16097_);
  and g_43037_(_16092_, _16096_, _16098_);
  or g_43038_(_16091_, _16097_, _16099_);
  and g_43039_(_16035_, _16048_, _16100_);
  or g_43040_(_16034_, _16047_, _16101_);
  and g_43041_(_16099_, _16100_, _16102_);
  or g_43042_(_16098_, _16101_, _16103_);
  and g_43043_(_16014_, _16022_, _16105_);
  or g_43044_(_16015_, _16021_, _16106_);
  and g_43045_(_16025_, _16033_, _16107_);
  or g_43046_(_16026_, _16032_, _16108_);
  and g_43047_(_16106_, _16108_, _16109_);
  or g_43048_(_16105_, _16107_, _16110_);
  and g_43049_(_16103_, _16109_, _16111_);
  or g_43050_(_16102_, _16110_, _16112_);
  and g_43051_(_16024_, _16112_, _16113_);
  or g_43052_(_16023_, _16111_, _16114_);
  and g_43053_(_16013_, _16114_, _16116_);
  or g_43054_(_16012_, _16113_, _16117_);
  and g_43055_(_15989_, _16000_, _16118_);
  or g_43056_(_15990_, _15999_, _16119_);
  and g_43057_(_16003_, _16010_, _16120_);
  or g_43058_(_16004_, _16011_, _16121_);
  and g_43059_(_16119_, _16121_, _16122_);
  or g_43060_(_16118_, _16120_, _16123_);
  and g_43061_(_16117_, _16122_, _16124_);
  or g_43062_(_16116_, _16123_, _16125_);
  and g_43063_(_16002_, _16125_, _16127_);
  or g_43064_(_16001_, _16124_, _16128_);
  and g_43065_(out[200], _15998_, _16129_);
  or g_43066_(out[201], _16129_, _16130_);
  not g_43067_(_16130_, _16131_);
  and g_43068_(out[202], _16130_, _16132_);
  xor g_43069_(out[202], _16130_, _16133_);
  xor g_43070_(out[202], _16131_, _16134_);
  and g_43071_(_15966_, _15984_, _16135_);
  or g_43072_(_15965_, _15982_, _16136_);
  and g_43073_(_15964_, _15982_, _16138_);
  or g_43074_(_15963_, _15984_, _16139_);
  and g_43075_(_16136_, _16139_, _16140_);
  or g_43076_(_16135_, _16138_, _16141_);
  and g_43077_(_16133_, _16141_, _16142_);
  or g_43078_(_16134_, _16140_, _16143_);
  and g_43079_(_15825_, _15839_, _16144_);
  or g_43080_(_15826_, _15841_, _16145_);
  xor g_43081_(out[203], _16132_, _16146_);
  xor g_43082_(_18848_, _16132_, _16147_);
  and g_43083_(_16144_, _16147_, _16149_);
  or g_43084_(_16145_, _16146_, _16150_);
  and g_43085_(_16145_, _16146_, _16151_);
  or g_43086_(_16144_, _16147_, _16152_);
  and g_43087_(out[201], _16129_, _16153_);
  xor g_43088_(out[201], _16129_, _16154_);
  or g_43089_(_16131_, _16153_, _16155_);
  and g_43090_(_15947_, _15984_, _16156_);
  or g_43091_(_15948_, _15982_, _16157_);
  and g_43092_(_15949_, _15982_, _16158_);
  or g_43093_(_15951_, _15984_, _16160_);
  and g_43094_(_16157_, _16160_, _16161_);
  or g_43095_(_16156_, _16158_, _16162_);
  and g_43096_(_16154_, _16161_, _16163_);
  or g_43097_(_16155_, _16162_, _16164_);
  and g_43098_(_16134_, _16140_, _16165_);
  or g_43099_(_16133_, _16141_, _16166_);
  and g_43100_(_16152_, _16166_, _16167_);
  or g_43101_(_16151_, _16165_, _16168_);
  and g_43102_(_16143_, _16164_, _16169_);
  or g_43103_(_16142_, _16163_, _16171_);
  and g_43104_(_16150_, _16169_, _16172_);
  or g_43105_(_16149_, _16171_, _16173_);
  and g_43106_(_16167_, _16172_, _16174_);
  or g_43107_(_16168_, _16173_, _16175_);
  xor g_43108_(out[200], _15998_, _16176_);
  xor g_43109_(_18947_, _15998_, _16177_);
  and g_43110_(_15934_, _15984_, _16178_);
  or g_43111_(_15935_, _15982_, _16179_);
  and g_43112_(_15936_, _15982_, _16180_);
  or g_43113_(_15937_, _15984_, _16182_);
  and g_43114_(_16179_, _16182_, _16183_);
  or g_43115_(_16178_, _16180_, _16184_);
  and g_43116_(_16176_, _16183_, _16185_);
  or g_43117_(_16177_, _16184_, _16186_);
  and g_43118_(_16155_, _16162_, _16187_);
  or g_43119_(_16154_, _16161_, _16188_);
  and g_43120_(_16186_, _16188_, _16189_);
  or g_43121_(_16185_, _16187_, _16190_);
  and g_43122_(_16177_, _16184_, _16191_);
  or g_43123_(_16176_, _16183_, _16193_);
  and g_43124_(_16189_, _16193_, _16194_);
  or g_43125_(_16190_, _16191_, _16195_);
  and g_43126_(_16174_, _16194_, _16196_);
  or g_43127_(_16175_, _16195_, _16197_);
  and g_43128_(_16128_, _16196_, _16198_);
  or g_43129_(_16127_, _16197_, _16199_);
  and g_43130_(_16174_, _16190_, _16200_);
  or g_43131_(_16175_, _16189_, _16201_);
  and g_43132_(_16143_, _16152_, _16202_);
  or g_43133_(_16142_, _16151_, _16204_);
  and g_43134_(_16150_, _16204_, _16205_);
  or g_43135_(_16149_, _16202_, _16206_);
  and g_43136_(_16201_, _16206_, _16207_);
  or g_43137_(_16200_, _16205_, _16208_);
  and g_43138_(_16199_, _16207_, _16209_);
  or g_43139_(_16198_, _16208_, _16210_);
  and g_43140_(_15990_, _16210_, _16211_);
  or g_43141_(_15989_, _16209_, _16212_);
  and g_43142_(_16000_, _16209_, _16213_);
  or g_43143_(_15999_, _16210_, _16215_);
  and g_43144_(_16212_, _16215_, _16216_);
  or g_43145_(_16211_, _16213_, _16217_);
  and g_43146_(out[192], _16209_, _16218_);
  or g_43147_(_18914_, _16210_, _16219_);
  and g_43148_(_16084_, _16210_, _16220_);
  or g_43149_(_16083_, _16209_, _16221_);
  and g_43150_(_16219_, _16221_, _16222_);
  or g_43151_(_16218_, _16220_, _16223_);
  and g_43152_(out[208], _16222_, _16224_);
  or g_43153_(_19024_, _16223_, _16226_);
  and g_43154_(_16074_, _16209_, _16227_);
  or g_43155_(_16075_, _16210_, _16228_);
  and g_43156_(_16070_, _16210_, _16229_);
  or g_43157_(_16069_, _16209_, _16230_);
  and g_43158_(_16228_, _16230_, _16231_);
  or g_43159_(_16227_, _16229_, _16232_);
  and g_43160_(out[209], _16232_, _16233_);
  or g_43161_(_19013_, _16231_, _16234_);
  or g_43162_(out[209], out[208], _16235_);
  xor g_43163_(out[209], out[208], _16237_);
  xor g_43164_(_19013_, out[208], _16238_);
  and g_43165_(_16224_, _16234_, _16239_);
  or g_43166_(_16226_, _16233_, _16240_);
  or g_43167_(out[208], _18849_, _16241_);
  xor g_43168_(out[210], _16235_, _16242_);
  xor g_43169_(_19035_, _16235_, _16243_);
  and g_43170_(_16050_, _16209_, _16244_);
  or g_43171_(_16051_, _16210_, _16245_);
  and g_43172_(_16057_, _16210_, _16246_);
  or g_43173_(_16056_, _16209_, _16248_);
  and g_43174_(_16245_, _16248_, _16249_);
  or g_43175_(_16244_, _16246_, _16250_);
  and g_43176_(_16242_, _16249_, _16251_);
  or g_43177_(_16243_, _16250_, _16252_);
  and g_43178_(_16231_, _16237_, _16253_);
  or g_43179_(_16232_, _16238_, _16254_);
  and g_43180_(_16252_, _16254_, _16255_);
  or g_43181_(_16251_, _16253_, _16256_);
  and g_43182_(_16240_, _16255_, _16257_);
  or g_43183_(_16239_, _16256_, _16259_);
  and g_43184_(out[211], _16241_, _16260_);
  xor g_43185_(out[211], _16241_, _16261_);
  xor g_43186_(_19046_, _16241_, _16262_);
  and g_43187_(_16037_, _16209_, _16263_);
  or g_43188_(_16036_, _16210_, _16264_);
  and g_43189_(_16044_, _16210_, _16265_);
  or g_43190_(_16043_, _16209_, _16266_);
  and g_43191_(_16264_, _16266_, _16267_);
  or g_43192_(_16263_, _16265_, _16268_);
  and g_43193_(_16261_, _16268_, _16270_);
  or g_43194_(_16262_, _16267_, _16271_);
  and g_43195_(_16243_, _16250_, _16272_);
  or g_43196_(_16242_, _16249_, _16273_);
  and g_43197_(_16271_, _16273_, _16274_);
  or g_43198_(_16270_, _16272_, _16275_);
  and g_43199_(_16259_, _16274_, _16276_);
  or g_43200_(_16257_, _16275_, _16277_);
  and g_43201_(_26601_, _16241_, _16278_);
  xor g_43202_(out[212], _16260_, _16279_);
  xor g_43203_(_19002_, _16260_, _16281_);
  and g_43204_(_16033_, _16210_, _16282_);
  or g_43205_(_16032_, _16209_, _16283_);
  and g_43206_(_16026_, _16209_, _16284_);
  or g_43207_(_16025_, _16210_, _16285_);
  and g_43208_(_16283_, _16285_, _16286_);
  or g_43209_(_16282_, _16284_, _16287_);
  and g_43210_(_16281_, _16286_, _16288_);
  or g_43211_(_16279_, _16287_, _16289_);
  and g_43212_(_16262_, _16267_, _16290_);
  or g_43213_(_16261_, _16268_, _16292_);
  and g_43214_(_16289_, _16292_, _16293_);
  or g_43215_(_16288_, _16290_, _16294_);
  and g_43216_(_16277_, _16293_, _16295_);
  or g_43217_(_16276_, _16294_, _16296_);
  and g_43218_(out[213], _16278_, _16297_);
  xor g_43219_(out[213], _16278_, _16298_);
  xor g_43220_(_18991_, _16278_, _16299_);
  and g_43221_(_16015_, _16209_, _16300_);
  or g_43222_(_16014_, _16210_, _16301_);
  and g_43223_(_16022_, _16210_, _16303_);
  or g_43224_(_16021_, _16209_, _16304_);
  and g_43225_(_16301_, _16304_, _16305_);
  or g_43226_(_16300_, _16303_, _16306_);
  and g_43227_(_16298_, _16306_, _16307_);
  or g_43228_(_16299_, _16305_, _16308_);
  and g_43229_(_16279_, _16287_, _16309_);
  or g_43230_(_16281_, _16286_, _16310_);
  and g_43231_(_16308_, _16310_, _16311_);
  or g_43232_(_16307_, _16309_, _16312_);
  and g_43233_(_16296_, _16311_, _16314_);
  or g_43234_(_16295_, _16312_, _16315_);
  or g_43235_(out[214], _16297_, _16316_);
  xor g_43236_(out[214], _16297_, _16317_);
  xor g_43237_(_18980_, _16297_, _16318_);
  and g_43238_(_16011_, _16210_, _16319_);
  or g_43239_(_16010_, _16209_, _16320_);
  and g_43240_(_16003_, _16209_, _16321_);
  or g_43241_(_16004_, _16210_, _16322_);
  and g_43242_(_16320_, _16322_, _16323_);
  or g_43243_(_16319_, _16321_, _16325_);
  and g_43244_(_16317_, _16323_, _16326_);
  or g_43245_(_16318_, _16325_, _16327_);
  and g_43246_(_16299_, _16305_, _16328_);
  or g_43247_(_16298_, _16306_, _16329_);
  and g_43248_(_16327_, _16329_, _16330_);
  or g_43249_(_16326_, _16328_, _16331_);
  and g_43250_(_16315_, _16330_, _16332_);
  or g_43251_(_16314_, _16331_, _16333_);
  and g_43252_(out[215], _16316_, _16334_);
  xor g_43253_(out[215], _16316_, _16336_);
  xor g_43254_(_18969_, _16316_, _16337_);
  and g_43255_(_16217_, _16336_, _16338_);
  or g_43256_(_16216_, _16337_, _16339_);
  and g_43257_(_16318_, _16325_, _16340_);
  or g_43258_(_16317_, _16323_, _16341_);
  and g_43259_(_16339_, _16341_, _16342_);
  or g_43260_(_16338_, _16340_, _16343_);
  and g_43261_(_16333_, _16342_, _16344_);
  or g_43262_(_16332_, _16343_, _16345_);
  and g_43263_(out[216], _16334_, _16347_);
  or g_43264_(out[217], _16347_, _16348_);
  xor g_43265_(out[217], _16347_, _16349_);
  xor g_43266_(_19068_, _16347_, _16350_);
  and g_43267_(_16162_, _16210_, _16351_);
  or g_43268_(_16161_, _16209_, _16352_);
  and g_43269_(_16154_, _16209_, _16353_);
  or g_43270_(_16155_, _16210_, _16354_);
  and g_43271_(_16352_, _16354_, _16355_);
  or g_43272_(_16351_, _16353_, _16356_);
  and g_43273_(_16349_, _16355_, _16358_);
  or g_43274_(_16350_, _16356_, _16359_);
  xor g_43275_(out[216], _16334_, _16360_);
  xor g_43276_(_19057_, _16334_, _16361_);
  and g_43277_(_16184_, _16210_, _16362_);
  or g_43278_(_16183_, _16209_, _16363_);
  and g_43279_(_16176_, _16209_, _16364_);
  or g_43280_(_16177_, _16210_, _16365_);
  and g_43281_(_16363_, _16365_, _16366_);
  or g_43282_(_16362_, _16364_, _16367_);
  and g_43283_(_16361_, _16367_, _16369_);
  or g_43284_(_16360_, _16366_, _16370_);
  and g_43285_(_16359_, _16370_, _16371_);
  or g_43286_(_16358_, _16369_, _16372_);
  and g_43287_(_16216_, _16337_, _16373_);
  or g_43288_(_16217_, _16336_, _16374_);
  and g_43289_(_16371_, _16374_, _16375_);
  or g_43290_(_16372_, _16373_, _16376_);
  and g_43291_(out[218], _16348_, _16377_);
  xor g_43292_(out[218], _16348_, _16378_);
  xor g_43293_(_19079_, _16348_, _16380_);
  and g_43294_(_16141_, _16210_, _16381_);
  or g_43295_(_16140_, _16209_, _16382_);
  and g_43296_(_16134_, _16209_, _16383_);
  or g_43297_(_16133_, _16210_, _16384_);
  and g_43298_(_16382_, _16384_, _16385_);
  or g_43299_(_16381_, _16383_, _16386_);
  and g_43300_(_16378_, _16386_, _16387_);
  or g_43301_(_16380_, _16385_, _16388_);
  and g_43302_(_16144_, _16146_, _16389_);
  or g_43303_(_16145_, _16147_, _16391_);
  xor g_43304_(out[219], _16377_, _16392_);
  xor g_43305_(_18958_, _16377_, _16393_);
  and g_43306_(_16391_, _16392_, _16394_);
  or g_43307_(_16389_, _16393_, _16395_);
  and g_43308_(_16388_, _16395_, _16396_);
  or g_43309_(_16387_, _16394_, _16397_);
  and g_43310_(_16389_, _16393_, _16398_);
  or g_43311_(_16391_, _16392_, _16399_);
  and g_43312_(_16380_, _16385_, _16400_);
  or g_43313_(_16378_, _16386_, _16402_);
  and g_43314_(_16399_, _16402_, _16403_);
  or g_43315_(_16398_, _16400_, _16404_);
  and g_43316_(_16360_, _16366_, _16405_);
  or g_43317_(_16361_, _16367_, _16406_);
  and g_43318_(_16350_, _16356_, _16407_);
  or g_43319_(_16349_, _16355_, _16408_);
  and g_43320_(_16406_, _16408_, _16409_);
  or g_43321_(_16405_, _16407_, _16410_);
  and g_43322_(_16403_, _16409_, _16411_);
  or g_43323_(_16404_, _16410_, _16413_);
  and g_43324_(_16396_, _16411_, _16414_);
  or g_43325_(_16397_, _16413_, _16415_);
  and g_43326_(_16375_, _16414_, _16416_);
  or g_43327_(_16376_, _16415_, _16417_);
  and g_43328_(_16345_, _16416_, _16418_);
  or g_43329_(_16344_, _16417_, _16419_);
  and g_43330_(_16397_, _16399_, _16420_);
  or g_43331_(_16396_, _16398_, _16421_);
  and g_43332_(_16403_, _16410_, _16422_);
  or g_43333_(_16404_, _16409_, _16424_);
  and g_43334_(_16359_, _16422_, _16425_);
  or g_43335_(_16358_, _16424_, _16426_);
  and g_43336_(_16421_, _16426_, _16427_);
  or g_43337_(_16420_, _16425_, _16428_);
  and g_43338_(_16419_, _16427_, _16429_);
  or g_43339_(_16418_, _16428_, _16430_);
  and g_43340_(_16217_, _16430_, _16431_);
  or g_43341_(_16216_, _16429_, _16432_);
  and g_43342_(_16337_, _16429_, _16433_);
  or g_43343_(_16336_, _16430_, _16435_);
  and g_43344_(_16432_, _16435_, _16436_);
  or g_43345_(_16431_, _16433_, _16437_);
  and g_43346_(out[208], _16429_, _16438_);
  or g_43347_(_19024_, _16430_, _16439_);
  and g_43348_(_16223_, _16430_, _16440_);
  or g_43349_(_16222_, _16429_, _16441_);
  and g_43350_(_16439_, _16441_, _16442_);
  or g_43351_(_16438_, _16440_, _16443_);
  and g_43352_(out[224], _16442_, _16444_);
  or g_43353_(_19156_, _16443_, _16446_);
  and g_43354_(_16237_, _16429_, _16447_);
  or g_43355_(_16238_, _16430_, _16448_);
  and g_43356_(_16232_, _16430_, _16449_);
  or g_43357_(_16231_, _16429_, _16450_);
  and g_43358_(_16448_, _16450_, _16451_);
  or g_43359_(_16447_, _16449_, _16452_);
  and g_43360_(out[225], _16452_, _16453_);
  or g_43361_(_19145_, _16451_, _16454_);
  or g_43362_(out[225], out[224], _16455_);
  xor g_43363_(out[225], out[224], _16457_);
  xor g_43364_(_19145_, out[224], _16458_);
  and g_43365_(_16444_, _16454_, _16459_);
  or g_43366_(_16446_, _16453_, _16460_);
  or g_43367_(out[224], _19229_, _16461_);
  xor g_43368_(out[226], _16455_, _16462_);
  xor g_43369_(_19167_, _16455_, _16463_);
  and g_43370_(_16250_, _16430_, _16464_);
  or g_43371_(_16249_, _16429_, _16465_);
  and g_43372_(_16242_, _16429_, _16466_);
  or g_43373_(_16243_, _16430_, _16468_);
  and g_43374_(_16465_, _16468_, _16469_);
  or g_43375_(_16464_, _16466_, _16470_);
  and g_43376_(_16462_, _16469_, _16471_);
  or g_43377_(_16463_, _16470_, _16472_);
  and g_43378_(_16451_, _16457_, _16473_);
  or g_43379_(_16452_, _16458_, _16474_);
  and g_43380_(_16472_, _16474_, _16475_);
  or g_43381_(_16471_, _16473_, _16476_);
  and g_43382_(_16460_, _16475_, _16477_);
  or g_43383_(_16459_, _16476_, _16479_);
  and g_43384_(out[227], _16461_, _16480_);
  xor g_43385_(out[227], _16461_, _16481_);
  xor g_43386_(_19178_, _16461_, _16482_);
  and g_43387_(_16262_, _16429_, _16483_);
  or g_43388_(_16261_, _16430_, _16484_);
  and g_43389_(_16268_, _16430_, _16485_);
  or g_43390_(_16267_, _16429_, _16486_);
  and g_43391_(_16484_, _16486_, _16487_);
  or g_43392_(_16483_, _16485_, _16488_);
  and g_43393_(_16481_, _16488_, _16490_);
  or g_43394_(_16482_, _16487_, _16491_);
  and g_43395_(_16463_, _16470_, _16492_);
  or g_43396_(_16462_, _16469_, _16493_);
  and g_43397_(_16491_, _16493_, _16494_);
  or g_43398_(_16490_, _16492_, _16495_);
  and g_43399_(_16479_, _16494_, _16496_);
  or g_43400_(_16477_, _16495_, _16497_);
  and g_43401_(_09300_, _16461_, _16498_);
  xor g_43402_(out[228], _16480_, _16499_);
  xor g_43403_(_19134_, _16480_, _16501_);
  and g_43404_(_16281_, _16429_, _16502_);
  or g_43405_(_16279_, _16430_, _16503_);
  and g_43406_(_16287_, _16430_, _16504_);
  or g_43407_(_16286_, _16429_, _16505_);
  and g_43408_(_16503_, _16505_, _16506_);
  or g_43409_(_16502_, _16504_, _16507_);
  and g_43410_(_16501_, _16506_, _16508_);
  or g_43411_(_16499_, _16507_, _16509_);
  and g_43412_(_16482_, _16487_, _16510_);
  or g_43413_(_16481_, _16488_, _16512_);
  and g_43414_(_16509_, _16512_, _16513_);
  or g_43415_(_16508_, _16510_, _16514_);
  and g_43416_(_16497_, _16513_, _16515_);
  or g_43417_(_16496_, _16514_, _16516_);
  and g_43418_(out[229], _16498_, _16517_);
  xor g_43419_(out[229], _16498_, _16518_);
  xor g_43420_(_19123_, _16498_, _16519_);
  and g_43421_(_16306_, _16430_, _16520_);
  or g_43422_(_16305_, _16429_, _16521_);
  and g_43423_(_16299_, _16429_, _16523_);
  or g_43424_(_16298_, _16430_, _16524_);
  and g_43425_(_16521_, _16524_, _16525_);
  or g_43426_(_16520_, _16523_, _16526_);
  and g_43427_(_16518_, _16526_, _16527_);
  or g_43428_(_16519_, _16525_, _16528_);
  and g_43429_(_16499_, _16507_, _16529_);
  or g_43430_(_16501_, _16506_, _16530_);
  and g_43431_(_16528_, _16530_, _16531_);
  or g_43432_(_16527_, _16529_, _16532_);
  and g_43433_(_16516_, _16531_, _16534_);
  or g_43434_(_16515_, _16532_, _16535_);
  or g_43435_(out[230], _16517_, _16536_);
  xor g_43436_(out[230], _16517_, _16537_);
  xor g_43437_(_19112_, _16517_, _16538_);
  and g_43438_(_16325_, _16430_, _16539_);
  or g_43439_(_16323_, _16429_, _16540_);
  and g_43440_(_16317_, _16429_, _16541_);
  or g_43441_(_16318_, _16430_, _16542_);
  and g_43442_(_16540_, _16542_, _16543_);
  or g_43443_(_16539_, _16541_, _16545_);
  and g_43444_(_16537_, _16543_, _16546_);
  or g_43445_(_16538_, _16545_, _16547_);
  and g_43446_(_16519_, _16525_, _16548_);
  or g_43447_(_16518_, _16526_, _16549_);
  and g_43448_(_16547_, _16549_, _16550_);
  or g_43449_(_16546_, _16548_, _16551_);
  and g_43450_(_16535_, _16550_, _16552_);
  or g_43451_(_16534_, _16551_, _16553_);
  and g_43452_(out[231], _16536_, _16554_);
  xor g_43453_(out[231], _16536_, _16556_);
  xor g_43454_(_19101_, _16536_, _16557_);
  and g_43455_(_16437_, _16556_, _16558_);
  or g_43456_(_16436_, _16557_, _16559_);
  and g_43457_(_16538_, _16545_, _16560_);
  or g_43458_(_16537_, _16543_, _16561_);
  and g_43459_(_16559_, _16561_, _16562_);
  or g_43460_(_16558_, _16560_, _16563_);
  and g_43461_(_16553_, _16562_, _16564_);
  or g_43462_(_16552_, _16563_, _16565_);
  and g_43463_(out[232], _16554_, _16567_);
  or g_43464_(out[233], _16567_, _16568_);
  and g_43465_(out[234], _16568_, _16569_);
  xor g_43466_(out[234], _16568_, _16570_);
  xor g_43467_(_19211_, _16568_, _16571_);
  and g_43468_(_16386_, _16430_, _16572_);
  or g_43469_(_16385_, _16429_, _16573_);
  and g_43470_(_16380_, _16429_, _16574_);
  or g_43471_(_16378_, _16430_, _16575_);
  and g_43472_(_16573_, _16575_, _16576_);
  or g_43473_(_16572_, _16574_, _16578_);
  and g_43474_(_16570_, _16578_, _16579_);
  or g_43475_(_16571_, _16576_, _16580_);
  and g_43476_(_16389_, _16392_, _16581_);
  or g_43477_(_16391_, _16393_, _16582_);
  xor g_43478_(out[235], _16569_, _16583_);
  xor g_43479_(_19090_, _16569_, _16584_);
  and g_43480_(_16582_, _16583_, _16585_);
  or g_43481_(_16581_, _16584_, _16586_);
  and g_43482_(_16580_, _16586_, _16587_);
  or g_43483_(_16579_, _16585_, _16589_);
  and g_43484_(_16571_, _16576_, _16590_);
  or g_43485_(_16570_, _16578_, _16591_);
  and g_43486_(_16581_, _16584_, _16592_);
  or g_43487_(_16582_, _16583_, _16593_);
  and g_43488_(_16591_, _16593_, _16594_);
  or g_43489_(_16590_, _16592_, _16595_);
  and g_43490_(_16587_, _16594_, _16596_);
  or g_43491_(_16589_, _16595_, _16597_);
  xor g_43492_(out[232], _16554_, _16598_);
  xor g_43493_(_19189_, _16554_, _16600_);
  and g_43494_(_16367_, _16430_, _16601_);
  or g_43495_(_16366_, _16429_, _16602_);
  and g_43496_(_16360_, _16429_, _16603_);
  or g_43497_(_16361_, _16430_, _16604_);
  and g_43498_(_16602_, _16604_, _16605_);
  or g_43499_(_16601_, _16603_, _16606_);
  and g_43500_(_16598_, _16605_, _16607_);
  or g_43501_(_16600_, _16606_, _16608_);
  xor g_43502_(out[233], _16567_, _16609_);
  xor g_43503_(_19200_, _16567_, _16611_);
  and g_43504_(_16356_, _16430_, _16612_);
  or g_43505_(_16355_, _16429_, _16613_);
  and g_43506_(_16349_, _16429_, _16614_);
  or g_43507_(_16350_, _16430_, _16615_);
  and g_43508_(_16613_, _16615_, _16616_);
  or g_43509_(_16612_, _16614_, _16617_);
  and g_43510_(_16611_, _16617_, _16618_);
  or g_43511_(_16609_, _16616_, _16619_);
  and g_43512_(_16608_, _16619_, _16620_);
  or g_43513_(_16607_, _16618_, _16622_);
  and g_43514_(_16600_, _16606_, _16623_);
  or g_43515_(_16598_, _16605_, _16624_);
  and g_43516_(_16609_, _16616_, _16625_);
  or g_43517_(_16611_, _16617_, _16626_);
  and g_43518_(_16436_, _16557_, _16627_);
  or g_43519_(_16437_, _16556_, _16628_);
  and g_43520_(_16626_, _16628_, _16629_);
  or g_43521_(_16625_, _16627_, _16630_);
  and g_43522_(_16624_, _16629_, _16631_);
  or g_43523_(_16623_, _16630_, _16633_);
  and g_43524_(_16620_, _16631_, _16634_);
  or g_43525_(_16622_, _16633_, _16635_);
  and g_43526_(_16596_, _16634_, _16636_);
  or g_43527_(_16597_, _16635_, _16637_);
  and g_43528_(_16565_, _16636_, _16638_);
  or g_43529_(_16564_, _16637_, _16639_);
  and g_43530_(_16622_, _16626_, _16640_);
  or g_43531_(_16620_, _16625_, _16641_);
  and g_43532_(_16596_, _16640_, _16642_);
  or g_43533_(_16597_, _16641_, _16644_);
  and g_43534_(_16589_, _16593_, _16645_);
  or g_43535_(_16587_, _16592_, _16646_);
  and g_43536_(_16644_, _16646_, _16647_);
  or g_43537_(_16642_, _16645_, _16648_);
  and g_43538_(_16639_, _16647_, _16649_);
  or g_43539_(_16638_, _16648_, _16650_);
  and g_43540_(_16436_, _16650_, _16651_);
  or g_43541_(_16437_, _16649_, _16652_);
  and g_43542_(_16556_, _16649_, _16653_);
  or g_43543_(_16557_, _16650_, _16655_);
  and g_43544_(_16652_, _16655_, _16656_);
  or g_43545_(_16651_, _16653_, _16657_);
  and g_43546_(out[224], _16649_, _16658_);
  or g_43547_(_19156_, _16650_, _16659_);
  and g_43548_(_16443_, _16650_, _16660_);
  or g_43549_(_16442_, _16649_, _16661_);
  and g_43550_(_16659_, _16661_, _16662_);
  or g_43551_(_16658_, _16660_, _16663_);
  and g_43552_(out[240], _16662_, _16664_);
  or g_43553_(_19288_, _16663_, _16666_);
  and g_43554_(_16458_, _16649_, _16667_);
  or g_43555_(_16457_, _16650_, _16668_);
  and g_43556_(_16451_, _16650_, _16669_);
  or g_43557_(_16452_, _16649_, _16670_);
  and g_43558_(_16668_, _16670_, _16671_);
  or g_43559_(_16667_, _16669_, _16672_);
  and g_43560_(out[241], _16671_, _16673_);
  or g_43561_(_19277_, _16672_, _16674_);
  or g_43562_(out[241], out[240], _16675_);
  xor g_43563_(out[241], out[240], _16677_);
  xor g_43564_(_19277_, out[240], _16678_);
  and g_43565_(_16664_, _16674_, _16679_);
  or g_43566_(_16666_, _16673_, _16680_);
  or g_43567_(out[240], _19441_, _16681_);
  xor g_43568_(out[242], _16675_, _16682_);
  xor g_43569_(_19299_, _16675_, _16683_);
  and g_43570_(_16463_, _16649_, _16684_);
  or g_43571_(_16462_, _16650_, _16685_);
  and g_43572_(_16469_, _16650_, _16686_);
  or g_43573_(_16470_, _16649_, _16688_);
  and g_43574_(_16685_, _16688_, _16689_);
  or g_43575_(_16684_, _16686_, _16690_);
  and g_43576_(_16682_, _16690_, _16691_);
  or g_43577_(_16683_, _16689_, _16692_);
  and g_43578_(_16672_, _16677_, _16693_);
  or g_43579_(_16671_, _16678_, _16694_);
  and g_43580_(_16692_, _16694_, _16695_);
  or g_43581_(_16691_, _16693_, _16696_);
  and g_43582_(_16680_, _16695_, _16697_);
  or g_43583_(_16679_, _16696_, _16699_);
  and g_43584_(out[243], _16681_, _16700_);
  xor g_43585_(out[243], _16681_, _16701_);
  xor g_43586_(_19310_, _16681_, _16702_);
  and g_43587_(_16481_, _16649_, _16703_);
  or g_43588_(_16482_, _16650_, _16704_);
  and g_43589_(_16487_, _16650_, _16705_);
  or g_43590_(_16488_, _16649_, _16706_);
  and g_43591_(_16704_, _16706_, _16707_);
  or g_43592_(_16703_, _16705_, _16708_);
  and g_43593_(_16701_, _16707_, _16710_);
  or g_43594_(_16702_, _16708_, _16711_);
  and g_43595_(_16683_, _16689_, _16712_);
  or g_43596_(_16682_, _16690_, _16713_);
  and g_43597_(_16711_, _16713_, _16714_);
  or g_43598_(_16710_, _16712_, _16715_);
  and g_43599_(_16699_, _16714_, _16716_);
  or g_43600_(_16697_, _16715_, _16717_);
  and g_43601_(_09472_, _16681_, _16718_);
  xor g_43602_(out[244], _16700_, _16719_);
  xor g_43603_(_19266_, _16700_, _16721_);
  and g_43604_(_16506_, _16650_, _16722_);
  or g_43605_(_16507_, _16649_, _16723_);
  and g_43606_(_16499_, _16649_, _16724_);
  or g_43607_(_16501_, _16650_, _16725_);
  and g_43608_(_16723_, _16725_, _16726_);
  or g_43609_(_16722_, _16724_, _16727_);
  and g_43610_(_16721_, _16727_, _16728_);
  or g_43611_(_16719_, _16726_, _16729_);
  and g_43612_(_16702_, _16708_, _16730_);
  or g_43613_(_16701_, _16707_, _16732_);
  and g_43614_(_16729_, _16732_, _16733_);
  or g_43615_(_16728_, _16730_, _16734_);
  and g_43616_(_16717_, _16733_, _16735_);
  or g_43617_(_16716_, _16734_, _16736_);
  and g_43618_(out[245], _16718_, _16737_);
  xor g_43619_(out[245], _16718_, _16738_);
  xor g_43620_(_19255_, _16718_, _16739_);
  and g_43621_(_16518_, _16649_, _16740_);
  or g_43622_(_16519_, _16650_, _16741_);
  and g_43623_(_16525_, _16650_, _16743_);
  or g_43624_(_16526_, _16649_, _16744_);
  and g_43625_(_16741_, _16744_, _16745_);
  or g_43626_(_16740_, _16743_, _16746_);
  and g_43627_(_16738_, _16745_, _16747_);
  or g_43628_(_16739_, _16746_, _16748_);
  and g_43629_(_16719_, _16726_, _16749_);
  or g_43630_(_16721_, _16727_, _16750_);
  and g_43631_(_16748_, _16750_, _16751_);
  or g_43632_(_16747_, _16749_, _16752_);
  and g_43633_(_16736_, _16751_, _16754_);
  or g_43634_(_16735_, _16752_, _16755_);
  or g_43635_(out[246], _16737_, _16756_);
  xor g_43636_(out[246], _16737_, _16757_);
  xor g_43637_(_19244_, _16737_, _16758_);
  and g_43638_(_16543_, _16650_, _16759_);
  or g_43639_(_16545_, _16649_, _16760_);
  and g_43640_(_16538_, _16649_, _16761_);
  or g_43641_(_16537_, _16650_, _16762_);
  and g_43642_(_16760_, _16762_, _16763_);
  or g_43643_(_16759_, _16761_, _16765_);
  and g_43644_(_16757_, _16765_, _16766_);
  or g_43645_(_16758_, _16763_, _16767_);
  and g_43646_(_16739_, _16746_, _16768_);
  or g_43647_(_16738_, _16745_, _16769_);
  and g_43648_(_16767_, _16769_, _16770_);
  or g_43649_(_16766_, _16768_, _16771_);
  and g_43650_(_16755_, _16770_, _16772_);
  or g_43651_(_16754_, _16771_, _16773_);
  and g_43652_(out[247], _16756_, _16774_);
  xor g_43653_(out[247], _16756_, _16776_);
  xor g_43654_(_19233_, _16756_, _16777_);
  and g_43655_(_16656_, _16776_, _16778_);
  or g_43656_(_16657_, _16777_, _16779_);
  and g_43657_(_16758_, _16763_, _16780_);
  or g_43658_(_16757_, _16765_, _16781_);
  and g_43659_(_16779_, _16781_, _16782_);
  or g_43660_(_16778_, _16780_, _16783_);
  and g_43661_(_16773_, _16782_, _16784_);
  or g_43662_(_16772_, _16783_, _16785_);
  and g_43663_(out[248], _16774_, _16787_);
  or g_43664_(out[249], _16787_, _16788_);
  xor g_43665_(out[249], _16787_, _16789_);
  xor g_43666_(_19332_, _16787_, _16790_);
  and g_43667_(_16617_, _16650_, _16791_);
  or g_43668_(_16616_, _16649_, _16792_);
  and g_43669_(_16609_, _16649_, _16793_);
  or g_43670_(_16611_, _16650_, _16794_);
  and g_43671_(_16792_, _16794_, _16795_);
  or g_43672_(_16791_, _16793_, _16796_);
  and g_43673_(_16789_, _16795_, _16798_);
  or g_43674_(_16790_, _16796_, _16799_);
  and g_43675_(_16657_, _16777_, _16800_);
  or g_43676_(_16656_, _16776_, _16801_);
  xor g_43677_(out[248], _16774_, _16802_);
  xor g_43678_(_19321_, _16774_, _16803_);
  and g_43679_(_16606_, _16650_, _16804_);
  or g_43680_(_16605_, _16649_, _16805_);
  and g_43681_(_16598_, _16649_, _16806_);
  or g_43682_(_16600_, _16650_, _16807_);
  and g_43683_(_16805_, _16807_, _16809_);
  or g_43684_(_16804_, _16806_, _16810_);
  and g_43685_(_16803_, _16810_, _16811_);
  or g_43686_(_16802_, _16809_, _16812_);
  and g_43687_(_16801_, _16812_, _16813_);
  or g_43688_(_16800_, _16811_, _16814_);
  and g_43689_(_16799_, _16813_, _16815_);
  or g_43690_(_16798_, _16814_, _16816_);
  and g_43691_(out[250], _16788_, _16817_);
  xor g_43692_(out[250], _16788_, _16818_);
  xor g_43693_(_19343_, _16788_, _16820_);
  and g_43694_(_16576_, _16650_, _16821_);
  or g_43695_(_16578_, _16649_, _16822_);
  and g_43696_(_16570_, _16649_, _16823_);
  or g_43697_(_16571_, _16650_, _16824_);
  and g_43698_(_16822_, _16824_, _16825_);
  or g_43699_(_16821_, _16823_, _16826_);
  and g_43700_(_16818_, _16825_, _16827_);
  or g_43701_(_16820_, _16826_, _16828_);
  and g_43702_(_16581_, _16583_, _16829_);
  or g_43703_(_16582_, _16584_, _16831_);
  xor g_43704_(out[251], _16817_, _16832_);
  xor g_43705_(_19222_, _16817_, _16833_);
  and g_43706_(_16831_, _16832_, _16834_);
  or g_43707_(_16829_, _16833_, _16835_);
  and g_43708_(_16828_, _16835_, _16836_);
  or g_43709_(_16827_, _16834_, _16837_);
  and g_43710_(_16802_, _16809_, _16838_);
  or g_43711_(_16803_, _16810_, _16839_);
  and g_43712_(_16790_, _16796_, _16840_);
  or g_43713_(_16789_, _16795_, _16842_);
  and g_43714_(_16839_, _16842_, _16843_);
  or g_43715_(_16838_, _16840_, _16844_);
  and g_43716_(_16829_, _16833_, _16845_);
  or g_43717_(_16831_, _16832_, _16846_);
  and g_43718_(_16820_, _16826_, _16847_);
  or g_43719_(_16818_, _16825_, _16848_);
  and g_43720_(_16846_, _16848_, _16849_);
  or g_43721_(_16845_, _16847_, _16850_);
  and g_43722_(_16836_, _16849_, _16851_);
  or g_43723_(_16837_, _16850_, _16853_);
  and g_43724_(_16843_, _16851_, _16854_);
  or g_43725_(_16844_, _16853_, _16855_);
  and g_43726_(_16815_, _16854_, _16856_);
  or g_43727_(_16816_, _16855_, _16857_);
  and g_43728_(_16785_, _16856_, _16858_);
  or g_43729_(_16784_, _16857_, _16859_);
  and g_43730_(_16837_, _16846_, _16860_);
  or g_43731_(_16836_, _16845_, _16861_);
  and g_43732_(_16844_, _16849_, _16862_);
  or g_43733_(_16843_, _16850_, _16864_);
  and g_43734_(_16799_, _16862_, _16865_);
  or g_43735_(_16798_, _16864_, _16866_);
  and g_43736_(_16861_, _16866_, _16867_);
  or g_43737_(_16860_, _16865_, _16868_);
  and g_43738_(_16859_, _16867_, _16869_);
  or g_43739_(_16858_, _16868_, _16870_);
  and g_43740_(_16657_, _16870_, _16871_);
  or g_43741_(_16656_, _16869_, _16872_);
  and g_43742_(_16776_, _16869_, _16873_);
  or g_43743_(_16777_, _16870_, _16875_);
  and g_43744_(_16872_, _16875_, _16876_);
  or g_43745_(_16871_, _16873_, _16877_);
  and g_43746_(_15810_, _16876_, _16878_);
  or g_43747_(_15811_, _16877_, _16879_);
  xor g_43748_(out[261], _15805_, _16880_);
  xor g_43749_(_19387_, _15805_, _16881_);
  and g_43750_(_16746_, _16870_, _16882_);
  or g_43751_(_16745_, _16869_, _16883_);
  and g_43752_(_16738_, _16869_, _16884_);
  or g_43753_(_16739_, _16870_, _16886_);
  and g_43754_(_16883_, _16886_, _16887_);
  or g_43755_(_16882_, _16884_, _16888_);
  and g_43756_(_16881_, _16888_, _16889_);
  or g_43757_(_16880_, _16887_, _16890_);
  xor g_43758_(out[260], _15802_, _16891_);
  xor g_43759_(_19398_, _15802_, _16892_);
  and g_43760_(_16719_, _16869_, _16893_);
  or g_43761_(_16721_, _16870_, _16894_);
  and g_43762_(_16727_, _16870_, _16895_);
  or g_43763_(_16726_, _16869_, _16897_);
  and g_43764_(_16894_, _16897_, _16898_);
  or g_43765_(_16893_, _16895_, _16899_);
  and g_43766_(_16891_, _16898_, _16900_);
  or g_43767_(_16892_, _16899_, _16901_);
  and g_43768_(out[240], _16869_, _16902_);
  or g_43769_(_19288_, _16870_, _16903_);
  and g_43770_(_16663_, _16870_, _16904_);
  or g_43771_(_16662_, _16869_, _16905_);
  and g_43772_(_16903_, _16905_, _16906_);
  or g_43773_(_16902_, _16904_, _16908_);
  and g_43774_(out[256], _16906_, _16909_);
  or g_43775_(_19420_, _16908_, _16910_);
  and g_43776_(_16678_, _16869_, _16911_);
  or g_43777_(_16677_, _16870_, _16912_);
  and g_43778_(_16672_, _16870_, _16913_);
  or g_43779_(_16671_, _16869_, _16914_);
  and g_43780_(_16912_, _16914_, _16915_);
  or g_43781_(_16911_, _16913_, _16916_);
  and g_43782_(out[257], _16915_, _16917_);
  or g_43783_(_19409_, _16916_, _16919_);
  xor g_43784_(out[257], out[256], _16920_);
  xor g_43785_(_19409_, out[256], _16921_);
  and g_43786_(_16909_, _16919_, _16922_);
  or g_43787_(_16910_, _16917_, _16923_);
  xor g_43788_(out[258], _15800_, _16924_);
  xor g_43789_(_19431_, _15800_, _16925_);
  and g_43790_(_16683_, _16869_, _16926_);
  or g_43791_(_16682_, _16870_, _16927_);
  and g_43792_(_16690_, _16870_, _16928_);
  or g_43793_(_16689_, _16869_, _16930_);
  and g_43794_(_16927_, _16930_, _16931_);
  or g_43795_(_16926_, _16928_, _16932_);
  and g_43796_(_16924_, _16932_, _16933_);
  or g_43797_(_16925_, _16931_, _16934_);
  and g_43798_(_16916_, _16920_, _16935_);
  or g_43799_(_16915_, _16921_, _16936_);
  and g_43800_(_16934_, _16936_, _16937_);
  or g_43801_(_16933_, _16935_, _16938_);
  and g_43802_(_16923_, _16937_, _16939_);
  or g_43803_(_16922_, _16938_, _16941_);
  and g_43804_(_16701_, _16869_, _16942_);
  or g_43805_(_16702_, _16870_, _16943_);
  and g_43806_(_16708_, _16870_, _16944_);
  or g_43807_(_16707_, _16869_, _16945_);
  and g_43808_(_16943_, _16945_, _16946_);
  or g_43809_(_16942_, _16944_, _16947_);
  and g_43810_(_15803_, _16946_, _16948_);
  or g_43811_(_15804_, _16947_, _16949_);
  and g_43812_(_16925_, _16931_, _16950_);
  or g_43813_(_16924_, _16932_, _16952_);
  and g_43814_(_16949_, _16952_, _16953_);
  or g_43815_(_16948_, _16950_, _16954_);
  and g_43816_(_16941_, _16953_, _16955_);
  or g_43817_(_16939_, _16954_, _16956_);
  and g_43818_(_16892_, _16899_, _16957_);
  or g_43819_(_16891_, _16898_, _16958_);
  and g_43820_(_15804_, _16947_, _16959_);
  or g_43821_(_15803_, _16946_, _16960_);
  and g_43822_(_16958_, _16960_, _16961_);
  or g_43823_(_16957_, _16959_, _16963_);
  and g_43824_(_16956_, _16961_, _16964_);
  or g_43825_(_16955_, _16963_, _16965_);
  and g_43826_(_16901_, _16965_, _16966_);
  or g_43827_(_16900_, _16964_, _16967_);
  and g_43828_(_16890_, _16967_, _16968_);
  or g_43829_(_16889_, _16966_, _16969_);
  xor g_43830_(out[262], _15806_, _16970_);
  xor g_43831_(_19376_, _15806_, _16971_);
  and g_43832_(_16765_, _16870_, _16972_);
  or g_43833_(_16763_, _16869_, _16974_);
  and g_43834_(_16758_, _16869_, _16975_);
  or g_43835_(_16757_, _16870_, _16976_);
  and g_43836_(_16974_, _16976_, _16977_);
  or g_43837_(_16972_, _16975_, _16978_);
  and g_43838_(_16971_, _16977_, _16979_);
  or g_43839_(_16970_, _16978_, _16980_);
  and g_43840_(_16880_, _16887_, _16981_);
  or g_43841_(_16881_, _16888_, _16982_);
  and g_43842_(_16980_, _16982_, _16983_);
  or g_43843_(_16979_, _16981_, _16985_);
  and g_43844_(_16969_, _16983_, _16986_);
  or g_43845_(_16968_, _16985_, _16987_);
  and g_43846_(_15811_, _16877_, _16988_);
  or g_43847_(_15810_, _16876_, _16989_);
  and g_43848_(_16970_, _16978_, _16990_);
  or g_43849_(_16971_, _16977_, _16991_);
  and g_43850_(_16989_, _16991_, _16992_);
  or g_43851_(_16988_, _16990_, _16993_);
  and g_43852_(_16987_, _16992_, _16994_);
  or g_43853_(_16986_, _16993_, _16996_);
  and g_43854_(_16879_, _16996_, _16997_);
  or g_43855_(_16878_, _16994_, _16998_);
  and g_43856_(_16826_, _16870_, _16999_);
  or g_43857_(_16825_, _16869_, _17000_);
  and g_43858_(_16818_, _16869_, _17001_);
  or g_43859_(_16820_, _16870_, _17002_);
  and g_43860_(_17000_, _17002_, _17003_);
  or g_43861_(_16999_, _17001_, _17004_);
  and g_43862_(out[264], _15809_, _17005_);
  or g_43863_(out[265], _17005_, _17007_);
  and g_43864_(out[266], _17007_, _17008_);
  xor g_43865_(out[266], _17007_, _17009_);
  xor g_43866_(_19475_, _17007_, _17010_);
  and g_43867_(_17003_, _17009_, _17011_);
  or g_43868_(_17004_, _17010_, _17012_);
  and g_43869_(_16829_, _16832_, _17013_);
  or g_43870_(_16831_, _16833_, _17014_);
  xor g_43871_(out[267], _17008_, _17015_);
  xor g_43872_(_19354_, _17008_, _17016_);
  and g_43873_(_17014_, _17015_, _17018_);
  or g_43874_(_17013_, _17016_, _17019_);
  and g_43875_(_17012_, _17019_, _17020_);
  or g_43876_(_17011_, _17018_, _17021_);
  and g_43877_(_17013_, _17016_, _17022_);
  or g_43878_(_17014_, _17015_, _17023_);
  and g_43879_(_17004_, _17010_, _17024_);
  or g_43880_(_17003_, _17009_, _17025_);
  and g_43881_(_17023_, _17025_, _17026_);
  or g_43882_(_17022_, _17024_, _17027_);
  and g_43883_(_17020_, _17026_, _17029_);
  or g_43884_(_17021_, _17027_, _17030_);
  xor g_43885_(out[264], _15809_, _17031_);
  not g_43886_(_17031_, _17032_);
  and g_43887_(_16810_, _16870_, _17033_);
  or g_43888_(_16809_, _16869_, _17034_);
  and g_43889_(_16802_, _16869_, _17035_);
  or g_43890_(_16803_, _16870_, _17036_);
  and g_43891_(_17034_, _17036_, _17037_);
  or g_43892_(_17033_, _17035_, _17038_);
  and g_43893_(_17032_, _17038_, _17040_);
  or g_43894_(_17031_, _17037_, _17041_);
  xor g_43895_(out[265], _17005_, _17042_);
  not g_43896_(_17042_, _17043_);
  and g_43897_(_16796_, _16870_, _17044_);
  or g_43898_(_16795_, _16869_, _17045_);
  and g_43899_(_16789_, _16869_, _17046_);
  or g_43900_(_16790_, _16870_, _17047_);
  and g_43901_(_17045_, _17047_, _17048_);
  or g_43902_(_17044_, _17046_, _17049_);
  and g_43903_(_17042_, _17048_, _17051_);
  or g_43904_(_17043_, _17049_, _17052_);
  and g_43905_(_17041_, _17052_, _17053_);
  or g_43906_(_17040_, _17051_, _17054_);
  and g_43907_(_17031_, _17037_, _17055_);
  or g_43908_(_17032_, _17038_, _17056_);
  and g_43909_(_17043_, _17049_, _17057_);
  or g_43910_(_17042_, _17048_, _17058_);
  and g_43911_(_17056_, _17058_, _17059_);
  or g_43912_(_17055_, _17057_, _17060_);
  and g_43913_(_17053_, _17059_, _17062_);
  or g_43914_(_17054_, _17060_, _17063_);
  and g_43915_(_17029_, _17062_, _17064_);
  or g_43916_(_17030_, _17063_, _17065_);
  and g_43917_(_16998_, _17064_, _17066_);
  or g_43918_(_16997_, _17065_, _17067_);
  and g_43919_(_17052_, _17060_, _17068_);
  or g_43920_(_17051_, _17059_, _17069_);
  and g_43921_(_17029_, _17068_, _17070_);
  or g_43922_(_17030_, _17069_, _17071_);
  and g_43923_(_17021_, _17023_, _17073_);
  or g_43924_(_17020_, _17022_, _17074_);
  and g_43925_(_17071_, _17074_, _17075_);
  or g_43926_(_17070_, _17073_, _17076_);
  and g_43927_(_17067_, _17075_, _17077_);
  or g_43928_(_17066_, _17076_, _17078_);
  and g_43929_(_15803_, _17077_, _17079_);
  or g_43930_(_15804_, _17078_, _17080_);
  and g_43931_(_16947_, _17078_, _17081_);
  or g_43932_(_16946_, _17077_, _17082_);
  and g_43933_(_17080_, _17082_, _17084_);
  or g_43934_(_17079_, _17081_, _17085_);
  and g_43935_(_15798_, _17084_, _17086_);
  or g_43936_(_15799_, _17085_, _17087_);
  xor g_43937_(out[274], _15788_, _17088_);
  xor g_43938_(_19563_, _15788_, _17089_);
  and g_43939_(_16924_, _17077_, _17090_);
  or g_43940_(_16925_, _17078_, _17091_);
  and g_43941_(_16931_, _17078_, _17092_);
  or g_43942_(_16932_, _17077_, _17093_);
  and g_43943_(_17091_, _17093_, _17095_);
  or g_43944_(_17090_, _17092_, _17096_);
  and g_43945_(_17088_, _17095_, _17097_);
  or g_43946_(_17089_, _17096_, _17098_);
  and g_43947_(_15799_, _17085_, _17099_);
  or g_43948_(_15798_, _17084_, _17100_);
  and g_43949_(_17098_, _17100_, _17101_);
  or g_43950_(_17097_, _17099_, _17102_);
  and g_43951_(_17087_, _17102_, _17103_);
  or g_43952_(_17086_, _17101_, _17104_);
  xor g_43953_(out[273], out[272], _17106_);
  not g_43954_(_17106_, _17107_);
  and g_43955_(_16920_, _17077_, _17108_);
  or g_43956_(_16921_, _17078_, _17109_);
  and g_43957_(_16915_, _17078_, _17110_);
  or g_43958_(_16916_, _17077_, _17111_);
  and g_43959_(_17109_, _17111_, _17112_);
  or g_43960_(_17108_, _17110_, _17113_);
  and g_43961_(_17106_, _17112_, _17114_);
  or g_43962_(_17107_, _17113_, _17115_);
  and g_43963_(out[256], _17077_, _17117_);
  or g_43964_(_19420_, _17078_, _17118_);
  and g_43965_(_16908_, _17078_, _17119_);
  not g_43966_(_17119_, _17120_);
  and g_43967_(_17118_, _17120_, _17121_);
  or g_43968_(_17117_, _17119_, _17122_);
  and g_43969_(_19552_, _17122_, _17123_);
  or g_43970_(out[272], _17121_, _17124_);
  xor g_43971_(_17106_, _17112_, _17125_);
  xor g_43972_(_17107_, _17112_, _17126_);
  and g_43973_(_17124_, _17125_, _17128_);
  or g_43974_(_17123_, _17126_, _17129_);
  and g_43975_(_17115_, _17129_, _17130_);
  or g_43976_(_17114_, _17128_, _17131_);
  and g_43977_(_17089_, _17096_, _17132_);
  or g_43978_(_17088_, _17095_, _17133_);
  and g_43979_(_17087_, _17133_, _17134_);
  or g_43980_(_17086_, _17132_, _17135_);
  and g_43981_(_17131_, _17134_, _17136_);
  or g_43982_(_17130_, _17135_, _17137_);
  and g_43983_(_17104_, _17137_, _17139_);
  or g_43984_(_17103_, _17136_, _17140_);
  and g_43985_(_17010_, _17077_, _17141_);
  or g_43986_(_17009_, _17078_, _17142_);
  and g_43987_(_17003_, _17078_, _17143_);
  or g_43988_(_17004_, _17077_, _17144_);
  and g_43989_(_17142_, _17144_, _17145_);
  or g_43990_(_17141_, _17143_, _17146_);
  and g_43991_(out[280], _15794_, _17147_);
  or g_43992_(out[281], _17147_, _17148_);
  and g_43993_(out[282], _17148_, _17150_);
  xor g_43994_(out[282], _17148_, _17151_);
  xor g_43995_(_19607_, _17148_, _17152_);
  and g_43996_(_17146_, _17151_, _17153_);
  or g_43997_(_17145_, _17152_, _17154_);
  xor g_43998_(out[281], _17147_, _17155_);
  xor g_43999_(_19596_, _17147_, _17156_);
  and g_44000_(_17042_, _17077_, _17157_);
  or g_44001_(_17043_, _17078_, _17158_);
  and g_44002_(_17049_, _17078_, _17159_);
  or g_44003_(_17048_, _17077_, _17161_);
  and g_44004_(_17158_, _17161_, _17162_);
  or g_44005_(_17157_, _17159_, _17163_);
  and g_44006_(_17156_, _17163_, _17164_);
  or g_44007_(_17155_, _17162_, _17165_);
  and g_44008_(_17154_, _17165_, _17166_);
  or g_44009_(_17153_, _17164_, _17167_);
  and g_44010_(_17013_, _17015_, _17168_);
  or g_44011_(_17014_, _17016_, _17169_);
  xor g_44012_(out[283], _17150_, _17170_);
  xor g_44013_(_19486_, _17150_, _17172_);
  and g_44014_(_17169_, _17170_, _17173_);
  or g_44015_(_17168_, _17172_, _17174_);
  xor g_44016_(out[280], _15794_, _17175_);
  xor g_44017_(_19585_, _15794_, _17176_);
  and g_44018_(_17031_, _17077_, _17177_);
  or g_44019_(_17032_, _17078_, _17178_);
  and g_44020_(_17038_, _17078_, _17179_);
  or g_44021_(_17037_, _17077_, _17180_);
  and g_44022_(_17178_, _17180_, _17181_);
  or g_44023_(_17177_, _17179_, _17183_);
  and g_44024_(_17175_, _17181_, _17184_);
  or g_44025_(_17176_, _17183_, _17185_);
  and g_44026_(_17174_, _17185_, _17186_);
  or g_44027_(_17173_, _17184_, _17187_);
  and g_44028_(_17166_, _17186_, _17188_);
  or g_44029_(_17167_, _17187_, _17189_);
  and g_44030_(_17145_, _17152_, _17190_);
  or g_44031_(_17146_, _17151_, _17191_);
  and g_44032_(_17168_, _17172_, _17192_);
  or g_44033_(_17169_, _17170_, _17194_);
  and g_44034_(_17191_, _17194_, _17195_);
  or g_44035_(_17190_, _17192_, _17196_);
  and g_44036_(_17176_, _17183_, _17197_);
  or g_44037_(_17175_, _17181_, _17198_);
  and g_44038_(_17155_, _17162_, _17199_);
  or g_44039_(_17156_, _17163_, _17200_);
  and g_44040_(_17198_, _17200_, _17201_);
  or g_44041_(_17197_, _17199_, _17202_);
  and g_44042_(_17195_, _17201_, _17203_);
  or g_44043_(_17196_, _17202_, _17205_);
  and g_44044_(_17188_, _17203_, _17206_);
  or g_44045_(_17189_, _17205_, _17207_);
  xor g_44046_(out[278], _15792_, _17208_);
  xor g_44047_(_19508_, _15792_, _17209_);
  or g_44048_(_16971_, _17078_, _17210_);
  or g_44049_(_16978_, _17077_, _17211_);
  and g_44050_(_17210_, _17211_, _17212_);
  not g_44051_(_17212_, _17213_);
  and g_44052_(_17208_, _17212_, _17214_);
  or g_44053_(_17209_, _17213_, _17216_);
  or g_44054_(_15811_, _17078_, _17217_);
  or g_44055_(_16876_, _17077_, _17218_);
  and g_44056_(_17217_, _17218_, _17219_);
  not g_44057_(_17219_, _17220_);
  and g_44058_(_15797_, _17220_, _17221_);
  or g_44059_(_15795_, _17219_, _17222_);
  and g_44060_(_17216_, _17222_, _17223_);
  or g_44061_(_17214_, _17221_, _17224_);
  and g_44062_(_15795_, _17219_, _17225_);
  or g_44063_(_15797_, _17220_, _17227_);
  and g_44064_(_17209_, _17213_, _17228_);
  or g_44065_(_17208_, _17212_, _17229_);
  and g_44066_(_17227_, _17229_, _17230_);
  or g_44067_(_17225_, _17228_, _17231_);
  and g_44068_(_17223_, _17230_, _17232_);
  or g_44069_(_17224_, _17231_, _17233_);
  xor g_44070_(out[277], _15791_, _17234_);
  xor g_44071_(_19519_, _15791_, _17235_);
  and g_44072_(_16880_, _17077_, _17236_);
  or g_44073_(_16881_, _17078_, _17238_);
  and g_44074_(_16888_, _17078_, _17239_);
  or g_44075_(_16887_, _17077_, _17240_);
  and g_44076_(_17238_, _17240_, _17241_);
  or g_44077_(_17236_, _17239_, _17242_);
  and g_44078_(_17235_, _17242_, _17243_);
  or g_44079_(_17234_, _17241_, _17244_);
  xor g_44080_(out[276], _15790_, _17245_);
  xor g_44081_(_19530_, _15790_, _17246_);
  and g_44082_(_16891_, _17077_, _17247_);
  or g_44083_(_16892_, _17078_, _17249_);
  and g_44084_(_16899_, _17078_, _17250_);
  or g_44085_(_16898_, _17077_, _17251_);
  and g_44086_(_17249_, _17251_, _17252_);
  or g_44087_(_17247_, _17250_, _17253_);
  and g_44088_(_17246_, _17253_, _17254_);
  or g_44089_(_17245_, _17252_, _17255_);
  and g_44090_(_17244_, _17255_, _17256_);
  or g_44091_(_17243_, _17254_, _17257_);
  and g_44092_(_17234_, _17241_, _17258_);
  or g_44093_(_17235_, _17242_, _17260_);
  and g_44094_(_17245_, _17252_, _17261_);
  or g_44095_(_17246_, _17253_, _17262_);
  and g_44096_(_17260_, _17262_, _17263_);
  or g_44097_(_17258_, _17261_, _17264_);
  and g_44098_(_17256_, _17263_, _17265_);
  or g_44099_(_17257_, _17264_, _17266_);
  and g_44100_(_17206_, _17265_, _17267_);
  or g_44101_(_17207_, _17266_, _17268_);
  and g_44102_(_17232_, _17267_, _17269_);
  or g_44103_(_17233_, _17268_, _17271_);
  and g_44104_(_17140_, _17269_, _17272_);
  or g_44105_(_17139_, _17271_, _17273_);
  and g_44106_(_17224_, _17227_, _17274_);
  or g_44107_(_17223_, _17225_, _17275_);
  and g_44108_(_17257_, _17260_, _17276_);
  or g_44109_(_17256_, _17258_, _17277_);
  and g_44110_(_17230_, _17276_, _17278_);
  or g_44111_(_17231_, _17277_, _17279_);
  and g_44112_(_17275_, _17279_, _17280_);
  or g_44113_(_17274_, _17278_, _17282_);
  and g_44114_(_17206_, _17282_, _17283_);
  or g_44115_(_17207_, _17280_, _17284_);
  and g_44116_(_17166_, _17202_, _17285_);
  or g_44117_(_17167_, _17201_, _17286_);
  and g_44118_(_17195_, _17286_, _17287_);
  or g_44119_(_17196_, _17285_, _17288_);
  and g_44120_(_17174_, _17288_, _17289_);
  or g_44121_(_17173_, _17287_, _17290_);
  and g_44122_(_17284_, _17290_, _17291_);
  or g_44123_(_17283_, _17289_, _17293_);
  and g_44124_(_17273_, _17291_, _17294_);
  or g_44125_(_17272_, _17293_, _17295_);
  and g_44126_(out[272], _17121_, _17296_);
  or g_44127_(_19552_, _17122_, _17297_);
  and g_44128_(_17101_, _17134_, _17298_);
  or g_44129_(_17102_, _17135_, _17299_);
  and g_44130_(_17297_, _17298_, _17300_);
  or g_44131_(_17296_, _17299_, _17301_);
  and g_44132_(_17128_, _17300_, _17302_);
  or g_44133_(_17129_, _17301_, _17304_);
  and g_44134_(_17269_, _17302_, _17305_);
  or g_44135_(_17271_, _17304_, _17306_);
  and g_44136_(_17295_, _17306_, _17307_);
  or g_44137_(_17294_, _17305_, _17308_);
  or g_44138_(_15797_, _17308_, _17309_);
  or g_44139_(_17219_, _17307_, _17310_);
  and g_44140_(_17309_, _17310_, _17311_);
  not g_44141_(_17311_, _17312_);
  and g_44142_(_15786_, _17311_, _17313_);
  or g_44143_(_15787_, _17312_, _17315_);
  xor g_44144_(out[294], _15782_, _17316_);
  xor g_44145_(_19640_, _15782_, _17317_);
  or g_44146_(_17209_, _17308_, _17318_);
  or g_44147_(_17212_, _17307_, _17319_);
  and g_44148_(_17318_, _17319_, _17320_);
  not g_44149_(_17320_, _17321_);
  and g_44150_(_17317_, _17321_, _17322_);
  or g_44151_(_17316_, _17320_, _17323_);
  xor g_44152_(out[293], _15781_, _17324_);
  xor g_44153_(_19651_, _15781_, _17326_);
  and g_44154_(_17234_, _17307_, _17327_);
  or g_44155_(_17235_, _17308_, _17328_);
  and g_44156_(_17242_, _17308_, _17329_);
  or g_44157_(_17241_, _17307_, _17330_);
  and g_44158_(_17328_, _17330_, _17331_);
  or g_44159_(_17327_, _17329_, _17332_);
  and g_44160_(_17326_, _17332_, _17333_);
  or g_44161_(_17324_, _17331_, _17334_);
  and g_44162_(out[272], _17307_, _17335_);
  or g_44163_(_19552_, _17308_, _17337_);
  and g_44164_(_17122_, _17308_, _17338_);
  or g_44165_(_17121_, _17307_, _17339_);
  and g_44166_(_17337_, _17339_, _17340_);
  or g_44167_(_17335_, _17338_, _17341_);
  and g_44168_(out[288], _17340_, _17342_);
  or g_44169_(_18573_, _17341_, _17343_);
  and g_44170_(_17107_, _17307_, _17344_);
  or g_44171_(_17106_, _17308_, _17345_);
  and g_44172_(_17112_, _17308_, _17346_);
  or g_44173_(_17113_, _17307_, _17348_);
  and g_44174_(_17345_, _17348_, _17349_);
  or g_44175_(_17344_, _17346_, _17350_);
  and g_44176_(out[289], _17349_, _17351_);
  or g_44177_(_19673_, _17350_, _17352_);
  xor g_44178_(out[288], out[289], _17353_);
  xor g_44179_(_18573_, out[289], _17354_);
  and g_44180_(_17342_, _17352_, _17355_);
  or g_44181_(_17343_, _17351_, _17356_);
  and g_44182_(_17088_, _17307_, _17357_);
  or g_44183_(_17089_, _17308_, _17359_);
  and g_44184_(_17096_, _17308_, _17360_);
  or g_44185_(_17095_, _17307_, _17361_);
  and g_44186_(_17359_, _17361_, _17362_);
  or g_44187_(_17357_, _17360_, _17363_);
  and g_44188_(_15778_, _17362_, _17364_);
  or g_44189_(_15779_, _17363_, _17365_);
  and g_44190_(_17350_, _17353_, _17366_);
  or g_44191_(_17349_, _17354_, _17367_);
  and g_44192_(_17365_, _17367_, _17368_);
  or g_44193_(_17364_, _17366_, _17370_);
  and g_44194_(_17356_, _17368_, _17371_);
  or g_44195_(_17355_, _17370_, _17372_);
  xor g_44196_(out[291], _15777_, _17373_);
  not g_44197_(_17373_, _17374_);
  and g_44198_(_15798_, _17307_, _17375_);
  and g_44199_(_17085_, _17308_, _17376_);
  or g_44200_(_17375_, _17376_, _17377_);
  not g_44201_(_17377_, _17378_);
  and g_44202_(_17373_, _17378_, _17379_);
  or g_44203_(_17374_, _17377_, _17381_);
  and g_44204_(_15779_, _17363_, _17382_);
  or g_44205_(_15778_, _17362_, _17383_);
  and g_44206_(_17381_, _17383_, _17384_);
  or g_44207_(_17379_, _17382_, _17385_);
  and g_44208_(_17372_, _17384_, _17386_);
  or g_44209_(_17371_, _17385_, _17387_);
  xor g_44210_(out[292], _15780_, _17388_);
  xor g_44211_(_19662_, _15780_, _17389_);
  and g_44212_(_17246_, _17307_, _17390_);
  or g_44213_(_17245_, _17308_, _17392_);
  and g_44214_(_17252_, _17308_, _17393_);
  or g_44215_(_17253_, _17307_, _17394_);
  and g_44216_(_17392_, _17394_, _17395_);
  or g_44217_(_17390_, _17393_, _17396_);
  and g_44218_(_17389_, _17395_, _17397_);
  or g_44219_(_17388_, _17396_, _17398_);
  and g_44220_(_17374_, _17377_, _17399_);
  or g_44221_(_17373_, _17378_, _17400_);
  and g_44222_(_17398_, _17400_, _17401_);
  or g_44223_(_17397_, _17399_, _17403_);
  and g_44224_(_17387_, _17401_, _17404_);
  or g_44225_(_17386_, _17403_, _17405_);
  and g_44226_(_17324_, _17331_, _17406_);
  or g_44227_(_17326_, _17332_, _17407_);
  and g_44228_(_17388_, _17396_, _17408_);
  or g_44229_(_17389_, _17395_, _17409_);
  and g_44230_(_17407_, _17409_, _17410_);
  or g_44231_(_17406_, _17408_, _17411_);
  and g_44232_(_17405_, _17410_, _17412_);
  or g_44233_(_17404_, _17411_, _17414_);
  and g_44234_(_17334_, _17414_, _17415_);
  or g_44235_(_17333_, _17412_, _17416_);
  and g_44236_(_17323_, _17416_, _17417_);
  or g_44237_(_17322_, _17415_, _17418_);
  and g_44238_(_15787_, _17312_, _17419_);
  or g_44239_(_15786_, _17311_, _17420_);
  and g_44240_(_17316_, _17320_, _17421_);
  or g_44241_(_17317_, _17321_, _17422_);
  and g_44242_(_17420_, _17422_, _17423_);
  or g_44243_(_17419_, _17421_, _17425_);
  and g_44244_(_17418_, _17423_, _17426_);
  or g_44245_(_17417_, _17425_, _17427_);
  and g_44246_(_17315_, _17427_, _17428_);
  or g_44247_(_17313_, _17426_, _17429_);
  or g_44248_(_17151_, _17308_, _17430_);
  or g_44249_(_17145_, _17307_, _17431_);
  and g_44250_(_17430_, _17431_, _17432_);
  not g_44251_(_17432_, _17433_);
  and g_44252_(out[296], _15784_, _17434_);
  or g_44253_(out[297], _17434_, _17436_);
  and g_44254_(out[298], _17436_, _17437_);
  xor g_44255_(out[298], _17436_, _17438_);
  not g_44256_(_17438_, _17439_);
  and g_44257_(_17433_, _17438_, _17440_);
  or g_44258_(_17432_, _17439_, _17441_);
  and g_44259_(_17432_, _17439_, _17442_);
  and g_44260_(_17168_, _17170_, _17443_);
  not g_44261_(_17443_, _17444_);
  xor g_44262_(out[299], _17437_, _17445_);
  not g_44263_(_17445_, _17447_);
  and g_44264_(_17444_, _17445_, _17448_);
  or g_44265_(_17443_, _17447_, _17449_);
  and g_44266_(_17443_, _17447_, _17450_);
  or g_44267_(_17444_, _17445_, _17451_);
  or g_44268_(_17442_, _17448_, _17452_);
  or g_44269_(_17440_, _17450_, _17453_);
  or g_44270_(_17452_, _17453_, _17454_);
  xor g_44271_(out[297], _17434_, _17455_);
  xor g_44272_(_19717_, _17434_, _17456_);
  or g_44273_(_17156_, _17308_, _17458_);
  or g_44274_(_17162_, _17307_, _17459_);
  and g_44275_(_17458_, _17459_, _17460_);
  or g_44276_(_17455_, _17460_, _17461_);
  xor g_44277_(out[296], _15784_, _17462_);
  not g_44278_(_17462_, _17463_);
  or g_44279_(_17175_, _17308_, _17464_);
  or g_44280_(_17183_, _17307_, _17465_);
  and g_44281_(_17464_, _17465_, _17466_);
  or g_44282_(_17463_, _17466_, _17467_);
  and g_44283_(_17461_, _17467_, _17469_);
  and g_44284_(_17455_, _17460_, _17470_);
  xor g_44285_(_17455_, _17460_, _17471_);
  xor g_44286_(_17456_, _17460_, _17472_);
  xor g_44287_(_17462_, _17466_, _17473_);
  or g_44288_(_17454_, _17473_, _17474_);
  not g_44289_(_17474_, _17475_);
  and g_44290_(_17471_, _17475_, _17476_);
  or g_44291_(_17472_, _17474_, _17477_);
  and g_44292_(_17429_, _17476_, _17478_);
  or g_44293_(_17428_, _17477_, _17480_);
  or g_44294_(_17469_, _17470_, _17481_);
  or g_44295_(_17454_, _17481_, _17482_);
  not g_44296_(_17482_, _17483_);
  and g_44297_(_17441_, _17449_, _17484_);
  or g_44298_(_17440_, _17448_, _17485_);
  and g_44299_(_17451_, _17485_, _17486_);
  or g_44300_(_17450_, _17484_, _17487_);
  and g_44301_(_17482_, _17487_, _17488_);
  or g_44302_(_17483_, _17486_, _17489_);
  and g_44303_(_17480_, _17488_, _17491_);
  or g_44304_(_17478_, _17489_, _17492_);
  or g_44305_(_15779_, _17492_, _17493_);
  or g_44306_(_17362_, _17491_, _17494_);
  and g_44307_(_17493_, _17494_, _17495_);
  not g_44308_(_17495_, _17496_);
  and g_44309_(_15773_, _17495_, _17497_);
  xor g_44310_(out[307], _15765_, _17498_);
  xor g_44311_(_19816_, _15765_, _17499_);
  and g_44312_(_17373_, _17491_, _17500_);
  and g_44313_(_17377_, _17492_, _17502_);
  or g_44314_(_17500_, _17502_, _17503_);
  and g_44315_(_17499_, _17503_, _17504_);
  or g_44316_(_17497_, _17504_, _17505_);
  or g_44317_(_17499_, _17503_, _17506_);
  xor g_44318_(_15773_, _17495_, _17507_);
  xor g_44319_(_15775_, _17495_, _17508_);
  xor g_44320_(_17499_, _17503_, _17509_);
  xor g_44321_(_17498_, _17503_, _17510_);
  and g_44322_(_17507_, _17509_, _17511_);
  or g_44323_(_17508_, _17510_, _17513_);
  xor g_44324_(out[304], out[305], _17514_);
  not g_44325_(_17514_, _17515_);
  or g_44326_(_17354_, _17492_, _17516_);
  not g_44327_(_17516_, _17517_);
  and g_44328_(_17349_, _17492_, _17518_);
  not g_44329_(_17518_, _17519_);
  and g_44330_(_17516_, _17519_, _17520_);
  or g_44331_(_17517_, _17518_, _17521_);
  and g_44332_(_17514_, _17520_, _17522_);
  or g_44333_(_17515_, _17521_, _17524_);
  and g_44334_(_17340_, _17492_, _17525_);
  not g_44335_(_17525_, _17526_);
  or g_44336_(out[288], _17492_, _17527_);
  not g_44337_(_17527_, _17528_);
  and g_44338_(_17526_, _17527_, _17529_);
  or g_44339_(_17525_, _17528_, _17530_);
  and g_44340_(_18562_, _17529_, _17531_);
  or g_44341_(out[304], _17530_, _17532_);
  xor g_44342_(_17514_, _17520_, _17533_);
  xor g_44343_(_17515_, _17520_, _17535_);
  and g_44344_(_17532_, _17533_, _17536_);
  or g_44345_(_17531_, _17535_, _17537_);
  and g_44346_(_17524_, _17537_, _17538_);
  or g_44347_(_17522_, _17536_, _17539_);
  and g_44348_(_17511_, _17539_, _17540_);
  or g_44349_(_17513_, _17538_, _17541_);
  and g_44350_(_17505_, _17506_, _17542_);
  not g_44351_(_17542_, _17543_);
  and g_44352_(_17541_, _17543_, _17544_);
  or g_44353_(_17540_, _17542_, _17546_);
  or g_44354_(out[313], _15771_, _17547_);
  xor g_44355_(out[313], _15771_, _17548_);
  not g_44356_(_17548_, _17549_);
  or g_44357_(_17456_, _17492_, _17550_);
  or g_44358_(_17460_, _17491_, _17551_);
  and g_44359_(_17550_, _17551_, _17552_);
  and g_44360_(_17548_, _17552_, _17553_);
  not g_44361_(_17553_, _17554_);
  or g_44362_(_17462_, _17492_, _17555_);
  or g_44363_(_17466_, _17491_, _17557_);
  and g_44364_(_17555_, _17557_, _17558_);
  or g_44365_(_15772_, _17558_, _17559_);
  not g_44366_(_17559_, _17560_);
  and g_44367_(_17554_, _17559_, _17561_);
  or g_44368_(_17553_, _17560_, _17562_);
  and g_44369_(out[314], _17547_, _17563_);
  xor g_44370_(out[314], _17547_, _17564_);
  xor g_44371_(_19849_, _17547_, _17565_);
  or g_44372_(_17438_, _17492_, _17566_);
  or g_44373_(_17432_, _17491_, _17568_);
  and g_44374_(_17566_, _17568_, _17569_);
  or g_44375_(_17565_, _17569_, _17570_);
  or g_44376_(_17548_, _17552_, _17571_);
  and g_44377_(_17570_, _17571_, _17572_);
  not g_44378_(_17572_, _17573_);
  and g_44379_(_17561_, _17572_, _17574_);
  or g_44380_(_17562_, _17573_, _17575_);
  and g_44381_(_17565_, _17569_, _17576_);
  and g_44382_(_17443_, _17445_, _17577_);
  not g_44383_(_17577_, _17579_);
  xor g_44384_(out[315], _17563_, _17580_);
  not g_44385_(_17580_, _17581_);
  and g_44386_(_17577_, _17581_, _17582_);
  or g_44387_(_17576_, _17582_, _17583_);
  and g_44388_(_17579_, _17580_, _17584_);
  not g_44389_(_17584_, _17585_);
  and g_44390_(_15772_, _17558_, _17586_);
  or g_44391_(_17584_, _17586_, _17587_);
  or g_44392_(_17583_, _17587_, _17588_);
  not g_44393_(_17588_, _17590_);
  and g_44394_(_17574_, _17590_, _17591_);
  or g_44395_(_17575_, _17588_, _17592_);
  xor g_44396_(out[311], _15769_, _17593_);
  not g_44397_(_17593_, _17594_);
  or g_44398_(_15787_, _17492_, _17595_);
  or g_44399_(_17311_, _17491_, _17596_);
  and g_44400_(_17595_, _17596_, _17597_);
  or g_44401_(_17593_, _17597_, _17598_);
  not g_44402_(_17598_, _17599_);
  xor g_44403_(out[310], _15768_, _17601_);
  not g_44404_(_17601_, _17602_);
  or g_44405_(_17317_, _17492_, _17603_);
  or g_44406_(_17320_, _17491_, _17604_);
  and g_44407_(_17603_, _17604_, _17605_);
  not g_44408_(_17605_, _17606_);
  and g_44409_(_17601_, _17605_, _17607_);
  not g_44410_(_17607_, _17608_);
  and g_44411_(_17598_, _17608_, _17609_);
  or g_44412_(_17599_, _17607_, _17610_);
  and g_44413_(_17593_, _17597_, _17612_);
  not g_44414_(_17612_, _17613_);
  xor g_44415_(_17593_, _17597_, _17614_);
  xor g_44416_(_17594_, _17597_, _17615_);
  xor g_44417_(_17601_, _17605_, _17616_);
  xor g_44418_(_17602_, _17605_, _17617_);
  and g_44419_(_17614_, _17616_, _17618_);
  or g_44420_(_17615_, _17617_, _17619_);
  xor g_44421_(out[309], _15767_, _17620_);
  xor g_44422_(_19783_, _15767_, _17621_);
  and g_44423_(_17324_, _17491_, _17623_);
  or g_44424_(_17326_, _17492_, _17624_);
  and g_44425_(_17332_, _17492_, _17625_);
  or g_44426_(_17331_, _17491_, _17626_);
  and g_44427_(_17624_, _17626_, _17627_);
  or g_44428_(_17623_, _17625_, _17628_);
  and g_44429_(_17621_, _17628_, _17629_);
  or g_44430_(_17620_, _17627_, _17630_);
  xor g_44431_(out[308], _15766_, _17631_);
  xor g_44432_(_19772_, _15766_, _17632_);
  and g_44433_(_17396_, _17492_, _17634_);
  or g_44434_(_17395_, _17491_, _17635_);
  and g_44435_(_17389_, _17491_, _17636_);
  or g_44436_(_17388_, _17492_, _17637_);
  and g_44437_(_17635_, _17637_, _17638_);
  or g_44438_(_17634_, _17636_, _17639_);
  and g_44439_(_17632_, _17638_, _17640_);
  or g_44440_(_17631_, _17639_, _17641_);
  and g_44441_(_17630_, _17641_, _17642_);
  or g_44442_(_17629_, _17640_, _17643_);
  and g_44443_(_17620_, _17627_, _17645_);
  or g_44444_(_17621_, _17628_, _17646_);
  or g_44445_(_17632_, _17638_, _17647_);
  not g_44446_(_17647_, _17648_);
  and g_44447_(_17646_, _17647_, _17649_);
  and g_44448_(_17642_, _17649_, _17650_);
  or g_44449_(_17643_, _17645_, _17651_);
  or g_44450_(_17619_, _17648_, _17652_);
  and g_44451_(_17618_, _17650_, _17653_);
  or g_44452_(_17651_, _17652_, _17654_);
  and g_44453_(_17591_, _17653_, _17656_);
  or g_44454_(_17592_, _17654_, _17657_);
  and g_44455_(_17546_, _17656_, _17658_);
  or g_44456_(_17544_, _17657_, _17659_);
  and g_44457_(_17618_, _17643_, _17660_);
  or g_44458_(_17619_, _17642_, _17661_);
  and g_44459_(_17646_, _17660_, _17662_);
  or g_44460_(_17645_, _17661_, _17663_);
  and g_44461_(_17610_, _17613_, _17664_);
  or g_44462_(_17609_, _17612_, _17665_);
  and g_44463_(_17663_, _17665_, _17667_);
  or g_44464_(_17662_, _17664_, _17668_);
  and g_44465_(_17591_, _17668_, _17669_);
  or g_44466_(_17592_, _17667_, _17670_);
  or g_44467_(_17553_, _17586_, _17671_);
  and g_44468_(_17572_, _17671_, _17672_);
  or g_44469_(_17583_, _17672_, _17673_);
  not g_44470_(_17673_, _17674_);
  and g_44471_(_17585_, _17673_, _17675_);
  or g_44472_(_17584_, _17674_, _17676_);
  and g_44473_(_17670_, _17676_, _17678_);
  or g_44474_(_17669_, _17675_, _17679_);
  and g_44475_(_17659_, _17678_, _17680_);
  or g_44476_(_17658_, _17679_, _17681_);
  and g_44477_(out[304], _17530_, _17682_);
  or g_44478_(_18562_, _17529_, _17683_);
  and g_44479_(_17511_, _17536_, _17684_);
  not g_44480_(_17684_, _17685_);
  and g_44481_(_17656_, _17684_, _17686_);
  or g_44482_(_17657_, _17685_, _17687_);
  and g_44483_(_17683_, _17686_, _17689_);
  or g_44484_(_17682_, _17687_, _17690_);
  and g_44485_(_17681_, _17690_, _17691_);
  or g_44486_(_17680_, _17689_, _17692_);
  or g_44487_(_17558_, _17691_, _17693_);
  and g_44488_(_15772_, _17691_, _17694_);
  not g_44489_(_17694_, _17695_);
  and g_44490_(_17693_, _17695_, _17696_);
  or g_44491_(_15716_, _15718_, _17697_);
  and g_44492_(_17577_, _17580_, _17698_);
  xor g_44493_(_17697_, _17698_, _17700_);
  and g_44494_(_15651_, _15757_, _17701_);
  or g_44495_(_15652_, _15758_, _17702_);
  and g_44496_(_15659_, _15758_, _17703_);
  or g_44497_(_15658_, _15757_, _17704_);
  and g_44498_(_17702_, _17704_, _17705_);
  or g_44499_(_17701_, _17703_, _17706_);
  and g_44500_(_17496_, _17692_, _17707_);
  or g_44501_(_17495_, _17691_, _17708_);
  and g_44502_(_15773_, _17691_, _17709_);
  or g_44503_(_15775_, _17692_, _17711_);
  and g_44504_(_17708_, _17711_, _17712_);
  or g_44505_(_17707_, _17709_, _17713_);
  or g_44506_(_17706_, _17712_, _17714_);
  or g_44507_(_15709_, _15758_, _17715_);
  not g_44508_(_17715_, _17716_);
  and g_44509_(_15712_, _15758_, _17717_);
  or g_44510_(_17716_, _17717_, _17718_);
  and g_44511_(_17564_, _17691_, _17719_);
  and g_44512_(_17569_, _17692_, _17720_);
  or g_44513_(_17719_, _17720_, _17722_);
  xor g_44514_(_17718_, _17722_, _17723_);
  or g_44515_(_21114_, _15758_, _17724_);
  or g_44516_(_15635_, _15757_, _17725_);
  and g_44517_(_17724_, _17725_, _17726_);
  or g_44518_(_17529_, _17691_, _17727_);
  or g_44519_(out[304], _17692_, _17728_);
  and g_44520_(_17727_, _17728_, _17729_);
  xor g_44521_(_17726_, _17729_, _17730_);
  and g_44522_(_15733_, _15757_, _17731_);
  or g_44523_(_15734_, _15758_, _17733_);
  and g_44524_(_15737_, _15758_, _17734_);
  not g_44525_(_17734_, _17735_);
  and g_44526_(_17733_, _17735_, _17736_);
  or g_44527_(_17731_, _17734_, _17737_);
  or g_44528_(_17552_, _17691_, _17738_);
  not g_44529_(_17738_, _17739_);
  and g_44530_(_17548_, _17691_, _17740_);
  or g_44531_(_17549_, _17692_, _17741_);
  and g_44532_(_17738_, _17741_, _17742_);
  or g_44533_(_17739_, _17740_, _17744_);
  or g_44534_(_17737_, _17742_, _17745_);
  or g_44535_(_15648_, _15758_, _17746_);
  not g_44536_(_17746_, _17747_);
  and g_44537_(_15645_, _15758_, _17748_);
  or g_44538_(_15644_, _15757_, _17749_);
  and g_44539_(_17746_, _17749_, _17750_);
  or g_44540_(_17747_, _17748_, _17751_);
  and g_44541_(_17514_, _17691_, _17752_);
  not g_44542_(_17752_, _17753_);
  and g_44543_(_17521_, _17692_, _17755_);
  or g_44544_(_17520_, _17691_, _17756_);
  and g_44545_(_17753_, _17756_, _17757_);
  or g_44546_(_17752_, _17755_, _17758_);
  or g_44547_(_17751_, _17757_, _17759_);
  or g_44548_(_15624_, _15758_, _17760_);
  not g_44549_(_17760_, _17761_);
  and g_44550_(_15627_, _15758_, _17762_);
  not g_44551_(_17762_, _17763_);
  and g_44552_(_17760_, _17763_, _17764_);
  or g_44553_(_17761_, _17762_, _17766_);
  or g_44554_(_17638_, _17691_, _17767_);
  not g_44555_(_17767_, _17768_);
  and g_44556_(_17632_, _17691_, _17769_);
  not g_44557_(_17769_, _17770_);
  and g_44558_(_17767_, _17770_, _17771_);
  or g_44559_(_17768_, _17769_, _17772_);
  or g_44560_(_17764_, _17772_, _17773_);
  or g_44561_(_17705_, _17713_, _17774_);
  or g_44562_(_15603_, _15758_, _17775_);
  not g_44563_(_17775_, _17777_);
  and g_44564_(_15610_, _15758_, _17778_);
  or g_44565_(_15608_, _15757_, _17779_);
  and g_44566_(_17775_, _17779_, _17780_);
  or g_44567_(_17777_, _17778_, _17781_);
  and g_44568_(_17606_, _17692_, _17782_);
  or g_44569_(_17605_, _17691_, _17783_);
  and g_44570_(_17601_, _17691_, _17784_);
  not g_44571_(_17784_, _17785_);
  and g_44572_(_17783_, _17785_, _17786_);
  or g_44573_(_17782_, _17784_, _17788_);
  or g_44574_(_17780_, _17788_, _17789_);
  or g_44575_(_17736_, _17744_, _17790_);
  or g_44576_(_15669_, _15758_, _17791_);
  not g_44577_(_17791_, _17792_);
  and g_44578_(_15672_, _15758_, _17793_);
  or g_44579_(_17792_, _17793_, _17794_);
  and g_44580_(_17503_, _17692_, _17795_);
  and g_44581_(_17498_, _17691_, _17796_);
  or g_44582_(_17795_, _17796_, _17797_);
  or g_44583_(_17766_, _17771_, _17799_);
  or g_44584_(_17781_, _17786_, _17800_);
  and g_44585_(_15621_, _15758_, _17801_);
  or g_44586_(_15619_, _15757_, _17802_);
  and g_44587_(_15614_, _15757_, _17803_);
  or g_44588_(_15613_, _15758_, _17804_);
  and g_44589_(_17802_, _17804_, _17805_);
  or g_44590_(_17801_, _17803_, _17806_);
  and g_44591_(_17628_, _17692_, _17807_);
  or g_44592_(_17627_, _17691_, _17808_);
  and g_44593_(_17620_, _17691_, _17810_);
  or g_44594_(_17621_, _17692_, _17811_);
  and g_44595_(_17808_, _17811_, _17812_);
  or g_44596_(_17807_, _17810_, _17813_);
  or g_44597_(_17806_, _17813_, _17814_);
  or g_44598_(_13848_, _15758_, _17815_);
  not g_44599_(_17815_, _17816_);
  and g_44600_(_15599_, _15758_, _17817_);
  or g_44601_(_17816_, _17817_, _17818_);
  or g_44602_(_17597_, _17691_, _17819_);
  not g_44603_(_17819_, _17821_);
  and g_44604_(_17593_, _17691_, _17822_);
  or g_44605_(_17821_, _17822_, _17823_);
  xor g_44606_(_17818_, _17823_, _17824_);
  or g_44607_(_17805_, _17812_, _17825_);
  or g_44608_(_17750_, _17758_, _17826_);
  and g_44609_(_17790_, _17799_, _17827_);
  xor g_44610_(_15762_, _17696_, _17828_);
  and g_44611_(_17714_, _17789_, _17829_);
  and g_44612_(_17773_, _17800_, _17830_);
  xor g_44613_(_17794_, _17797_, _17832_);
  and g_44614_(_17829_, _17832_, _17833_);
  and g_44615_(_17830_, _17833_, _17834_);
  and g_44616_(_17745_, _17825_, _17835_);
  and g_44617_(_17774_, _17814_, _17836_);
  and g_44618_(_17835_, _17836_, _17837_);
  and g_44619_(_17723_, _17837_, _17838_);
  and g_44620_(_17834_, _17838_, _17839_);
  and g_44621_(_17827_, _17828_, _17840_);
  and g_44622_(_17700_, _17826_, _17841_);
  and g_44623_(_17730_, _17841_, _17843_);
  and g_44624_(_17759_, _17824_, _17844_);
  and g_44625_(_17843_, _17844_, _17845_);
  and g_44626_(_17840_, _17845_, _17846_);
  and g_44627_(_17839_, _17846_, _17847_);
  or g_44628_(_13837_, _17847_, _17848_);
  and g_44629_(_13837_, _17847_, _17849_);
  xor g_44630_(_13836_, _17847_, _17850_);
  xor g_44631_(_10622_, _17850_, _17851_);
  xor g_44632_(_10621_, _17850_, _17852_);
  and g_44633_(_24416_, _17852_, _17854_);
  not g_44634_(_17854_, _17855_);
  and g_44635_(_24415_, _17851_, _17856_);
  xor g_44636_(_24415_, _17851_, _17857_);
  xor g_44637_(_20522_, _17857_, out[320]);
  or g_44638_(_10621_, _17849_, _17858_);
  and g_44639_(_17848_, _17858_, _17859_);
  or g_44640_(_20522_, _17856_, _17860_);
  and g_44641_(_17855_, _17860_, _17861_);
  and g_44642_(_17859_, _17861_, out[322]);
  xor g_44643_(_17859_, _17861_, out[321]);
  czero b_0_(out[334]);
  czero b_1_(out[333]);
  czero b_2_(out[332]);
  czero b_3_(out[331]);
  czero b_4_(out[330]);
  czero b_5_(out[329]);
  czero b_6_(out[328]);
  czero b_7_(out[327]);
  czero b_8_(out[326]);
  czero b_9_(out[325]);
  czero b_10_(out[326]);
  buf b_11_(set1[42], out[202]);
  buf b_12_(set1[67], out[227]);
  buf b_13_(set1[52], out[212]);
  buf b_14_(set2[15], out[15]);
  czero b_15_(out[335]);
  buf b_16_(set1[44], out[204]);
  buf b_17_(set1[80], out[240]);
  buf b_18_(set1[82], out[242]);
  buf b_19_(set2[10], out[10]);
  buf b_20_(set1[144], out[304]);
  buf b_21_(set1[50], out[210]);
  buf b_22_(set2[141], out[141]);
  buf b_23_(set2[42], out[42]);
  buf b_24_(set1[99], out[259]);
  buf b_25_(set1[17], out[177]);
  buf b_26_(set1[138], out[298]);
  buf b_27_(set1[30], out[190]);
  buf b_28_(set1[111], out[271]);
  buf b_29_(set1[130], out[290]);
  buf b_30_(set1[108], out[268]);
  buf b_31_(set2[126], out[126]);
  buf b_32_(set1[73], out[233]);
  buf b_33_(set2[36], out[36]);
  buf b_34_(set1[31], out[191]);
  buf b_35_(set1[95], out[255]);
  buf b_36_(set1[110], out[270]);
  buf b_37_(set1[76], out[236]);
  buf b_38_(set1[153], out[313]);
  buf b_39_(set2[155], out[155]);
  buf b_40_(set1[148], out[308]);
  buf b_41_(set2[79], out[79]);
  buf b_42_(set1[53], out[213]);
  buf b_43_(set1[77], out[237]);
  buf b_44_(set2[11], out[11]);
  czero b_45_(out[330]);
  buf b_46_(set2[8], out[8]);
  czero b_47_(out[335]);
  buf b_48_(set1[119], out[279]);
  buf b_49_(set1[102], out[262]);
  buf b_50_(set1[121], out[281]);
  buf b_51_(set2[110], out[110]);
  buf b_52_(set2[76], out[76]);
  buf b_53_(set1[114], out[274]);
  buf b_54_(set1[147], out[307]);
  buf b_55_(set2[24], out[24]);
  buf b_56_(set2[14], out[14]);
  buf b_57_(set1[3], out[163]);
  buf b_58_(set1[132], out[292]);
  buf b_59_(set1[113], out[273]);
  buf b_60_(set1[51], out[211]);
  buf b_61_(set2[105], out[105]);
  buf b_62_(set2[46], out[46]);
  buf b_63_(set2[56], out[56]);
  buf b_64_(set2[64], out[64]);
  buf b_65_(set2[39], out[39]);
  buf b_66_(set1[5], out[165]);
  czero b_67_(out[333]);
  buf b_68_(set1[70], out[230]);
  buf b_69_(set2[80], out[80]);
  buf b_70_(set1[140], out[300]);
  czero b_71_(out[323]);
  buf b_72_(set2[5], out[5]);
  buf b_73_(set2[147], out[147]);
  buf b_74_(set2[33], out[33]);
  buf b_75_(set1[21], out[181]);
  buf b_76_(set1[12], out[172]);
  buf b_77_(set2[124], out[124]);
  buf b_78_(set2[21], out[21]);
  buf b_79_(set2[43], out[43]);
  buf b_80_(set2[99], out[99]);
  buf b_81_(set2[145], out[145]);
  buf b_82_(set1[117], out[277]);
  buf b_83_(set1[124], out[284]);
  buf b_84_(set1[9], out[169]);
  buf b_85_(set2[35], out[35]);
  buf b_86_(set1[136], out[296]);
  buf b_87_(set2[152], out[152]);
  buf b_88_(set2[72], out[72]);
  buf b_89_(set1[101], out[261]);
  buf b_90_(set1[29], out[189]);
  buf b_91_(set2[116], out[116]);
  buf b_92_(set1[156], out[316]);
  buf b_93_(set2[101], out[101]);
  buf b_94_(set2[134], out[134]);
  buf b_95_(set1[109], out[269]);
  buf b_96_(set1[149], out[309]);
  buf b_97_(set1[134], out[294]);
  buf b_98_(set2[143], out[143]);
  buf b_99_(set2[19], out[19]);
  buf b_100_(set2[55], out[55]);
  czero b_101_(out[331]);
  buf b_102_(set2[13], out[13]);
  buf b_103_(set1[98], out[258]);
  buf b_104_(set1[48], out[208]);
  buf b_105_(set1[152], out[312]);
  buf b_106_(set1[56], out[216]);
  buf b_107_(set1[115], out[275]);
  buf b_108_(set1[157], out[317]);
  buf b_109_(set1[125], out[285]);
  buf b_110_(set2[130], out[130]);
  buf b_111_(set2[29], out[29]);
  buf b_112_(set2[107], out[107]);
  buf b_113_(set2[25], out[25]);
  buf b_114_(set1[69], out[229]);
  buf b_115_(set2[104], out[104]);
  buf b_116_(set1[66], out[226]);
  buf b_117_(set1[154], out[314]);
  buf b_118_(set1[61], out[221]);
  buf b_119_(set1[47], out[207]);
  buf b_120_(set1[0], out[160]);
  buf b_121_(set1[8], out[168]);
  buf b_122_(set2[142], out[142]);
  buf b_123_(set2[133], out[133]);
  buf b_124_(set2[61], out[61]);
  czero b_125_(out[325]);
  buf b_126_(set2[157], out[157]);
  buf b_127_(set1[46], out[206]);
  buf b_128_(set2[154], out[154]);
  buf b_129_(set2[81], out[81]);
  buf b_130_(set2[90], out[90]);
  buf b_131_(set2[122], out[122]);
  buf b_132_(set2[75], out[75]);
  buf b_133_(set2[118], out[118]);
  buf b_134_(set1[116], out[276]);
  buf b_135_(set2[26], out[26]);
  buf b_136_(set2[7], out[7]);
  buf b_137_(set1[71], out[231]);
  buf b_138_(set2[149], out[149]);
  buf b_139_(set1[16], out[176]);
  czero b_140_(out[334]);
  buf b_141_(set2[139], out[139]);
  buf b_142_(set2[103], out[103]);
  buf b_143_(set2[112], out[112]);
  buf b_144_(set1[120], out[280]);
  buf b_145_(set1[62], out[222]);
  buf b_146_(set1[93], out[253]);
  buf b_147_(set2[114], out[114]);
  buf b_148_(set1[100], out[260]);
  buf b_149_(set1[13], out[173]);
  buf b_150_(set1[6], out[166]);
  buf b_151_(set1[55], out[215]);
  czero b_152_(_26838_);
  buf b_153_(set1[25], out[185]);
  buf b_154_(set2[121], out[121]);
  buf b_155_(set1[10], out[170]);
  buf b_156_(set2[88], out[88]);
  buf b_157_(set2[70], out[70]);
  buf b_158_(set2[94], out[94]);
  czero b_159_(out[327]);
  buf b_160_(set2[20], out[20]);
  buf b_161_(set2[97], out[97]);
  buf b_162_(set1[90], out[250]);
  buf b_163_(set2[138], out[138]);
  buf b_164_(set1[38], out[198]);
  buf b_165_(set2[41], out[41]);
  buf b_166_(set1[107], out[267]);
  buf b_167_(set2[95], out[95]);
  buf b_168_(set1[143], out[303]);
  buf b_169_(set1[43], out[203]);
  buf b_170_(set1[106], out[266]);
  buf b_171_(set1[84], out[244]);
  buf b_172_(set2[6], out[6]);
  buf b_173_(set1[129], out[289]);
  czero b_174_(out[328]);
  buf b_175_(set1[81], out[241]);
  czero b_176_(out[324]);
  buf b_177_(set2[48], out[48]);
  buf b_178_(set1[20], out[180]);
  buf b_179_(set2[127], out[127]);
  buf b_180_(set1[64], out[224]);
  buf b_181_(set1[28], out[188]);
  buf b_182_(set2[45], out[45]);
  buf b_183_(set2[12], out[12]);
  buf b_184_(set2[84], out[84]);
  buf b_185_(set2[17], out[17]);
  buf b_186_(set1[141], out[301]);
  buf b_187_(set2[60], out[60]);
  buf b_188_(set2[63], out[63]);
  buf b_189_(set1[27], out[187]);
  buf b_190_(set2[120], out[120]);
  buf b_191_(set2[93], out[93]);
  buf b_192_(set1[105], out[265]);
  buf b_193_(set2[73], out[73]);
  buf b_194_(set1[54], out[214]);
  buf b_195_(set2[38], out[38]);
  buf b_196_(set2[54], out[54]);
  buf b_197_(set1[49], out[209]);
  buf b_198_(set2[58], out[58]);
  buf b_199_(set1[45], out[205]);
  buf b_200_(set2[52], out[52]);
  buf b_201_(set1[72], out[232]);
  buf b_202_(set2[22], out[22]);
  buf b_203_(set2[40], out[40]);
  buf b_204_(set2[111], out[111]);
  buf b_205_(set2[4], out[4]);
  buf b_206_(set2[66], out[66]);
  buf b_207_(set1[127], out[287]);
  buf b_208_(set2[146], out[146]);
  buf b_209_(set2[159], out[159]);
  buf b_210_(set1[59], out[219]);
  buf b_211_(set2[16], out[16]);
  buf b_212_(set1[7], out[167]);
  buf b_213_(set2[28], out[28]);
  buf b_214_(set2[69], out[69]);
  buf b_215_(set2[108], out[108]);
  buf b_216_(set2[87], out[87]);
  buf b_217_(set2[91], out[91]);
  buf b_218_(set1[126], out[286]);
  czero b_219_(out[329]);
  buf b_220_(set1[135], out[295]);
  buf b_221_(set1[40], out[200]);
  buf b_222_(set1[35], out[195]);
  buf b_223_(set2[119], out[119]);
  buf b_224_(set2[131], out[131]);
  buf b_225_(set1[92], out[252]);
  buf b_226_(set2[100], out[100]);
  buf b_227_(set2[77], out[77]);
  buf b_228_(set2[78], out[78]);
  buf b_229_(set2[115], out[115]);
  buf b_230_(set1[131], out[291]);
  buf b_231_(set1[128], out[288]);
  buf b_232_(set2[1], out[1]);
  buf b_233_(set2[86], out[86]);
  buf b_234_(set2[123], out[123]);
  buf b_235_(set1[96], out[256]);
  buf b_236_(set2[27], out[27]);
  buf b_237_(set2[50], out[50]);
  buf b_238_(set1[85], out[245]);
  buf b_239_(set1[151], out[311]);
  buf b_240_(set1[133], out[293]);
  buf b_241_(set2[62], out[62]);
  buf b_242_(set1[88], out[248]);
  buf b_243_(set2[125], out[125]);
  buf b_244_(set1[34], out[194]);
  buf b_245_(set2[37], out[37]);
  buf b_246_(set2[82], out[82]);
  buf b_247_(set1[63], out[223]);
  buf b_248_(set1[112], out[272]);
  buf b_249_(set1[37], out[197]);
  buf b_250_(set1[94], out[254]);
  buf b_251_(set2[51], out[51]);
  buf b_252_(set2[140], out[140]);
  buf b_253_(set2[117], out[117]);
  buf b_254_(set2[98], out[98]);
  buf b_255_(set2[67], out[67]);
  buf b_256_(set2[0], out[0]);
  buf b_257_(set1[33], out[193]);
  buf b_258_(set1[139], out[299]);
  buf b_259_(set1[158], out[318]);
  buf b_260_(set2[9], out[9]);
  buf b_261_(set1[65], out[225]);
  buf b_262_(set1[103], out[263]);
  buf b_263_(set1[1], out[161]);
  buf b_264_(set1[68], out[228]);
  buf b_265_(set1[123], out[283]);
  buf b_266_(set2[30], out[30]);
  buf b_267_(set1[145], out[305]);
  buf b_268_(set2[59], out[59]);
  buf b_269_(set1[41], out[201]);
  buf b_270_(set2[49], out[49]);
  buf b_271_(set2[83], out[83]);
  buf b_272_(set2[135], out[135]);
  buf b_273_(set2[68], out[68]);
  buf b_274_(set1[32], out[192]);
  buf b_275_(set2[132], out[132]);
  buf b_276_(set2[148], out[148]);
  buf b_277_(set2[129], out[129]);
  buf b_278_(set1[79], out[239]);
  buf b_279_(set1[18], out[178]);
  buf b_280_(set1[104], out[264]);
  buf b_281_(set1[97], out[257]);
  buf b_282_(set1[150], out[310]);
  buf b_283_(set1[2], out[162]);
  buf b_284_(set1[159], out[319]);
  buf b_285_(set1[89], out[249]);
  buf b_286_(set1[137], out[297]);
  buf b_287_(set2[137], out[137]);
  buf b_288_(set2[156], out[156]);
  buf b_289_(set2[158], out[158]);
  buf b_290_(set2[71], out[71]);
  buf b_291_(set2[106], out[106]);
  buf b_292_(set1[22], out[182]);
  buf b_293_(set2[18], out[18]);
  buf b_294_(set1[75], out[235]);
  buf b_295_(set2[102], out[102]);
  buf b_296_(set1[86], out[246]);
  buf b_297_(set1[122], out[282]);
  buf b_298_(set1[36], out[196]);
  buf b_299_(set2[74], out[74]);
  buf b_300_(set1[24], out[184]);
  buf b_301_(set1[142], out[302]);
  buf b_302_(set2[89], out[89]);
  buf b_303_(set2[96], out[96]);
  buf b_304_(set2[92], out[92]);
  buf b_305_(set2[32], out[32]);
  buf b_306_(set1[26], out[186]);
  buf b_307_(set1[87], out[247]);
  buf b_308_(set2[113], out[113]);
  buf b_309_(set1[58], out[218]);
  buf b_310_(set1[19], out[179]);
  buf b_311_(set2[3], out[3]);
  buf b_312_(set2[31], out[31]);
  buf b_313_(set2[144], out[144]);
  buf b_314_(set2[85], out[85]);
  buf b_315_(set2[65], out[65]);
  buf b_316_(set2[23], out[23]);
  czero b_317_(_26839_);
  buf b_318_(set1[4], out[164]);
  buf b_319_(set2[53], out[53]);
  buf b_320_(set2[57], out[57]);
  buf b_321_(set1[23], out[183]);
  czero b_322_(out[332]);
  buf b_323_(set2[128], out[128]);
  buf b_324_(set1[57], out[217]);
  buf b_325_(set2[44], out[44]);
  buf b_326_(set2[150], out[150]);
  buf b_327_(set1[155], out[315]);
  buf b_328_(set2[136], out[136]);
  buf b_329_(set2[47], out[47]);
  buf b_330_(set2[109], out[109]);
  buf b_331_(set1[14], out[174]);
  buf b_332_(set1[15], out[175]);
  buf b_333_(set1[91], out[251]);
  buf b_334_(set1[60], out[220]);
  buf b_335_(set2[34], out[34]);
  buf b_336_(set1[74], out[234]);
  buf b_337_(set1[118], out[278]);
  buf b_338_(set1[11], out[171]);
  czero b_339_(out[324]);
  buf b_340_(set1[39], out[199]);
  buf b_341_(set2[2], out[2]);
  buf b_342_(set1[83], out[243]);
  buf b_343_(set1[78], out[238]);
  buf b_344_(set1[146], out[306]);
  buf b_345_(set2[151], out[151]);
  buf b_346_(set2[153], out[153]);

endmodule
