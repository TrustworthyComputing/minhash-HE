module min_hash(
  input wire [1199:0] set1,
  input wire [1199:0] set2,
  output wire [2415:0] out
);
  wire [15:0] set1_unflattened[75];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  assign set1_unflattened[50] = set1[815:800];
  assign set1_unflattened[51] = set1[831:816];
  assign set1_unflattened[52] = set1[847:832];
  assign set1_unflattened[53] = set1[863:848];
  assign set1_unflattened[54] = set1[879:864];
  assign set1_unflattened[55] = set1[895:880];
  assign set1_unflattened[56] = set1[911:896];
  assign set1_unflattened[57] = set1[927:912];
  assign set1_unflattened[58] = set1[943:928];
  assign set1_unflattened[59] = set1[959:944];
  assign set1_unflattened[60] = set1[975:960];
  assign set1_unflattened[61] = set1[991:976];
  assign set1_unflattened[62] = set1[1007:992];
  assign set1_unflattened[63] = set1[1023:1008];
  assign set1_unflattened[64] = set1[1039:1024];
  assign set1_unflattened[65] = set1[1055:1040];
  assign set1_unflattened[66] = set1[1071:1056];
  assign set1_unflattened[67] = set1[1087:1072];
  assign set1_unflattened[68] = set1[1103:1088];
  assign set1_unflattened[69] = set1[1119:1104];
  assign set1_unflattened[70] = set1[1135:1120];
  assign set1_unflattened[71] = set1[1151:1136];
  assign set1_unflattened[72] = set1[1167:1152];
  assign set1_unflattened[73] = set1[1183:1168];
  assign set1_unflattened[74] = set1[1199:1184];
  wire [15:0] set2_unflattened[75];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  assign set2_unflattened[50] = set2[815:800];
  assign set2_unflattened[51] = set2[831:816];
  assign set2_unflattened[52] = set2[847:832];
  assign set2_unflattened[53] = set2[863:848];
  assign set2_unflattened[54] = set2[879:864];
  assign set2_unflattened[55] = set2[895:880];
  assign set2_unflattened[56] = set2[911:896];
  assign set2_unflattened[57] = set2[927:912];
  assign set2_unflattened[58] = set2[943:928];
  assign set2_unflattened[59] = set2[959:944];
  assign set2_unflattened[60] = set2[975:960];
  assign set2_unflattened[61] = set2[991:976];
  assign set2_unflattened[62] = set2[1007:992];
  assign set2_unflattened[63] = set2[1023:1008];
  assign set2_unflattened[64] = set2[1039:1024];
  assign set2_unflattened[65] = set2[1055:1040];
  assign set2_unflattened[66] = set2[1071:1056];
  assign set2_unflattened[67] = set2[1087:1072];
  assign set2_unflattened[68] = set2[1103:1088];
  assign set2_unflattened[69] = set2[1119:1104];
  assign set2_unflattened[70] = set2[1135:1120];
  assign set2_unflattened[71] = set2[1151:1136];
  assign set2_unflattened[72] = set2[1167:1152];
  assign set2_unflattened[73] = set2[1183:1168];
  assign set2_unflattened[74] = set2[1199:1184];
  wire [15:0] array_index_130213;
  wire [15:0] array_index_130214;
  wire [11:0] add_130221;
  wire [11:0] add_130224;
  wire [15:0] array_index_130229;
  wire [15:0] array_index_130232;
  wire [10:0] add_130236;
  wire [10:0] add_130239;
  wire [11:0] add_130255;
  wire [11:0] sel_130257;
  wire [11:0] add_130260;
  wire [11:0] sel_130262;
  wire [15:0] array_index_130277;
  wire [15:0] array_index_130280;
  wire [8:0] add_130284;
  wire [8:0] add_130287;
  wire [10:0] add_130290;
  wire [11:0] sel_130293;
  wire [10:0] add_130295;
  wire [11:0] sel_130298;
  wire [11:0] add_130315;
  wire [11:0] sel_130317;
  wire [11:0] add_130320;
  wire [11:0] sel_130322;
  wire [15:0] array_index_130343;
  wire [15:0] array_index_130346;
  wire [10:0] add_130350;
  wire [10:0] add_130352;
  wire [8:0] add_130354;
  wire [11:0] sel_130357;
  wire [8:0] add_130359;
  wire [11:0] sel_130362;
  wire [10:0] add_130364;
  wire [11:0] sel_130367;
  wire [10:0] add_130369;
  wire [11:0] sel_130372;
  wire [11:0] add_130393;
  wire [11:0] sel_130395;
  wire [11:0] add_130398;
  wire [11:0] sel_130400;
  wire [15:0] array_index_130427;
  wire [15:0] array_index_130430;
  wire [10:0] add_130434;
  wire [10:0] add_130436;
  wire [10:0] add_130438;
  wire [11:0] sel_130440;
  wire [10:0] add_130442;
  wire [11:0] sel_130444;
  wire [8:0] add_130446;
  wire [11:0] sel_130449;
  wire [8:0] add_130451;
  wire [11:0] sel_130454;
  wire [10:0] add_130456;
  wire [11:0] sel_130459;
  wire [10:0] add_130461;
  wire [11:0] sel_130464;
  wire [11:0] add_130489;
  wire [11:0] sel_130491;
  wire [11:0] add_130494;
  wire [11:0] sel_130496;
  wire [15:0] array_index_130527;
  wire [15:0] array_index_130530;
  wire [10:0] add_130534;
  wire [11:0] sel_130536;
  wire [10:0] add_130538;
  wire [11:0] sel_130540;
  wire [10:0] add_130542;
  wire [11:0] sel_130544;
  wire [10:0] add_130546;
  wire [11:0] sel_130548;
  wire [8:0] add_130550;
  wire [11:0] sel_130553;
  wire [8:0] add_130555;
  wire [11:0] sel_130558;
  wire [10:0] add_130560;
  wire [11:0] sel_130563;
  wire [10:0] add_130565;
  wire [11:0] sel_130568;
  wire [11:0] add_130593;
  wire [11:0] sel_130595;
  wire [11:0] add_130598;
  wire [11:0] sel_130600;
  wire [15:0] array_index_130629;
  wire [15:0] array_index_130632;
  wire [10:0] add_130636;
  wire [11:0] sel_130638;
  wire [10:0] add_130640;
  wire [11:0] sel_130642;
  wire [10:0] add_130644;
  wire [11:0] sel_130646;
  wire [10:0] add_130648;
  wire [11:0] sel_130650;
  wire [8:0] add_130652;
  wire [11:0] sel_130655;
  wire [8:0] add_130657;
  wire [11:0] sel_130660;
  wire [10:0] add_130662;
  wire [11:0] sel_130665;
  wire [10:0] add_130667;
  wire [11:0] sel_130670;
  wire [11:0] add_130695;
  wire [11:0] sel_130697;
  wire [11:0] add_130700;
  wire [11:0] sel_130702;
  wire [15:0] array_index_130731;
  wire [15:0] array_index_130734;
  wire [10:0] add_130738;
  wire [11:0] sel_130740;
  wire [10:0] add_130742;
  wire [11:0] sel_130744;
  wire [10:0] add_130746;
  wire [11:0] sel_130748;
  wire [10:0] add_130750;
  wire [11:0] sel_130752;
  wire [8:0] add_130754;
  wire [11:0] sel_130757;
  wire [8:0] add_130759;
  wire [11:0] sel_130762;
  wire [10:0] add_130764;
  wire [11:0] sel_130767;
  wire [10:0] add_130769;
  wire [11:0] sel_130772;
  wire [11:0] add_130797;
  wire [11:0] sel_130799;
  wire [11:0] add_130802;
  wire [11:0] sel_130804;
  wire [15:0] array_index_130833;
  wire [15:0] array_index_130836;
  wire [10:0] add_130840;
  wire [11:0] sel_130842;
  wire [10:0] add_130844;
  wire [11:0] sel_130846;
  wire [10:0] add_130848;
  wire [11:0] sel_130850;
  wire [10:0] add_130852;
  wire [11:0] sel_130854;
  wire [8:0] add_130856;
  wire [11:0] sel_130859;
  wire [8:0] add_130861;
  wire [11:0] sel_130864;
  wire [10:0] add_130866;
  wire [11:0] sel_130869;
  wire [10:0] add_130871;
  wire [11:0] sel_130874;
  wire [11:0] add_130899;
  wire [11:0] sel_130901;
  wire [11:0] add_130904;
  wire [11:0] sel_130906;
  wire [15:0] array_index_130935;
  wire [15:0] array_index_130938;
  wire [10:0] add_130942;
  wire [11:0] sel_130944;
  wire [10:0] add_130946;
  wire [11:0] sel_130948;
  wire [10:0] add_130950;
  wire [11:0] sel_130952;
  wire [10:0] add_130954;
  wire [11:0] sel_130956;
  wire [8:0] add_130958;
  wire [11:0] sel_130961;
  wire [8:0] add_130963;
  wire [11:0] sel_130966;
  wire [10:0] add_130968;
  wire [11:0] sel_130971;
  wire [10:0] add_130973;
  wire [11:0] sel_130976;
  wire [11:0] add_131001;
  wire [11:0] sel_131003;
  wire [11:0] add_131006;
  wire [11:0] sel_131008;
  wire [15:0] array_index_131037;
  wire [15:0] array_index_131040;
  wire [10:0] add_131044;
  wire [11:0] sel_131046;
  wire [10:0] add_131048;
  wire [11:0] sel_131050;
  wire [10:0] add_131052;
  wire [11:0] sel_131054;
  wire [10:0] add_131056;
  wire [11:0] sel_131058;
  wire [8:0] add_131060;
  wire [11:0] sel_131063;
  wire [8:0] add_131065;
  wire [11:0] sel_131068;
  wire [10:0] add_131070;
  wire [11:0] sel_131073;
  wire [10:0] add_131075;
  wire [11:0] sel_131078;
  wire [11:0] add_131103;
  wire [11:0] sel_131105;
  wire [11:0] add_131108;
  wire [11:0] sel_131110;
  wire [15:0] array_index_131139;
  wire [15:0] array_index_131142;
  wire [10:0] add_131146;
  wire [11:0] sel_131148;
  wire [10:0] add_131150;
  wire [11:0] sel_131152;
  wire [10:0] add_131154;
  wire [11:0] sel_131156;
  wire [10:0] add_131158;
  wire [11:0] sel_131160;
  wire [8:0] add_131162;
  wire [11:0] sel_131165;
  wire [8:0] add_131167;
  wire [11:0] sel_131170;
  wire [10:0] add_131172;
  wire [11:0] sel_131175;
  wire [10:0] add_131177;
  wire [11:0] sel_131180;
  wire [11:0] add_131205;
  wire [11:0] sel_131207;
  wire [11:0] add_131210;
  wire [11:0] sel_131212;
  wire [15:0] array_index_131241;
  wire [15:0] array_index_131244;
  wire [10:0] add_131248;
  wire [11:0] sel_131250;
  wire [10:0] add_131252;
  wire [11:0] sel_131254;
  wire [10:0] add_131256;
  wire [11:0] sel_131258;
  wire [10:0] add_131260;
  wire [11:0] sel_131262;
  wire [8:0] add_131264;
  wire [11:0] sel_131267;
  wire [8:0] add_131269;
  wire [11:0] sel_131272;
  wire [10:0] add_131274;
  wire [11:0] sel_131277;
  wire [10:0] add_131279;
  wire [11:0] sel_131282;
  wire [11:0] add_131307;
  wire [11:0] sel_131309;
  wire [11:0] add_131312;
  wire [11:0] sel_131314;
  wire [15:0] array_index_131343;
  wire [15:0] array_index_131346;
  wire [10:0] add_131350;
  wire [11:0] sel_131352;
  wire [10:0] add_131354;
  wire [11:0] sel_131356;
  wire [10:0] add_131358;
  wire [11:0] sel_131360;
  wire [10:0] add_131362;
  wire [11:0] sel_131364;
  wire [8:0] add_131366;
  wire [11:0] sel_131369;
  wire [8:0] add_131371;
  wire [11:0] sel_131374;
  wire [10:0] add_131376;
  wire [11:0] sel_131379;
  wire [10:0] add_131381;
  wire [11:0] sel_131384;
  wire [11:0] add_131409;
  wire [11:0] sel_131411;
  wire [11:0] add_131414;
  wire [11:0] sel_131416;
  wire [15:0] array_index_131445;
  wire [15:0] array_index_131448;
  wire [10:0] add_131452;
  wire [11:0] sel_131454;
  wire [10:0] add_131456;
  wire [11:0] sel_131458;
  wire [10:0] add_131460;
  wire [11:0] sel_131462;
  wire [10:0] add_131464;
  wire [11:0] sel_131466;
  wire [8:0] add_131468;
  wire [11:0] sel_131471;
  wire [8:0] add_131473;
  wire [11:0] sel_131476;
  wire [10:0] add_131478;
  wire [11:0] sel_131481;
  wire [10:0] add_131483;
  wire [11:0] sel_131486;
  wire [11:0] add_131511;
  wire [11:0] sel_131513;
  wire [11:0] add_131516;
  wire [11:0] sel_131518;
  wire [15:0] array_index_131547;
  wire [15:0] array_index_131550;
  wire [10:0] add_131554;
  wire [11:0] sel_131556;
  wire [10:0] add_131558;
  wire [11:0] sel_131560;
  wire [10:0] add_131562;
  wire [11:0] sel_131564;
  wire [10:0] add_131566;
  wire [11:0] sel_131568;
  wire [8:0] add_131570;
  wire [11:0] sel_131573;
  wire [8:0] add_131575;
  wire [11:0] sel_131578;
  wire [10:0] add_131580;
  wire [11:0] sel_131583;
  wire [10:0] add_131585;
  wire [11:0] sel_131588;
  wire [11:0] add_131613;
  wire [11:0] sel_131615;
  wire [11:0] add_131618;
  wire [11:0] sel_131620;
  wire [15:0] array_index_131649;
  wire [15:0] array_index_131652;
  wire [10:0] add_131656;
  wire [11:0] sel_131658;
  wire [10:0] add_131660;
  wire [11:0] sel_131662;
  wire [10:0] add_131664;
  wire [11:0] sel_131666;
  wire [10:0] add_131668;
  wire [11:0] sel_131670;
  wire [8:0] add_131672;
  wire [11:0] sel_131675;
  wire [8:0] add_131677;
  wire [11:0] sel_131680;
  wire [10:0] add_131682;
  wire [11:0] sel_131685;
  wire [10:0] add_131687;
  wire [11:0] sel_131690;
  wire [11:0] add_131715;
  wire [11:0] sel_131717;
  wire [11:0] add_131720;
  wire [11:0] sel_131722;
  wire [15:0] array_index_131751;
  wire [15:0] array_index_131754;
  wire [10:0] add_131758;
  wire [11:0] sel_131760;
  wire [10:0] add_131762;
  wire [11:0] sel_131764;
  wire [10:0] add_131766;
  wire [11:0] sel_131768;
  wire [10:0] add_131770;
  wire [11:0] sel_131772;
  wire [8:0] add_131774;
  wire [11:0] sel_131777;
  wire [8:0] add_131779;
  wire [11:0] sel_131782;
  wire [10:0] add_131784;
  wire [11:0] sel_131787;
  wire [10:0] add_131789;
  wire [11:0] sel_131792;
  wire [11:0] add_131817;
  wire [11:0] sel_131819;
  wire [11:0] add_131822;
  wire [11:0] sel_131824;
  wire [15:0] array_index_131853;
  wire [15:0] array_index_131856;
  wire [10:0] add_131860;
  wire [11:0] sel_131862;
  wire [10:0] add_131864;
  wire [11:0] sel_131866;
  wire [10:0] add_131868;
  wire [11:0] sel_131870;
  wire [10:0] add_131872;
  wire [11:0] sel_131874;
  wire [8:0] add_131876;
  wire [11:0] sel_131879;
  wire [8:0] add_131881;
  wire [11:0] sel_131884;
  wire [10:0] add_131886;
  wire [11:0] sel_131889;
  wire [10:0] add_131891;
  wire [11:0] sel_131894;
  wire [11:0] add_131919;
  wire [11:0] sel_131921;
  wire [11:0] add_131924;
  wire [11:0] sel_131926;
  wire [15:0] array_index_131955;
  wire [15:0] array_index_131958;
  wire [10:0] add_131962;
  wire [11:0] sel_131964;
  wire [10:0] add_131966;
  wire [11:0] sel_131968;
  wire [10:0] add_131970;
  wire [11:0] sel_131972;
  wire [10:0] add_131974;
  wire [11:0] sel_131976;
  wire [8:0] add_131978;
  wire [11:0] sel_131981;
  wire [8:0] add_131983;
  wire [11:0] sel_131986;
  wire [10:0] add_131988;
  wire [11:0] sel_131991;
  wire [10:0] add_131993;
  wire [11:0] sel_131996;
  wire [11:0] add_132021;
  wire [11:0] sel_132023;
  wire [11:0] add_132026;
  wire [11:0] sel_132028;
  wire [15:0] array_index_132057;
  wire [15:0] array_index_132060;
  wire [10:0] add_132064;
  wire [11:0] sel_132066;
  wire [10:0] add_132068;
  wire [11:0] sel_132070;
  wire [10:0] add_132072;
  wire [11:0] sel_132074;
  wire [10:0] add_132076;
  wire [11:0] sel_132078;
  wire [8:0] add_132080;
  wire [11:0] sel_132083;
  wire [8:0] add_132085;
  wire [11:0] sel_132088;
  wire [10:0] add_132090;
  wire [11:0] sel_132093;
  wire [10:0] add_132095;
  wire [11:0] sel_132098;
  wire [11:0] add_132123;
  wire [11:0] sel_132125;
  wire [11:0] add_132128;
  wire [11:0] sel_132130;
  wire [15:0] array_index_132159;
  wire [15:0] array_index_132162;
  wire [10:0] add_132166;
  wire [11:0] sel_132168;
  wire [10:0] add_132170;
  wire [11:0] sel_132172;
  wire [10:0] add_132174;
  wire [11:0] sel_132176;
  wire [10:0] add_132178;
  wire [11:0] sel_132180;
  wire [8:0] add_132182;
  wire [11:0] sel_132185;
  wire [8:0] add_132187;
  wire [11:0] sel_132190;
  wire [10:0] add_132192;
  wire [11:0] sel_132195;
  wire [10:0] add_132197;
  wire [11:0] sel_132200;
  wire [11:0] add_132225;
  wire [11:0] sel_132227;
  wire [11:0] add_132230;
  wire [11:0] sel_132232;
  wire [15:0] array_index_132261;
  wire [15:0] array_index_132264;
  wire [10:0] add_132268;
  wire [11:0] sel_132270;
  wire [10:0] add_132272;
  wire [11:0] sel_132274;
  wire [10:0] add_132276;
  wire [11:0] sel_132278;
  wire [10:0] add_132280;
  wire [11:0] sel_132282;
  wire [8:0] add_132284;
  wire [11:0] sel_132287;
  wire [8:0] add_132289;
  wire [11:0] sel_132292;
  wire [10:0] add_132294;
  wire [11:0] sel_132297;
  wire [10:0] add_132299;
  wire [11:0] sel_132302;
  wire [11:0] add_132327;
  wire [11:0] sel_132329;
  wire [11:0] add_132332;
  wire [11:0] sel_132334;
  wire [15:0] array_index_132363;
  wire [15:0] array_index_132366;
  wire [10:0] add_132370;
  wire [11:0] sel_132372;
  wire [10:0] add_132374;
  wire [11:0] sel_132376;
  wire [10:0] add_132378;
  wire [11:0] sel_132380;
  wire [10:0] add_132382;
  wire [11:0] sel_132384;
  wire [8:0] add_132386;
  wire [11:0] sel_132389;
  wire [8:0] add_132391;
  wire [11:0] sel_132394;
  wire [10:0] add_132396;
  wire [11:0] sel_132399;
  wire [10:0] add_132401;
  wire [11:0] sel_132404;
  wire [11:0] add_132429;
  wire [11:0] sel_132431;
  wire [11:0] add_132434;
  wire [11:0] sel_132436;
  wire [15:0] array_index_132465;
  wire [15:0] array_index_132468;
  wire [10:0] add_132472;
  wire [11:0] sel_132474;
  wire [10:0] add_132476;
  wire [11:0] sel_132478;
  wire [10:0] add_132480;
  wire [11:0] sel_132482;
  wire [10:0] add_132484;
  wire [11:0] sel_132486;
  wire [8:0] add_132488;
  wire [11:0] sel_132491;
  wire [8:0] add_132493;
  wire [11:0] sel_132496;
  wire [10:0] add_132498;
  wire [11:0] sel_132501;
  wire [10:0] add_132503;
  wire [11:0] sel_132506;
  wire [11:0] add_132531;
  wire [11:0] sel_132533;
  wire [11:0] add_132536;
  wire [11:0] sel_132538;
  wire [15:0] array_index_132567;
  wire [15:0] array_index_132570;
  wire [10:0] add_132574;
  wire [11:0] sel_132576;
  wire [10:0] add_132578;
  wire [11:0] sel_132580;
  wire [10:0] add_132582;
  wire [11:0] sel_132584;
  wire [10:0] add_132586;
  wire [11:0] sel_132588;
  wire [8:0] add_132590;
  wire [11:0] sel_132593;
  wire [8:0] add_132595;
  wire [11:0] sel_132598;
  wire [10:0] add_132600;
  wire [11:0] sel_132603;
  wire [10:0] add_132605;
  wire [11:0] sel_132608;
  wire [11:0] add_132633;
  wire [11:0] sel_132635;
  wire [11:0] add_132638;
  wire [11:0] sel_132640;
  wire [15:0] array_index_132669;
  wire [15:0] array_index_132672;
  wire [10:0] add_132676;
  wire [11:0] sel_132678;
  wire [10:0] add_132680;
  wire [11:0] sel_132682;
  wire [10:0] add_132684;
  wire [11:0] sel_132686;
  wire [10:0] add_132688;
  wire [11:0] sel_132690;
  wire [8:0] add_132692;
  wire [11:0] sel_132695;
  wire [8:0] add_132697;
  wire [11:0] sel_132700;
  wire [10:0] add_132702;
  wire [11:0] sel_132705;
  wire [10:0] add_132707;
  wire [11:0] sel_132710;
  wire [11:0] add_132735;
  wire [11:0] sel_132737;
  wire [11:0] add_132740;
  wire [11:0] sel_132742;
  wire [15:0] array_index_132771;
  wire [15:0] array_index_132774;
  wire [10:0] add_132778;
  wire [11:0] sel_132780;
  wire [10:0] add_132782;
  wire [11:0] sel_132784;
  wire [10:0] add_132786;
  wire [11:0] sel_132788;
  wire [10:0] add_132790;
  wire [11:0] sel_132792;
  wire [8:0] add_132794;
  wire [11:0] sel_132797;
  wire [8:0] add_132799;
  wire [11:0] sel_132802;
  wire [10:0] add_132804;
  wire [11:0] sel_132807;
  wire [10:0] add_132809;
  wire [11:0] sel_132812;
  wire [11:0] add_132837;
  wire [11:0] sel_132839;
  wire [11:0] add_132842;
  wire [11:0] sel_132844;
  wire [15:0] array_index_132873;
  wire [15:0] array_index_132876;
  wire [10:0] add_132880;
  wire [11:0] sel_132882;
  wire [10:0] add_132884;
  wire [11:0] sel_132886;
  wire [10:0] add_132888;
  wire [11:0] sel_132890;
  wire [10:0] add_132892;
  wire [11:0] sel_132894;
  wire [8:0] add_132896;
  wire [11:0] sel_132899;
  wire [8:0] add_132901;
  wire [11:0] sel_132904;
  wire [10:0] add_132906;
  wire [11:0] sel_132909;
  wire [10:0] add_132911;
  wire [11:0] sel_132914;
  wire [11:0] add_132939;
  wire [11:0] sel_132941;
  wire [11:0] add_132944;
  wire [11:0] sel_132946;
  wire [15:0] array_index_132975;
  wire [15:0] array_index_132978;
  wire [10:0] add_132982;
  wire [11:0] sel_132984;
  wire [10:0] add_132986;
  wire [11:0] sel_132988;
  wire [10:0] add_132990;
  wire [11:0] sel_132992;
  wire [10:0] add_132994;
  wire [11:0] sel_132996;
  wire [8:0] add_132998;
  wire [11:0] sel_133001;
  wire [8:0] add_133003;
  wire [11:0] sel_133006;
  wire [10:0] add_133008;
  wire [11:0] sel_133011;
  wire [10:0] add_133013;
  wire [11:0] sel_133016;
  wire [11:0] add_133041;
  wire [11:0] sel_133043;
  wire [11:0] add_133046;
  wire [11:0] sel_133048;
  wire [15:0] array_index_133077;
  wire [15:0] array_index_133080;
  wire [10:0] add_133084;
  wire [11:0] sel_133086;
  wire [10:0] add_133088;
  wire [11:0] sel_133090;
  wire [10:0] add_133092;
  wire [11:0] sel_133094;
  wire [10:0] add_133096;
  wire [11:0] sel_133098;
  wire [8:0] add_133100;
  wire [11:0] sel_133103;
  wire [8:0] add_133105;
  wire [11:0] sel_133108;
  wire [10:0] add_133110;
  wire [11:0] sel_133113;
  wire [10:0] add_133115;
  wire [11:0] sel_133118;
  wire [11:0] add_133143;
  wire [11:0] sel_133145;
  wire [11:0] add_133148;
  wire [11:0] sel_133150;
  wire [15:0] array_index_133179;
  wire [15:0] array_index_133182;
  wire [10:0] add_133186;
  wire [11:0] sel_133188;
  wire [10:0] add_133190;
  wire [11:0] sel_133192;
  wire [10:0] add_133194;
  wire [11:0] sel_133196;
  wire [10:0] add_133198;
  wire [11:0] sel_133200;
  wire [8:0] add_133202;
  wire [11:0] sel_133205;
  wire [8:0] add_133207;
  wire [11:0] sel_133210;
  wire [10:0] add_133212;
  wire [11:0] sel_133215;
  wire [10:0] add_133217;
  wire [11:0] sel_133220;
  wire [11:0] add_133245;
  wire [11:0] sel_133247;
  wire [11:0] add_133250;
  wire [11:0] sel_133252;
  wire [15:0] array_index_133281;
  wire [15:0] array_index_133284;
  wire [10:0] add_133288;
  wire [11:0] sel_133290;
  wire [10:0] add_133292;
  wire [11:0] sel_133294;
  wire [10:0] add_133296;
  wire [11:0] sel_133298;
  wire [10:0] add_133300;
  wire [11:0] sel_133302;
  wire [8:0] add_133304;
  wire [11:0] sel_133307;
  wire [8:0] add_133309;
  wire [11:0] sel_133312;
  wire [10:0] add_133314;
  wire [11:0] sel_133317;
  wire [10:0] add_133319;
  wire [11:0] sel_133322;
  wire [11:0] add_133347;
  wire [11:0] sel_133349;
  wire [11:0] add_133352;
  wire [11:0] sel_133354;
  wire [15:0] array_index_133383;
  wire [15:0] array_index_133386;
  wire [10:0] add_133390;
  wire [11:0] sel_133392;
  wire [10:0] add_133394;
  wire [11:0] sel_133396;
  wire [10:0] add_133398;
  wire [11:0] sel_133400;
  wire [10:0] add_133402;
  wire [11:0] sel_133404;
  wire [8:0] add_133406;
  wire [11:0] sel_133409;
  wire [8:0] add_133411;
  wire [11:0] sel_133414;
  wire [10:0] add_133416;
  wire [11:0] sel_133419;
  wire [10:0] add_133421;
  wire [11:0] sel_133424;
  wire [11:0] add_133449;
  wire [11:0] sel_133451;
  wire [11:0] add_133454;
  wire [11:0] sel_133456;
  wire [15:0] array_index_133485;
  wire [15:0] array_index_133488;
  wire [10:0] add_133492;
  wire [11:0] sel_133494;
  wire [10:0] add_133496;
  wire [11:0] sel_133498;
  wire [10:0] add_133500;
  wire [11:0] sel_133502;
  wire [10:0] add_133504;
  wire [11:0] sel_133506;
  wire [8:0] add_133508;
  wire [11:0] sel_133511;
  wire [8:0] add_133513;
  wire [11:0] sel_133516;
  wire [10:0] add_133518;
  wire [11:0] sel_133521;
  wire [10:0] add_133523;
  wire [11:0] sel_133526;
  wire [11:0] add_133551;
  wire [11:0] sel_133553;
  wire [11:0] add_133556;
  wire [11:0] sel_133558;
  wire [15:0] array_index_133587;
  wire [15:0] array_index_133590;
  wire [10:0] add_133594;
  wire [11:0] sel_133596;
  wire [10:0] add_133598;
  wire [11:0] sel_133600;
  wire [10:0] add_133602;
  wire [11:0] sel_133604;
  wire [10:0] add_133606;
  wire [11:0] sel_133608;
  wire [8:0] add_133610;
  wire [11:0] sel_133613;
  wire [8:0] add_133615;
  wire [11:0] sel_133618;
  wire [10:0] add_133620;
  wire [11:0] sel_133623;
  wire [10:0] add_133625;
  wire [11:0] sel_133628;
  wire [11:0] add_133653;
  wire [11:0] sel_133655;
  wire [11:0] add_133658;
  wire [11:0] sel_133660;
  wire [15:0] array_index_133689;
  wire [15:0] array_index_133692;
  wire [10:0] add_133696;
  wire [11:0] sel_133698;
  wire [10:0] add_133700;
  wire [11:0] sel_133702;
  wire [10:0] add_133704;
  wire [11:0] sel_133706;
  wire [10:0] add_133708;
  wire [11:0] sel_133710;
  wire [8:0] add_133712;
  wire [11:0] sel_133715;
  wire [8:0] add_133717;
  wire [11:0] sel_133720;
  wire [10:0] add_133722;
  wire [11:0] sel_133725;
  wire [10:0] add_133727;
  wire [11:0] sel_133730;
  wire [11:0] add_133755;
  wire [11:0] sel_133757;
  wire [11:0] add_133760;
  wire [11:0] sel_133762;
  wire [15:0] array_index_133791;
  wire [15:0] array_index_133794;
  wire [10:0] add_133798;
  wire [11:0] sel_133800;
  wire [10:0] add_133802;
  wire [11:0] sel_133804;
  wire [10:0] add_133806;
  wire [11:0] sel_133808;
  wire [10:0] add_133810;
  wire [11:0] sel_133812;
  wire [8:0] add_133814;
  wire [11:0] sel_133817;
  wire [8:0] add_133819;
  wire [11:0] sel_133822;
  wire [10:0] add_133824;
  wire [11:0] sel_133827;
  wire [10:0] add_133829;
  wire [11:0] sel_133832;
  wire [11:0] add_133857;
  wire [11:0] sel_133859;
  wire [11:0] add_133862;
  wire [11:0] sel_133864;
  wire [15:0] array_index_133893;
  wire [15:0] array_index_133896;
  wire [10:0] add_133900;
  wire [11:0] sel_133902;
  wire [10:0] add_133904;
  wire [11:0] sel_133906;
  wire [10:0] add_133908;
  wire [11:0] sel_133910;
  wire [10:0] add_133912;
  wire [11:0] sel_133914;
  wire [8:0] add_133916;
  wire [11:0] sel_133919;
  wire [8:0] add_133921;
  wire [11:0] sel_133924;
  wire [10:0] add_133926;
  wire [11:0] sel_133929;
  wire [10:0] add_133931;
  wire [11:0] sel_133934;
  wire [11:0] add_133959;
  wire [11:0] sel_133961;
  wire [11:0] add_133964;
  wire [11:0] sel_133966;
  wire [15:0] array_index_133995;
  wire [15:0] array_index_133998;
  wire [10:0] add_134002;
  wire [11:0] sel_134004;
  wire [10:0] add_134006;
  wire [11:0] sel_134008;
  wire [10:0] add_134010;
  wire [11:0] sel_134012;
  wire [10:0] add_134014;
  wire [11:0] sel_134016;
  wire [8:0] add_134018;
  wire [11:0] sel_134021;
  wire [8:0] add_134023;
  wire [11:0] sel_134026;
  wire [10:0] add_134028;
  wire [11:0] sel_134031;
  wire [10:0] add_134033;
  wire [11:0] sel_134036;
  wire [11:0] add_134061;
  wire [11:0] sel_134063;
  wire [11:0] add_134066;
  wire [11:0] sel_134068;
  wire [15:0] array_index_134097;
  wire [15:0] array_index_134100;
  wire [10:0] add_134104;
  wire [11:0] sel_134106;
  wire [10:0] add_134108;
  wire [11:0] sel_134110;
  wire [10:0] add_134112;
  wire [11:0] sel_134114;
  wire [10:0] add_134116;
  wire [11:0] sel_134118;
  wire [8:0] add_134120;
  wire [11:0] sel_134123;
  wire [8:0] add_134125;
  wire [11:0] sel_134128;
  wire [10:0] add_134130;
  wire [11:0] sel_134133;
  wire [10:0] add_134135;
  wire [11:0] sel_134138;
  wire [11:0] add_134163;
  wire [11:0] sel_134165;
  wire [11:0] add_134168;
  wire [11:0] sel_134170;
  wire [15:0] array_index_134199;
  wire [15:0] array_index_134202;
  wire [10:0] add_134206;
  wire [11:0] sel_134208;
  wire [10:0] add_134210;
  wire [11:0] sel_134212;
  wire [10:0] add_134214;
  wire [11:0] sel_134216;
  wire [10:0] add_134218;
  wire [11:0] sel_134220;
  wire [8:0] add_134222;
  wire [11:0] sel_134225;
  wire [8:0] add_134227;
  wire [11:0] sel_134230;
  wire [10:0] add_134232;
  wire [11:0] sel_134235;
  wire [10:0] add_134237;
  wire [11:0] sel_134240;
  wire [11:0] add_134265;
  wire [11:0] sel_134267;
  wire [11:0] add_134270;
  wire [11:0] sel_134272;
  wire [15:0] array_index_134301;
  wire [15:0] array_index_134304;
  wire [10:0] add_134308;
  wire [11:0] sel_134310;
  wire [10:0] add_134312;
  wire [11:0] sel_134314;
  wire [10:0] add_134316;
  wire [11:0] sel_134318;
  wire [10:0] add_134320;
  wire [11:0] sel_134322;
  wire [8:0] add_134324;
  wire [11:0] sel_134327;
  wire [8:0] add_134329;
  wire [11:0] sel_134332;
  wire [10:0] add_134334;
  wire [11:0] sel_134337;
  wire [10:0] add_134339;
  wire [11:0] sel_134342;
  wire [11:0] add_134367;
  wire [11:0] sel_134369;
  wire [11:0] add_134372;
  wire [11:0] sel_134374;
  wire [15:0] array_index_134403;
  wire [15:0] array_index_134406;
  wire [10:0] add_134410;
  wire [11:0] sel_134412;
  wire [10:0] add_134414;
  wire [11:0] sel_134416;
  wire [10:0] add_134418;
  wire [11:0] sel_134420;
  wire [10:0] add_134422;
  wire [11:0] sel_134424;
  wire [8:0] add_134426;
  wire [11:0] sel_134429;
  wire [8:0] add_134431;
  wire [11:0] sel_134434;
  wire [10:0] add_134436;
  wire [11:0] sel_134439;
  wire [10:0] add_134441;
  wire [11:0] sel_134444;
  wire [11:0] add_134469;
  wire [11:0] sel_134471;
  wire [11:0] add_134474;
  wire [11:0] sel_134476;
  wire [15:0] array_index_134505;
  wire [15:0] array_index_134508;
  wire [10:0] add_134512;
  wire [11:0] sel_134514;
  wire [10:0] add_134516;
  wire [11:0] sel_134518;
  wire [10:0] add_134520;
  wire [11:0] sel_134522;
  wire [10:0] add_134524;
  wire [11:0] sel_134526;
  wire [8:0] add_134528;
  wire [11:0] sel_134531;
  wire [8:0] add_134533;
  wire [11:0] sel_134536;
  wire [10:0] add_134538;
  wire [11:0] sel_134541;
  wire [10:0] add_134543;
  wire [11:0] sel_134546;
  wire [11:0] add_134571;
  wire [11:0] sel_134573;
  wire [11:0] add_134576;
  wire [11:0] sel_134578;
  wire [15:0] array_index_134607;
  wire [15:0] array_index_134610;
  wire [10:0] add_134614;
  wire [11:0] sel_134616;
  wire [10:0] add_134618;
  wire [11:0] sel_134620;
  wire [10:0] add_134622;
  wire [11:0] sel_134624;
  wire [10:0] add_134626;
  wire [11:0] sel_134628;
  wire [8:0] add_134630;
  wire [11:0] sel_134633;
  wire [8:0] add_134635;
  wire [11:0] sel_134638;
  wire [10:0] add_134640;
  wire [11:0] sel_134643;
  wire [10:0] add_134645;
  wire [11:0] sel_134648;
  wire [11:0] add_134673;
  wire [11:0] sel_134675;
  wire [11:0] add_134678;
  wire [11:0] sel_134680;
  wire [15:0] array_index_134709;
  wire [15:0] array_index_134712;
  wire [10:0] add_134716;
  wire [11:0] sel_134718;
  wire [10:0] add_134720;
  wire [11:0] sel_134722;
  wire [10:0] add_134724;
  wire [11:0] sel_134726;
  wire [10:0] add_134728;
  wire [11:0] sel_134730;
  wire [8:0] add_134732;
  wire [11:0] sel_134735;
  wire [8:0] add_134737;
  wire [11:0] sel_134740;
  wire [10:0] add_134742;
  wire [11:0] sel_134745;
  wire [10:0] add_134747;
  wire [11:0] sel_134750;
  wire [11:0] add_134775;
  wire [11:0] sel_134777;
  wire [11:0] add_134780;
  wire [11:0] sel_134782;
  wire [15:0] array_index_134811;
  wire [15:0] array_index_134814;
  wire [10:0] add_134818;
  wire [11:0] sel_134820;
  wire [10:0] add_134822;
  wire [11:0] sel_134824;
  wire [10:0] add_134826;
  wire [11:0] sel_134828;
  wire [10:0] add_134830;
  wire [11:0] sel_134832;
  wire [8:0] add_134834;
  wire [11:0] sel_134837;
  wire [8:0] add_134839;
  wire [11:0] sel_134842;
  wire [10:0] add_134844;
  wire [11:0] sel_134847;
  wire [10:0] add_134849;
  wire [11:0] sel_134852;
  wire [11:0] add_134877;
  wire [11:0] sel_134879;
  wire [11:0] add_134882;
  wire [11:0] sel_134884;
  wire [15:0] array_index_134913;
  wire [15:0] array_index_134916;
  wire [10:0] add_134920;
  wire [11:0] sel_134922;
  wire [10:0] add_134924;
  wire [11:0] sel_134926;
  wire [10:0] add_134928;
  wire [11:0] sel_134930;
  wire [10:0] add_134932;
  wire [11:0] sel_134934;
  wire [8:0] add_134936;
  wire [11:0] sel_134939;
  wire [8:0] add_134941;
  wire [11:0] sel_134944;
  wire [10:0] add_134946;
  wire [11:0] sel_134949;
  wire [10:0] add_134951;
  wire [11:0] sel_134954;
  wire [11:0] add_134979;
  wire [11:0] sel_134981;
  wire [11:0] add_134984;
  wire [11:0] sel_134986;
  wire [15:0] array_index_135015;
  wire [15:0] array_index_135018;
  wire [10:0] add_135022;
  wire [11:0] sel_135024;
  wire [10:0] add_135026;
  wire [11:0] sel_135028;
  wire [10:0] add_135030;
  wire [11:0] sel_135032;
  wire [10:0] add_135034;
  wire [11:0] sel_135036;
  wire [8:0] add_135038;
  wire [11:0] sel_135041;
  wire [8:0] add_135043;
  wire [11:0] sel_135046;
  wire [10:0] add_135048;
  wire [11:0] sel_135051;
  wire [10:0] add_135053;
  wire [11:0] sel_135056;
  wire [11:0] add_135081;
  wire [11:0] sel_135083;
  wire [11:0] add_135086;
  wire [11:0] sel_135088;
  wire [15:0] array_index_135117;
  wire [15:0] array_index_135120;
  wire [10:0] add_135124;
  wire [11:0] sel_135126;
  wire [10:0] add_135128;
  wire [11:0] sel_135130;
  wire [10:0] add_135132;
  wire [11:0] sel_135134;
  wire [10:0] add_135136;
  wire [11:0] sel_135138;
  wire [8:0] add_135140;
  wire [11:0] sel_135143;
  wire [8:0] add_135145;
  wire [11:0] sel_135148;
  wire [10:0] add_135150;
  wire [11:0] sel_135153;
  wire [10:0] add_135155;
  wire [11:0] sel_135158;
  wire [11:0] add_135183;
  wire [11:0] sel_135185;
  wire [11:0] add_135188;
  wire [11:0] sel_135190;
  wire [15:0] array_index_135219;
  wire [15:0] array_index_135222;
  wire [10:0] add_135226;
  wire [11:0] sel_135228;
  wire [10:0] add_135230;
  wire [11:0] sel_135232;
  wire [10:0] add_135234;
  wire [11:0] sel_135236;
  wire [10:0] add_135238;
  wire [11:0] sel_135240;
  wire [8:0] add_135242;
  wire [11:0] sel_135245;
  wire [8:0] add_135247;
  wire [11:0] sel_135250;
  wire [10:0] add_135252;
  wire [11:0] sel_135255;
  wire [10:0] add_135257;
  wire [11:0] sel_135260;
  wire [11:0] add_135285;
  wire [11:0] sel_135287;
  wire [11:0] add_135290;
  wire [11:0] sel_135292;
  wire [15:0] array_index_135321;
  wire [15:0] array_index_135324;
  wire [10:0] add_135328;
  wire [11:0] sel_135330;
  wire [10:0] add_135332;
  wire [11:0] sel_135334;
  wire [10:0] add_135336;
  wire [11:0] sel_135338;
  wire [10:0] add_135340;
  wire [11:0] sel_135342;
  wire [8:0] add_135344;
  wire [11:0] sel_135347;
  wire [8:0] add_135349;
  wire [11:0] sel_135352;
  wire [10:0] add_135354;
  wire [11:0] sel_135357;
  wire [10:0] add_135359;
  wire [11:0] sel_135362;
  wire [11:0] add_135387;
  wire [11:0] sel_135389;
  wire [11:0] add_135392;
  wire [11:0] sel_135394;
  wire [15:0] array_index_135423;
  wire [15:0] array_index_135426;
  wire [10:0] add_135430;
  wire [11:0] sel_135432;
  wire [10:0] add_135434;
  wire [11:0] sel_135436;
  wire [10:0] add_135438;
  wire [11:0] sel_135440;
  wire [10:0] add_135442;
  wire [11:0] sel_135444;
  wire [8:0] add_135446;
  wire [11:0] sel_135449;
  wire [8:0] add_135451;
  wire [11:0] sel_135454;
  wire [10:0] add_135456;
  wire [11:0] sel_135459;
  wire [10:0] add_135461;
  wire [11:0] sel_135464;
  wire [11:0] add_135489;
  wire [11:0] sel_135491;
  wire [11:0] add_135494;
  wire [11:0] sel_135496;
  wire [15:0] array_index_135525;
  wire [15:0] array_index_135528;
  wire [10:0] add_135532;
  wire [11:0] sel_135534;
  wire [10:0] add_135536;
  wire [11:0] sel_135538;
  wire [10:0] add_135540;
  wire [11:0] sel_135542;
  wire [10:0] add_135544;
  wire [11:0] sel_135546;
  wire [8:0] add_135548;
  wire [11:0] sel_135551;
  wire [8:0] add_135553;
  wire [11:0] sel_135556;
  wire [10:0] add_135558;
  wire [11:0] sel_135561;
  wire [10:0] add_135563;
  wire [11:0] sel_135566;
  wire [11:0] add_135591;
  wire [11:0] sel_135593;
  wire [11:0] add_135596;
  wire [11:0] sel_135598;
  wire [15:0] array_index_135627;
  wire [15:0] array_index_135630;
  wire [10:0] add_135634;
  wire [11:0] sel_135636;
  wire [10:0] add_135638;
  wire [11:0] sel_135640;
  wire [10:0] add_135642;
  wire [11:0] sel_135644;
  wire [10:0] add_135646;
  wire [11:0] sel_135648;
  wire [8:0] add_135650;
  wire [11:0] sel_135653;
  wire [8:0] add_135655;
  wire [11:0] sel_135658;
  wire [10:0] add_135660;
  wire [11:0] sel_135663;
  wire [10:0] add_135665;
  wire [11:0] sel_135668;
  wire [11:0] add_135693;
  wire [11:0] sel_135695;
  wire [11:0] add_135698;
  wire [11:0] sel_135700;
  wire [15:0] array_index_135729;
  wire [15:0] array_index_135732;
  wire [10:0] add_135736;
  wire [11:0] sel_135738;
  wire [10:0] add_135740;
  wire [11:0] sel_135742;
  wire [10:0] add_135744;
  wire [11:0] sel_135746;
  wire [10:0] add_135748;
  wire [11:0] sel_135750;
  wire [8:0] add_135752;
  wire [11:0] sel_135755;
  wire [8:0] add_135757;
  wire [11:0] sel_135760;
  wire [10:0] add_135762;
  wire [11:0] sel_135765;
  wire [10:0] add_135767;
  wire [11:0] sel_135770;
  wire [11:0] add_135795;
  wire [11:0] sel_135797;
  wire [11:0] add_135800;
  wire [11:0] sel_135802;
  wire [15:0] array_index_135831;
  wire [15:0] array_index_135834;
  wire [10:0] add_135838;
  wire [11:0] sel_135840;
  wire [10:0] add_135842;
  wire [11:0] sel_135844;
  wire [10:0] add_135846;
  wire [11:0] sel_135848;
  wire [10:0] add_135850;
  wire [11:0] sel_135852;
  wire [8:0] add_135854;
  wire [11:0] sel_135857;
  wire [8:0] add_135859;
  wire [11:0] sel_135862;
  wire [10:0] add_135864;
  wire [11:0] sel_135867;
  wire [10:0] add_135869;
  wire [11:0] sel_135872;
  wire [11:0] add_135897;
  wire [11:0] sel_135899;
  wire [11:0] add_135902;
  wire [11:0] sel_135904;
  wire [15:0] array_index_135933;
  wire [15:0] array_index_135936;
  wire [10:0] add_135940;
  wire [11:0] sel_135942;
  wire [10:0] add_135944;
  wire [11:0] sel_135946;
  wire [10:0] add_135948;
  wire [11:0] sel_135950;
  wire [10:0] add_135952;
  wire [11:0] sel_135954;
  wire [8:0] add_135956;
  wire [11:0] sel_135959;
  wire [8:0] add_135961;
  wire [11:0] sel_135964;
  wire [10:0] add_135966;
  wire [11:0] sel_135969;
  wire [10:0] add_135971;
  wire [11:0] sel_135974;
  wire [11:0] add_135999;
  wire [11:0] sel_136001;
  wire [11:0] add_136004;
  wire [11:0] sel_136006;
  wire [15:0] array_index_136035;
  wire [15:0] array_index_136038;
  wire [10:0] add_136042;
  wire [11:0] sel_136044;
  wire [10:0] add_136046;
  wire [11:0] sel_136048;
  wire [10:0] add_136050;
  wire [11:0] sel_136052;
  wire [10:0] add_136054;
  wire [11:0] sel_136056;
  wire [8:0] add_136058;
  wire [11:0] sel_136061;
  wire [8:0] add_136063;
  wire [11:0] sel_136066;
  wire [10:0] add_136068;
  wire [11:0] sel_136071;
  wire [10:0] add_136073;
  wire [11:0] sel_136076;
  wire [11:0] add_136101;
  wire [11:0] sel_136103;
  wire [11:0] add_136106;
  wire [11:0] sel_136108;
  wire [15:0] array_index_136137;
  wire [15:0] array_index_136140;
  wire [10:0] add_136144;
  wire [11:0] sel_136146;
  wire [10:0] add_136148;
  wire [11:0] sel_136150;
  wire [10:0] add_136152;
  wire [11:0] sel_136154;
  wire [10:0] add_136156;
  wire [11:0] sel_136158;
  wire [8:0] add_136160;
  wire [11:0] sel_136163;
  wire [8:0] add_136165;
  wire [11:0] sel_136168;
  wire [10:0] add_136170;
  wire [11:0] sel_136173;
  wire [10:0] add_136175;
  wire [11:0] sel_136178;
  wire [11:0] add_136203;
  wire [11:0] sel_136205;
  wire [11:0] add_136208;
  wire [11:0] sel_136210;
  wire [15:0] array_index_136239;
  wire [15:0] array_index_136242;
  wire [10:0] add_136246;
  wire [11:0] sel_136248;
  wire [10:0] add_136250;
  wire [11:0] sel_136252;
  wire [10:0] add_136254;
  wire [11:0] sel_136256;
  wire [10:0] add_136258;
  wire [11:0] sel_136260;
  wire [8:0] add_136262;
  wire [11:0] sel_136265;
  wire [8:0] add_136267;
  wire [11:0] sel_136270;
  wire [10:0] add_136272;
  wire [11:0] sel_136275;
  wire [10:0] add_136277;
  wire [11:0] sel_136280;
  wire [11:0] add_136305;
  wire [11:0] sel_136307;
  wire [11:0] add_136310;
  wire [11:0] sel_136312;
  wire [15:0] array_index_136341;
  wire [15:0] array_index_136344;
  wire [10:0] add_136348;
  wire [11:0] sel_136350;
  wire [10:0] add_136352;
  wire [11:0] sel_136354;
  wire [10:0] add_136356;
  wire [11:0] sel_136358;
  wire [10:0] add_136360;
  wire [11:0] sel_136362;
  wire [8:0] add_136364;
  wire [11:0] sel_136367;
  wire [8:0] add_136369;
  wire [11:0] sel_136372;
  wire [10:0] add_136374;
  wire [11:0] sel_136377;
  wire [10:0] add_136379;
  wire [11:0] sel_136382;
  wire [11:0] add_136407;
  wire [11:0] sel_136409;
  wire [11:0] add_136412;
  wire [11:0] sel_136414;
  wire [15:0] array_index_136443;
  wire [15:0] array_index_136446;
  wire [10:0] add_136450;
  wire [11:0] sel_136452;
  wire [10:0] add_136454;
  wire [11:0] sel_136456;
  wire [10:0] add_136458;
  wire [11:0] sel_136460;
  wire [10:0] add_136462;
  wire [11:0] sel_136464;
  wire [8:0] add_136466;
  wire [11:0] sel_136469;
  wire [8:0] add_136471;
  wire [11:0] sel_136474;
  wire [10:0] add_136476;
  wire [11:0] sel_136479;
  wire [10:0] add_136481;
  wire [11:0] sel_136484;
  wire [11:0] add_136509;
  wire [11:0] sel_136511;
  wire [11:0] add_136514;
  wire [11:0] sel_136516;
  wire [15:0] array_index_136545;
  wire [15:0] array_index_136548;
  wire [10:0] add_136552;
  wire [11:0] sel_136554;
  wire [10:0] add_136556;
  wire [11:0] sel_136558;
  wire [10:0] add_136560;
  wire [11:0] sel_136562;
  wire [10:0] add_136564;
  wire [11:0] sel_136566;
  wire [8:0] add_136568;
  wire [11:0] sel_136571;
  wire [8:0] add_136573;
  wire [11:0] sel_136576;
  wire [10:0] add_136578;
  wire [11:0] sel_136581;
  wire [10:0] add_136583;
  wire [11:0] sel_136586;
  wire [11:0] add_136611;
  wire [11:0] sel_136613;
  wire [11:0] add_136616;
  wire [11:0] sel_136618;
  wire [15:0] array_index_136647;
  wire [15:0] array_index_136650;
  wire [10:0] add_136654;
  wire [11:0] sel_136656;
  wire [10:0] add_136658;
  wire [11:0] sel_136660;
  wire [10:0] add_136662;
  wire [11:0] sel_136664;
  wire [10:0] add_136666;
  wire [11:0] sel_136668;
  wire [8:0] add_136670;
  wire [11:0] sel_136673;
  wire [8:0] add_136675;
  wire [11:0] sel_136678;
  wire [10:0] add_136680;
  wire [11:0] sel_136683;
  wire [10:0] add_136685;
  wire [11:0] sel_136688;
  wire [11:0] add_136713;
  wire [11:0] sel_136715;
  wire [11:0] add_136718;
  wire [11:0] sel_136720;
  wire [15:0] array_index_136749;
  wire [15:0] array_index_136752;
  wire [10:0] add_136756;
  wire [11:0] sel_136758;
  wire [10:0] add_136760;
  wire [11:0] sel_136762;
  wire [10:0] add_136764;
  wire [11:0] sel_136766;
  wire [10:0] add_136768;
  wire [11:0] sel_136770;
  wire [8:0] add_136772;
  wire [11:0] sel_136775;
  wire [8:0] add_136777;
  wire [11:0] sel_136780;
  wire [10:0] add_136782;
  wire [11:0] sel_136785;
  wire [10:0] add_136787;
  wire [11:0] sel_136790;
  wire [11:0] add_136815;
  wire [11:0] sel_136817;
  wire [11:0] add_136820;
  wire [11:0] sel_136822;
  wire [15:0] array_index_136851;
  wire [15:0] array_index_136854;
  wire [10:0] add_136858;
  wire [11:0] sel_136860;
  wire [10:0] add_136862;
  wire [11:0] sel_136864;
  wire [10:0] add_136866;
  wire [11:0] sel_136868;
  wire [10:0] add_136870;
  wire [11:0] sel_136872;
  wire [8:0] add_136874;
  wire [11:0] sel_136877;
  wire [8:0] add_136879;
  wire [11:0] sel_136882;
  wire [10:0] add_136884;
  wire [11:0] sel_136887;
  wire [10:0] add_136889;
  wire [11:0] sel_136892;
  wire [11:0] add_136917;
  wire [11:0] sel_136919;
  wire [11:0] add_136922;
  wire [11:0] sel_136924;
  wire [15:0] array_index_136953;
  wire [15:0] array_index_136956;
  wire [10:0] add_136960;
  wire [11:0] sel_136962;
  wire [10:0] add_136964;
  wire [11:0] sel_136966;
  wire [10:0] add_136968;
  wire [11:0] sel_136970;
  wire [10:0] add_136972;
  wire [11:0] sel_136974;
  wire [8:0] add_136976;
  wire [11:0] sel_136979;
  wire [8:0] add_136981;
  wire [11:0] sel_136984;
  wire [10:0] add_136986;
  wire [11:0] sel_136989;
  wire [10:0] add_136991;
  wire [11:0] sel_136994;
  wire [11:0] add_137019;
  wire [11:0] sel_137021;
  wire [11:0] add_137024;
  wire [11:0] sel_137026;
  wire [15:0] array_index_137055;
  wire [15:0] array_index_137058;
  wire [10:0] add_137062;
  wire [11:0] sel_137064;
  wire [10:0] add_137066;
  wire [11:0] sel_137068;
  wire [10:0] add_137070;
  wire [11:0] sel_137072;
  wire [10:0] add_137074;
  wire [11:0] sel_137076;
  wire [8:0] add_137078;
  wire [11:0] sel_137081;
  wire [8:0] add_137083;
  wire [11:0] sel_137086;
  wire [10:0] add_137088;
  wire [11:0] sel_137091;
  wire [10:0] add_137093;
  wire [11:0] sel_137096;
  wire [11:0] add_137121;
  wire [11:0] sel_137123;
  wire [11:0] add_137126;
  wire [11:0] sel_137128;
  wire [15:0] array_index_137157;
  wire [15:0] array_index_137160;
  wire [10:0] add_137164;
  wire [11:0] sel_137166;
  wire [10:0] add_137168;
  wire [11:0] sel_137170;
  wire [10:0] add_137172;
  wire [11:0] sel_137174;
  wire [10:0] add_137176;
  wire [11:0] sel_137178;
  wire [8:0] add_137180;
  wire [11:0] sel_137183;
  wire [8:0] add_137185;
  wire [11:0] sel_137188;
  wire [10:0] add_137190;
  wire [11:0] sel_137193;
  wire [10:0] add_137195;
  wire [11:0] sel_137198;
  wire [11:0] add_137223;
  wire [11:0] sel_137225;
  wire [11:0] add_137228;
  wire [11:0] sel_137230;
  wire [15:0] array_index_137259;
  wire [15:0] array_index_137262;
  wire [10:0] add_137266;
  wire [11:0] sel_137268;
  wire [10:0] add_137270;
  wire [11:0] sel_137272;
  wire [10:0] add_137274;
  wire [11:0] sel_137276;
  wire [10:0] add_137278;
  wire [11:0] sel_137280;
  wire [8:0] add_137282;
  wire [11:0] sel_137285;
  wire [8:0] add_137287;
  wire [11:0] sel_137290;
  wire [10:0] add_137292;
  wire [11:0] sel_137295;
  wire [10:0] add_137297;
  wire [11:0] sel_137300;
  wire [11:0] add_137325;
  wire [11:0] sel_137327;
  wire [11:0] add_137330;
  wire [11:0] sel_137332;
  wire [15:0] array_index_137361;
  wire [15:0] array_index_137364;
  wire [10:0] add_137368;
  wire [11:0] sel_137370;
  wire [10:0] add_137372;
  wire [11:0] sel_137374;
  wire [10:0] add_137376;
  wire [11:0] sel_137378;
  wire [10:0] add_137380;
  wire [11:0] sel_137382;
  wire [8:0] add_137384;
  wire [11:0] sel_137387;
  wire [8:0] add_137389;
  wire [11:0] sel_137392;
  wire [10:0] add_137394;
  wire [11:0] sel_137397;
  wire [10:0] add_137399;
  wire [11:0] sel_137402;
  wire [11:0] add_137427;
  wire [11:0] sel_137429;
  wire [11:0] add_137432;
  wire [11:0] sel_137434;
  wire [15:0] array_index_137463;
  wire [15:0] array_index_137466;
  wire [10:0] add_137470;
  wire [11:0] sel_137472;
  wire [10:0] add_137474;
  wire [11:0] sel_137476;
  wire [10:0] add_137478;
  wire [11:0] sel_137480;
  wire [10:0] add_137482;
  wire [11:0] sel_137484;
  wire [8:0] add_137486;
  wire [11:0] sel_137489;
  wire [8:0] add_137491;
  wire [11:0] sel_137494;
  wire [10:0] add_137496;
  wire [11:0] sel_137499;
  wire [10:0] add_137501;
  wire [11:0] sel_137504;
  wire [11:0] add_137529;
  wire [11:0] sel_137531;
  wire [11:0] add_137534;
  wire [11:0] sel_137536;
  wire [15:0] array_index_137565;
  wire [15:0] array_index_137568;
  wire [10:0] add_137572;
  wire [11:0] sel_137574;
  wire [10:0] add_137576;
  wire [11:0] sel_137578;
  wire [10:0] add_137580;
  wire [11:0] sel_137582;
  wire [10:0] add_137584;
  wire [11:0] sel_137586;
  wire [8:0] add_137588;
  wire [11:0] sel_137591;
  wire [8:0] add_137593;
  wire [11:0] sel_137596;
  wire [10:0] add_137598;
  wire [11:0] sel_137601;
  wire [10:0] add_137603;
  wire [11:0] sel_137606;
  wire [11:0] add_137630;
  wire [11:0] sel_137632;
  wire [11:0] add_137634;
  wire [11:0] sel_137636;
  wire [10:0] add_137670;
  wire [11:0] sel_137672;
  wire [10:0] add_137674;
  wire [11:0] sel_137676;
  wire [10:0] add_137678;
  wire [11:0] sel_137680;
  wire [10:0] add_137682;
  wire [11:0] sel_137684;
  wire [8:0] add_137686;
  wire [11:0] sel_137689;
  wire [8:0] add_137691;
  wire [11:0] sel_137694;
  wire [10:0] add_137696;
  wire [11:0] sel_137699;
  wire [10:0] add_137701;
  wire [11:0] sel_137704;
  wire [10:0] add_137752;
  wire [11:0] sel_137754;
  wire [10:0] add_137756;
  wire [11:0] sel_137758;
  wire [10:0] add_137760;
  wire [11:0] sel_137762;
  wire [10:0] add_137764;
  wire [11:0] sel_137766;
  wire [8:0] add_137768;
  wire [11:0] sel_137771;
  wire [8:0] add_137773;
  wire [11:0] sel_137776;
  wire [1:0] concat_137779;
  wire [1:0] add_137794;
  wire [10:0] add_137814;
  wire [11:0] sel_137816;
  wire [10:0] add_137818;
  wire [11:0] sel_137820;
  wire [10:0] add_137822;
  wire [11:0] sel_137824;
  wire [10:0] add_137826;
  wire [11:0] sel_137828;
  wire [2:0] concat_137831;
  wire [2:0] add_137842;
  wire [10:0] add_137856;
  wire [11:0] sel_137858;
  wire [10:0] add_137860;
  wire [11:0] sel_137862;
  wire [3:0] concat_137865;
  wire [3:0] add_137872;
  wire [4:0] concat_137881;
  wire [4:0] add_137884;
  assign array_index_130213 = set1_unflattened[7'h00];
  assign array_index_130214 = set2_unflattened[7'h00];
  assign add_130221 = array_index_130213[11:0] + 12'h247;
  assign add_130224 = array_index_130214[11:0] + 12'h247;
  assign array_index_130229 = set1_unflattened[7'h01];
  assign array_index_130232 = set2_unflattened[7'h01];
  assign add_130236 = array_index_130213[11:1] + 11'h247;
  assign add_130239 = array_index_130214[11:1] + 11'h247;
  assign add_130255 = array_index_130229[11:0] + 12'h247;
  assign sel_130257 = $signed({1'h0, add_130221}) < $signed(13'h0fff) ? add_130221 : 12'hfff;
  assign add_130260 = array_index_130232[11:0] + 12'h247;
  assign sel_130262 = $signed({1'h0, add_130224}) < $signed(13'h0fff) ? add_130224 : 12'hfff;
  assign array_index_130277 = set1_unflattened[7'h02];
  assign array_index_130280 = set2_unflattened[7'h02];
  assign add_130284 = array_index_130213[11:3] + 9'h0bd;
  assign add_130287 = array_index_130214[11:3] + 9'h0bd;
  assign add_130290 = array_index_130229[11:1] + 11'h247;
  assign sel_130293 = $signed({1'h0, add_130236, array_index_130213[0]}) < $signed(13'h0fff) ? {add_130236, array_index_130213[0]} : 12'hfff;
  assign add_130295 = array_index_130232[11:1] + 11'h247;
  assign sel_130298 = $signed({1'h0, add_130239, array_index_130214[0]}) < $signed(13'h0fff) ? {add_130239, array_index_130214[0]} : 12'hfff;
  assign add_130315 = array_index_130277[11:0] + 12'h247;
  assign sel_130317 = $signed({1'h0, add_130255}) < $signed({1'h0, sel_130257}) ? add_130255 : sel_130257;
  assign add_130320 = array_index_130280[11:0] + 12'h247;
  assign sel_130322 = $signed({1'h0, add_130260}) < $signed({1'h0, sel_130262}) ? add_130260 : sel_130262;
  assign array_index_130343 = set1_unflattened[7'h03];
  assign array_index_130346 = set2_unflattened[7'h03];
  assign add_130350 = array_index_130213[11:1] + 11'h347;
  assign add_130352 = array_index_130214[11:1] + 11'h347;
  assign add_130354 = array_index_130229[11:3] + 9'h0bd;
  assign sel_130357 = $signed({1'h0, add_130284, array_index_130213[2:0]}) < $signed(13'h0fff) ? {add_130284, array_index_130213[2:0]} : 12'hfff;
  assign add_130359 = array_index_130232[11:3] + 9'h0bd;
  assign sel_130362 = $signed({1'h0, add_130287, array_index_130214[2:0]}) < $signed(13'h0fff) ? {add_130287, array_index_130214[2:0]} : 12'hfff;
  assign add_130364 = array_index_130277[11:1] + 11'h247;
  assign sel_130367 = $signed({1'h0, add_130290, array_index_130229[0]}) < $signed({1'h0, sel_130293}) ? {add_130290, array_index_130229[0]} : sel_130293;
  assign add_130369 = array_index_130280[11:1] + 11'h247;
  assign sel_130372 = $signed({1'h0, add_130295, array_index_130232[0]}) < $signed({1'h0, sel_130298}) ? {add_130295, array_index_130232[0]} : sel_130298;
  assign add_130393 = array_index_130343[11:0] + 12'h247;
  assign sel_130395 = $signed({1'h0, add_130315}) < $signed({1'h0, sel_130317}) ? add_130315 : sel_130317;
  assign add_130398 = array_index_130346[11:0] + 12'h247;
  assign sel_130400 = $signed({1'h0, add_130320}) < $signed({1'h0, sel_130322}) ? add_130320 : sel_130322;
  assign array_index_130427 = set1_unflattened[7'h04];
  assign array_index_130430 = set2_unflattened[7'h04];
  assign add_130434 = array_index_130213[11:1] + 11'h79d;
  assign add_130436 = array_index_130214[11:1] + 11'h79d;
  assign add_130438 = array_index_130229[11:1] + 11'h347;
  assign sel_130440 = $signed({1'h0, add_130350, array_index_130213[0]}) < $signed(13'h0fff) ? {add_130350, array_index_130213[0]} : 12'hfff;
  assign add_130442 = array_index_130232[11:1] + 11'h347;
  assign sel_130444 = $signed({1'h0, add_130352, array_index_130214[0]}) < $signed(13'h0fff) ? {add_130352, array_index_130214[0]} : 12'hfff;
  assign add_130446 = array_index_130277[11:3] + 9'h0bd;
  assign sel_130449 = $signed({1'h0, add_130354, array_index_130229[2:0]}) < $signed({1'h0, sel_130357}) ? {add_130354, array_index_130229[2:0]} : sel_130357;
  assign add_130451 = array_index_130280[11:3] + 9'h0bd;
  assign sel_130454 = $signed({1'h0, add_130359, array_index_130232[2:0]}) < $signed({1'h0, sel_130362}) ? {add_130359, array_index_130232[2:0]} : sel_130362;
  assign add_130456 = array_index_130343[11:1] + 11'h247;
  assign sel_130459 = $signed({1'h0, add_130364, array_index_130277[0]}) < $signed({1'h0, sel_130367}) ? {add_130364, array_index_130277[0]} : sel_130367;
  assign add_130461 = array_index_130346[11:1] + 11'h247;
  assign sel_130464 = $signed({1'h0, add_130369, array_index_130280[0]}) < $signed({1'h0, sel_130372}) ? {add_130369, array_index_130280[0]} : sel_130372;
  assign add_130489 = array_index_130427[11:0] + 12'h247;
  assign sel_130491 = $signed({1'h0, add_130393}) < $signed({1'h0, sel_130395}) ? add_130393 : sel_130395;
  assign add_130494 = array_index_130430[11:0] + 12'h247;
  assign sel_130496 = $signed({1'h0, add_130398}) < $signed({1'h0, sel_130400}) ? add_130398 : sel_130400;
  assign array_index_130527 = set1_unflattened[7'h05];
  assign array_index_130530 = set2_unflattened[7'h05];
  assign add_130534 = array_index_130229[11:1] + 11'h79d;
  assign sel_130536 = $signed({1'h0, add_130434, array_index_130213[0]}) < $signed(13'h0fff) ? {add_130434, array_index_130213[0]} : 12'hfff;
  assign add_130538 = array_index_130232[11:1] + 11'h79d;
  assign sel_130540 = $signed({1'h0, add_130436, array_index_130214[0]}) < $signed(13'h0fff) ? {add_130436, array_index_130214[0]} : 12'hfff;
  assign add_130542 = array_index_130277[11:1] + 11'h347;
  assign sel_130544 = $signed({1'h0, add_130438, array_index_130229[0]}) < $signed({1'h0, sel_130440}) ? {add_130438, array_index_130229[0]} : sel_130440;
  assign add_130546 = array_index_130280[11:1] + 11'h347;
  assign sel_130548 = $signed({1'h0, add_130442, array_index_130232[0]}) < $signed({1'h0, sel_130444}) ? {add_130442, array_index_130232[0]} : sel_130444;
  assign add_130550 = array_index_130343[11:3] + 9'h0bd;
  assign sel_130553 = $signed({1'h0, add_130446, array_index_130277[2:0]}) < $signed({1'h0, sel_130449}) ? {add_130446, array_index_130277[2:0]} : sel_130449;
  assign add_130555 = array_index_130346[11:3] + 9'h0bd;
  assign sel_130558 = $signed({1'h0, add_130451, array_index_130280[2:0]}) < $signed({1'h0, sel_130454}) ? {add_130451, array_index_130280[2:0]} : sel_130454;
  assign add_130560 = array_index_130427[11:1] + 11'h247;
  assign sel_130563 = $signed({1'h0, add_130456, array_index_130343[0]}) < $signed({1'h0, sel_130459}) ? {add_130456, array_index_130343[0]} : sel_130459;
  assign add_130565 = array_index_130430[11:1] + 11'h247;
  assign sel_130568 = $signed({1'h0, add_130461, array_index_130346[0]}) < $signed({1'h0, sel_130464}) ? {add_130461, array_index_130346[0]} : sel_130464;
  assign add_130593 = array_index_130527[11:0] + 12'h247;
  assign sel_130595 = $signed({1'h0, add_130489}) < $signed({1'h0, sel_130491}) ? add_130489 : sel_130491;
  assign add_130598 = array_index_130530[11:0] + 12'h247;
  assign sel_130600 = $signed({1'h0, add_130494}) < $signed({1'h0, sel_130496}) ? add_130494 : sel_130496;
  assign array_index_130629 = set1_unflattened[7'h06];
  assign array_index_130632 = set2_unflattened[7'h06];
  assign add_130636 = array_index_130277[11:1] + 11'h79d;
  assign sel_130638 = $signed({1'h0, add_130534, array_index_130229[0]}) < $signed({1'h0, sel_130536}) ? {add_130534, array_index_130229[0]} : sel_130536;
  assign add_130640 = array_index_130280[11:1] + 11'h79d;
  assign sel_130642 = $signed({1'h0, add_130538, array_index_130232[0]}) < $signed({1'h0, sel_130540}) ? {add_130538, array_index_130232[0]} : sel_130540;
  assign add_130644 = array_index_130343[11:1] + 11'h347;
  assign sel_130646 = $signed({1'h0, add_130542, array_index_130277[0]}) < $signed({1'h0, sel_130544}) ? {add_130542, array_index_130277[0]} : sel_130544;
  assign add_130648 = array_index_130346[11:1] + 11'h347;
  assign sel_130650 = $signed({1'h0, add_130546, array_index_130280[0]}) < $signed({1'h0, sel_130548}) ? {add_130546, array_index_130280[0]} : sel_130548;
  assign add_130652 = array_index_130427[11:3] + 9'h0bd;
  assign sel_130655 = $signed({1'h0, add_130550, array_index_130343[2:0]}) < $signed({1'h0, sel_130553}) ? {add_130550, array_index_130343[2:0]} : sel_130553;
  assign add_130657 = array_index_130430[11:3] + 9'h0bd;
  assign sel_130660 = $signed({1'h0, add_130555, array_index_130346[2:0]}) < $signed({1'h0, sel_130558}) ? {add_130555, array_index_130346[2:0]} : sel_130558;
  assign add_130662 = array_index_130527[11:1] + 11'h247;
  assign sel_130665 = $signed({1'h0, add_130560, array_index_130427[0]}) < $signed({1'h0, sel_130563}) ? {add_130560, array_index_130427[0]} : sel_130563;
  assign add_130667 = array_index_130530[11:1] + 11'h247;
  assign sel_130670 = $signed({1'h0, add_130565, array_index_130430[0]}) < $signed({1'h0, sel_130568}) ? {add_130565, array_index_130430[0]} : sel_130568;
  assign add_130695 = array_index_130629[11:0] + 12'h247;
  assign sel_130697 = $signed({1'h0, add_130593}) < $signed({1'h0, sel_130595}) ? add_130593 : sel_130595;
  assign add_130700 = array_index_130632[11:0] + 12'h247;
  assign sel_130702 = $signed({1'h0, add_130598}) < $signed({1'h0, sel_130600}) ? add_130598 : sel_130600;
  assign array_index_130731 = set1_unflattened[7'h07];
  assign array_index_130734 = set2_unflattened[7'h07];
  assign add_130738 = array_index_130343[11:1] + 11'h79d;
  assign sel_130740 = $signed({1'h0, add_130636, array_index_130277[0]}) < $signed({1'h0, sel_130638}) ? {add_130636, array_index_130277[0]} : sel_130638;
  assign add_130742 = array_index_130346[11:1] + 11'h79d;
  assign sel_130744 = $signed({1'h0, add_130640, array_index_130280[0]}) < $signed({1'h0, sel_130642}) ? {add_130640, array_index_130280[0]} : sel_130642;
  assign add_130746 = array_index_130427[11:1] + 11'h347;
  assign sel_130748 = $signed({1'h0, add_130644, array_index_130343[0]}) < $signed({1'h0, sel_130646}) ? {add_130644, array_index_130343[0]} : sel_130646;
  assign add_130750 = array_index_130430[11:1] + 11'h347;
  assign sel_130752 = $signed({1'h0, add_130648, array_index_130346[0]}) < $signed({1'h0, sel_130650}) ? {add_130648, array_index_130346[0]} : sel_130650;
  assign add_130754 = array_index_130527[11:3] + 9'h0bd;
  assign sel_130757 = $signed({1'h0, add_130652, array_index_130427[2:0]}) < $signed({1'h0, sel_130655}) ? {add_130652, array_index_130427[2:0]} : sel_130655;
  assign add_130759 = array_index_130530[11:3] + 9'h0bd;
  assign sel_130762 = $signed({1'h0, add_130657, array_index_130430[2:0]}) < $signed({1'h0, sel_130660}) ? {add_130657, array_index_130430[2:0]} : sel_130660;
  assign add_130764 = array_index_130629[11:1] + 11'h247;
  assign sel_130767 = $signed({1'h0, add_130662, array_index_130527[0]}) < $signed({1'h0, sel_130665}) ? {add_130662, array_index_130527[0]} : sel_130665;
  assign add_130769 = array_index_130632[11:1] + 11'h247;
  assign sel_130772 = $signed({1'h0, add_130667, array_index_130530[0]}) < $signed({1'h0, sel_130670}) ? {add_130667, array_index_130530[0]} : sel_130670;
  assign add_130797 = array_index_130731[11:0] + 12'h247;
  assign sel_130799 = $signed({1'h0, add_130695}) < $signed({1'h0, sel_130697}) ? add_130695 : sel_130697;
  assign add_130802 = array_index_130734[11:0] + 12'h247;
  assign sel_130804 = $signed({1'h0, add_130700}) < $signed({1'h0, sel_130702}) ? add_130700 : sel_130702;
  assign array_index_130833 = set1_unflattened[7'h08];
  assign array_index_130836 = set2_unflattened[7'h08];
  assign add_130840 = array_index_130427[11:1] + 11'h79d;
  assign sel_130842 = $signed({1'h0, add_130738, array_index_130343[0]}) < $signed({1'h0, sel_130740}) ? {add_130738, array_index_130343[0]} : sel_130740;
  assign add_130844 = array_index_130430[11:1] + 11'h79d;
  assign sel_130846 = $signed({1'h0, add_130742, array_index_130346[0]}) < $signed({1'h0, sel_130744}) ? {add_130742, array_index_130346[0]} : sel_130744;
  assign add_130848 = array_index_130527[11:1] + 11'h347;
  assign sel_130850 = $signed({1'h0, add_130746, array_index_130427[0]}) < $signed({1'h0, sel_130748}) ? {add_130746, array_index_130427[0]} : sel_130748;
  assign add_130852 = array_index_130530[11:1] + 11'h347;
  assign sel_130854 = $signed({1'h0, add_130750, array_index_130430[0]}) < $signed({1'h0, sel_130752}) ? {add_130750, array_index_130430[0]} : sel_130752;
  assign add_130856 = array_index_130629[11:3] + 9'h0bd;
  assign sel_130859 = $signed({1'h0, add_130754, array_index_130527[2:0]}) < $signed({1'h0, sel_130757}) ? {add_130754, array_index_130527[2:0]} : sel_130757;
  assign add_130861 = array_index_130632[11:3] + 9'h0bd;
  assign sel_130864 = $signed({1'h0, add_130759, array_index_130530[2:0]}) < $signed({1'h0, sel_130762}) ? {add_130759, array_index_130530[2:0]} : sel_130762;
  assign add_130866 = array_index_130731[11:1] + 11'h247;
  assign sel_130869 = $signed({1'h0, add_130764, array_index_130629[0]}) < $signed({1'h0, sel_130767}) ? {add_130764, array_index_130629[0]} : sel_130767;
  assign add_130871 = array_index_130734[11:1] + 11'h247;
  assign sel_130874 = $signed({1'h0, add_130769, array_index_130632[0]}) < $signed({1'h0, sel_130772}) ? {add_130769, array_index_130632[0]} : sel_130772;
  assign add_130899 = array_index_130833[11:0] + 12'h247;
  assign sel_130901 = $signed({1'h0, add_130797}) < $signed({1'h0, sel_130799}) ? add_130797 : sel_130799;
  assign add_130904 = array_index_130836[11:0] + 12'h247;
  assign sel_130906 = $signed({1'h0, add_130802}) < $signed({1'h0, sel_130804}) ? add_130802 : sel_130804;
  assign array_index_130935 = set1_unflattened[7'h09];
  assign array_index_130938 = set2_unflattened[7'h09];
  assign add_130942 = array_index_130527[11:1] + 11'h79d;
  assign sel_130944 = $signed({1'h0, add_130840, array_index_130427[0]}) < $signed({1'h0, sel_130842}) ? {add_130840, array_index_130427[0]} : sel_130842;
  assign add_130946 = array_index_130530[11:1] + 11'h79d;
  assign sel_130948 = $signed({1'h0, add_130844, array_index_130430[0]}) < $signed({1'h0, sel_130846}) ? {add_130844, array_index_130430[0]} : sel_130846;
  assign add_130950 = array_index_130629[11:1] + 11'h347;
  assign sel_130952 = $signed({1'h0, add_130848, array_index_130527[0]}) < $signed({1'h0, sel_130850}) ? {add_130848, array_index_130527[0]} : sel_130850;
  assign add_130954 = array_index_130632[11:1] + 11'h347;
  assign sel_130956 = $signed({1'h0, add_130852, array_index_130530[0]}) < $signed({1'h0, sel_130854}) ? {add_130852, array_index_130530[0]} : sel_130854;
  assign add_130958 = array_index_130731[11:3] + 9'h0bd;
  assign sel_130961 = $signed({1'h0, add_130856, array_index_130629[2:0]}) < $signed({1'h0, sel_130859}) ? {add_130856, array_index_130629[2:0]} : sel_130859;
  assign add_130963 = array_index_130734[11:3] + 9'h0bd;
  assign sel_130966 = $signed({1'h0, add_130861, array_index_130632[2:0]}) < $signed({1'h0, sel_130864}) ? {add_130861, array_index_130632[2:0]} : sel_130864;
  assign add_130968 = array_index_130833[11:1] + 11'h247;
  assign sel_130971 = $signed({1'h0, add_130866, array_index_130731[0]}) < $signed({1'h0, sel_130869}) ? {add_130866, array_index_130731[0]} : sel_130869;
  assign add_130973 = array_index_130836[11:1] + 11'h247;
  assign sel_130976 = $signed({1'h0, add_130871, array_index_130734[0]}) < $signed({1'h0, sel_130874}) ? {add_130871, array_index_130734[0]} : sel_130874;
  assign add_131001 = array_index_130935[11:0] + 12'h247;
  assign sel_131003 = $signed({1'h0, add_130899}) < $signed({1'h0, sel_130901}) ? add_130899 : sel_130901;
  assign add_131006 = array_index_130938[11:0] + 12'h247;
  assign sel_131008 = $signed({1'h0, add_130904}) < $signed({1'h0, sel_130906}) ? add_130904 : sel_130906;
  assign array_index_131037 = set1_unflattened[7'h0a];
  assign array_index_131040 = set2_unflattened[7'h0a];
  assign add_131044 = array_index_130629[11:1] + 11'h79d;
  assign sel_131046 = $signed({1'h0, add_130942, array_index_130527[0]}) < $signed({1'h0, sel_130944}) ? {add_130942, array_index_130527[0]} : sel_130944;
  assign add_131048 = array_index_130632[11:1] + 11'h79d;
  assign sel_131050 = $signed({1'h0, add_130946, array_index_130530[0]}) < $signed({1'h0, sel_130948}) ? {add_130946, array_index_130530[0]} : sel_130948;
  assign add_131052 = array_index_130731[11:1] + 11'h347;
  assign sel_131054 = $signed({1'h0, add_130950, array_index_130629[0]}) < $signed({1'h0, sel_130952}) ? {add_130950, array_index_130629[0]} : sel_130952;
  assign add_131056 = array_index_130734[11:1] + 11'h347;
  assign sel_131058 = $signed({1'h0, add_130954, array_index_130632[0]}) < $signed({1'h0, sel_130956}) ? {add_130954, array_index_130632[0]} : sel_130956;
  assign add_131060 = array_index_130833[11:3] + 9'h0bd;
  assign sel_131063 = $signed({1'h0, add_130958, array_index_130731[2:0]}) < $signed({1'h0, sel_130961}) ? {add_130958, array_index_130731[2:0]} : sel_130961;
  assign add_131065 = array_index_130836[11:3] + 9'h0bd;
  assign sel_131068 = $signed({1'h0, add_130963, array_index_130734[2:0]}) < $signed({1'h0, sel_130966}) ? {add_130963, array_index_130734[2:0]} : sel_130966;
  assign add_131070 = array_index_130935[11:1] + 11'h247;
  assign sel_131073 = $signed({1'h0, add_130968, array_index_130833[0]}) < $signed({1'h0, sel_130971}) ? {add_130968, array_index_130833[0]} : sel_130971;
  assign add_131075 = array_index_130938[11:1] + 11'h247;
  assign sel_131078 = $signed({1'h0, add_130973, array_index_130836[0]}) < $signed({1'h0, sel_130976}) ? {add_130973, array_index_130836[0]} : sel_130976;
  assign add_131103 = array_index_131037[11:0] + 12'h247;
  assign sel_131105 = $signed({1'h0, add_131001}) < $signed({1'h0, sel_131003}) ? add_131001 : sel_131003;
  assign add_131108 = array_index_131040[11:0] + 12'h247;
  assign sel_131110 = $signed({1'h0, add_131006}) < $signed({1'h0, sel_131008}) ? add_131006 : sel_131008;
  assign array_index_131139 = set1_unflattened[7'h0b];
  assign array_index_131142 = set2_unflattened[7'h0b];
  assign add_131146 = array_index_130731[11:1] + 11'h79d;
  assign sel_131148 = $signed({1'h0, add_131044, array_index_130629[0]}) < $signed({1'h0, sel_131046}) ? {add_131044, array_index_130629[0]} : sel_131046;
  assign add_131150 = array_index_130734[11:1] + 11'h79d;
  assign sel_131152 = $signed({1'h0, add_131048, array_index_130632[0]}) < $signed({1'h0, sel_131050}) ? {add_131048, array_index_130632[0]} : sel_131050;
  assign add_131154 = array_index_130833[11:1] + 11'h347;
  assign sel_131156 = $signed({1'h0, add_131052, array_index_130731[0]}) < $signed({1'h0, sel_131054}) ? {add_131052, array_index_130731[0]} : sel_131054;
  assign add_131158 = array_index_130836[11:1] + 11'h347;
  assign sel_131160 = $signed({1'h0, add_131056, array_index_130734[0]}) < $signed({1'h0, sel_131058}) ? {add_131056, array_index_130734[0]} : sel_131058;
  assign add_131162 = array_index_130935[11:3] + 9'h0bd;
  assign sel_131165 = $signed({1'h0, add_131060, array_index_130833[2:0]}) < $signed({1'h0, sel_131063}) ? {add_131060, array_index_130833[2:0]} : sel_131063;
  assign add_131167 = array_index_130938[11:3] + 9'h0bd;
  assign sel_131170 = $signed({1'h0, add_131065, array_index_130836[2:0]}) < $signed({1'h0, sel_131068}) ? {add_131065, array_index_130836[2:0]} : sel_131068;
  assign add_131172 = array_index_131037[11:1] + 11'h247;
  assign sel_131175 = $signed({1'h0, add_131070, array_index_130935[0]}) < $signed({1'h0, sel_131073}) ? {add_131070, array_index_130935[0]} : sel_131073;
  assign add_131177 = array_index_131040[11:1] + 11'h247;
  assign sel_131180 = $signed({1'h0, add_131075, array_index_130938[0]}) < $signed({1'h0, sel_131078}) ? {add_131075, array_index_130938[0]} : sel_131078;
  assign add_131205 = array_index_131139[11:0] + 12'h247;
  assign sel_131207 = $signed({1'h0, add_131103}) < $signed({1'h0, sel_131105}) ? add_131103 : sel_131105;
  assign add_131210 = array_index_131142[11:0] + 12'h247;
  assign sel_131212 = $signed({1'h0, add_131108}) < $signed({1'h0, sel_131110}) ? add_131108 : sel_131110;
  assign array_index_131241 = set1_unflattened[7'h0c];
  assign array_index_131244 = set2_unflattened[7'h0c];
  assign add_131248 = array_index_130833[11:1] + 11'h79d;
  assign sel_131250 = $signed({1'h0, add_131146, array_index_130731[0]}) < $signed({1'h0, sel_131148}) ? {add_131146, array_index_130731[0]} : sel_131148;
  assign add_131252 = array_index_130836[11:1] + 11'h79d;
  assign sel_131254 = $signed({1'h0, add_131150, array_index_130734[0]}) < $signed({1'h0, sel_131152}) ? {add_131150, array_index_130734[0]} : sel_131152;
  assign add_131256 = array_index_130935[11:1] + 11'h347;
  assign sel_131258 = $signed({1'h0, add_131154, array_index_130833[0]}) < $signed({1'h0, sel_131156}) ? {add_131154, array_index_130833[0]} : sel_131156;
  assign add_131260 = array_index_130938[11:1] + 11'h347;
  assign sel_131262 = $signed({1'h0, add_131158, array_index_130836[0]}) < $signed({1'h0, sel_131160}) ? {add_131158, array_index_130836[0]} : sel_131160;
  assign add_131264 = array_index_131037[11:3] + 9'h0bd;
  assign sel_131267 = $signed({1'h0, add_131162, array_index_130935[2:0]}) < $signed({1'h0, sel_131165}) ? {add_131162, array_index_130935[2:0]} : sel_131165;
  assign add_131269 = array_index_131040[11:3] + 9'h0bd;
  assign sel_131272 = $signed({1'h0, add_131167, array_index_130938[2:0]}) < $signed({1'h0, sel_131170}) ? {add_131167, array_index_130938[2:0]} : sel_131170;
  assign add_131274 = array_index_131139[11:1] + 11'h247;
  assign sel_131277 = $signed({1'h0, add_131172, array_index_131037[0]}) < $signed({1'h0, sel_131175}) ? {add_131172, array_index_131037[0]} : sel_131175;
  assign add_131279 = array_index_131142[11:1] + 11'h247;
  assign sel_131282 = $signed({1'h0, add_131177, array_index_131040[0]}) < $signed({1'h0, sel_131180}) ? {add_131177, array_index_131040[0]} : sel_131180;
  assign add_131307 = array_index_131241[11:0] + 12'h247;
  assign sel_131309 = $signed({1'h0, add_131205}) < $signed({1'h0, sel_131207}) ? add_131205 : sel_131207;
  assign add_131312 = array_index_131244[11:0] + 12'h247;
  assign sel_131314 = $signed({1'h0, add_131210}) < $signed({1'h0, sel_131212}) ? add_131210 : sel_131212;
  assign array_index_131343 = set1_unflattened[7'h0d];
  assign array_index_131346 = set2_unflattened[7'h0d];
  assign add_131350 = array_index_130935[11:1] + 11'h79d;
  assign sel_131352 = $signed({1'h0, add_131248, array_index_130833[0]}) < $signed({1'h0, sel_131250}) ? {add_131248, array_index_130833[0]} : sel_131250;
  assign add_131354 = array_index_130938[11:1] + 11'h79d;
  assign sel_131356 = $signed({1'h0, add_131252, array_index_130836[0]}) < $signed({1'h0, sel_131254}) ? {add_131252, array_index_130836[0]} : sel_131254;
  assign add_131358 = array_index_131037[11:1] + 11'h347;
  assign sel_131360 = $signed({1'h0, add_131256, array_index_130935[0]}) < $signed({1'h0, sel_131258}) ? {add_131256, array_index_130935[0]} : sel_131258;
  assign add_131362 = array_index_131040[11:1] + 11'h347;
  assign sel_131364 = $signed({1'h0, add_131260, array_index_130938[0]}) < $signed({1'h0, sel_131262}) ? {add_131260, array_index_130938[0]} : sel_131262;
  assign add_131366 = array_index_131139[11:3] + 9'h0bd;
  assign sel_131369 = $signed({1'h0, add_131264, array_index_131037[2:0]}) < $signed({1'h0, sel_131267}) ? {add_131264, array_index_131037[2:0]} : sel_131267;
  assign add_131371 = array_index_131142[11:3] + 9'h0bd;
  assign sel_131374 = $signed({1'h0, add_131269, array_index_131040[2:0]}) < $signed({1'h0, sel_131272}) ? {add_131269, array_index_131040[2:0]} : sel_131272;
  assign add_131376 = array_index_131241[11:1] + 11'h247;
  assign sel_131379 = $signed({1'h0, add_131274, array_index_131139[0]}) < $signed({1'h0, sel_131277}) ? {add_131274, array_index_131139[0]} : sel_131277;
  assign add_131381 = array_index_131244[11:1] + 11'h247;
  assign sel_131384 = $signed({1'h0, add_131279, array_index_131142[0]}) < $signed({1'h0, sel_131282}) ? {add_131279, array_index_131142[0]} : sel_131282;
  assign add_131409 = array_index_131343[11:0] + 12'h247;
  assign sel_131411 = $signed({1'h0, add_131307}) < $signed({1'h0, sel_131309}) ? add_131307 : sel_131309;
  assign add_131414 = array_index_131346[11:0] + 12'h247;
  assign sel_131416 = $signed({1'h0, add_131312}) < $signed({1'h0, sel_131314}) ? add_131312 : sel_131314;
  assign array_index_131445 = set1_unflattened[7'h0e];
  assign array_index_131448 = set2_unflattened[7'h0e];
  assign add_131452 = array_index_131037[11:1] + 11'h79d;
  assign sel_131454 = $signed({1'h0, add_131350, array_index_130935[0]}) < $signed({1'h0, sel_131352}) ? {add_131350, array_index_130935[0]} : sel_131352;
  assign add_131456 = array_index_131040[11:1] + 11'h79d;
  assign sel_131458 = $signed({1'h0, add_131354, array_index_130938[0]}) < $signed({1'h0, sel_131356}) ? {add_131354, array_index_130938[0]} : sel_131356;
  assign add_131460 = array_index_131139[11:1] + 11'h347;
  assign sel_131462 = $signed({1'h0, add_131358, array_index_131037[0]}) < $signed({1'h0, sel_131360}) ? {add_131358, array_index_131037[0]} : sel_131360;
  assign add_131464 = array_index_131142[11:1] + 11'h347;
  assign sel_131466 = $signed({1'h0, add_131362, array_index_131040[0]}) < $signed({1'h0, sel_131364}) ? {add_131362, array_index_131040[0]} : sel_131364;
  assign add_131468 = array_index_131241[11:3] + 9'h0bd;
  assign sel_131471 = $signed({1'h0, add_131366, array_index_131139[2:0]}) < $signed({1'h0, sel_131369}) ? {add_131366, array_index_131139[2:0]} : sel_131369;
  assign add_131473 = array_index_131244[11:3] + 9'h0bd;
  assign sel_131476 = $signed({1'h0, add_131371, array_index_131142[2:0]}) < $signed({1'h0, sel_131374}) ? {add_131371, array_index_131142[2:0]} : sel_131374;
  assign add_131478 = array_index_131343[11:1] + 11'h247;
  assign sel_131481 = $signed({1'h0, add_131376, array_index_131241[0]}) < $signed({1'h0, sel_131379}) ? {add_131376, array_index_131241[0]} : sel_131379;
  assign add_131483 = array_index_131346[11:1] + 11'h247;
  assign sel_131486 = $signed({1'h0, add_131381, array_index_131244[0]}) < $signed({1'h0, sel_131384}) ? {add_131381, array_index_131244[0]} : sel_131384;
  assign add_131511 = array_index_131445[11:0] + 12'h247;
  assign sel_131513 = $signed({1'h0, add_131409}) < $signed({1'h0, sel_131411}) ? add_131409 : sel_131411;
  assign add_131516 = array_index_131448[11:0] + 12'h247;
  assign sel_131518 = $signed({1'h0, add_131414}) < $signed({1'h0, sel_131416}) ? add_131414 : sel_131416;
  assign array_index_131547 = set1_unflattened[7'h0f];
  assign array_index_131550 = set2_unflattened[7'h0f];
  assign add_131554 = array_index_131139[11:1] + 11'h79d;
  assign sel_131556 = $signed({1'h0, add_131452, array_index_131037[0]}) < $signed({1'h0, sel_131454}) ? {add_131452, array_index_131037[0]} : sel_131454;
  assign add_131558 = array_index_131142[11:1] + 11'h79d;
  assign sel_131560 = $signed({1'h0, add_131456, array_index_131040[0]}) < $signed({1'h0, sel_131458}) ? {add_131456, array_index_131040[0]} : sel_131458;
  assign add_131562 = array_index_131241[11:1] + 11'h347;
  assign sel_131564 = $signed({1'h0, add_131460, array_index_131139[0]}) < $signed({1'h0, sel_131462}) ? {add_131460, array_index_131139[0]} : sel_131462;
  assign add_131566 = array_index_131244[11:1] + 11'h347;
  assign sel_131568 = $signed({1'h0, add_131464, array_index_131142[0]}) < $signed({1'h0, sel_131466}) ? {add_131464, array_index_131142[0]} : sel_131466;
  assign add_131570 = array_index_131343[11:3] + 9'h0bd;
  assign sel_131573 = $signed({1'h0, add_131468, array_index_131241[2:0]}) < $signed({1'h0, sel_131471}) ? {add_131468, array_index_131241[2:0]} : sel_131471;
  assign add_131575 = array_index_131346[11:3] + 9'h0bd;
  assign sel_131578 = $signed({1'h0, add_131473, array_index_131244[2:0]}) < $signed({1'h0, sel_131476}) ? {add_131473, array_index_131244[2:0]} : sel_131476;
  assign add_131580 = array_index_131445[11:1] + 11'h247;
  assign sel_131583 = $signed({1'h0, add_131478, array_index_131343[0]}) < $signed({1'h0, sel_131481}) ? {add_131478, array_index_131343[0]} : sel_131481;
  assign add_131585 = array_index_131448[11:1] + 11'h247;
  assign sel_131588 = $signed({1'h0, add_131483, array_index_131346[0]}) < $signed({1'h0, sel_131486}) ? {add_131483, array_index_131346[0]} : sel_131486;
  assign add_131613 = array_index_131547[11:0] + 12'h247;
  assign sel_131615 = $signed({1'h0, add_131511}) < $signed({1'h0, sel_131513}) ? add_131511 : sel_131513;
  assign add_131618 = array_index_131550[11:0] + 12'h247;
  assign sel_131620 = $signed({1'h0, add_131516}) < $signed({1'h0, sel_131518}) ? add_131516 : sel_131518;
  assign array_index_131649 = set1_unflattened[7'h10];
  assign array_index_131652 = set2_unflattened[7'h10];
  assign add_131656 = array_index_131241[11:1] + 11'h79d;
  assign sel_131658 = $signed({1'h0, add_131554, array_index_131139[0]}) < $signed({1'h0, sel_131556}) ? {add_131554, array_index_131139[0]} : sel_131556;
  assign add_131660 = array_index_131244[11:1] + 11'h79d;
  assign sel_131662 = $signed({1'h0, add_131558, array_index_131142[0]}) < $signed({1'h0, sel_131560}) ? {add_131558, array_index_131142[0]} : sel_131560;
  assign add_131664 = array_index_131343[11:1] + 11'h347;
  assign sel_131666 = $signed({1'h0, add_131562, array_index_131241[0]}) < $signed({1'h0, sel_131564}) ? {add_131562, array_index_131241[0]} : sel_131564;
  assign add_131668 = array_index_131346[11:1] + 11'h347;
  assign sel_131670 = $signed({1'h0, add_131566, array_index_131244[0]}) < $signed({1'h0, sel_131568}) ? {add_131566, array_index_131244[0]} : sel_131568;
  assign add_131672 = array_index_131445[11:3] + 9'h0bd;
  assign sel_131675 = $signed({1'h0, add_131570, array_index_131343[2:0]}) < $signed({1'h0, sel_131573}) ? {add_131570, array_index_131343[2:0]} : sel_131573;
  assign add_131677 = array_index_131448[11:3] + 9'h0bd;
  assign sel_131680 = $signed({1'h0, add_131575, array_index_131346[2:0]}) < $signed({1'h0, sel_131578}) ? {add_131575, array_index_131346[2:0]} : sel_131578;
  assign add_131682 = array_index_131547[11:1] + 11'h247;
  assign sel_131685 = $signed({1'h0, add_131580, array_index_131445[0]}) < $signed({1'h0, sel_131583}) ? {add_131580, array_index_131445[0]} : sel_131583;
  assign add_131687 = array_index_131550[11:1] + 11'h247;
  assign sel_131690 = $signed({1'h0, add_131585, array_index_131448[0]}) < $signed({1'h0, sel_131588}) ? {add_131585, array_index_131448[0]} : sel_131588;
  assign add_131715 = array_index_131649[11:0] + 12'h247;
  assign sel_131717 = $signed({1'h0, add_131613}) < $signed({1'h0, sel_131615}) ? add_131613 : sel_131615;
  assign add_131720 = array_index_131652[11:0] + 12'h247;
  assign sel_131722 = $signed({1'h0, add_131618}) < $signed({1'h0, sel_131620}) ? add_131618 : sel_131620;
  assign array_index_131751 = set1_unflattened[7'h11];
  assign array_index_131754 = set2_unflattened[7'h11];
  assign add_131758 = array_index_131343[11:1] + 11'h79d;
  assign sel_131760 = $signed({1'h0, add_131656, array_index_131241[0]}) < $signed({1'h0, sel_131658}) ? {add_131656, array_index_131241[0]} : sel_131658;
  assign add_131762 = array_index_131346[11:1] + 11'h79d;
  assign sel_131764 = $signed({1'h0, add_131660, array_index_131244[0]}) < $signed({1'h0, sel_131662}) ? {add_131660, array_index_131244[0]} : sel_131662;
  assign add_131766 = array_index_131445[11:1] + 11'h347;
  assign sel_131768 = $signed({1'h0, add_131664, array_index_131343[0]}) < $signed({1'h0, sel_131666}) ? {add_131664, array_index_131343[0]} : sel_131666;
  assign add_131770 = array_index_131448[11:1] + 11'h347;
  assign sel_131772 = $signed({1'h0, add_131668, array_index_131346[0]}) < $signed({1'h0, sel_131670}) ? {add_131668, array_index_131346[0]} : sel_131670;
  assign add_131774 = array_index_131547[11:3] + 9'h0bd;
  assign sel_131777 = $signed({1'h0, add_131672, array_index_131445[2:0]}) < $signed({1'h0, sel_131675}) ? {add_131672, array_index_131445[2:0]} : sel_131675;
  assign add_131779 = array_index_131550[11:3] + 9'h0bd;
  assign sel_131782 = $signed({1'h0, add_131677, array_index_131448[2:0]}) < $signed({1'h0, sel_131680}) ? {add_131677, array_index_131448[2:0]} : sel_131680;
  assign add_131784 = array_index_131649[11:1] + 11'h247;
  assign sel_131787 = $signed({1'h0, add_131682, array_index_131547[0]}) < $signed({1'h0, sel_131685}) ? {add_131682, array_index_131547[0]} : sel_131685;
  assign add_131789 = array_index_131652[11:1] + 11'h247;
  assign sel_131792 = $signed({1'h0, add_131687, array_index_131550[0]}) < $signed({1'h0, sel_131690}) ? {add_131687, array_index_131550[0]} : sel_131690;
  assign add_131817 = array_index_131751[11:0] + 12'h247;
  assign sel_131819 = $signed({1'h0, add_131715}) < $signed({1'h0, sel_131717}) ? add_131715 : sel_131717;
  assign add_131822 = array_index_131754[11:0] + 12'h247;
  assign sel_131824 = $signed({1'h0, add_131720}) < $signed({1'h0, sel_131722}) ? add_131720 : sel_131722;
  assign array_index_131853 = set1_unflattened[7'h12];
  assign array_index_131856 = set2_unflattened[7'h12];
  assign add_131860 = array_index_131445[11:1] + 11'h79d;
  assign sel_131862 = $signed({1'h0, add_131758, array_index_131343[0]}) < $signed({1'h0, sel_131760}) ? {add_131758, array_index_131343[0]} : sel_131760;
  assign add_131864 = array_index_131448[11:1] + 11'h79d;
  assign sel_131866 = $signed({1'h0, add_131762, array_index_131346[0]}) < $signed({1'h0, sel_131764}) ? {add_131762, array_index_131346[0]} : sel_131764;
  assign add_131868 = array_index_131547[11:1] + 11'h347;
  assign sel_131870 = $signed({1'h0, add_131766, array_index_131445[0]}) < $signed({1'h0, sel_131768}) ? {add_131766, array_index_131445[0]} : sel_131768;
  assign add_131872 = array_index_131550[11:1] + 11'h347;
  assign sel_131874 = $signed({1'h0, add_131770, array_index_131448[0]}) < $signed({1'h0, sel_131772}) ? {add_131770, array_index_131448[0]} : sel_131772;
  assign add_131876 = array_index_131649[11:3] + 9'h0bd;
  assign sel_131879 = $signed({1'h0, add_131774, array_index_131547[2:0]}) < $signed({1'h0, sel_131777}) ? {add_131774, array_index_131547[2:0]} : sel_131777;
  assign add_131881 = array_index_131652[11:3] + 9'h0bd;
  assign sel_131884 = $signed({1'h0, add_131779, array_index_131550[2:0]}) < $signed({1'h0, sel_131782}) ? {add_131779, array_index_131550[2:0]} : sel_131782;
  assign add_131886 = array_index_131751[11:1] + 11'h247;
  assign sel_131889 = $signed({1'h0, add_131784, array_index_131649[0]}) < $signed({1'h0, sel_131787}) ? {add_131784, array_index_131649[0]} : sel_131787;
  assign add_131891 = array_index_131754[11:1] + 11'h247;
  assign sel_131894 = $signed({1'h0, add_131789, array_index_131652[0]}) < $signed({1'h0, sel_131792}) ? {add_131789, array_index_131652[0]} : sel_131792;
  assign add_131919 = array_index_131853[11:0] + 12'h247;
  assign sel_131921 = $signed({1'h0, add_131817}) < $signed({1'h0, sel_131819}) ? add_131817 : sel_131819;
  assign add_131924 = array_index_131856[11:0] + 12'h247;
  assign sel_131926 = $signed({1'h0, add_131822}) < $signed({1'h0, sel_131824}) ? add_131822 : sel_131824;
  assign array_index_131955 = set1_unflattened[7'h13];
  assign array_index_131958 = set2_unflattened[7'h13];
  assign add_131962 = array_index_131547[11:1] + 11'h79d;
  assign sel_131964 = $signed({1'h0, add_131860, array_index_131445[0]}) < $signed({1'h0, sel_131862}) ? {add_131860, array_index_131445[0]} : sel_131862;
  assign add_131966 = array_index_131550[11:1] + 11'h79d;
  assign sel_131968 = $signed({1'h0, add_131864, array_index_131448[0]}) < $signed({1'h0, sel_131866}) ? {add_131864, array_index_131448[0]} : sel_131866;
  assign add_131970 = array_index_131649[11:1] + 11'h347;
  assign sel_131972 = $signed({1'h0, add_131868, array_index_131547[0]}) < $signed({1'h0, sel_131870}) ? {add_131868, array_index_131547[0]} : sel_131870;
  assign add_131974 = array_index_131652[11:1] + 11'h347;
  assign sel_131976 = $signed({1'h0, add_131872, array_index_131550[0]}) < $signed({1'h0, sel_131874}) ? {add_131872, array_index_131550[0]} : sel_131874;
  assign add_131978 = array_index_131751[11:3] + 9'h0bd;
  assign sel_131981 = $signed({1'h0, add_131876, array_index_131649[2:0]}) < $signed({1'h0, sel_131879}) ? {add_131876, array_index_131649[2:0]} : sel_131879;
  assign add_131983 = array_index_131754[11:3] + 9'h0bd;
  assign sel_131986 = $signed({1'h0, add_131881, array_index_131652[2:0]}) < $signed({1'h0, sel_131884}) ? {add_131881, array_index_131652[2:0]} : sel_131884;
  assign add_131988 = array_index_131853[11:1] + 11'h247;
  assign sel_131991 = $signed({1'h0, add_131886, array_index_131751[0]}) < $signed({1'h0, sel_131889}) ? {add_131886, array_index_131751[0]} : sel_131889;
  assign add_131993 = array_index_131856[11:1] + 11'h247;
  assign sel_131996 = $signed({1'h0, add_131891, array_index_131754[0]}) < $signed({1'h0, sel_131894}) ? {add_131891, array_index_131754[0]} : sel_131894;
  assign add_132021 = array_index_131955[11:0] + 12'h247;
  assign sel_132023 = $signed({1'h0, add_131919}) < $signed({1'h0, sel_131921}) ? add_131919 : sel_131921;
  assign add_132026 = array_index_131958[11:0] + 12'h247;
  assign sel_132028 = $signed({1'h0, add_131924}) < $signed({1'h0, sel_131926}) ? add_131924 : sel_131926;
  assign array_index_132057 = set1_unflattened[7'h14];
  assign array_index_132060 = set2_unflattened[7'h14];
  assign add_132064 = array_index_131649[11:1] + 11'h79d;
  assign sel_132066 = $signed({1'h0, add_131962, array_index_131547[0]}) < $signed({1'h0, sel_131964}) ? {add_131962, array_index_131547[0]} : sel_131964;
  assign add_132068 = array_index_131652[11:1] + 11'h79d;
  assign sel_132070 = $signed({1'h0, add_131966, array_index_131550[0]}) < $signed({1'h0, sel_131968}) ? {add_131966, array_index_131550[0]} : sel_131968;
  assign add_132072 = array_index_131751[11:1] + 11'h347;
  assign sel_132074 = $signed({1'h0, add_131970, array_index_131649[0]}) < $signed({1'h0, sel_131972}) ? {add_131970, array_index_131649[0]} : sel_131972;
  assign add_132076 = array_index_131754[11:1] + 11'h347;
  assign sel_132078 = $signed({1'h0, add_131974, array_index_131652[0]}) < $signed({1'h0, sel_131976}) ? {add_131974, array_index_131652[0]} : sel_131976;
  assign add_132080 = array_index_131853[11:3] + 9'h0bd;
  assign sel_132083 = $signed({1'h0, add_131978, array_index_131751[2:0]}) < $signed({1'h0, sel_131981}) ? {add_131978, array_index_131751[2:0]} : sel_131981;
  assign add_132085 = array_index_131856[11:3] + 9'h0bd;
  assign sel_132088 = $signed({1'h0, add_131983, array_index_131754[2:0]}) < $signed({1'h0, sel_131986}) ? {add_131983, array_index_131754[2:0]} : sel_131986;
  assign add_132090 = array_index_131955[11:1] + 11'h247;
  assign sel_132093 = $signed({1'h0, add_131988, array_index_131853[0]}) < $signed({1'h0, sel_131991}) ? {add_131988, array_index_131853[0]} : sel_131991;
  assign add_132095 = array_index_131958[11:1] + 11'h247;
  assign sel_132098 = $signed({1'h0, add_131993, array_index_131856[0]}) < $signed({1'h0, sel_131996}) ? {add_131993, array_index_131856[0]} : sel_131996;
  assign add_132123 = array_index_132057[11:0] + 12'h247;
  assign sel_132125 = $signed({1'h0, add_132021}) < $signed({1'h0, sel_132023}) ? add_132021 : sel_132023;
  assign add_132128 = array_index_132060[11:0] + 12'h247;
  assign sel_132130 = $signed({1'h0, add_132026}) < $signed({1'h0, sel_132028}) ? add_132026 : sel_132028;
  assign array_index_132159 = set1_unflattened[7'h15];
  assign array_index_132162 = set2_unflattened[7'h15];
  assign add_132166 = array_index_131751[11:1] + 11'h79d;
  assign sel_132168 = $signed({1'h0, add_132064, array_index_131649[0]}) < $signed({1'h0, sel_132066}) ? {add_132064, array_index_131649[0]} : sel_132066;
  assign add_132170 = array_index_131754[11:1] + 11'h79d;
  assign sel_132172 = $signed({1'h0, add_132068, array_index_131652[0]}) < $signed({1'h0, sel_132070}) ? {add_132068, array_index_131652[0]} : sel_132070;
  assign add_132174 = array_index_131853[11:1] + 11'h347;
  assign sel_132176 = $signed({1'h0, add_132072, array_index_131751[0]}) < $signed({1'h0, sel_132074}) ? {add_132072, array_index_131751[0]} : sel_132074;
  assign add_132178 = array_index_131856[11:1] + 11'h347;
  assign sel_132180 = $signed({1'h0, add_132076, array_index_131754[0]}) < $signed({1'h0, sel_132078}) ? {add_132076, array_index_131754[0]} : sel_132078;
  assign add_132182 = array_index_131955[11:3] + 9'h0bd;
  assign sel_132185 = $signed({1'h0, add_132080, array_index_131853[2:0]}) < $signed({1'h0, sel_132083}) ? {add_132080, array_index_131853[2:0]} : sel_132083;
  assign add_132187 = array_index_131958[11:3] + 9'h0bd;
  assign sel_132190 = $signed({1'h0, add_132085, array_index_131856[2:0]}) < $signed({1'h0, sel_132088}) ? {add_132085, array_index_131856[2:0]} : sel_132088;
  assign add_132192 = array_index_132057[11:1] + 11'h247;
  assign sel_132195 = $signed({1'h0, add_132090, array_index_131955[0]}) < $signed({1'h0, sel_132093}) ? {add_132090, array_index_131955[0]} : sel_132093;
  assign add_132197 = array_index_132060[11:1] + 11'h247;
  assign sel_132200 = $signed({1'h0, add_132095, array_index_131958[0]}) < $signed({1'h0, sel_132098}) ? {add_132095, array_index_131958[0]} : sel_132098;
  assign add_132225 = array_index_132159[11:0] + 12'h247;
  assign sel_132227 = $signed({1'h0, add_132123}) < $signed({1'h0, sel_132125}) ? add_132123 : sel_132125;
  assign add_132230 = array_index_132162[11:0] + 12'h247;
  assign sel_132232 = $signed({1'h0, add_132128}) < $signed({1'h0, sel_132130}) ? add_132128 : sel_132130;
  assign array_index_132261 = set1_unflattened[7'h16];
  assign array_index_132264 = set2_unflattened[7'h16];
  assign add_132268 = array_index_131853[11:1] + 11'h79d;
  assign sel_132270 = $signed({1'h0, add_132166, array_index_131751[0]}) < $signed({1'h0, sel_132168}) ? {add_132166, array_index_131751[0]} : sel_132168;
  assign add_132272 = array_index_131856[11:1] + 11'h79d;
  assign sel_132274 = $signed({1'h0, add_132170, array_index_131754[0]}) < $signed({1'h0, sel_132172}) ? {add_132170, array_index_131754[0]} : sel_132172;
  assign add_132276 = array_index_131955[11:1] + 11'h347;
  assign sel_132278 = $signed({1'h0, add_132174, array_index_131853[0]}) < $signed({1'h0, sel_132176}) ? {add_132174, array_index_131853[0]} : sel_132176;
  assign add_132280 = array_index_131958[11:1] + 11'h347;
  assign sel_132282 = $signed({1'h0, add_132178, array_index_131856[0]}) < $signed({1'h0, sel_132180}) ? {add_132178, array_index_131856[0]} : sel_132180;
  assign add_132284 = array_index_132057[11:3] + 9'h0bd;
  assign sel_132287 = $signed({1'h0, add_132182, array_index_131955[2:0]}) < $signed({1'h0, sel_132185}) ? {add_132182, array_index_131955[2:0]} : sel_132185;
  assign add_132289 = array_index_132060[11:3] + 9'h0bd;
  assign sel_132292 = $signed({1'h0, add_132187, array_index_131958[2:0]}) < $signed({1'h0, sel_132190}) ? {add_132187, array_index_131958[2:0]} : sel_132190;
  assign add_132294 = array_index_132159[11:1] + 11'h247;
  assign sel_132297 = $signed({1'h0, add_132192, array_index_132057[0]}) < $signed({1'h0, sel_132195}) ? {add_132192, array_index_132057[0]} : sel_132195;
  assign add_132299 = array_index_132162[11:1] + 11'h247;
  assign sel_132302 = $signed({1'h0, add_132197, array_index_132060[0]}) < $signed({1'h0, sel_132200}) ? {add_132197, array_index_132060[0]} : sel_132200;
  assign add_132327 = array_index_132261[11:0] + 12'h247;
  assign sel_132329 = $signed({1'h0, add_132225}) < $signed({1'h0, sel_132227}) ? add_132225 : sel_132227;
  assign add_132332 = array_index_132264[11:0] + 12'h247;
  assign sel_132334 = $signed({1'h0, add_132230}) < $signed({1'h0, sel_132232}) ? add_132230 : sel_132232;
  assign array_index_132363 = set1_unflattened[7'h17];
  assign array_index_132366 = set2_unflattened[7'h17];
  assign add_132370 = array_index_131955[11:1] + 11'h79d;
  assign sel_132372 = $signed({1'h0, add_132268, array_index_131853[0]}) < $signed({1'h0, sel_132270}) ? {add_132268, array_index_131853[0]} : sel_132270;
  assign add_132374 = array_index_131958[11:1] + 11'h79d;
  assign sel_132376 = $signed({1'h0, add_132272, array_index_131856[0]}) < $signed({1'h0, sel_132274}) ? {add_132272, array_index_131856[0]} : sel_132274;
  assign add_132378 = array_index_132057[11:1] + 11'h347;
  assign sel_132380 = $signed({1'h0, add_132276, array_index_131955[0]}) < $signed({1'h0, sel_132278}) ? {add_132276, array_index_131955[0]} : sel_132278;
  assign add_132382 = array_index_132060[11:1] + 11'h347;
  assign sel_132384 = $signed({1'h0, add_132280, array_index_131958[0]}) < $signed({1'h0, sel_132282}) ? {add_132280, array_index_131958[0]} : sel_132282;
  assign add_132386 = array_index_132159[11:3] + 9'h0bd;
  assign sel_132389 = $signed({1'h0, add_132284, array_index_132057[2:0]}) < $signed({1'h0, sel_132287}) ? {add_132284, array_index_132057[2:0]} : sel_132287;
  assign add_132391 = array_index_132162[11:3] + 9'h0bd;
  assign sel_132394 = $signed({1'h0, add_132289, array_index_132060[2:0]}) < $signed({1'h0, sel_132292}) ? {add_132289, array_index_132060[2:0]} : sel_132292;
  assign add_132396 = array_index_132261[11:1] + 11'h247;
  assign sel_132399 = $signed({1'h0, add_132294, array_index_132159[0]}) < $signed({1'h0, sel_132297}) ? {add_132294, array_index_132159[0]} : sel_132297;
  assign add_132401 = array_index_132264[11:1] + 11'h247;
  assign sel_132404 = $signed({1'h0, add_132299, array_index_132162[0]}) < $signed({1'h0, sel_132302}) ? {add_132299, array_index_132162[0]} : sel_132302;
  assign add_132429 = array_index_132363[11:0] + 12'h247;
  assign sel_132431 = $signed({1'h0, add_132327}) < $signed({1'h0, sel_132329}) ? add_132327 : sel_132329;
  assign add_132434 = array_index_132366[11:0] + 12'h247;
  assign sel_132436 = $signed({1'h0, add_132332}) < $signed({1'h0, sel_132334}) ? add_132332 : sel_132334;
  assign array_index_132465 = set1_unflattened[7'h18];
  assign array_index_132468 = set2_unflattened[7'h18];
  assign add_132472 = array_index_132057[11:1] + 11'h79d;
  assign sel_132474 = $signed({1'h0, add_132370, array_index_131955[0]}) < $signed({1'h0, sel_132372}) ? {add_132370, array_index_131955[0]} : sel_132372;
  assign add_132476 = array_index_132060[11:1] + 11'h79d;
  assign sel_132478 = $signed({1'h0, add_132374, array_index_131958[0]}) < $signed({1'h0, sel_132376}) ? {add_132374, array_index_131958[0]} : sel_132376;
  assign add_132480 = array_index_132159[11:1] + 11'h347;
  assign sel_132482 = $signed({1'h0, add_132378, array_index_132057[0]}) < $signed({1'h0, sel_132380}) ? {add_132378, array_index_132057[0]} : sel_132380;
  assign add_132484 = array_index_132162[11:1] + 11'h347;
  assign sel_132486 = $signed({1'h0, add_132382, array_index_132060[0]}) < $signed({1'h0, sel_132384}) ? {add_132382, array_index_132060[0]} : sel_132384;
  assign add_132488 = array_index_132261[11:3] + 9'h0bd;
  assign sel_132491 = $signed({1'h0, add_132386, array_index_132159[2:0]}) < $signed({1'h0, sel_132389}) ? {add_132386, array_index_132159[2:0]} : sel_132389;
  assign add_132493 = array_index_132264[11:3] + 9'h0bd;
  assign sel_132496 = $signed({1'h0, add_132391, array_index_132162[2:0]}) < $signed({1'h0, sel_132394}) ? {add_132391, array_index_132162[2:0]} : sel_132394;
  assign add_132498 = array_index_132363[11:1] + 11'h247;
  assign sel_132501 = $signed({1'h0, add_132396, array_index_132261[0]}) < $signed({1'h0, sel_132399}) ? {add_132396, array_index_132261[0]} : sel_132399;
  assign add_132503 = array_index_132366[11:1] + 11'h247;
  assign sel_132506 = $signed({1'h0, add_132401, array_index_132264[0]}) < $signed({1'h0, sel_132404}) ? {add_132401, array_index_132264[0]} : sel_132404;
  assign add_132531 = array_index_132465[11:0] + 12'h247;
  assign sel_132533 = $signed({1'h0, add_132429}) < $signed({1'h0, sel_132431}) ? add_132429 : sel_132431;
  assign add_132536 = array_index_132468[11:0] + 12'h247;
  assign sel_132538 = $signed({1'h0, add_132434}) < $signed({1'h0, sel_132436}) ? add_132434 : sel_132436;
  assign array_index_132567 = set1_unflattened[7'h19];
  assign array_index_132570 = set2_unflattened[7'h19];
  assign add_132574 = array_index_132159[11:1] + 11'h79d;
  assign sel_132576 = $signed({1'h0, add_132472, array_index_132057[0]}) < $signed({1'h0, sel_132474}) ? {add_132472, array_index_132057[0]} : sel_132474;
  assign add_132578 = array_index_132162[11:1] + 11'h79d;
  assign sel_132580 = $signed({1'h0, add_132476, array_index_132060[0]}) < $signed({1'h0, sel_132478}) ? {add_132476, array_index_132060[0]} : sel_132478;
  assign add_132582 = array_index_132261[11:1] + 11'h347;
  assign sel_132584 = $signed({1'h0, add_132480, array_index_132159[0]}) < $signed({1'h0, sel_132482}) ? {add_132480, array_index_132159[0]} : sel_132482;
  assign add_132586 = array_index_132264[11:1] + 11'h347;
  assign sel_132588 = $signed({1'h0, add_132484, array_index_132162[0]}) < $signed({1'h0, sel_132486}) ? {add_132484, array_index_132162[0]} : sel_132486;
  assign add_132590 = array_index_132363[11:3] + 9'h0bd;
  assign sel_132593 = $signed({1'h0, add_132488, array_index_132261[2:0]}) < $signed({1'h0, sel_132491}) ? {add_132488, array_index_132261[2:0]} : sel_132491;
  assign add_132595 = array_index_132366[11:3] + 9'h0bd;
  assign sel_132598 = $signed({1'h0, add_132493, array_index_132264[2:0]}) < $signed({1'h0, sel_132496}) ? {add_132493, array_index_132264[2:0]} : sel_132496;
  assign add_132600 = array_index_132465[11:1] + 11'h247;
  assign sel_132603 = $signed({1'h0, add_132498, array_index_132363[0]}) < $signed({1'h0, sel_132501}) ? {add_132498, array_index_132363[0]} : sel_132501;
  assign add_132605 = array_index_132468[11:1] + 11'h247;
  assign sel_132608 = $signed({1'h0, add_132503, array_index_132366[0]}) < $signed({1'h0, sel_132506}) ? {add_132503, array_index_132366[0]} : sel_132506;
  assign add_132633 = array_index_132567[11:0] + 12'h247;
  assign sel_132635 = $signed({1'h0, add_132531}) < $signed({1'h0, sel_132533}) ? add_132531 : sel_132533;
  assign add_132638 = array_index_132570[11:0] + 12'h247;
  assign sel_132640 = $signed({1'h0, add_132536}) < $signed({1'h0, sel_132538}) ? add_132536 : sel_132538;
  assign array_index_132669 = set1_unflattened[7'h1a];
  assign array_index_132672 = set2_unflattened[7'h1a];
  assign add_132676 = array_index_132261[11:1] + 11'h79d;
  assign sel_132678 = $signed({1'h0, add_132574, array_index_132159[0]}) < $signed({1'h0, sel_132576}) ? {add_132574, array_index_132159[0]} : sel_132576;
  assign add_132680 = array_index_132264[11:1] + 11'h79d;
  assign sel_132682 = $signed({1'h0, add_132578, array_index_132162[0]}) < $signed({1'h0, sel_132580}) ? {add_132578, array_index_132162[0]} : sel_132580;
  assign add_132684 = array_index_132363[11:1] + 11'h347;
  assign sel_132686 = $signed({1'h0, add_132582, array_index_132261[0]}) < $signed({1'h0, sel_132584}) ? {add_132582, array_index_132261[0]} : sel_132584;
  assign add_132688 = array_index_132366[11:1] + 11'h347;
  assign sel_132690 = $signed({1'h0, add_132586, array_index_132264[0]}) < $signed({1'h0, sel_132588}) ? {add_132586, array_index_132264[0]} : sel_132588;
  assign add_132692 = array_index_132465[11:3] + 9'h0bd;
  assign sel_132695 = $signed({1'h0, add_132590, array_index_132363[2:0]}) < $signed({1'h0, sel_132593}) ? {add_132590, array_index_132363[2:0]} : sel_132593;
  assign add_132697 = array_index_132468[11:3] + 9'h0bd;
  assign sel_132700 = $signed({1'h0, add_132595, array_index_132366[2:0]}) < $signed({1'h0, sel_132598}) ? {add_132595, array_index_132366[2:0]} : sel_132598;
  assign add_132702 = array_index_132567[11:1] + 11'h247;
  assign sel_132705 = $signed({1'h0, add_132600, array_index_132465[0]}) < $signed({1'h0, sel_132603}) ? {add_132600, array_index_132465[0]} : sel_132603;
  assign add_132707 = array_index_132570[11:1] + 11'h247;
  assign sel_132710 = $signed({1'h0, add_132605, array_index_132468[0]}) < $signed({1'h0, sel_132608}) ? {add_132605, array_index_132468[0]} : sel_132608;
  assign add_132735 = array_index_132669[11:0] + 12'h247;
  assign sel_132737 = $signed({1'h0, add_132633}) < $signed({1'h0, sel_132635}) ? add_132633 : sel_132635;
  assign add_132740 = array_index_132672[11:0] + 12'h247;
  assign sel_132742 = $signed({1'h0, add_132638}) < $signed({1'h0, sel_132640}) ? add_132638 : sel_132640;
  assign array_index_132771 = set1_unflattened[7'h1b];
  assign array_index_132774 = set2_unflattened[7'h1b];
  assign add_132778 = array_index_132363[11:1] + 11'h79d;
  assign sel_132780 = $signed({1'h0, add_132676, array_index_132261[0]}) < $signed({1'h0, sel_132678}) ? {add_132676, array_index_132261[0]} : sel_132678;
  assign add_132782 = array_index_132366[11:1] + 11'h79d;
  assign sel_132784 = $signed({1'h0, add_132680, array_index_132264[0]}) < $signed({1'h0, sel_132682}) ? {add_132680, array_index_132264[0]} : sel_132682;
  assign add_132786 = array_index_132465[11:1] + 11'h347;
  assign sel_132788 = $signed({1'h0, add_132684, array_index_132363[0]}) < $signed({1'h0, sel_132686}) ? {add_132684, array_index_132363[0]} : sel_132686;
  assign add_132790 = array_index_132468[11:1] + 11'h347;
  assign sel_132792 = $signed({1'h0, add_132688, array_index_132366[0]}) < $signed({1'h0, sel_132690}) ? {add_132688, array_index_132366[0]} : sel_132690;
  assign add_132794 = array_index_132567[11:3] + 9'h0bd;
  assign sel_132797 = $signed({1'h0, add_132692, array_index_132465[2:0]}) < $signed({1'h0, sel_132695}) ? {add_132692, array_index_132465[2:0]} : sel_132695;
  assign add_132799 = array_index_132570[11:3] + 9'h0bd;
  assign sel_132802 = $signed({1'h0, add_132697, array_index_132468[2:0]}) < $signed({1'h0, sel_132700}) ? {add_132697, array_index_132468[2:0]} : sel_132700;
  assign add_132804 = array_index_132669[11:1] + 11'h247;
  assign sel_132807 = $signed({1'h0, add_132702, array_index_132567[0]}) < $signed({1'h0, sel_132705}) ? {add_132702, array_index_132567[0]} : sel_132705;
  assign add_132809 = array_index_132672[11:1] + 11'h247;
  assign sel_132812 = $signed({1'h0, add_132707, array_index_132570[0]}) < $signed({1'h0, sel_132710}) ? {add_132707, array_index_132570[0]} : sel_132710;
  assign add_132837 = array_index_132771[11:0] + 12'h247;
  assign sel_132839 = $signed({1'h0, add_132735}) < $signed({1'h0, sel_132737}) ? add_132735 : sel_132737;
  assign add_132842 = array_index_132774[11:0] + 12'h247;
  assign sel_132844 = $signed({1'h0, add_132740}) < $signed({1'h0, sel_132742}) ? add_132740 : sel_132742;
  assign array_index_132873 = set1_unflattened[7'h1c];
  assign array_index_132876 = set2_unflattened[7'h1c];
  assign add_132880 = array_index_132465[11:1] + 11'h79d;
  assign sel_132882 = $signed({1'h0, add_132778, array_index_132363[0]}) < $signed({1'h0, sel_132780}) ? {add_132778, array_index_132363[0]} : sel_132780;
  assign add_132884 = array_index_132468[11:1] + 11'h79d;
  assign sel_132886 = $signed({1'h0, add_132782, array_index_132366[0]}) < $signed({1'h0, sel_132784}) ? {add_132782, array_index_132366[0]} : sel_132784;
  assign add_132888 = array_index_132567[11:1] + 11'h347;
  assign sel_132890 = $signed({1'h0, add_132786, array_index_132465[0]}) < $signed({1'h0, sel_132788}) ? {add_132786, array_index_132465[0]} : sel_132788;
  assign add_132892 = array_index_132570[11:1] + 11'h347;
  assign sel_132894 = $signed({1'h0, add_132790, array_index_132468[0]}) < $signed({1'h0, sel_132792}) ? {add_132790, array_index_132468[0]} : sel_132792;
  assign add_132896 = array_index_132669[11:3] + 9'h0bd;
  assign sel_132899 = $signed({1'h0, add_132794, array_index_132567[2:0]}) < $signed({1'h0, sel_132797}) ? {add_132794, array_index_132567[2:0]} : sel_132797;
  assign add_132901 = array_index_132672[11:3] + 9'h0bd;
  assign sel_132904 = $signed({1'h0, add_132799, array_index_132570[2:0]}) < $signed({1'h0, sel_132802}) ? {add_132799, array_index_132570[2:0]} : sel_132802;
  assign add_132906 = array_index_132771[11:1] + 11'h247;
  assign sel_132909 = $signed({1'h0, add_132804, array_index_132669[0]}) < $signed({1'h0, sel_132807}) ? {add_132804, array_index_132669[0]} : sel_132807;
  assign add_132911 = array_index_132774[11:1] + 11'h247;
  assign sel_132914 = $signed({1'h0, add_132809, array_index_132672[0]}) < $signed({1'h0, sel_132812}) ? {add_132809, array_index_132672[0]} : sel_132812;
  assign add_132939 = array_index_132873[11:0] + 12'h247;
  assign sel_132941 = $signed({1'h0, add_132837}) < $signed({1'h0, sel_132839}) ? add_132837 : sel_132839;
  assign add_132944 = array_index_132876[11:0] + 12'h247;
  assign sel_132946 = $signed({1'h0, add_132842}) < $signed({1'h0, sel_132844}) ? add_132842 : sel_132844;
  assign array_index_132975 = set1_unflattened[7'h1d];
  assign array_index_132978 = set2_unflattened[7'h1d];
  assign add_132982 = array_index_132567[11:1] + 11'h79d;
  assign sel_132984 = $signed({1'h0, add_132880, array_index_132465[0]}) < $signed({1'h0, sel_132882}) ? {add_132880, array_index_132465[0]} : sel_132882;
  assign add_132986 = array_index_132570[11:1] + 11'h79d;
  assign sel_132988 = $signed({1'h0, add_132884, array_index_132468[0]}) < $signed({1'h0, sel_132886}) ? {add_132884, array_index_132468[0]} : sel_132886;
  assign add_132990 = array_index_132669[11:1] + 11'h347;
  assign sel_132992 = $signed({1'h0, add_132888, array_index_132567[0]}) < $signed({1'h0, sel_132890}) ? {add_132888, array_index_132567[0]} : sel_132890;
  assign add_132994 = array_index_132672[11:1] + 11'h347;
  assign sel_132996 = $signed({1'h0, add_132892, array_index_132570[0]}) < $signed({1'h0, sel_132894}) ? {add_132892, array_index_132570[0]} : sel_132894;
  assign add_132998 = array_index_132771[11:3] + 9'h0bd;
  assign sel_133001 = $signed({1'h0, add_132896, array_index_132669[2:0]}) < $signed({1'h0, sel_132899}) ? {add_132896, array_index_132669[2:0]} : sel_132899;
  assign add_133003 = array_index_132774[11:3] + 9'h0bd;
  assign sel_133006 = $signed({1'h0, add_132901, array_index_132672[2:0]}) < $signed({1'h0, sel_132904}) ? {add_132901, array_index_132672[2:0]} : sel_132904;
  assign add_133008 = array_index_132873[11:1] + 11'h247;
  assign sel_133011 = $signed({1'h0, add_132906, array_index_132771[0]}) < $signed({1'h0, sel_132909}) ? {add_132906, array_index_132771[0]} : sel_132909;
  assign add_133013 = array_index_132876[11:1] + 11'h247;
  assign sel_133016 = $signed({1'h0, add_132911, array_index_132774[0]}) < $signed({1'h0, sel_132914}) ? {add_132911, array_index_132774[0]} : sel_132914;
  assign add_133041 = array_index_132975[11:0] + 12'h247;
  assign sel_133043 = $signed({1'h0, add_132939}) < $signed({1'h0, sel_132941}) ? add_132939 : sel_132941;
  assign add_133046 = array_index_132978[11:0] + 12'h247;
  assign sel_133048 = $signed({1'h0, add_132944}) < $signed({1'h0, sel_132946}) ? add_132944 : sel_132946;
  assign array_index_133077 = set1_unflattened[7'h1e];
  assign array_index_133080 = set2_unflattened[7'h1e];
  assign add_133084 = array_index_132669[11:1] + 11'h79d;
  assign sel_133086 = $signed({1'h0, add_132982, array_index_132567[0]}) < $signed({1'h0, sel_132984}) ? {add_132982, array_index_132567[0]} : sel_132984;
  assign add_133088 = array_index_132672[11:1] + 11'h79d;
  assign sel_133090 = $signed({1'h0, add_132986, array_index_132570[0]}) < $signed({1'h0, sel_132988}) ? {add_132986, array_index_132570[0]} : sel_132988;
  assign add_133092 = array_index_132771[11:1] + 11'h347;
  assign sel_133094 = $signed({1'h0, add_132990, array_index_132669[0]}) < $signed({1'h0, sel_132992}) ? {add_132990, array_index_132669[0]} : sel_132992;
  assign add_133096 = array_index_132774[11:1] + 11'h347;
  assign sel_133098 = $signed({1'h0, add_132994, array_index_132672[0]}) < $signed({1'h0, sel_132996}) ? {add_132994, array_index_132672[0]} : sel_132996;
  assign add_133100 = array_index_132873[11:3] + 9'h0bd;
  assign sel_133103 = $signed({1'h0, add_132998, array_index_132771[2:0]}) < $signed({1'h0, sel_133001}) ? {add_132998, array_index_132771[2:0]} : sel_133001;
  assign add_133105 = array_index_132876[11:3] + 9'h0bd;
  assign sel_133108 = $signed({1'h0, add_133003, array_index_132774[2:0]}) < $signed({1'h0, sel_133006}) ? {add_133003, array_index_132774[2:0]} : sel_133006;
  assign add_133110 = array_index_132975[11:1] + 11'h247;
  assign sel_133113 = $signed({1'h0, add_133008, array_index_132873[0]}) < $signed({1'h0, sel_133011}) ? {add_133008, array_index_132873[0]} : sel_133011;
  assign add_133115 = array_index_132978[11:1] + 11'h247;
  assign sel_133118 = $signed({1'h0, add_133013, array_index_132876[0]}) < $signed({1'h0, sel_133016}) ? {add_133013, array_index_132876[0]} : sel_133016;
  assign add_133143 = array_index_133077[11:0] + 12'h247;
  assign sel_133145 = $signed({1'h0, add_133041}) < $signed({1'h0, sel_133043}) ? add_133041 : sel_133043;
  assign add_133148 = array_index_133080[11:0] + 12'h247;
  assign sel_133150 = $signed({1'h0, add_133046}) < $signed({1'h0, sel_133048}) ? add_133046 : sel_133048;
  assign array_index_133179 = set1_unflattened[7'h1f];
  assign array_index_133182 = set2_unflattened[7'h1f];
  assign add_133186 = array_index_132771[11:1] + 11'h79d;
  assign sel_133188 = $signed({1'h0, add_133084, array_index_132669[0]}) < $signed({1'h0, sel_133086}) ? {add_133084, array_index_132669[0]} : sel_133086;
  assign add_133190 = array_index_132774[11:1] + 11'h79d;
  assign sel_133192 = $signed({1'h0, add_133088, array_index_132672[0]}) < $signed({1'h0, sel_133090}) ? {add_133088, array_index_132672[0]} : sel_133090;
  assign add_133194 = array_index_132873[11:1] + 11'h347;
  assign sel_133196 = $signed({1'h0, add_133092, array_index_132771[0]}) < $signed({1'h0, sel_133094}) ? {add_133092, array_index_132771[0]} : sel_133094;
  assign add_133198 = array_index_132876[11:1] + 11'h347;
  assign sel_133200 = $signed({1'h0, add_133096, array_index_132774[0]}) < $signed({1'h0, sel_133098}) ? {add_133096, array_index_132774[0]} : sel_133098;
  assign add_133202 = array_index_132975[11:3] + 9'h0bd;
  assign sel_133205 = $signed({1'h0, add_133100, array_index_132873[2:0]}) < $signed({1'h0, sel_133103}) ? {add_133100, array_index_132873[2:0]} : sel_133103;
  assign add_133207 = array_index_132978[11:3] + 9'h0bd;
  assign sel_133210 = $signed({1'h0, add_133105, array_index_132876[2:0]}) < $signed({1'h0, sel_133108}) ? {add_133105, array_index_132876[2:0]} : sel_133108;
  assign add_133212 = array_index_133077[11:1] + 11'h247;
  assign sel_133215 = $signed({1'h0, add_133110, array_index_132975[0]}) < $signed({1'h0, sel_133113}) ? {add_133110, array_index_132975[0]} : sel_133113;
  assign add_133217 = array_index_133080[11:1] + 11'h247;
  assign sel_133220 = $signed({1'h0, add_133115, array_index_132978[0]}) < $signed({1'h0, sel_133118}) ? {add_133115, array_index_132978[0]} : sel_133118;
  assign add_133245 = array_index_133179[11:0] + 12'h247;
  assign sel_133247 = $signed({1'h0, add_133143}) < $signed({1'h0, sel_133145}) ? add_133143 : sel_133145;
  assign add_133250 = array_index_133182[11:0] + 12'h247;
  assign sel_133252 = $signed({1'h0, add_133148}) < $signed({1'h0, sel_133150}) ? add_133148 : sel_133150;
  assign array_index_133281 = set1_unflattened[7'h20];
  assign array_index_133284 = set2_unflattened[7'h20];
  assign add_133288 = array_index_132873[11:1] + 11'h79d;
  assign sel_133290 = $signed({1'h0, add_133186, array_index_132771[0]}) < $signed({1'h0, sel_133188}) ? {add_133186, array_index_132771[0]} : sel_133188;
  assign add_133292 = array_index_132876[11:1] + 11'h79d;
  assign sel_133294 = $signed({1'h0, add_133190, array_index_132774[0]}) < $signed({1'h0, sel_133192}) ? {add_133190, array_index_132774[0]} : sel_133192;
  assign add_133296 = array_index_132975[11:1] + 11'h347;
  assign sel_133298 = $signed({1'h0, add_133194, array_index_132873[0]}) < $signed({1'h0, sel_133196}) ? {add_133194, array_index_132873[0]} : sel_133196;
  assign add_133300 = array_index_132978[11:1] + 11'h347;
  assign sel_133302 = $signed({1'h0, add_133198, array_index_132876[0]}) < $signed({1'h0, sel_133200}) ? {add_133198, array_index_132876[0]} : sel_133200;
  assign add_133304 = array_index_133077[11:3] + 9'h0bd;
  assign sel_133307 = $signed({1'h0, add_133202, array_index_132975[2:0]}) < $signed({1'h0, sel_133205}) ? {add_133202, array_index_132975[2:0]} : sel_133205;
  assign add_133309 = array_index_133080[11:3] + 9'h0bd;
  assign sel_133312 = $signed({1'h0, add_133207, array_index_132978[2:0]}) < $signed({1'h0, sel_133210}) ? {add_133207, array_index_132978[2:0]} : sel_133210;
  assign add_133314 = array_index_133179[11:1] + 11'h247;
  assign sel_133317 = $signed({1'h0, add_133212, array_index_133077[0]}) < $signed({1'h0, sel_133215}) ? {add_133212, array_index_133077[0]} : sel_133215;
  assign add_133319 = array_index_133182[11:1] + 11'h247;
  assign sel_133322 = $signed({1'h0, add_133217, array_index_133080[0]}) < $signed({1'h0, sel_133220}) ? {add_133217, array_index_133080[0]} : sel_133220;
  assign add_133347 = array_index_133281[11:0] + 12'h247;
  assign sel_133349 = $signed({1'h0, add_133245}) < $signed({1'h0, sel_133247}) ? add_133245 : sel_133247;
  assign add_133352 = array_index_133284[11:0] + 12'h247;
  assign sel_133354 = $signed({1'h0, add_133250}) < $signed({1'h0, sel_133252}) ? add_133250 : sel_133252;
  assign array_index_133383 = set1_unflattened[7'h21];
  assign array_index_133386 = set2_unflattened[7'h21];
  assign add_133390 = array_index_132975[11:1] + 11'h79d;
  assign sel_133392 = $signed({1'h0, add_133288, array_index_132873[0]}) < $signed({1'h0, sel_133290}) ? {add_133288, array_index_132873[0]} : sel_133290;
  assign add_133394 = array_index_132978[11:1] + 11'h79d;
  assign sel_133396 = $signed({1'h0, add_133292, array_index_132876[0]}) < $signed({1'h0, sel_133294}) ? {add_133292, array_index_132876[0]} : sel_133294;
  assign add_133398 = array_index_133077[11:1] + 11'h347;
  assign sel_133400 = $signed({1'h0, add_133296, array_index_132975[0]}) < $signed({1'h0, sel_133298}) ? {add_133296, array_index_132975[0]} : sel_133298;
  assign add_133402 = array_index_133080[11:1] + 11'h347;
  assign sel_133404 = $signed({1'h0, add_133300, array_index_132978[0]}) < $signed({1'h0, sel_133302}) ? {add_133300, array_index_132978[0]} : sel_133302;
  assign add_133406 = array_index_133179[11:3] + 9'h0bd;
  assign sel_133409 = $signed({1'h0, add_133304, array_index_133077[2:0]}) < $signed({1'h0, sel_133307}) ? {add_133304, array_index_133077[2:0]} : sel_133307;
  assign add_133411 = array_index_133182[11:3] + 9'h0bd;
  assign sel_133414 = $signed({1'h0, add_133309, array_index_133080[2:0]}) < $signed({1'h0, sel_133312}) ? {add_133309, array_index_133080[2:0]} : sel_133312;
  assign add_133416 = array_index_133281[11:1] + 11'h247;
  assign sel_133419 = $signed({1'h0, add_133314, array_index_133179[0]}) < $signed({1'h0, sel_133317}) ? {add_133314, array_index_133179[0]} : sel_133317;
  assign add_133421 = array_index_133284[11:1] + 11'h247;
  assign sel_133424 = $signed({1'h0, add_133319, array_index_133182[0]}) < $signed({1'h0, sel_133322}) ? {add_133319, array_index_133182[0]} : sel_133322;
  assign add_133449 = array_index_133383[11:0] + 12'h247;
  assign sel_133451 = $signed({1'h0, add_133347}) < $signed({1'h0, sel_133349}) ? add_133347 : sel_133349;
  assign add_133454 = array_index_133386[11:0] + 12'h247;
  assign sel_133456 = $signed({1'h0, add_133352}) < $signed({1'h0, sel_133354}) ? add_133352 : sel_133354;
  assign array_index_133485 = set1_unflattened[7'h22];
  assign array_index_133488 = set2_unflattened[7'h22];
  assign add_133492 = array_index_133077[11:1] + 11'h79d;
  assign sel_133494 = $signed({1'h0, add_133390, array_index_132975[0]}) < $signed({1'h0, sel_133392}) ? {add_133390, array_index_132975[0]} : sel_133392;
  assign add_133496 = array_index_133080[11:1] + 11'h79d;
  assign sel_133498 = $signed({1'h0, add_133394, array_index_132978[0]}) < $signed({1'h0, sel_133396}) ? {add_133394, array_index_132978[0]} : sel_133396;
  assign add_133500 = array_index_133179[11:1] + 11'h347;
  assign sel_133502 = $signed({1'h0, add_133398, array_index_133077[0]}) < $signed({1'h0, sel_133400}) ? {add_133398, array_index_133077[0]} : sel_133400;
  assign add_133504 = array_index_133182[11:1] + 11'h347;
  assign sel_133506 = $signed({1'h0, add_133402, array_index_133080[0]}) < $signed({1'h0, sel_133404}) ? {add_133402, array_index_133080[0]} : sel_133404;
  assign add_133508 = array_index_133281[11:3] + 9'h0bd;
  assign sel_133511 = $signed({1'h0, add_133406, array_index_133179[2:0]}) < $signed({1'h0, sel_133409}) ? {add_133406, array_index_133179[2:0]} : sel_133409;
  assign add_133513 = array_index_133284[11:3] + 9'h0bd;
  assign sel_133516 = $signed({1'h0, add_133411, array_index_133182[2:0]}) < $signed({1'h0, sel_133414}) ? {add_133411, array_index_133182[2:0]} : sel_133414;
  assign add_133518 = array_index_133383[11:1] + 11'h247;
  assign sel_133521 = $signed({1'h0, add_133416, array_index_133281[0]}) < $signed({1'h0, sel_133419}) ? {add_133416, array_index_133281[0]} : sel_133419;
  assign add_133523 = array_index_133386[11:1] + 11'h247;
  assign sel_133526 = $signed({1'h0, add_133421, array_index_133284[0]}) < $signed({1'h0, sel_133424}) ? {add_133421, array_index_133284[0]} : sel_133424;
  assign add_133551 = array_index_133485[11:0] + 12'h247;
  assign sel_133553 = $signed({1'h0, add_133449}) < $signed({1'h0, sel_133451}) ? add_133449 : sel_133451;
  assign add_133556 = array_index_133488[11:0] + 12'h247;
  assign sel_133558 = $signed({1'h0, add_133454}) < $signed({1'h0, sel_133456}) ? add_133454 : sel_133456;
  assign array_index_133587 = set1_unflattened[7'h23];
  assign array_index_133590 = set2_unflattened[7'h23];
  assign add_133594 = array_index_133179[11:1] + 11'h79d;
  assign sel_133596 = $signed({1'h0, add_133492, array_index_133077[0]}) < $signed({1'h0, sel_133494}) ? {add_133492, array_index_133077[0]} : sel_133494;
  assign add_133598 = array_index_133182[11:1] + 11'h79d;
  assign sel_133600 = $signed({1'h0, add_133496, array_index_133080[0]}) < $signed({1'h0, sel_133498}) ? {add_133496, array_index_133080[0]} : sel_133498;
  assign add_133602 = array_index_133281[11:1] + 11'h347;
  assign sel_133604 = $signed({1'h0, add_133500, array_index_133179[0]}) < $signed({1'h0, sel_133502}) ? {add_133500, array_index_133179[0]} : sel_133502;
  assign add_133606 = array_index_133284[11:1] + 11'h347;
  assign sel_133608 = $signed({1'h0, add_133504, array_index_133182[0]}) < $signed({1'h0, sel_133506}) ? {add_133504, array_index_133182[0]} : sel_133506;
  assign add_133610 = array_index_133383[11:3] + 9'h0bd;
  assign sel_133613 = $signed({1'h0, add_133508, array_index_133281[2:0]}) < $signed({1'h0, sel_133511}) ? {add_133508, array_index_133281[2:0]} : sel_133511;
  assign add_133615 = array_index_133386[11:3] + 9'h0bd;
  assign sel_133618 = $signed({1'h0, add_133513, array_index_133284[2:0]}) < $signed({1'h0, sel_133516}) ? {add_133513, array_index_133284[2:0]} : sel_133516;
  assign add_133620 = array_index_133485[11:1] + 11'h247;
  assign sel_133623 = $signed({1'h0, add_133518, array_index_133383[0]}) < $signed({1'h0, sel_133521}) ? {add_133518, array_index_133383[0]} : sel_133521;
  assign add_133625 = array_index_133488[11:1] + 11'h247;
  assign sel_133628 = $signed({1'h0, add_133523, array_index_133386[0]}) < $signed({1'h0, sel_133526}) ? {add_133523, array_index_133386[0]} : sel_133526;
  assign add_133653 = array_index_133587[11:0] + 12'h247;
  assign sel_133655 = $signed({1'h0, add_133551}) < $signed({1'h0, sel_133553}) ? add_133551 : sel_133553;
  assign add_133658 = array_index_133590[11:0] + 12'h247;
  assign sel_133660 = $signed({1'h0, add_133556}) < $signed({1'h0, sel_133558}) ? add_133556 : sel_133558;
  assign array_index_133689 = set1_unflattened[7'h24];
  assign array_index_133692 = set2_unflattened[7'h24];
  assign add_133696 = array_index_133281[11:1] + 11'h79d;
  assign sel_133698 = $signed({1'h0, add_133594, array_index_133179[0]}) < $signed({1'h0, sel_133596}) ? {add_133594, array_index_133179[0]} : sel_133596;
  assign add_133700 = array_index_133284[11:1] + 11'h79d;
  assign sel_133702 = $signed({1'h0, add_133598, array_index_133182[0]}) < $signed({1'h0, sel_133600}) ? {add_133598, array_index_133182[0]} : sel_133600;
  assign add_133704 = array_index_133383[11:1] + 11'h347;
  assign sel_133706 = $signed({1'h0, add_133602, array_index_133281[0]}) < $signed({1'h0, sel_133604}) ? {add_133602, array_index_133281[0]} : sel_133604;
  assign add_133708 = array_index_133386[11:1] + 11'h347;
  assign sel_133710 = $signed({1'h0, add_133606, array_index_133284[0]}) < $signed({1'h0, sel_133608}) ? {add_133606, array_index_133284[0]} : sel_133608;
  assign add_133712 = array_index_133485[11:3] + 9'h0bd;
  assign sel_133715 = $signed({1'h0, add_133610, array_index_133383[2:0]}) < $signed({1'h0, sel_133613}) ? {add_133610, array_index_133383[2:0]} : sel_133613;
  assign add_133717 = array_index_133488[11:3] + 9'h0bd;
  assign sel_133720 = $signed({1'h0, add_133615, array_index_133386[2:0]}) < $signed({1'h0, sel_133618}) ? {add_133615, array_index_133386[2:0]} : sel_133618;
  assign add_133722 = array_index_133587[11:1] + 11'h247;
  assign sel_133725 = $signed({1'h0, add_133620, array_index_133485[0]}) < $signed({1'h0, sel_133623}) ? {add_133620, array_index_133485[0]} : sel_133623;
  assign add_133727 = array_index_133590[11:1] + 11'h247;
  assign sel_133730 = $signed({1'h0, add_133625, array_index_133488[0]}) < $signed({1'h0, sel_133628}) ? {add_133625, array_index_133488[0]} : sel_133628;
  assign add_133755 = array_index_133689[11:0] + 12'h247;
  assign sel_133757 = $signed({1'h0, add_133653}) < $signed({1'h0, sel_133655}) ? add_133653 : sel_133655;
  assign add_133760 = array_index_133692[11:0] + 12'h247;
  assign sel_133762 = $signed({1'h0, add_133658}) < $signed({1'h0, sel_133660}) ? add_133658 : sel_133660;
  assign array_index_133791 = set1_unflattened[7'h25];
  assign array_index_133794 = set2_unflattened[7'h25];
  assign add_133798 = array_index_133383[11:1] + 11'h79d;
  assign sel_133800 = $signed({1'h0, add_133696, array_index_133281[0]}) < $signed({1'h0, sel_133698}) ? {add_133696, array_index_133281[0]} : sel_133698;
  assign add_133802 = array_index_133386[11:1] + 11'h79d;
  assign sel_133804 = $signed({1'h0, add_133700, array_index_133284[0]}) < $signed({1'h0, sel_133702}) ? {add_133700, array_index_133284[0]} : sel_133702;
  assign add_133806 = array_index_133485[11:1] + 11'h347;
  assign sel_133808 = $signed({1'h0, add_133704, array_index_133383[0]}) < $signed({1'h0, sel_133706}) ? {add_133704, array_index_133383[0]} : sel_133706;
  assign add_133810 = array_index_133488[11:1] + 11'h347;
  assign sel_133812 = $signed({1'h0, add_133708, array_index_133386[0]}) < $signed({1'h0, sel_133710}) ? {add_133708, array_index_133386[0]} : sel_133710;
  assign add_133814 = array_index_133587[11:3] + 9'h0bd;
  assign sel_133817 = $signed({1'h0, add_133712, array_index_133485[2:0]}) < $signed({1'h0, sel_133715}) ? {add_133712, array_index_133485[2:0]} : sel_133715;
  assign add_133819 = array_index_133590[11:3] + 9'h0bd;
  assign sel_133822 = $signed({1'h0, add_133717, array_index_133488[2:0]}) < $signed({1'h0, sel_133720}) ? {add_133717, array_index_133488[2:0]} : sel_133720;
  assign add_133824 = array_index_133689[11:1] + 11'h247;
  assign sel_133827 = $signed({1'h0, add_133722, array_index_133587[0]}) < $signed({1'h0, sel_133725}) ? {add_133722, array_index_133587[0]} : sel_133725;
  assign add_133829 = array_index_133692[11:1] + 11'h247;
  assign sel_133832 = $signed({1'h0, add_133727, array_index_133590[0]}) < $signed({1'h0, sel_133730}) ? {add_133727, array_index_133590[0]} : sel_133730;
  assign add_133857 = array_index_133791[11:0] + 12'h247;
  assign sel_133859 = $signed({1'h0, add_133755}) < $signed({1'h0, sel_133757}) ? add_133755 : sel_133757;
  assign add_133862 = array_index_133794[11:0] + 12'h247;
  assign sel_133864 = $signed({1'h0, add_133760}) < $signed({1'h0, sel_133762}) ? add_133760 : sel_133762;
  assign array_index_133893 = set1_unflattened[7'h26];
  assign array_index_133896 = set2_unflattened[7'h26];
  assign add_133900 = array_index_133485[11:1] + 11'h79d;
  assign sel_133902 = $signed({1'h0, add_133798, array_index_133383[0]}) < $signed({1'h0, sel_133800}) ? {add_133798, array_index_133383[0]} : sel_133800;
  assign add_133904 = array_index_133488[11:1] + 11'h79d;
  assign sel_133906 = $signed({1'h0, add_133802, array_index_133386[0]}) < $signed({1'h0, sel_133804}) ? {add_133802, array_index_133386[0]} : sel_133804;
  assign add_133908 = array_index_133587[11:1] + 11'h347;
  assign sel_133910 = $signed({1'h0, add_133806, array_index_133485[0]}) < $signed({1'h0, sel_133808}) ? {add_133806, array_index_133485[0]} : sel_133808;
  assign add_133912 = array_index_133590[11:1] + 11'h347;
  assign sel_133914 = $signed({1'h0, add_133810, array_index_133488[0]}) < $signed({1'h0, sel_133812}) ? {add_133810, array_index_133488[0]} : sel_133812;
  assign add_133916 = array_index_133689[11:3] + 9'h0bd;
  assign sel_133919 = $signed({1'h0, add_133814, array_index_133587[2:0]}) < $signed({1'h0, sel_133817}) ? {add_133814, array_index_133587[2:0]} : sel_133817;
  assign add_133921 = array_index_133692[11:3] + 9'h0bd;
  assign sel_133924 = $signed({1'h0, add_133819, array_index_133590[2:0]}) < $signed({1'h0, sel_133822}) ? {add_133819, array_index_133590[2:0]} : sel_133822;
  assign add_133926 = array_index_133791[11:1] + 11'h247;
  assign sel_133929 = $signed({1'h0, add_133824, array_index_133689[0]}) < $signed({1'h0, sel_133827}) ? {add_133824, array_index_133689[0]} : sel_133827;
  assign add_133931 = array_index_133794[11:1] + 11'h247;
  assign sel_133934 = $signed({1'h0, add_133829, array_index_133692[0]}) < $signed({1'h0, sel_133832}) ? {add_133829, array_index_133692[0]} : sel_133832;
  assign add_133959 = array_index_133893[11:0] + 12'h247;
  assign sel_133961 = $signed({1'h0, add_133857}) < $signed({1'h0, sel_133859}) ? add_133857 : sel_133859;
  assign add_133964 = array_index_133896[11:0] + 12'h247;
  assign sel_133966 = $signed({1'h0, add_133862}) < $signed({1'h0, sel_133864}) ? add_133862 : sel_133864;
  assign array_index_133995 = set1_unflattened[7'h27];
  assign array_index_133998 = set2_unflattened[7'h27];
  assign add_134002 = array_index_133587[11:1] + 11'h79d;
  assign sel_134004 = $signed({1'h0, add_133900, array_index_133485[0]}) < $signed({1'h0, sel_133902}) ? {add_133900, array_index_133485[0]} : sel_133902;
  assign add_134006 = array_index_133590[11:1] + 11'h79d;
  assign sel_134008 = $signed({1'h0, add_133904, array_index_133488[0]}) < $signed({1'h0, sel_133906}) ? {add_133904, array_index_133488[0]} : sel_133906;
  assign add_134010 = array_index_133689[11:1] + 11'h347;
  assign sel_134012 = $signed({1'h0, add_133908, array_index_133587[0]}) < $signed({1'h0, sel_133910}) ? {add_133908, array_index_133587[0]} : sel_133910;
  assign add_134014 = array_index_133692[11:1] + 11'h347;
  assign sel_134016 = $signed({1'h0, add_133912, array_index_133590[0]}) < $signed({1'h0, sel_133914}) ? {add_133912, array_index_133590[0]} : sel_133914;
  assign add_134018 = array_index_133791[11:3] + 9'h0bd;
  assign sel_134021 = $signed({1'h0, add_133916, array_index_133689[2:0]}) < $signed({1'h0, sel_133919}) ? {add_133916, array_index_133689[2:0]} : sel_133919;
  assign add_134023 = array_index_133794[11:3] + 9'h0bd;
  assign sel_134026 = $signed({1'h0, add_133921, array_index_133692[2:0]}) < $signed({1'h0, sel_133924}) ? {add_133921, array_index_133692[2:0]} : sel_133924;
  assign add_134028 = array_index_133893[11:1] + 11'h247;
  assign sel_134031 = $signed({1'h0, add_133926, array_index_133791[0]}) < $signed({1'h0, sel_133929}) ? {add_133926, array_index_133791[0]} : sel_133929;
  assign add_134033 = array_index_133896[11:1] + 11'h247;
  assign sel_134036 = $signed({1'h0, add_133931, array_index_133794[0]}) < $signed({1'h0, sel_133934}) ? {add_133931, array_index_133794[0]} : sel_133934;
  assign add_134061 = array_index_133995[11:0] + 12'h247;
  assign sel_134063 = $signed({1'h0, add_133959}) < $signed({1'h0, sel_133961}) ? add_133959 : sel_133961;
  assign add_134066 = array_index_133998[11:0] + 12'h247;
  assign sel_134068 = $signed({1'h0, add_133964}) < $signed({1'h0, sel_133966}) ? add_133964 : sel_133966;
  assign array_index_134097 = set1_unflattened[7'h28];
  assign array_index_134100 = set2_unflattened[7'h28];
  assign add_134104 = array_index_133689[11:1] + 11'h79d;
  assign sel_134106 = $signed({1'h0, add_134002, array_index_133587[0]}) < $signed({1'h0, sel_134004}) ? {add_134002, array_index_133587[0]} : sel_134004;
  assign add_134108 = array_index_133692[11:1] + 11'h79d;
  assign sel_134110 = $signed({1'h0, add_134006, array_index_133590[0]}) < $signed({1'h0, sel_134008}) ? {add_134006, array_index_133590[0]} : sel_134008;
  assign add_134112 = array_index_133791[11:1] + 11'h347;
  assign sel_134114 = $signed({1'h0, add_134010, array_index_133689[0]}) < $signed({1'h0, sel_134012}) ? {add_134010, array_index_133689[0]} : sel_134012;
  assign add_134116 = array_index_133794[11:1] + 11'h347;
  assign sel_134118 = $signed({1'h0, add_134014, array_index_133692[0]}) < $signed({1'h0, sel_134016}) ? {add_134014, array_index_133692[0]} : sel_134016;
  assign add_134120 = array_index_133893[11:3] + 9'h0bd;
  assign sel_134123 = $signed({1'h0, add_134018, array_index_133791[2:0]}) < $signed({1'h0, sel_134021}) ? {add_134018, array_index_133791[2:0]} : sel_134021;
  assign add_134125 = array_index_133896[11:3] + 9'h0bd;
  assign sel_134128 = $signed({1'h0, add_134023, array_index_133794[2:0]}) < $signed({1'h0, sel_134026}) ? {add_134023, array_index_133794[2:0]} : sel_134026;
  assign add_134130 = array_index_133995[11:1] + 11'h247;
  assign sel_134133 = $signed({1'h0, add_134028, array_index_133893[0]}) < $signed({1'h0, sel_134031}) ? {add_134028, array_index_133893[0]} : sel_134031;
  assign add_134135 = array_index_133998[11:1] + 11'h247;
  assign sel_134138 = $signed({1'h0, add_134033, array_index_133896[0]}) < $signed({1'h0, sel_134036}) ? {add_134033, array_index_133896[0]} : sel_134036;
  assign add_134163 = array_index_134097[11:0] + 12'h247;
  assign sel_134165 = $signed({1'h0, add_134061}) < $signed({1'h0, sel_134063}) ? add_134061 : sel_134063;
  assign add_134168 = array_index_134100[11:0] + 12'h247;
  assign sel_134170 = $signed({1'h0, add_134066}) < $signed({1'h0, sel_134068}) ? add_134066 : sel_134068;
  assign array_index_134199 = set1_unflattened[7'h29];
  assign array_index_134202 = set2_unflattened[7'h29];
  assign add_134206 = array_index_133791[11:1] + 11'h79d;
  assign sel_134208 = $signed({1'h0, add_134104, array_index_133689[0]}) < $signed({1'h0, sel_134106}) ? {add_134104, array_index_133689[0]} : sel_134106;
  assign add_134210 = array_index_133794[11:1] + 11'h79d;
  assign sel_134212 = $signed({1'h0, add_134108, array_index_133692[0]}) < $signed({1'h0, sel_134110}) ? {add_134108, array_index_133692[0]} : sel_134110;
  assign add_134214 = array_index_133893[11:1] + 11'h347;
  assign sel_134216 = $signed({1'h0, add_134112, array_index_133791[0]}) < $signed({1'h0, sel_134114}) ? {add_134112, array_index_133791[0]} : sel_134114;
  assign add_134218 = array_index_133896[11:1] + 11'h347;
  assign sel_134220 = $signed({1'h0, add_134116, array_index_133794[0]}) < $signed({1'h0, sel_134118}) ? {add_134116, array_index_133794[0]} : sel_134118;
  assign add_134222 = array_index_133995[11:3] + 9'h0bd;
  assign sel_134225 = $signed({1'h0, add_134120, array_index_133893[2:0]}) < $signed({1'h0, sel_134123}) ? {add_134120, array_index_133893[2:0]} : sel_134123;
  assign add_134227 = array_index_133998[11:3] + 9'h0bd;
  assign sel_134230 = $signed({1'h0, add_134125, array_index_133896[2:0]}) < $signed({1'h0, sel_134128}) ? {add_134125, array_index_133896[2:0]} : sel_134128;
  assign add_134232 = array_index_134097[11:1] + 11'h247;
  assign sel_134235 = $signed({1'h0, add_134130, array_index_133995[0]}) < $signed({1'h0, sel_134133}) ? {add_134130, array_index_133995[0]} : sel_134133;
  assign add_134237 = array_index_134100[11:1] + 11'h247;
  assign sel_134240 = $signed({1'h0, add_134135, array_index_133998[0]}) < $signed({1'h0, sel_134138}) ? {add_134135, array_index_133998[0]} : sel_134138;
  assign add_134265 = array_index_134199[11:0] + 12'h247;
  assign sel_134267 = $signed({1'h0, add_134163}) < $signed({1'h0, sel_134165}) ? add_134163 : sel_134165;
  assign add_134270 = array_index_134202[11:0] + 12'h247;
  assign sel_134272 = $signed({1'h0, add_134168}) < $signed({1'h0, sel_134170}) ? add_134168 : sel_134170;
  assign array_index_134301 = set1_unflattened[7'h2a];
  assign array_index_134304 = set2_unflattened[7'h2a];
  assign add_134308 = array_index_133893[11:1] + 11'h79d;
  assign sel_134310 = $signed({1'h0, add_134206, array_index_133791[0]}) < $signed({1'h0, sel_134208}) ? {add_134206, array_index_133791[0]} : sel_134208;
  assign add_134312 = array_index_133896[11:1] + 11'h79d;
  assign sel_134314 = $signed({1'h0, add_134210, array_index_133794[0]}) < $signed({1'h0, sel_134212}) ? {add_134210, array_index_133794[0]} : sel_134212;
  assign add_134316 = array_index_133995[11:1] + 11'h347;
  assign sel_134318 = $signed({1'h0, add_134214, array_index_133893[0]}) < $signed({1'h0, sel_134216}) ? {add_134214, array_index_133893[0]} : sel_134216;
  assign add_134320 = array_index_133998[11:1] + 11'h347;
  assign sel_134322 = $signed({1'h0, add_134218, array_index_133896[0]}) < $signed({1'h0, sel_134220}) ? {add_134218, array_index_133896[0]} : sel_134220;
  assign add_134324 = array_index_134097[11:3] + 9'h0bd;
  assign sel_134327 = $signed({1'h0, add_134222, array_index_133995[2:0]}) < $signed({1'h0, sel_134225}) ? {add_134222, array_index_133995[2:0]} : sel_134225;
  assign add_134329 = array_index_134100[11:3] + 9'h0bd;
  assign sel_134332 = $signed({1'h0, add_134227, array_index_133998[2:0]}) < $signed({1'h0, sel_134230}) ? {add_134227, array_index_133998[2:0]} : sel_134230;
  assign add_134334 = array_index_134199[11:1] + 11'h247;
  assign sel_134337 = $signed({1'h0, add_134232, array_index_134097[0]}) < $signed({1'h0, sel_134235}) ? {add_134232, array_index_134097[0]} : sel_134235;
  assign add_134339 = array_index_134202[11:1] + 11'h247;
  assign sel_134342 = $signed({1'h0, add_134237, array_index_134100[0]}) < $signed({1'h0, sel_134240}) ? {add_134237, array_index_134100[0]} : sel_134240;
  assign add_134367 = array_index_134301[11:0] + 12'h247;
  assign sel_134369 = $signed({1'h0, add_134265}) < $signed({1'h0, sel_134267}) ? add_134265 : sel_134267;
  assign add_134372 = array_index_134304[11:0] + 12'h247;
  assign sel_134374 = $signed({1'h0, add_134270}) < $signed({1'h0, sel_134272}) ? add_134270 : sel_134272;
  assign array_index_134403 = set1_unflattened[7'h2b];
  assign array_index_134406 = set2_unflattened[7'h2b];
  assign add_134410 = array_index_133995[11:1] + 11'h79d;
  assign sel_134412 = $signed({1'h0, add_134308, array_index_133893[0]}) < $signed({1'h0, sel_134310}) ? {add_134308, array_index_133893[0]} : sel_134310;
  assign add_134414 = array_index_133998[11:1] + 11'h79d;
  assign sel_134416 = $signed({1'h0, add_134312, array_index_133896[0]}) < $signed({1'h0, sel_134314}) ? {add_134312, array_index_133896[0]} : sel_134314;
  assign add_134418 = array_index_134097[11:1] + 11'h347;
  assign sel_134420 = $signed({1'h0, add_134316, array_index_133995[0]}) < $signed({1'h0, sel_134318}) ? {add_134316, array_index_133995[0]} : sel_134318;
  assign add_134422 = array_index_134100[11:1] + 11'h347;
  assign sel_134424 = $signed({1'h0, add_134320, array_index_133998[0]}) < $signed({1'h0, sel_134322}) ? {add_134320, array_index_133998[0]} : sel_134322;
  assign add_134426 = array_index_134199[11:3] + 9'h0bd;
  assign sel_134429 = $signed({1'h0, add_134324, array_index_134097[2:0]}) < $signed({1'h0, sel_134327}) ? {add_134324, array_index_134097[2:0]} : sel_134327;
  assign add_134431 = array_index_134202[11:3] + 9'h0bd;
  assign sel_134434 = $signed({1'h0, add_134329, array_index_134100[2:0]}) < $signed({1'h0, sel_134332}) ? {add_134329, array_index_134100[2:0]} : sel_134332;
  assign add_134436 = array_index_134301[11:1] + 11'h247;
  assign sel_134439 = $signed({1'h0, add_134334, array_index_134199[0]}) < $signed({1'h0, sel_134337}) ? {add_134334, array_index_134199[0]} : sel_134337;
  assign add_134441 = array_index_134304[11:1] + 11'h247;
  assign sel_134444 = $signed({1'h0, add_134339, array_index_134202[0]}) < $signed({1'h0, sel_134342}) ? {add_134339, array_index_134202[0]} : sel_134342;
  assign add_134469 = array_index_134403[11:0] + 12'h247;
  assign sel_134471 = $signed({1'h0, add_134367}) < $signed({1'h0, sel_134369}) ? add_134367 : sel_134369;
  assign add_134474 = array_index_134406[11:0] + 12'h247;
  assign sel_134476 = $signed({1'h0, add_134372}) < $signed({1'h0, sel_134374}) ? add_134372 : sel_134374;
  assign array_index_134505 = set1_unflattened[7'h2c];
  assign array_index_134508 = set2_unflattened[7'h2c];
  assign add_134512 = array_index_134097[11:1] + 11'h79d;
  assign sel_134514 = $signed({1'h0, add_134410, array_index_133995[0]}) < $signed({1'h0, sel_134412}) ? {add_134410, array_index_133995[0]} : sel_134412;
  assign add_134516 = array_index_134100[11:1] + 11'h79d;
  assign sel_134518 = $signed({1'h0, add_134414, array_index_133998[0]}) < $signed({1'h0, sel_134416}) ? {add_134414, array_index_133998[0]} : sel_134416;
  assign add_134520 = array_index_134199[11:1] + 11'h347;
  assign sel_134522 = $signed({1'h0, add_134418, array_index_134097[0]}) < $signed({1'h0, sel_134420}) ? {add_134418, array_index_134097[0]} : sel_134420;
  assign add_134524 = array_index_134202[11:1] + 11'h347;
  assign sel_134526 = $signed({1'h0, add_134422, array_index_134100[0]}) < $signed({1'h0, sel_134424}) ? {add_134422, array_index_134100[0]} : sel_134424;
  assign add_134528 = array_index_134301[11:3] + 9'h0bd;
  assign sel_134531 = $signed({1'h0, add_134426, array_index_134199[2:0]}) < $signed({1'h0, sel_134429}) ? {add_134426, array_index_134199[2:0]} : sel_134429;
  assign add_134533 = array_index_134304[11:3] + 9'h0bd;
  assign sel_134536 = $signed({1'h0, add_134431, array_index_134202[2:0]}) < $signed({1'h0, sel_134434}) ? {add_134431, array_index_134202[2:0]} : sel_134434;
  assign add_134538 = array_index_134403[11:1] + 11'h247;
  assign sel_134541 = $signed({1'h0, add_134436, array_index_134301[0]}) < $signed({1'h0, sel_134439}) ? {add_134436, array_index_134301[0]} : sel_134439;
  assign add_134543 = array_index_134406[11:1] + 11'h247;
  assign sel_134546 = $signed({1'h0, add_134441, array_index_134304[0]}) < $signed({1'h0, sel_134444}) ? {add_134441, array_index_134304[0]} : sel_134444;
  assign add_134571 = array_index_134505[11:0] + 12'h247;
  assign sel_134573 = $signed({1'h0, add_134469}) < $signed({1'h0, sel_134471}) ? add_134469 : sel_134471;
  assign add_134576 = array_index_134508[11:0] + 12'h247;
  assign sel_134578 = $signed({1'h0, add_134474}) < $signed({1'h0, sel_134476}) ? add_134474 : sel_134476;
  assign array_index_134607 = set1_unflattened[7'h2d];
  assign array_index_134610 = set2_unflattened[7'h2d];
  assign add_134614 = array_index_134199[11:1] + 11'h79d;
  assign sel_134616 = $signed({1'h0, add_134512, array_index_134097[0]}) < $signed({1'h0, sel_134514}) ? {add_134512, array_index_134097[0]} : sel_134514;
  assign add_134618 = array_index_134202[11:1] + 11'h79d;
  assign sel_134620 = $signed({1'h0, add_134516, array_index_134100[0]}) < $signed({1'h0, sel_134518}) ? {add_134516, array_index_134100[0]} : sel_134518;
  assign add_134622 = array_index_134301[11:1] + 11'h347;
  assign sel_134624 = $signed({1'h0, add_134520, array_index_134199[0]}) < $signed({1'h0, sel_134522}) ? {add_134520, array_index_134199[0]} : sel_134522;
  assign add_134626 = array_index_134304[11:1] + 11'h347;
  assign sel_134628 = $signed({1'h0, add_134524, array_index_134202[0]}) < $signed({1'h0, sel_134526}) ? {add_134524, array_index_134202[0]} : sel_134526;
  assign add_134630 = array_index_134403[11:3] + 9'h0bd;
  assign sel_134633 = $signed({1'h0, add_134528, array_index_134301[2:0]}) < $signed({1'h0, sel_134531}) ? {add_134528, array_index_134301[2:0]} : sel_134531;
  assign add_134635 = array_index_134406[11:3] + 9'h0bd;
  assign sel_134638 = $signed({1'h0, add_134533, array_index_134304[2:0]}) < $signed({1'h0, sel_134536}) ? {add_134533, array_index_134304[2:0]} : sel_134536;
  assign add_134640 = array_index_134505[11:1] + 11'h247;
  assign sel_134643 = $signed({1'h0, add_134538, array_index_134403[0]}) < $signed({1'h0, sel_134541}) ? {add_134538, array_index_134403[0]} : sel_134541;
  assign add_134645 = array_index_134508[11:1] + 11'h247;
  assign sel_134648 = $signed({1'h0, add_134543, array_index_134406[0]}) < $signed({1'h0, sel_134546}) ? {add_134543, array_index_134406[0]} : sel_134546;
  assign add_134673 = array_index_134607[11:0] + 12'h247;
  assign sel_134675 = $signed({1'h0, add_134571}) < $signed({1'h0, sel_134573}) ? add_134571 : sel_134573;
  assign add_134678 = array_index_134610[11:0] + 12'h247;
  assign sel_134680 = $signed({1'h0, add_134576}) < $signed({1'h0, sel_134578}) ? add_134576 : sel_134578;
  assign array_index_134709 = set1_unflattened[7'h2e];
  assign array_index_134712 = set2_unflattened[7'h2e];
  assign add_134716 = array_index_134301[11:1] + 11'h79d;
  assign sel_134718 = $signed({1'h0, add_134614, array_index_134199[0]}) < $signed({1'h0, sel_134616}) ? {add_134614, array_index_134199[0]} : sel_134616;
  assign add_134720 = array_index_134304[11:1] + 11'h79d;
  assign sel_134722 = $signed({1'h0, add_134618, array_index_134202[0]}) < $signed({1'h0, sel_134620}) ? {add_134618, array_index_134202[0]} : sel_134620;
  assign add_134724 = array_index_134403[11:1] + 11'h347;
  assign sel_134726 = $signed({1'h0, add_134622, array_index_134301[0]}) < $signed({1'h0, sel_134624}) ? {add_134622, array_index_134301[0]} : sel_134624;
  assign add_134728 = array_index_134406[11:1] + 11'h347;
  assign sel_134730 = $signed({1'h0, add_134626, array_index_134304[0]}) < $signed({1'h0, sel_134628}) ? {add_134626, array_index_134304[0]} : sel_134628;
  assign add_134732 = array_index_134505[11:3] + 9'h0bd;
  assign sel_134735 = $signed({1'h0, add_134630, array_index_134403[2:0]}) < $signed({1'h0, sel_134633}) ? {add_134630, array_index_134403[2:0]} : sel_134633;
  assign add_134737 = array_index_134508[11:3] + 9'h0bd;
  assign sel_134740 = $signed({1'h0, add_134635, array_index_134406[2:0]}) < $signed({1'h0, sel_134638}) ? {add_134635, array_index_134406[2:0]} : sel_134638;
  assign add_134742 = array_index_134607[11:1] + 11'h247;
  assign sel_134745 = $signed({1'h0, add_134640, array_index_134505[0]}) < $signed({1'h0, sel_134643}) ? {add_134640, array_index_134505[0]} : sel_134643;
  assign add_134747 = array_index_134610[11:1] + 11'h247;
  assign sel_134750 = $signed({1'h0, add_134645, array_index_134508[0]}) < $signed({1'h0, sel_134648}) ? {add_134645, array_index_134508[0]} : sel_134648;
  assign add_134775 = array_index_134709[11:0] + 12'h247;
  assign sel_134777 = $signed({1'h0, add_134673}) < $signed({1'h0, sel_134675}) ? add_134673 : sel_134675;
  assign add_134780 = array_index_134712[11:0] + 12'h247;
  assign sel_134782 = $signed({1'h0, add_134678}) < $signed({1'h0, sel_134680}) ? add_134678 : sel_134680;
  assign array_index_134811 = set1_unflattened[7'h2f];
  assign array_index_134814 = set2_unflattened[7'h2f];
  assign add_134818 = array_index_134403[11:1] + 11'h79d;
  assign sel_134820 = $signed({1'h0, add_134716, array_index_134301[0]}) < $signed({1'h0, sel_134718}) ? {add_134716, array_index_134301[0]} : sel_134718;
  assign add_134822 = array_index_134406[11:1] + 11'h79d;
  assign sel_134824 = $signed({1'h0, add_134720, array_index_134304[0]}) < $signed({1'h0, sel_134722}) ? {add_134720, array_index_134304[0]} : sel_134722;
  assign add_134826 = array_index_134505[11:1] + 11'h347;
  assign sel_134828 = $signed({1'h0, add_134724, array_index_134403[0]}) < $signed({1'h0, sel_134726}) ? {add_134724, array_index_134403[0]} : sel_134726;
  assign add_134830 = array_index_134508[11:1] + 11'h347;
  assign sel_134832 = $signed({1'h0, add_134728, array_index_134406[0]}) < $signed({1'h0, sel_134730}) ? {add_134728, array_index_134406[0]} : sel_134730;
  assign add_134834 = array_index_134607[11:3] + 9'h0bd;
  assign sel_134837 = $signed({1'h0, add_134732, array_index_134505[2:0]}) < $signed({1'h0, sel_134735}) ? {add_134732, array_index_134505[2:0]} : sel_134735;
  assign add_134839 = array_index_134610[11:3] + 9'h0bd;
  assign sel_134842 = $signed({1'h0, add_134737, array_index_134508[2:0]}) < $signed({1'h0, sel_134740}) ? {add_134737, array_index_134508[2:0]} : sel_134740;
  assign add_134844 = array_index_134709[11:1] + 11'h247;
  assign sel_134847 = $signed({1'h0, add_134742, array_index_134607[0]}) < $signed({1'h0, sel_134745}) ? {add_134742, array_index_134607[0]} : sel_134745;
  assign add_134849 = array_index_134712[11:1] + 11'h247;
  assign sel_134852 = $signed({1'h0, add_134747, array_index_134610[0]}) < $signed({1'h0, sel_134750}) ? {add_134747, array_index_134610[0]} : sel_134750;
  assign add_134877 = array_index_134811[11:0] + 12'h247;
  assign sel_134879 = $signed({1'h0, add_134775}) < $signed({1'h0, sel_134777}) ? add_134775 : sel_134777;
  assign add_134882 = array_index_134814[11:0] + 12'h247;
  assign sel_134884 = $signed({1'h0, add_134780}) < $signed({1'h0, sel_134782}) ? add_134780 : sel_134782;
  assign array_index_134913 = set1_unflattened[7'h30];
  assign array_index_134916 = set2_unflattened[7'h30];
  assign add_134920 = array_index_134505[11:1] + 11'h79d;
  assign sel_134922 = $signed({1'h0, add_134818, array_index_134403[0]}) < $signed({1'h0, sel_134820}) ? {add_134818, array_index_134403[0]} : sel_134820;
  assign add_134924 = array_index_134508[11:1] + 11'h79d;
  assign sel_134926 = $signed({1'h0, add_134822, array_index_134406[0]}) < $signed({1'h0, sel_134824}) ? {add_134822, array_index_134406[0]} : sel_134824;
  assign add_134928 = array_index_134607[11:1] + 11'h347;
  assign sel_134930 = $signed({1'h0, add_134826, array_index_134505[0]}) < $signed({1'h0, sel_134828}) ? {add_134826, array_index_134505[0]} : sel_134828;
  assign add_134932 = array_index_134610[11:1] + 11'h347;
  assign sel_134934 = $signed({1'h0, add_134830, array_index_134508[0]}) < $signed({1'h0, sel_134832}) ? {add_134830, array_index_134508[0]} : sel_134832;
  assign add_134936 = array_index_134709[11:3] + 9'h0bd;
  assign sel_134939 = $signed({1'h0, add_134834, array_index_134607[2:0]}) < $signed({1'h0, sel_134837}) ? {add_134834, array_index_134607[2:0]} : sel_134837;
  assign add_134941 = array_index_134712[11:3] + 9'h0bd;
  assign sel_134944 = $signed({1'h0, add_134839, array_index_134610[2:0]}) < $signed({1'h0, sel_134842}) ? {add_134839, array_index_134610[2:0]} : sel_134842;
  assign add_134946 = array_index_134811[11:1] + 11'h247;
  assign sel_134949 = $signed({1'h0, add_134844, array_index_134709[0]}) < $signed({1'h0, sel_134847}) ? {add_134844, array_index_134709[0]} : sel_134847;
  assign add_134951 = array_index_134814[11:1] + 11'h247;
  assign sel_134954 = $signed({1'h0, add_134849, array_index_134712[0]}) < $signed({1'h0, sel_134852}) ? {add_134849, array_index_134712[0]} : sel_134852;
  assign add_134979 = array_index_134913[11:0] + 12'h247;
  assign sel_134981 = $signed({1'h0, add_134877}) < $signed({1'h0, sel_134879}) ? add_134877 : sel_134879;
  assign add_134984 = array_index_134916[11:0] + 12'h247;
  assign sel_134986 = $signed({1'h0, add_134882}) < $signed({1'h0, sel_134884}) ? add_134882 : sel_134884;
  assign array_index_135015 = set1_unflattened[7'h31];
  assign array_index_135018 = set2_unflattened[7'h31];
  assign add_135022 = array_index_134607[11:1] + 11'h79d;
  assign sel_135024 = $signed({1'h0, add_134920, array_index_134505[0]}) < $signed({1'h0, sel_134922}) ? {add_134920, array_index_134505[0]} : sel_134922;
  assign add_135026 = array_index_134610[11:1] + 11'h79d;
  assign sel_135028 = $signed({1'h0, add_134924, array_index_134508[0]}) < $signed({1'h0, sel_134926}) ? {add_134924, array_index_134508[0]} : sel_134926;
  assign add_135030 = array_index_134709[11:1] + 11'h347;
  assign sel_135032 = $signed({1'h0, add_134928, array_index_134607[0]}) < $signed({1'h0, sel_134930}) ? {add_134928, array_index_134607[0]} : sel_134930;
  assign add_135034 = array_index_134712[11:1] + 11'h347;
  assign sel_135036 = $signed({1'h0, add_134932, array_index_134610[0]}) < $signed({1'h0, sel_134934}) ? {add_134932, array_index_134610[0]} : sel_134934;
  assign add_135038 = array_index_134811[11:3] + 9'h0bd;
  assign sel_135041 = $signed({1'h0, add_134936, array_index_134709[2:0]}) < $signed({1'h0, sel_134939}) ? {add_134936, array_index_134709[2:0]} : sel_134939;
  assign add_135043 = array_index_134814[11:3] + 9'h0bd;
  assign sel_135046 = $signed({1'h0, add_134941, array_index_134712[2:0]}) < $signed({1'h0, sel_134944}) ? {add_134941, array_index_134712[2:0]} : sel_134944;
  assign add_135048 = array_index_134913[11:1] + 11'h247;
  assign sel_135051 = $signed({1'h0, add_134946, array_index_134811[0]}) < $signed({1'h0, sel_134949}) ? {add_134946, array_index_134811[0]} : sel_134949;
  assign add_135053 = array_index_134916[11:1] + 11'h247;
  assign sel_135056 = $signed({1'h0, add_134951, array_index_134814[0]}) < $signed({1'h0, sel_134954}) ? {add_134951, array_index_134814[0]} : sel_134954;
  assign add_135081 = array_index_135015[11:0] + 12'h247;
  assign sel_135083 = $signed({1'h0, add_134979}) < $signed({1'h0, sel_134981}) ? add_134979 : sel_134981;
  assign add_135086 = array_index_135018[11:0] + 12'h247;
  assign sel_135088 = $signed({1'h0, add_134984}) < $signed({1'h0, sel_134986}) ? add_134984 : sel_134986;
  assign array_index_135117 = set1_unflattened[7'h32];
  assign array_index_135120 = set2_unflattened[7'h32];
  assign add_135124 = array_index_134709[11:1] + 11'h79d;
  assign sel_135126 = $signed({1'h0, add_135022, array_index_134607[0]}) < $signed({1'h0, sel_135024}) ? {add_135022, array_index_134607[0]} : sel_135024;
  assign add_135128 = array_index_134712[11:1] + 11'h79d;
  assign sel_135130 = $signed({1'h0, add_135026, array_index_134610[0]}) < $signed({1'h0, sel_135028}) ? {add_135026, array_index_134610[0]} : sel_135028;
  assign add_135132 = array_index_134811[11:1] + 11'h347;
  assign sel_135134 = $signed({1'h0, add_135030, array_index_134709[0]}) < $signed({1'h0, sel_135032}) ? {add_135030, array_index_134709[0]} : sel_135032;
  assign add_135136 = array_index_134814[11:1] + 11'h347;
  assign sel_135138 = $signed({1'h0, add_135034, array_index_134712[0]}) < $signed({1'h0, sel_135036}) ? {add_135034, array_index_134712[0]} : sel_135036;
  assign add_135140 = array_index_134913[11:3] + 9'h0bd;
  assign sel_135143 = $signed({1'h0, add_135038, array_index_134811[2:0]}) < $signed({1'h0, sel_135041}) ? {add_135038, array_index_134811[2:0]} : sel_135041;
  assign add_135145 = array_index_134916[11:3] + 9'h0bd;
  assign sel_135148 = $signed({1'h0, add_135043, array_index_134814[2:0]}) < $signed({1'h0, sel_135046}) ? {add_135043, array_index_134814[2:0]} : sel_135046;
  assign add_135150 = array_index_135015[11:1] + 11'h247;
  assign sel_135153 = $signed({1'h0, add_135048, array_index_134913[0]}) < $signed({1'h0, sel_135051}) ? {add_135048, array_index_134913[0]} : sel_135051;
  assign add_135155 = array_index_135018[11:1] + 11'h247;
  assign sel_135158 = $signed({1'h0, add_135053, array_index_134916[0]}) < $signed({1'h0, sel_135056}) ? {add_135053, array_index_134916[0]} : sel_135056;
  assign add_135183 = array_index_135117[11:0] + 12'h247;
  assign sel_135185 = $signed({1'h0, add_135081}) < $signed({1'h0, sel_135083}) ? add_135081 : sel_135083;
  assign add_135188 = array_index_135120[11:0] + 12'h247;
  assign sel_135190 = $signed({1'h0, add_135086}) < $signed({1'h0, sel_135088}) ? add_135086 : sel_135088;
  assign array_index_135219 = set1_unflattened[7'h33];
  assign array_index_135222 = set2_unflattened[7'h33];
  assign add_135226 = array_index_134811[11:1] + 11'h79d;
  assign sel_135228 = $signed({1'h0, add_135124, array_index_134709[0]}) < $signed({1'h0, sel_135126}) ? {add_135124, array_index_134709[0]} : sel_135126;
  assign add_135230 = array_index_134814[11:1] + 11'h79d;
  assign sel_135232 = $signed({1'h0, add_135128, array_index_134712[0]}) < $signed({1'h0, sel_135130}) ? {add_135128, array_index_134712[0]} : sel_135130;
  assign add_135234 = array_index_134913[11:1] + 11'h347;
  assign sel_135236 = $signed({1'h0, add_135132, array_index_134811[0]}) < $signed({1'h0, sel_135134}) ? {add_135132, array_index_134811[0]} : sel_135134;
  assign add_135238 = array_index_134916[11:1] + 11'h347;
  assign sel_135240 = $signed({1'h0, add_135136, array_index_134814[0]}) < $signed({1'h0, sel_135138}) ? {add_135136, array_index_134814[0]} : sel_135138;
  assign add_135242 = array_index_135015[11:3] + 9'h0bd;
  assign sel_135245 = $signed({1'h0, add_135140, array_index_134913[2:0]}) < $signed({1'h0, sel_135143}) ? {add_135140, array_index_134913[2:0]} : sel_135143;
  assign add_135247 = array_index_135018[11:3] + 9'h0bd;
  assign sel_135250 = $signed({1'h0, add_135145, array_index_134916[2:0]}) < $signed({1'h0, sel_135148}) ? {add_135145, array_index_134916[2:0]} : sel_135148;
  assign add_135252 = array_index_135117[11:1] + 11'h247;
  assign sel_135255 = $signed({1'h0, add_135150, array_index_135015[0]}) < $signed({1'h0, sel_135153}) ? {add_135150, array_index_135015[0]} : sel_135153;
  assign add_135257 = array_index_135120[11:1] + 11'h247;
  assign sel_135260 = $signed({1'h0, add_135155, array_index_135018[0]}) < $signed({1'h0, sel_135158}) ? {add_135155, array_index_135018[0]} : sel_135158;
  assign add_135285 = array_index_135219[11:0] + 12'h247;
  assign sel_135287 = $signed({1'h0, add_135183}) < $signed({1'h0, sel_135185}) ? add_135183 : sel_135185;
  assign add_135290 = array_index_135222[11:0] + 12'h247;
  assign sel_135292 = $signed({1'h0, add_135188}) < $signed({1'h0, sel_135190}) ? add_135188 : sel_135190;
  assign array_index_135321 = set1_unflattened[7'h34];
  assign array_index_135324 = set2_unflattened[7'h34];
  assign add_135328 = array_index_134913[11:1] + 11'h79d;
  assign sel_135330 = $signed({1'h0, add_135226, array_index_134811[0]}) < $signed({1'h0, sel_135228}) ? {add_135226, array_index_134811[0]} : sel_135228;
  assign add_135332 = array_index_134916[11:1] + 11'h79d;
  assign sel_135334 = $signed({1'h0, add_135230, array_index_134814[0]}) < $signed({1'h0, sel_135232}) ? {add_135230, array_index_134814[0]} : sel_135232;
  assign add_135336 = array_index_135015[11:1] + 11'h347;
  assign sel_135338 = $signed({1'h0, add_135234, array_index_134913[0]}) < $signed({1'h0, sel_135236}) ? {add_135234, array_index_134913[0]} : sel_135236;
  assign add_135340 = array_index_135018[11:1] + 11'h347;
  assign sel_135342 = $signed({1'h0, add_135238, array_index_134916[0]}) < $signed({1'h0, sel_135240}) ? {add_135238, array_index_134916[0]} : sel_135240;
  assign add_135344 = array_index_135117[11:3] + 9'h0bd;
  assign sel_135347 = $signed({1'h0, add_135242, array_index_135015[2:0]}) < $signed({1'h0, sel_135245}) ? {add_135242, array_index_135015[2:0]} : sel_135245;
  assign add_135349 = array_index_135120[11:3] + 9'h0bd;
  assign sel_135352 = $signed({1'h0, add_135247, array_index_135018[2:0]}) < $signed({1'h0, sel_135250}) ? {add_135247, array_index_135018[2:0]} : sel_135250;
  assign add_135354 = array_index_135219[11:1] + 11'h247;
  assign sel_135357 = $signed({1'h0, add_135252, array_index_135117[0]}) < $signed({1'h0, sel_135255}) ? {add_135252, array_index_135117[0]} : sel_135255;
  assign add_135359 = array_index_135222[11:1] + 11'h247;
  assign sel_135362 = $signed({1'h0, add_135257, array_index_135120[0]}) < $signed({1'h0, sel_135260}) ? {add_135257, array_index_135120[0]} : sel_135260;
  assign add_135387 = array_index_135321[11:0] + 12'h247;
  assign sel_135389 = $signed({1'h0, add_135285}) < $signed({1'h0, sel_135287}) ? add_135285 : sel_135287;
  assign add_135392 = array_index_135324[11:0] + 12'h247;
  assign sel_135394 = $signed({1'h0, add_135290}) < $signed({1'h0, sel_135292}) ? add_135290 : sel_135292;
  assign array_index_135423 = set1_unflattened[7'h35];
  assign array_index_135426 = set2_unflattened[7'h35];
  assign add_135430 = array_index_135015[11:1] + 11'h79d;
  assign sel_135432 = $signed({1'h0, add_135328, array_index_134913[0]}) < $signed({1'h0, sel_135330}) ? {add_135328, array_index_134913[0]} : sel_135330;
  assign add_135434 = array_index_135018[11:1] + 11'h79d;
  assign sel_135436 = $signed({1'h0, add_135332, array_index_134916[0]}) < $signed({1'h0, sel_135334}) ? {add_135332, array_index_134916[0]} : sel_135334;
  assign add_135438 = array_index_135117[11:1] + 11'h347;
  assign sel_135440 = $signed({1'h0, add_135336, array_index_135015[0]}) < $signed({1'h0, sel_135338}) ? {add_135336, array_index_135015[0]} : sel_135338;
  assign add_135442 = array_index_135120[11:1] + 11'h347;
  assign sel_135444 = $signed({1'h0, add_135340, array_index_135018[0]}) < $signed({1'h0, sel_135342}) ? {add_135340, array_index_135018[0]} : sel_135342;
  assign add_135446 = array_index_135219[11:3] + 9'h0bd;
  assign sel_135449 = $signed({1'h0, add_135344, array_index_135117[2:0]}) < $signed({1'h0, sel_135347}) ? {add_135344, array_index_135117[2:0]} : sel_135347;
  assign add_135451 = array_index_135222[11:3] + 9'h0bd;
  assign sel_135454 = $signed({1'h0, add_135349, array_index_135120[2:0]}) < $signed({1'h0, sel_135352}) ? {add_135349, array_index_135120[2:0]} : sel_135352;
  assign add_135456 = array_index_135321[11:1] + 11'h247;
  assign sel_135459 = $signed({1'h0, add_135354, array_index_135219[0]}) < $signed({1'h0, sel_135357}) ? {add_135354, array_index_135219[0]} : sel_135357;
  assign add_135461 = array_index_135324[11:1] + 11'h247;
  assign sel_135464 = $signed({1'h0, add_135359, array_index_135222[0]}) < $signed({1'h0, sel_135362}) ? {add_135359, array_index_135222[0]} : sel_135362;
  assign add_135489 = array_index_135423[11:0] + 12'h247;
  assign sel_135491 = $signed({1'h0, add_135387}) < $signed({1'h0, sel_135389}) ? add_135387 : sel_135389;
  assign add_135494 = array_index_135426[11:0] + 12'h247;
  assign sel_135496 = $signed({1'h0, add_135392}) < $signed({1'h0, sel_135394}) ? add_135392 : sel_135394;
  assign array_index_135525 = set1_unflattened[7'h36];
  assign array_index_135528 = set2_unflattened[7'h36];
  assign add_135532 = array_index_135117[11:1] + 11'h79d;
  assign sel_135534 = $signed({1'h0, add_135430, array_index_135015[0]}) < $signed({1'h0, sel_135432}) ? {add_135430, array_index_135015[0]} : sel_135432;
  assign add_135536 = array_index_135120[11:1] + 11'h79d;
  assign sel_135538 = $signed({1'h0, add_135434, array_index_135018[0]}) < $signed({1'h0, sel_135436}) ? {add_135434, array_index_135018[0]} : sel_135436;
  assign add_135540 = array_index_135219[11:1] + 11'h347;
  assign sel_135542 = $signed({1'h0, add_135438, array_index_135117[0]}) < $signed({1'h0, sel_135440}) ? {add_135438, array_index_135117[0]} : sel_135440;
  assign add_135544 = array_index_135222[11:1] + 11'h347;
  assign sel_135546 = $signed({1'h0, add_135442, array_index_135120[0]}) < $signed({1'h0, sel_135444}) ? {add_135442, array_index_135120[0]} : sel_135444;
  assign add_135548 = array_index_135321[11:3] + 9'h0bd;
  assign sel_135551 = $signed({1'h0, add_135446, array_index_135219[2:0]}) < $signed({1'h0, sel_135449}) ? {add_135446, array_index_135219[2:0]} : sel_135449;
  assign add_135553 = array_index_135324[11:3] + 9'h0bd;
  assign sel_135556 = $signed({1'h0, add_135451, array_index_135222[2:0]}) < $signed({1'h0, sel_135454}) ? {add_135451, array_index_135222[2:0]} : sel_135454;
  assign add_135558 = array_index_135423[11:1] + 11'h247;
  assign sel_135561 = $signed({1'h0, add_135456, array_index_135321[0]}) < $signed({1'h0, sel_135459}) ? {add_135456, array_index_135321[0]} : sel_135459;
  assign add_135563 = array_index_135426[11:1] + 11'h247;
  assign sel_135566 = $signed({1'h0, add_135461, array_index_135324[0]}) < $signed({1'h0, sel_135464}) ? {add_135461, array_index_135324[0]} : sel_135464;
  assign add_135591 = array_index_135525[11:0] + 12'h247;
  assign sel_135593 = $signed({1'h0, add_135489}) < $signed({1'h0, sel_135491}) ? add_135489 : sel_135491;
  assign add_135596 = array_index_135528[11:0] + 12'h247;
  assign sel_135598 = $signed({1'h0, add_135494}) < $signed({1'h0, sel_135496}) ? add_135494 : sel_135496;
  assign array_index_135627 = set1_unflattened[7'h37];
  assign array_index_135630 = set2_unflattened[7'h37];
  assign add_135634 = array_index_135219[11:1] + 11'h79d;
  assign sel_135636 = $signed({1'h0, add_135532, array_index_135117[0]}) < $signed({1'h0, sel_135534}) ? {add_135532, array_index_135117[0]} : sel_135534;
  assign add_135638 = array_index_135222[11:1] + 11'h79d;
  assign sel_135640 = $signed({1'h0, add_135536, array_index_135120[0]}) < $signed({1'h0, sel_135538}) ? {add_135536, array_index_135120[0]} : sel_135538;
  assign add_135642 = array_index_135321[11:1] + 11'h347;
  assign sel_135644 = $signed({1'h0, add_135540, array_index_135219[0]}) < $signed({1'h0, sel_135542}) ? {add_135540, array_index_135219[0]} : sel_135542;
  assign add_135646 = array_index_135324[11:1] + 11'h347;
  assign sel_135648 = $signed({1'h0, add_135544, array_index_135222[0]}) < $signed({1'h0, sel_135546}) ? {add_135544, array_index_135222[0]} : sel_135546;
  assign add_135650 = array_index_135423[11:3] + 9'h0bd;
  assign sel_135653 = $signed({1'h0, add_135548, array_index_135321[2:0]}) < $signed({1'h0, sel_135551}) ? {add_135548, array_index_135321[2:0]} : sel_135551;
  assign add_135655 = array_index_135426[11:3] + 9'h0bd;
  assign sel_135658 = $signed({1'h0, add_135553, array_index_135324[2:0]}) < $signed({1'h0, sel_135556}) ? {add_135553, array_index_135324[2:0]} : sel_135556;
  assign add_135660 = array_index_135525[11:1] + 11'h247;
  assign sel_135663 = $signed({1'h0, add_135558, array_index_135423[0]}) < $signed({1'h0, sel_135561}) ? {add_135558, array_index_135423[0]} : sel_135561;
  assign add_135665 = array_index_135528[11:1] + 11'h247;
  assign sel_135668 = $signed({1'h0, add_135563, array_index_135426[0]}) < $signed({1'h0, sel_135566}) ? {add_135563, array_index_135426[0]} : sel_135566;
  assign add_135693 = array_index_135627[11:0] + 12'h247;
  assign sel_135695 = $signed({1'h0, add_135591}) < $signed({1'h0, sel_135593}) ? add_135591 : sel_135593;
  assign add_135698 = array_index_135630[11:0] + 12'h247;
  assign sel_135700 = $signed({1'h0, add_135596}) < $signed({1'h0, sel_135598}) ? add_135596 : sel_135598;
  assign array_index_135729 = set1_unflattened[7'h38];
  assign array_index_135732 = set2_unflattened[7'h38];
  assign add_135736 = array_index_135321[11:1] + 11'h79d;
  assign sel_135738 = $signed({1'h0, add_135634, array_index_135219[0]}) < $signed({1'h0, sel_135636}) ? {add_135634, array_index_135219[0]} : sel_135636;
  assign add_135740 = array_index_135324[11:1] + 11'h79d;
  assign sel_135742 = $signed({1'h0, add_135638, array_index_135222[0]}) < $signed({1'h0, sel_135640}) ? {add_135638, array_index_135222[0]} : sel_135640;
  assign add_135744 = array_index_135423[11:1] + 11'h347;
  assign sel_135746 = $signed({1'h0, add_135642, array_index_135321[0]}) < $signed({1'h0, sel_135644}) ? {add_135642, array_index_135321[0]} : sel_135644;
  assign add_135748 = array_index_135426[11:1] + 11'h347;
  assign sel_135750 = $signed({1'h0, add_135646, array_index_135324[0]}) < $signed({1'h0, sel_135648}) ? {add_135646, array_index_135324[0]} : sel_135648;
  assign add_135752 = array_index_135525[11:3] + 9'h0bd;
  assign sel_135755 = $signed({1'h0, add_135650, array_index_135423[2:0]}) < $signed({1'h0, sel_135653}) ? {add_135650, array_index_135423[2:0]} : sel_135653;
  assign add_135757 = array_index_135528[11:3] + 9'h0bd;
  assign sel_135760 = $signed({1'h0, add_135655, array_index_135426[2:0]}) < $signed({1'h0, sel_135658}) ? {add_135655, array_index_135426[2:0]} : sel_135658;
  assign add_135762 = array_index_135627[11:1] + 11'h247;
  assign sel_135765 = $signed({1'h0, add_135660, array_index_135525[0]}) < $signed({1'h0, sel_135663}) ? {add_135660, array_index_135525[0]} : sel_135663;
  assign add_135767 = array_index_135630[11:1] + 11'h247;
  assign sel_135770 = $signed({1'h0, add_135665, array_index_135528[0]}) < $signed({1'h0, sel_135668}) ? {add_135665, array_index_135528[0]} : sel_135668;
  assign add_135795 = array_index_135729[11:0] + 12'h247;
  assign sel_135797 = $signed({1'h0, add_135693}) < $signed({1'h0, sel_135695}) ? add_135693 : sel_135695;
  assign add_135800 = array_index_135732[11:0] + 12'h247;
  assign sel_135802 = $signed({1'h0, add_135698}) < $signed({1'h0, sel_135700}) ? add_135698 : sel_135700;
  assign array_index_135831 = set1_unflattened[7'h39];
  assign array_index_135834 = set2_unflattened[7'h39];
  assign add_135838 = array_index_135423[11:1] + 11'h79d;
  assign sel_135840 = $signed({1'h0, add_135736, array_index_135321[0]}) < $signed({1'h0, sel_135738}) ? {add_135736, array_index_135321[0]} : sel_135738;
  assign add_135842 = array_index_135426[11:1] + 11'h79d;
  assign sel_135844 = $signed({1'h0, add_135740, array_index_135324[0]}) < $signed({1'h0, sel_135742}) ? {add_135740, array_index_135324[0]} : sel_135742;
  assign add_135846 = array_index_135525[11:1] + 11'h347;
  assign sel_135848 = $signed({1'h0, add_135744, array_index_135423[0]}) < $signed({1'h0, sel_135746}) ? {add_135744, array_index_135423[0]} : sel_135746;
  assign add_135850 = array_index_135528[11:1] + 11'h347;
  assign sel_135852 = $signed({1'h0, add_135748, array_index_135426[0]}) < $signed({1'h0, sel_135750}) ? {add_135748, array_index_135426[0]} : sel_135750;
  assign add_135854 = array_index_135627[11:3] + 9'h0bd;
  assign sel_135857 = $signed({1'h0, add_135752, array_index_135525[2:0]}) < $signed({1'h0, sel_135755}) ? {add_135752, array_index_135525[2:0]} : sel_135755;
  assign add_135859 = array_index_135630[11:3] + 9'h0bd;
  assign sel_135862 = $signed({1'h0, add_135757, array_index_135528[2:0]}) < $signed({1'h0, sel_135760}) ? {add_135757, array_index_135528[2:0]} : sel_135760;
  assign add_135864 = array_index_135729[11:1] + 11'h247;
  assign sel_135867 = $signed({1'h0, add_135762, array_index_135627[0]}) < $signed({1'h0, sel_135765}) ? {add_135762, array_index_135627[0]} : sel_135765;
  assign add_135869 = array_index_135732[11:1] + 11'h247;
  assign sel_135872 = $signed({1'h0, add_135767, array_index_135630[0]}) < $signed({1'h0, sel_135770}) ? {add_135767, array_index_135630[0]} : sel_135770;
  assign add_135897 = array_index_135831[11:0] + 12'h247;
  assign sel_135899 = $signed({1'h0, add_135795}) < $signed({1'h0, sel_135797}) ? add_135795 : sel_135797;
  assign add_135902 = array_index_135834[11:0] + 12'h247;
  assign sel_135904 = $signed({1'h0, add_135800}) < $signed({1'h0, sel_135802}) ? add_135800 : sel_135802;
  assign array_index_135933 = set1_unflattened[7'h3a];
  assign array_index_135936 = set2_unflattened[7'h3a];
  assign add_135940 = array_index_135525[11:1] + 11'h79d;
  assign sel_135942 = $signed({1'h0, add_135838, array_index_135423[0]}) < $signed({1'h0, sel_135840}) ? {add_135838, array_index_135423[0]} : sel_135840;
  assign add_135944 = array_index_135528[11:1] + 11'h79d;
  assign sel_135946 = $signed({1'h0, add_135842, array_index_135426[0]}) < $signed({1'h0, sel_135844}) ? {add_135842, array_index_135426[0]} : sel_135844;
  assign add_135948 = array_index_135627[11:1] + 11'h347;
  assign sel_135950 = $signed({1'h0, add_135846, array_index_135525[0]}) < $signed({1'h0, sel_135848}) ? {add_135846, array_index_135525[0]} : sel_135848;
  assign add_135952 = array_index_135630[11:1] + 11'h347;
  assign sel_135954 = $signed({1'h0, add_135850, array_index_135528[0]}) < $signed({1'h0, sel_135852}) ? {add_135850, array_index_135528[0]} : sel_135852;
  assign add_135956 = array_index_135729[11:3] + 9'h0bd;
  assign sel_135959 = $signed({1'h0, add_135854, array_index_135627[2:0]}) < $signed({1'h0, sel_135857}) ? {add_135854, array_index_135627[2:0]} : sel_135857;
  assign add_135961 = array_index_135732[11:3] + 9'h0bd;
  assign sel_135964 = $signed({1'h0, add_135859, array_index_135630[2:0]}) < $signed({1'h0, sel_135862}) ? {add_135859, array_index_135630[2:0]} : sel_135862;
  assign add_135966 = array_index_135831[11:1] + 11'h247;
  assign sel_135969 = $signed({1'h0, add_135864, array_index_135729[0]}) < $signed({1'h0, sel_135867}) ? {add_135864, array_index_135729[0]} : sel_135867;
  assign add_135971 = array_index_135834[11:1] + 11'h247;
  assign sel_135974 = $signed({1'h0, add_135869, array_index_135732[0]}) < $signed({1'h0, sel_135872}) ? {add_135869, array_index_135732[0]} : sel_135872;
  assign add_135999 = array_index_135933[11:0] + 12'h247;
  assign sel_136001 = $signed({1'h0, add_135897}) < $signed({1'h0, sel_135899}) ? add_135897 : sel_135899;
  assign add_136004 = array_index_135936[11:0] + 12'h247;
  assign sel_136006 = $signed({1'h0, add_135902}) < $signed({1'h0, sel_135904}) ? add_135902 : sel_135904;
  assign array_index_136035 = set1_unflattened[7'h3b];
  assign array_index_136038 = set2_unflattened[7'h3b];
  assign add_136042 = array_index_135627[11:1] + 11'h79d;
  assign sel_136044 = $signed({1'h0, add_135940, array_index_135525[0]}) < $signed({1'h0, sel_135942}) ? {add_135940, array_index_135525[0]} : sel_135942;
  assign add_136046 = array_index_135630[11:1] + 11'h79d;
  assign sel_136048 = $signed({1'h0, add_135944, array_index_135528[0]}) < $signed({1'h0, sel_135946}) ? {add_135944, array_index_135528[0]} : sel_135946;
  assign add_136050 = array_index_135729[11:1] + 11'h347;
  assign sel_136052 = $signed({1'h0, add_135948, array_index_135627[0]}) < $signed({1'h0, sel_135950}) ? {add_135948, array_index_135627[0]} : sel_135950;
  assign add_136054 = array_index_135732[11:1] + 11'h347;
  assign sel_136056 = $signed({1'h0, add_135952, array_index_135630[0]}) < $signed({1'h0, sel_135954}) ? {add_135952, array_index_135630[0]} : sel_135954;
  assign add_136058 = array_index_135831[11:3] + 9'h0bd;
  assign sel_136061 = $signed({1'h0, add_135956, array_index_135729[2:0]}) < $signed({1'h0, sel_135959}) ? {add_135956, array_index_135729[2:0]} : sel_135959;
  assign add_136063 = array_index_135834[11:3] + 9'h0bd;
  assign sel_136066 = $signed({1'h0, add_135961, array_index_135732[2:0]}) < $signed({1'h0, sel_135964}) ? {add_135961, array_index_135732[2:0]} : sel_135964;
  assign add_136068 = array_index_135933[11:1] + 11'h247;
  assign sel_136071 = $signed({1'h0, add_135966, array_index_135831[0]}) < $signed({1'h0, sel_135969}) ? {add_135966, array_index_135831[0]} : sel_135969;
  assign add_136073 = array_index_135936[11:1] + 11'h247;
  assign sel_136076 = $signed({1'h0, add_135971, array_index_135834[0]}) < $signed({1'h0, sel_135974}) ? {add_135971, array_index_135834[0]} : sel_135974;
  assign add_136101 = array_index_136035[11:0] + 12'h247;
  assign sel_136103 = $signed({1'h0, add_135999}) < $signed({1'h0, sel_136001}) ? add_135999 : sel_136001;
  assign add_136106 = array_index_136038[11:0] + 12'h247;
  assign sel_136108 = $signed({1'h0, add_136004}) < $signed({1'h0, sel_136006}) ? add_136004 : sel_136006;
  assign array_index_136137 = set1_unflattened[7'h3c];
  assign array_index_136140 = set2_unflattened[7'h3c];
  assign add_136144 = array_index_135729[11:1] + 11'h79d;
  assign sel_136146 = $signed({1'h0, add_136042, array_index_135627[0]}) < $signed({1'h0, sel_136044}) ? {add_136042, array_index_135627[0]} : sel_136044;
  assign add_136148 = array_index_135732[11:1] + 11'h79d;
  assign sel_136150 = $signed({1'h0, add_136046, array_index_135630[0]}) < $signed({1'h0, sel_136048}) ? {add_136046, array_index_135630[0]} : sel_136048;
  assign add_136152 = array_index_135831[11:1] + 11'h347;
  assign sel_136154 = $signed({1'h0, add_136050, array_index_135729[0]}) < $signed({1'h0, sel_136052}) ? {add_136050, array_index_135729[0]} : sel_136052;
  assign add_136156 = array_index_135834[11:1] + 11'h347;
  assign sel_136158 = $signed({1'h0, add_136054, array_index_135732[0]}) < $signed({1'h0, sel_136056}) ? {add_136054, array_index_135732[0]} : sel_136056;
  assign add_136160 = array_index_135933[11:3] + 9'h0bd;
  assign sel_136163 = $signed({1'h0, add_136058, array_index_135831[2:0]}) < $signed({1'h0, sel_136061}) ? {add_136058, array_index_135831[2:0]} : sel_136061;
  assign add_136165 = array_index_135936[11:3] + 9'h0bd;
  assign sel_136168 = $signed({1'h0, add_136063, array_index_135834[2:0]}) < $signed({1'h0, sel_136066}) ? {add_136063, array_index_135834[2:0]} : sel_136066;
  assign add_136170 = array_index_136035[11:1] + 11'h247;
  assign sel_136173 = $signed({1'h0, add_136068, array_index_135933[0]}) < $signed({1'h0, sel_136071}) ? {add_136068, array_index_135933[0]} : sel_136071;
  assign add_136175 = array_index_136038[11:1] + 11'h247;
  assign sel_136178 = $signed({1'h0, add_136073, array_index_135936[0]}) < $signed({1'h0, sel_136076}) ? {add_136073, array_index_135936[0]} : sel_136076;
  assign add_136203 = array_index_136137[11:0] + 12'h247;
  assign sel_136205 = $signed({1'h0, add_136101}) < $signed({1'h0, sel_136103}) ? add_136101 : sel_136103;
  assign add_136208 = array_index_136140[11:0] + 12'h247;
  assign sel_136210 = $signed({1'h0, add_136106}) < $signed({1'h0, sel_136108}) ? add_136106 : sel_136108;
  assign array_index_136239 = set1_unflattened[7'h3d];
  assign array_index_136242 = set2_unflattened[7'h3d];
  assign add_136246 = array_index_135831[11:1] + 11'h79d;
  assign sel_136248 = $signed({1'h0, add_136144, array_index_135729[0]}) < $signed({1'h0, sel_136146}) ? {add_136144, array_index_135729[0]} : sel_136146;
  assign add_136250 = array_index_135834[11:1] + 11'h79d;
  assign sel_136252 = $signed({1'h0, add_136148, array_index_135732[0]}) < $signed({1'h0, sel_136150}) ? {add_136148, array_index_135732[0]} : sel_136150;
  assign add_136254 = array_index_135933[11:1] + 11'h347;
  assign sel_136256 = $signed({1'h0, add_136152, array_index_135831[0]}) < $signed({1'h0, sel_136154}) ? {add_136152, array_index_135831[0]} : sel_136154;
  assign add_136258 = array_index_135936[11:1] + 11'h347;
  assign sel_136260 = $signed({1'h0, add_136156, array_index_135834[0]}) < $signed({1'h0, sel_136158}) ? {add_136156, array_index_135834[0]} : sel_136158;
  assign add_136262 = array_index_136035[11:3] + 9'h0bd;
  assign sel_136265 = $signed({1'h0, add_136160, array_index_135933[2:0]}) < $signed({1'h0, sel_136163}) ? {add_136160, array_index_135933[2:0]} : sel_136163;
  assign add_136267 = array_index_136038[11:3] + 9'h0bd;
  assign sel_136270 = $signed({1'h0, add_136165, array_index_135936[2:0]}) < $signed({1'h0, sel_136168}) ? {add_136165, array_index_135936[2:0]} : sel_136168;
  assign add_136272 = array_index_136137[11:1] + 11'h247;
  assign sel_136275 = $signed({1'h0, add_136170, array_index_136035[0]}) < $signed({1'h0, sel_136173}) ? {add_136170, array_index_136035[0]} : sel_136173;
  assign add_136277 = array_index_136140[11:1] + 11'h247;
  assign sel_136280 = $signed({1'h0, add_136175, array_index_136038[0]}) < $signed({1'h0, sel_136178}) ? {add_136175, array_index_136038[0]} : sel_136178;
  assign add_136305 = array_index_136239[11:0] + 12'h247;
  assign sel_136307 = $signed({1'h0, add_136203}) < $signed({1'h0, sel_136205}) ? add_136203 : sel_136205;
  assign add_136310 = array_index_136242[11:0] + 12'h247;
  assign sel_136312 = $signed({1'h0, add_136208}) < $signed({1'h0, sel_136210}) ? add_136208 : sel_136210;
  assign array_index_136341 = set1_unflattened[7'h3e];
  assign array_index_136344 = set2_unflattened[7'h3e];
  assign add_136348 = array_index_135933[11:1] + 11'h79d;
  assign sel_136350 = $signed({1'h0, add_136246, array_index_135831[0]}) < $signed({1'h0, sel_136248}) ? {add_136246, array_index_135831[0]} : sel_136248;
  assign add_136352 = array_index_135936[11:1] + 11'h79d;
  assign sel_136354 = $signed({1'h0, add_136250, array_index_135834[0]}) < $signed({1'h0, sel_136252}) ? {add_136250, array_index_135834[0]} : sel_136252;
  assign add_136356 = array_index_136035[11:1] + 11'h347;
  assign sel_136358 = $signed({1'h0, add_136254, array_index_135933[0]}) < $signed({1'h0, sel_136256}) ? {add_136254, array_index_135933[0]} : sel_136256;
  assign add_136360 = array_index_136038[11:1] + 11'h347;
  assign sel_136362 = $signed({1'h0, add_136258, array_index_135936[0]}) < $signed({1'h0, sel_136260}) ? {add_136258, array_index_135936[0]} : sel_136260;
  assign add_136364 = array_index_136137[11:3] + 9'h0bd;
  assign sel_136367 = $signed({1'h0, add_136262, array_index_136035[2:0]}) < $signed({1'h0, sel_136265}) ? {add_136262, array_index_136035[2:0]} : sel_136265;
  assign add_136369 = array_index_136140[11:3] + 9'h0bd;
  assign sel_136372 = $signed({1'h0, add_136267, array_index_136038[2:0]}) < $signed({1'h0, sel_136270}) ? {add_136267, array_index_136038[2:0]} : sel_136270;
  assign add_136374 = array_index_136239[11:1] + 11'h247;
  assign sel_136377 = $signed({1'h0, add_136272, array_index_136137[0]}) < $signed({1'h0, sel_136275}) ? {add_136272, array_index_136137[0]} : sel_136275;
  assign add_136379 = array_index_136242[11:1] + 11'h247;
  assign sel_136382 = $signed({1'h0, add_136277, array_index_136140[0]}) < $signed({1'h0, sel_136280}) ? {add_136277, array_index_136140[0]} : sel_136280;
  assign add_136407 = array_index_136341[11:0] + 12'h247;
  assign sel_136409 = $signed({1'h0, add_136305}) < $signed({1'h0, sel_136307}) ? add_136305 : sel_136307;
  assign add_136412 = array_index_136344[11:0] + 12'h247;
  assign sel_136414 = $signed({1'h0, add_136310}) < $signed({1'h0, sel_136312}) ? add_136310 : sel_136312;
  assign array_index_136443 = set1_unflattened[7'h3f];
  assign array_index_136446 = set2_unflattened[7'h3f];
  assign add_136450 = array_index_136035[11:1] + 11'h79d;
  assign sel_136452 = $signed({1'h0, add_136348, array_index_135933[0]}) < $signed({1'h0, sel_136350}) ? {add_136348, array_index_135933[0]} : sel_136350;
  assign add_136454 = array_index_136038[11:1] + 11'h79d;
  assign sel_136456 = $signed({1'h0, add_136352, array_index_135936[0]}) < $signed({1'h0, sel_136354}) ? {add_136352, array_index_135936[0]} : sel_136354;
  assign add_136458 = array_index_136137[11:1] + 11'h347;
  assign sel_136460 = $signed({1'h0, add_136356, array_index_136035[0]}) < $signed({1'h0, sel_136358}) ? {add_136356, array_index_136035[0]} : sel_136358;
  assign add_136462 = array_index_136140[11:1] + 11'h347;
  assign sel_136464 = $signed({1'h0, add_136360, array_index_136038[0]}) < $signed({1'h0, sel_136362}) ? {add_136360, array_index_136038[0]} : sel_136362;
  assign add_136466 = array_index_136239[11:3] + 9'h0bd;
  assign sel_136469 = $signed({1'h0, add_136364, array_index_136137[2:0]}) < $signed({1'h0, sel_136367}) ? {add_136364, array_index_136137[2:0]} : sel_136367;
  assign add_136471 = array_index_136242[11:3] + 9'h0bd;
  assign sel_136474 = $signed({1'h0, add_136369, array_index_136140[2:0]}) < $signed({1'h0, sel_136372}) ? {add_136369, array_index_136140[2:0]} : sel_136372;
  assign add_136476 = array_index_136341[11:1] + 11'h247;
  assign sel_136479 = $signed({1'h0, add_136374, array_index_136239[0]}) < $signed({1'h0, sel_136377}) ? {add_136374, array_index_136239[0]} : sel_136377;
  assign add_136481 = array_index_136344[11:1] + 11'h247;
  assign sel_136484 = $signed({1'h0, add_136379, array_index_136242[0]}) < $signed({1'h0, sel_136382}) ? {add_136379, array_index_136242[0]} : sel_136382;
  assign add_136509 = array_index_136443[11:0] + 12'h247;
  assign sel_136511 = $signed({1'h0, add_136407}) < $signed({1'h0, sel_136409}) ? add_136407 : sel_136409;
  assign add_136514 = array_index_136446[11:0] + 12'h247;
  assign sel_136516 = $signed({1'h0, add_136412}) < $signed({1'h0, sel_136414}) ? add_136412 : sel_136414;
  assign array_index_136545 = set1_unflattened[7'h40];
  assign array_index_136548 = set2_unflattened[7'h40];
  assign add_136552 = array_index_136137[11:1] + 11'h79d;
  assign sel_136554 = $signed({1'h0, add_136450, array_index_136035[0]}) < $signed({1'h0, sel_136452}) ? {add_136450, array_index_136035[0]} : sel_136452;
  assign add_136556 = array_index_136140[11:1] + 11'h79d;
  assign sel_136558 = $signed({1'h0, add_136454, array_index_136038[0]}) < $signed({1'h0, sel_136456}) ? {add_136454, array_index_136038[0]} : sel_136456;
  assign add_136560 = array_index_136239[11:1] + 11'h347;
  assign sel_136562 = $signed({1'h0, add_136458, array_index_136137[0]}) < $signed({1'h0, sel_136460}) ? {add_136458, array_index_136137[0]} : sel_136460;
  assign add_136564 = array_index_136242[11:1] + 11'h347;
  assign sel_136566 = $signed({1'h0, add_136462, array_index_136140[0]}) < $signed({1'h0, sel_136464}) ? {add_136462, array_index_136140[0]} : sel_136464;
  assign add_136568 = array_index_136341[11:3] + 9'h0bd;
  assign sel_136571 = $signed({1'h0, add_136466, array_index_136239[2:0]}) < $signed({1'h0, sel_136469}) ? {add_136466, array_index_136239[2:0]} : sel_136469;
  assign add_136573 = array_index_136344[11:3] + 9'h0bd;
  assign sel_136576 = $signed({1'h0, add_136471, array_index_136242[2:0]}) < $signed({1'h0, sel_136474}) ? {add_136471, array_index_136242[2:0]} : sel_136474;
  assign add_136578 = array_index_136443[11:1] + 11'h247;
  assign sel_136581 = $signed({1'h0, add_136476, array_index_136341[0]}) < $signed({1'h0, sel_136479}) ? {add_136476, array_index_136341[0]} : sel_136479;
  assign add_136583 = array_index_136446[11:1] + 11'h247;
  assign sel_136586 = $signed({1'h0, add_136481, array_index_136344[0]}) < $signed({1'h0, sel_136484}) ? {add_136481, array_index_136344[0]} : sel_136484;
  assign add_136611 = array_index_136545[11:0] + 12'h247;
  assign sel_136613 = $signed({1'h0, add_136509}) < $signed({1'h0, sel_136511}) ? add_136509 : sel_136511;
  assign add_136616 = array_index_136548[11:0] + 12'h247;
  assign sel_136618 = $signed({1'h0, add_136514}) < $signed({1'h0, sel_136516}) ? add_136514 : sel_136516;
  assign array_index_136647 = set1_unflattened[7'h41];
  assign array_index_136650 = set2_unflattened[7'h41];
  assign add_136654 = array_index_136239[11:1] + 11'h79d;
  assign sel_136656 = $signed({1'h0, add_136552, array_index_136137[0]}) < $signed({1'h0, sel_136554}) ? {add_136552, array_index_136137[0]} : sel_136554;
  assign add_136658 = array_index_136242[11:1] + 11'h79d;
  assign sel_136660 = $signed({1'h0, add_136556, array_index_136140[0]}) < $signed({1'h0, sel_136558}) ? {add_136556, array_index_136140[0]} : sel_136558;
  assign add_136662 = array_index_136341[11:1] + 11'h347;
  assign sel_136664 = $signed({1'h0, add_136560, array_index_136239[0]}) < $signed({1'h0, sel_136562}) ? {add_136560, array_index_136239[0]} : sel_136562;
  assign add_136666 = array_index_136344[11:1] + 11'h347;
  assign sel_136668 = $signed({1'h0, add_136564, array_index_136242[0]}) < $signed({1'h0, sel_136566}) ? {add_136564, array_index_136242[0]} : sel_136566;
  assign add_136670 = array_index_136443[11:3] + 9'h0bd;
  assign sel_136673 = $signed({1'h0, add_136568, array_index_136341[2:0]}) < $signed({1'h0, sel_136571}) ? {add_136568, array_index_136341[2:0]} : sel_136571;
  assign add_136675 = array_index_136446[11:3] + 9'h0bd;
  assign sel_136678 = $signed({1'h0, add_136573, array_index_136344[2:0]}) < $signed({1'h0, sel_136576}) ? {add_136573, array_index_136344[2:0]} : sel_136576;
  assign add_136680 = array_index_136545[11:1] + 11'h247;
  assign sel_136683 = $signed({1'h0, add_136578, array_index_136443[0]}) < $signed({1'h0, sel_136581}) ? {add_136578, array_index_136443[0]} : sel_136581;
  assign add_136685 = array_index_136548[11:1] + 11'h247;
  assign sel_136688 = $signed({1'h0, add_136583, array_index_136446[0]}) < $signed({1'h0, sel_136586}) ? {add_136583, array_index_136446[0]} : sel_136586;
  assign add_136713 = array_index_136647[11:0] + 12'h247;
  assign sel_136715 = $signed({1'h0, add_136611}) < $signed({1'h0, sel_136613}) ? add_136611 : sel_136613;
  assign add_136718 = array_index_136650[11:0] + 12'h247;
  assign sel_136720 = $signed({1'h0, add_136616}) < $signed({1'h0, sel_136618}) ? add_136616 : sel_136618;
  assign array_index_136749 = set1_unflattened[7'h42];
  assign array_index_136752 = set2_unflattened[7'h42];
  assign add_136756 = array_index_136341[11:1] + 11'h79d;
  assign sel_136758 = $signed({1'h0, add_136654, array_index_136239[0]}) < $signed({1'h0, sel_136656}) ? {add_136654, array_index_136239[0]} : sel_136656;
  assign add_136760 = array_index_136344[11:1] + 11'h79d;
  assign sel_136762 = $signed({1'h0, add_136658, array_index_136242[0]}) < $signed({1'h0, sel_136660}) ? {add_136658, array_index_136242[0]} : sel_136660;
  assign add_136764 = array_index_136443[11:1] + 11'h347;
  assign sel_136766 = $signed({1'h0, add_136662, array_index_136341[0]}) < $signed({1'h0, sel_136664}) ? {add_136662, array_index_136341[0]} : sel_136664;
  assign add_136768 = array_index_136446[11:1] + 11'h347;
  assign sel_136770 = $signed({1'h0, add_136666, array_index_136344[0]}) < $signed({1'h0, sel_136668}) ? {add_136666, array_index_136344[0]} : sel_136668;
  assign add_136772 = array_index_136545[11:3] + 9'h0bd;
  assign sel_136775 = $signed({1'h0, add_136670, array_index_136443[2:0]}) < $signed({1'h0, sel_136673}) ? {add_136670, array_index_136443[2:0]} : sel_136673;
  assign add_136777 = array_index_136548[11:3] + 9'h0bd;
  assign sel_136780 = $signed({1'h0, add_136675, array_index_136446[2:0]}) < $signed({1'h0, sel_136678}) ? {add_136675, array_index_136446[2:0]} : sel_136678;
  assign add_136782 = array_index_136647[11:1] + 11'h247;
  assign sel_136785 = $signed({1'h0, add_136680, array_index_136545[0]}) < $signed({1'h0, sel_136683}) ? {add_136680, array_index_136545[0]} : sel_136683;
  assign add_136787 = array_index_136650[11:1] + 11'h247;
  assign sel_136790 = $signed({1'h0, add_136685, array_index_136548[0]}) < $signed({1'h0, sel_136688}) ? {add_136685, array_index_136548[0]} : sel_136688;
  assign add_136815 = array_index_136749[11:0] + 12'h247;
  assign sel_136817 = $signed({1'h0, add_136713}) < $signed({1'h0, sel_136715}) ? add_136713 : sel_136715;
  assign add_136820 = array_index_136752[11:0] + 12'h247;
  assign sel_136822 = $signed({1'h0, add_136718}) < $signed({1'h0, sel_136720}) ? add_136718 : sel_136720;
  assign array_index_136851 = set1_unflattened[7'h43];
  assign array_index_136854 = set2_unflattened[7'h43];
  assign add_136858 = array_index_136443[11:1] + 11'h79d;
  assign sel_136860 = $signed({1'h0, add_136756, array_index_136341[0]}) < $signed({1'h0, sel_136758}) ? {add_136756, array_index_136341[0]} : sel_136758;
  assign add_136862 = array_index_136446[11:1] + 11'h79d;
  assign sel_136864 = $signed({1'h0, add_136760, array_index_136344[0]}) < $signed({1'h0, sel_136762}) ? {add_136760, array_index_136344[0]} : sel_136762;
  assign add_136866 = array_index_136545[11:1] + 11'h347;
  assign sel_136868 = $signed({1'h0, add_136764, array_index_136443[0]}) < $signed({1'h0, sel_136766}) ? {add_136764, array_index_136443[0]} : sel_136766;
  assign add_136870 = array_index_136548[11:1] + 11'h347;
  assign sel_136872 = $signed({1'h0, add_136768, array_index_136446[0]}) < $signed({1'h0, sel_136770}) ? {add_136768, array_index_136446[0]} : sel_136770;
  assign add_136874 = array_index_136647[11:3] + 9'h0bd;
  assign sel_136877 = $signed({1'h0, add_136772, array_index_136545[2:0]}) < $signed({1'h0, sel_136775}) ? {add_136772, array_index_136545[2:0]} : sel_136775;
  assign add_136879 = array_index_136650[11:3] + 9'h0bd;
  assign sel_136882 = $signed({1'h0, add_136777, array_index_136548[2:0]}) < $signed({1'h0, sel_136780}) ? {add_136777, array_index_136548[2:0]} : sel_136780;
  assign add_136884 = array_index_136749[11:1] + 11'h247;
  assign sel_136887 = $signed({1'h0, add_136782, array_index_136647[0]}) < $signed({1'h0, sel_136785}) ? {add_136782, array_index_136647[0]} : sel_136785;
  assign add_136889 = array_index_136752[11:1] + 11'h247;
  assign sel_136892 = $signed({1'h0, add_136787, array_index_136650[0]}) < $signed({1'h0, sel_136790}) ? {add_136787, array_index_136650[0]} : sel_136790;
  assign add_136917 = array_index_136851[11:0] + 12'h247;
  assign sel_136919 = $signed({1'h0, add_136815}) < $signed({1'h0, sel_136817}) ? add_136815 : sel_136817;
  assign add_136922 = array_index_136854[11:0] + 12'h247;
  assign sel_136924 = $signed({1'h0, add_136820}) < $signed({1'h0, sel_136822}) ? add_136820 : sel_136822;
  assign array_index_136953 = set1_unflattened[7'h44];
  assign array_index_136956 = set2_unflattened[7'h44];
  assign add_136960 = array_index_136545[11:1] + 11'h79d;
  assign sel_136962 = $signed({1'h0, add_136858, array_index_136443[0]}) < $signed({1'h0, sel_136860}) ? {add_136858, array_index_136443[0]} : sel_136860;
  assign add_136964 = array_index_136548[11:1] + 11'h79d;
  assign sel_136966 = $signed({1'h0, add_136862, array_index_136446[0]}) < $signed({1'h0, sel_136864}) ? {add_136862, array_index_136446[0]} : sel_136864;
  assign add_136968 = array_index_136647[11:1] + 11'h347;
  assign sel_136970 = $signed({1'h0, add_136866, array_index_136545[0]}) < $signed({1'h0, sel_136868}) ? {add_136866, array_index_136545[0]} : sel_136868;
  assign add_136972 = array_index_136650[11:1] + 11'h347;
  assign sel_136974 = $signed({1'h0, add_136870, array_index_136548[0]}) < $signed({1'h0, sel_136872}) ? {add_136870, array_index_136548[0]} : sel_136872;
  assign add_136976 = array_index_136749[11:3] + 9'h0bd;
  assign sel_136979 = $signed({1'h0, add_136874, array_index_136647[2:0]}) < $signed({1'h0, sel_136877}) ? {add_136874, array_index_136647[2:0]} : sel_136877;
  assign add_136981 = array_index_136752[11:3] + 9'h0bd;
  assign sel_136984 = $signed({1'h0, add_136879, array_index_136650[2:0]}) < $signed({1'h0, sel_136882}) ? {add_136879, array_index_136650[2:0]} : sel_136882;
  assign add_136986 = array_index_136851[11:1] + 11'h247;
  assign sel_136989 = $signed({1'h0, add_136884, array_index_136749[0]}) < $signed({1'h0, sel_136887}) ? {add_136884, array_index_136749[0]} : sel_136887;
  assign add_136991 = array_index_136854[11:1] + 11'h247;
  assign sel_136994 = $signed({1'h0, add_136889, array_index_136752[0]}) < $signed({1'h0, sel_136892}) ? {add_136889, array_index_136752[0]} : sel_136892;
  assign add_137019 = array_index_136953[11:0] + 12'h247;
  assign sel_137021 = $signed({1'h0, add_136917}) < $signed({1'h0, sel_136919}) ? add_136917 : sel_136919;
  assign add_137024 = array_index_136956[11:0] + 12'h247;
  assign sel_137026 = $signed({1'h0, add_136922}) < $signed({1'h0, sel_136924}) ? add_136922 : sel_136924;
  assign array_index_137055 = set1_unflattened[7'h45];
  assign array_index_137058 = set2_unflattened[7'h45];
  assign add_137062 = array_index_136647[11:1] + 11'h79d;
  assign sel_137064 = $signed({1'h0, add_136960, array_index_136545[0]}) < $signed({1'h0, sel_136962}) ? {add_136960, array_index_136545[0]} : sel_136962;
  assign add_137066 = array_index_136650[11:1] + 11'h79d;
  assign sel_137068 = $signed({1'h0, add_136964, array_index_136548[0]}) < $signed({1'h0, sel_136966}) ? {add_136964, array_index_136548[0]} : sel_136966;
  assign add_137070 = array_index_136749[11:1] + 11'h347;
  assign sel_137072 = $signed({1'h0, add_136968, array_index_136647[0]}) < $signed({1'h0, sel_136970}) ? {add_136968, array_index_136647[0]} : sel_136970;
  assign add_137074 = array_index_136752[11:1] + 11'h347;
  assign sel_137076 = $signed({1'h0, add_136972, array_index_136650[0]}) < $signed({1'h0, sel_136974}) ? {add_136972, array_index_136650[0]} : sel_136974;
  assign add_137078 = array_index_136851[11:3] + 9'h0bd;
  assign sel_137081 = $signed({1'h0, add_136976, array_index_136749[2:0]}) < $signed({1'h0, sel_136979}) ? {add_136976, array_index_136749[2:0]} : sel_136979;
  assign add_137083 = array_index_136854[11:3] + 9'h0bd;
  assign sel_137086 = $signed({1'h0, add_136981, array_index_136752[2:0]}) < $signed({1'h0, sel_136984}) ? {add_136981, array_index_136752[2:0]} : sel_136984;
  assign add_137088 = array_index_136953[11:1] + 11'h247;
  assign sel_137091 = $signed({1'h0, add_136986, array_index_136851[0]}) < $signed({1'h0, sel_136989}) ? {add_136986, array_index_136851[0]} : sel_136989;
  assign add_137093 = array_index_136956[11:1] + 11'h247;
  assign sel_137096 = $signed({1'h0, add_136991, array_index_136854[0]}) < $signed({1'h0, sel_136994}) ? {add_136991, array_index_136854[0]} : sel_136994;
  assign add_137121 = array_index_137055[11:0] + 12'h247;
  assign sel_137123 = $signed({1'h0, add_137019}) < $signed({1'h0, sel_137021}) ? add_137019 : sel_137021;
  assign add_137126 = array_index_137058[11:0] + 12'h247;
  assign sel_137128 = $signed({1'h0, add_137024}) < $signed({1'h0, sel_137026}) ? add_137024 : sel_137026;
  assign array_index_137157 = set1_unflattened[7'h46];
  assign array_index_137160 = set2_unflattened[7'h46];
  assign add_137164 = array_index_136749[11:1] + 11'h79d;
  assign sel_137166 = $signed({1'h0, add_137062, array_index_136647[0]}) < $signed({1'h0, sel_137064}) ? {add_137062, array_index_136647[0]} : sel_137064;
  assign add_137168 = array_index_136752[11:1] + 11'h79d;
  assign sel_137170 = $signed({1'h0, add_137066, array_index_136650[0]}) < $signed({1'h0, sel_137068}) ? {add_137066, array_index_136650[0]} : sel_137068;
  assign add_137172 = array_index_136851[11:1] + 11'h347;
  assign sel_137174 = $signed({1'h0, add_137070, array_index_136749[0]}) < $signed({1'h0, sel_137072}) ? {add_137070, array_index_136749[0]} : sel_137072;
  assign add_137176 = array_index_136854[11:1] + 11'h347;
  assign sel_137178 = $signed({1'h0, add_137074, array_index_136752[0]}) < $signed({1'h0, sel_137076}) ? {add_137074, array_index_136752[0]} : sel_137076;
  assign add_137180 = array_index_136953[11:3] + 9'h0bd;
  assign sel_137183 = $signed({1'h0, add_137078, array_index_136851[2:0]}) < $signed({1'h0, sel_137081}) ? {add_137078, array_index_136851[2:0]} : sel_137081;
  assign add_137185 = array_index_136956[11:3] + 9'h0bd;
  assign sel_137188 = $signed({1'h0, add_137083, array_index_136854[2:0]}) < $signed({1'h0, sel_137086}) ? {add_137083, array_index_136854[2:0]} : sel_137086;
  assign add_137190 = array_index_137055[11:1] + 11'h247;
  assign sel_137193 = $signed({1'h0, add_137088, array_index_136953[0]}) < $signed({1'h0, sel_137091}) ? {add_137088, array_index_136953[0]} : sel_137091;
  assign add_137195 = array_index_137058[11:1] + 11'h247;
  assign sel_137198 = $signed({1'h0, add_137093, array_index_136956[0]}) < $signed({1'h0, sel_137096}) ? {add_137093, array_index_136956[0]} : sel_137096;
  assign add_137223 = array_index_137157[11:0] + 12'h247;
  assign sel_137225 = $signed({1'h0, add_137121}) < $signed({1'h0, sel_137123}) ? add_137121 : sel_137123;
  assign add_137228 = array_index_137160[11:0] + 12'h247;
  assign sel_137230 = $signed({1'h0, add_137126}) < $signed({1'h0, sel_137128}) ? add_137126 : sel_137128;
  assign array_index_137259 = set1_unflattened[7'h47];
  assign array_index_137262 = set2_unflattened[7'h47];
  assign add_137266 = array_index_136851[11:1] + 11'h79d;
  assign sel_137268 = $signed({1'h0, add_137164, array_index_136749[0]}) < $signed({1'h0, sel_137166}) ? {add_137164, array_index_136749[0]} : sel_137166;
  assign add_137270 = array_index_136854[11:1] + 11'h79d;
  assign sel_137272 = $signed({1'h0, add_137168, array_index_136752[0]}) < $signed({1'h0, sel_137170}) ? {add_137168, array_index_136752[0]} : sel_137170;
  assign add_137274 = array_index_136953[11:1] + 11'h347;
  assign sel_137276 = $signed({1'h0, add_137172, array_index_136851[0]}) < $signed({1'h0, sel_137174}) ? {add_137172, array_index_136851[0]} : sel_137174;
  assign add_137278 = array_index_136956[11:1] + 11'h347;
  assign sel_137280 = $signed({1'h0, add_137176, array_index_136854[0]}) < $signed({1'h0, sel_137178}) ? {add_137176, array_index_136854[0]} : sel_137178;
  assign add_137282 = array_index_137055[11:3] + 9'h0bd;
  assign sel_137285 = $signed({1'h0, add_137180, array_index_136953[2:0]}) < $signed({1'h0, sel_137183}) ? {add_137180, array_index_136953[2:0]} : sel_137183;
  assign add_137287 = array_index_137058[11:3] + 9'h0bd;
  assign sel_137290 = $signed({1'h0, add_137185, array_index_136956[2:0]}) < $signed({1'h0, sel_137188}) ? {add_137185, array_index_136956[2:0]} : sel_137188;
  assign add_137292 = array_index_137157[11:1] + 11'h247;
  assign sel_137295 = $signed({1'h0, add_137190, array_index_137055[0]}) < $signed({1'h0, sel_137193}) ? {add_137190, array_index_137055[0]} : sel_137193;
  assign add_137297 = array_index_137160[11:1] + 11'h247;
  assign sel_137300 = $signed({1'h0, add_137195, array_index_137058[0]}) < $signed({1'h0, sel_137198}) ? {add_137195, array_index_137058[0]} : sel_137198;
  assign add_137325 = array_index_137259[11:0] + 12'h247;
  assign sel_137327 = $signed({1'h0, add_137223}) < $signed({1'h0, sel_137225}) ? add_137223 : sel_137225;
  assign add_137330 = array_index_137262[11:0] + 12'h247;
  assign sel_137332 = $signed({1'h0, add_137228}) < $signed({1'h0, sel_137230}) ? add_137228 : sel_137230;
  assign array_index_137361 = set1_unflattened[7'h48];
  assign array_index_137364 = set2_unflattened[7'h48];
  assign add_137368 = array_index_136953[11:1] + 11'h79d;
  assign sel_137370 = $signed({1'h0, add_137266, array_index_136851[0]}) < $signed({1'h0, sel_137268}) ? {add_137266, array_index_136851[0]} : sel_137268;
  assign add_137372 = array_index_136956[11:1] + 11'h79d;
  assign sel_137374 = $signed({1'h0, add_137270, array_index_136854[0]}) < $signed({1'h0, sel_137272}) ? {add_137270, array_index_136854[0]} : sel_137272;
  assign add_137376 = array_index_137055[11:1] + 11'h347;
  assign sel_137378 = $signed({1'h0, add_137274, array_index_136953[0]}) < $signed({1'h0, sel_137276}) ? {add_137274, array_index_136953[0]} : sel_137276;
  assign add_137380 = array_index_137058[11:1] + 11'h347;
  assign sel_137382 = $signed({1'h0, add_137278, array_index_136956[0]}) < $signed({1'h0, sel_137280}) ? {add_137278, array_index_136956[0]} : sel_137280;
  assign add_137384 = array_index_137157[11:3] + 9'h0bd;
  assign sel_137387 = $signed({1'h0, add_137282, array_index_137055[2:0]}) < $signed({1'h0, sel_137285}) ? {add_137282, array_index_137055[2:0]} : sel_137285;
  assign add_137389 = array_index_137160[11:3] + 9'h0bd;
  assign sel_137392 = $signed({1'h0, add_137287, array_index_137058[2:0]}) < $signed({1'h0, sel_137290}) ? {add_137287, array_index_137058[2:0]} : sel_137290;
  assign add_137394 = array_index_137259[11:1] + 11'h247;
  assign sel_137397 = $signed({1'h0, add_137292, array_index_137157[0]}) < $signed({1'h0, sel_137295}) ? {add_137292, array_index_137157[0]} : sel_137295;
  assign add_137399 = array_index_137262[11:1] + 11'h247;
  assign sel_137402 = $signed({1'h0, add_137297, array_index_137160[0]}) < $signed({1'h0, sel_137300}) ? {add_137297, array_index_137160[0]} : sel_137300;
  assign add_137427 = array_index_137361[11:0] + 12'h247;
  assign sel_137429 = $signed({1'h0, add_137325}) < $signed({1'h0, sel_137327}) ? add_137325 : sel_137327;
  assign add_137432 = array_index_137364[11:0] + 12'h247;
  assign sel_137434 = $signed({1'h0, add_137330}) < $signed({1'h0, sel_137332}) ? add_137330 : sel_137332;
  assign array_index_137463 = set1_unflattened[7'h49];
  assign array_index_137466 = set2_unflattened[7'h49];
  assign add_137470 = array_index_137055[11:1] + 11'h79d;
  assign sel_137472 = $signed({1'h0, add_137368, array_index_136953[0]}) < $signed({1'h0, sel_137370}) ? {add_137368, array_index_136953[0]} : sel_137370;
  assign add_137474 = array_index_137058[11:1] + 11'h79d;
  assign sel_137476 = $signed({1'h0, add_137372, array_index_136956[0]}) < $signed({1'h0, sel_137374}) ? {add_137372, array_index_136956[0]} : sel_137374;
  assign add_137478 = array_index_137157[11:1] + 11'h347;
  assign sel_137480 = $signed({1'h0, add_137376, array_index_137055[0]}) < $signed({1'h0, sel_137378}) ? {add_137376, array_index_137055[0]} : sel_137378;
  assign add_137482 = array_index_137160[11:1] + 11'h347;
  assign sel_137484 = $signed({1'h0, add_137380, array_index_137058[0]}) < $signed({1'h0, sel_137382}) ? {add_137380, array_index_137058[0]} : sel_137382;
  assign add_137486 = array_index_137259[11:3] + 9'h0bd;
  assign sel_137489 = $signed({1'h0, add_137384, array_index_137157[2:0]}) < $signed({1'h0, sel_137387}) ? {add_137384, array_index_137157[2:0]} : sel_137387;
  assign add_137491 = array_index_137262[11:3] + 9'h0bd;
  assign sel_137494 = $signed({1'h0, add_137389, array_index_137160[2:0]}) < $signed({1'h0, sel_137392}) ? {add_137389, array_index_137160[2:0]} : sel_137392;
  assign add_137496 = array_index_137361[11:1] + 11'h247;
  assign sel_137499 = $signed({1'h0, add_137394, array_index_137259[0]}) < $signed({1'h0, sel_137397}) ? {add_137394, array_index_137259[0]} : sel_137397;
  assign add_137501 = array_index_137364[11:1] + 11'h247;
  assign sel_137504 = $signed({1'h0, add_137399, array_index_137262[0]}) < $signed({1'h0, sel_137402}) ? {add_137399, array_index_137262[0]} : sel_137402;
  assign add_137529 = array_index_137463[11:0] + 12'h247;
  assign sel_137531 = $signed({1'h0, add_137427}) < $signed({1'h0, sel_137429}) ? add_137427 : sel_137429;
  assign add_137534 = array_index_137466[11:0] + 12'h247;
  assign sel_137536 = $signed({1'h0, add_137432}) < $signed({1'h0, sel_137434}) ? add_137432 : sel_137434;
  assign array_index_137565 = set1_unflattened[7'h4a];
  assign array_index_137568 = set2_unflattened[7'h4a];
  assign add_137572 = array_index_137157[11:1] + 11'h79d;
  assign sel_137574 = $signed({1'h0, add_137470, array_index_137055[0]}) < $signed({1'h0, sel_137472}) ? {add_137470, array_index_137055[0]} : sel_137472;
  assign add_137576 = array_index_137160[11:1] + 11'h79d;
  assign sel_137578 = $signed({1'h0, add_137474, array_index_137058[0]}) < $signed({1'h0, sel_137476}) ? {add_137474, array_index_137058[0]} : sel_137476;
  assign add_137580 = array_index_137259[11:1] + 11'h347;
  assign sel_137582 = $signed({1'h0, add_137478, array_index_137157[0]}) < $signed({1'h0, sel_137480}) ? {add_137478, array_index_137157[0]} : sel_137480;
  assign add_137584 = array_index_137262[11:1] + 11'h347;
  assign sel_137586 = $signed({1'h0, add_137482, array_index_137160[0]}) < $signed({1'h0, sel_137484}) ? {add_137482, array_index_137160[0]} : sel_137484;
  assign add_137588 = array_index_137361[11:3] + 9'h0bd;
  assign sel_137591 = $signed({1'h0, add_137486, array_index_137259[2:0]}) < $signed({1'h0, sel_137489}) ? {add_137486, array_index_137259[2:0]} : sel_137489;
  assign add_137593 = array_index_137364[11:3] + 9'h0bd;
  assign sel_137596 = $signed({1'h0, add_137491, array_index_137262[2:0]}) < $signed({1'h0, sel_137494}) ? {add_137491, array_index_137262[2:0]} : sel_137494;
  assign add_137598 = array_index_137463[11:1] + 11'h247;
  assign sel_137601 = $signed({1'h0, add_137496, array_index_137361[0]}) < $signed({1'h0, sel_137499}) ? {add_137496, array_index_137361[0]} : sel_137499;
  assign add_137603 = array_index_137466[11:1] + 11'h247;
  assign sel_137606 = $signed({1'h0, add_137501, array_index_137364[0]}) < $signed({1'h0, sel_137504}) ? {add_137501, array_index_137364[0]} : sel_137504;
  assign add_137630 = array_index_137565[11:0] + 12'h247;
  assign sel_137632 = $signed({1'h0, add_137529}) < $signed({1'h0, sel_137531}) ? add_137529 : sel_137531;
  assign add_137634 = array_index_137568[11:0] + 12'h247;
  assign sel_137636 = $signed({1'h0, add_137534}) < $signed({1'h0, sel_137536}) ? add_137534 : sel_137536;
  assign add_137670 = array_index_137259[11:1] + 11'h79d;
  assign sel_137672 = $signed({1'h0, add_137572, array_index_137157[0]}) < $signed({1'h0, sel_137574}) ? {add_137572, array_index_137157[0]} : sel_137574;
  assign add_137674 = array_index_137262[11:1] + 11'h79d;
  assign sel_137676 = $signed({1'h0, add_137576, array_index_137160[0]}) < $signed({1'h0, sel_137578}) ? {add_137576, array_index_137160[0]} : sel_137578;
  assign add_137678 = array_index_137361[11:1] + 11'h347;
  assign sel_137680 = $signed({1'h0, add_137580, array_index_137259[0]}) < $signed({1'h0, sel_137582}) ? {add_137580, array_index_137259[0]} : sel_137582;
  assign add_137682 = array_index_137364[11:1] + 11'h347;
  assign sel_137684 = $signed({1'h0, add_137584, array_index_137262[0]}) < $signed({1'h0, sel_137586}) ? {add_137584, array_index_137262[0]} : sel_137586;
  assign add_137686 = array_index_137463[11:3] + 9'h0bd;
  assign sel_137689 = $signed({1'h0, add_137588, array_index_137361[2:0]}) < $signed({1'h0, sel_137591}) ? {add_137588, array_index_137361[2:0]} : sel_137591;
  assign add_137691 = array_index_137466[11:3] + 9'h0bd;
  assign sel_137694 = $signed({1'h0, add_137593, array_index_137364[2:0]}) < $signed({1'h0, sel_137596}) ? {add_137593, array_index_137364[2:0]} : sel_137596;
  assign add_137696 = array_index_137565[11:1] + 11'h247;
  assign sel_137699 = $signed({1'h0, add_137598, array_index_137463[0]}) < $signed({1'h0, sel_137601}) ? {add_137598, array_index_137463[0]} : sel_137601;
  assign add_137701 = array_index_137568[11:1] + 11'h247;
  assign sel_137704 = $signed({1'h0, add_137603, array_index_137466[0]}) < $signed({1'h0, sel_137606}) ? {add_137603, array_index_137466[0]} : sel_137606;
  assign add_137752 = array_index_137361[11:1] + 11'h79d;
  assign sel_137754 = $signed({1'h0, add_137670, array_index_137259[0]}) < $signed({1'h0, sel_137672}) ? {add_137670, array_index_137259[0]} : sel_137672;
  assign add_137756 = array_index_137364[11:1] + 11'h79d;
  assign sel_137758 = $signed({1'h0, add_137674, array_index_137262[0]}) < $signed({1'h0, sel_137676}) ? {add_137674, array_index_137262[0]} : sel_137676;
  assign add_137760 = array_index_137463[11:1] + 11'h347;
  assign sel_137762 = $signed({1'h0, add_137678, array_index_137361[0]}) < $signed({1'h0, sel_137680}) ? {add_137678, array_index_137361[0]} : sel_137680;
  assign add_137764 = array_index_137466[11:1] + 11'h347;
  assign sel_137766 = $signed({1'h0, add_137682, array_index_137364[0]}) < $signed({1'h0, sel_137684}) ? {add_137682, array_index_137364[0]} : sel_137684;
  assign add_137768 = array_index_137565[11:3] + 9'h0bd;
  assign sel_137771 = $signed({1'h0, add_137686, array_index_137463[2:0]}) < $signed({1'h0, sel_137689}) ? {add_137686, array_index_137463[2:0]} : sel_137689;
  assign add_137773 = array_index_137568[11:3] + 9'h0bd;
  assign sel_137776 = $signed({1'h0, add_137691, array_index_137466[2:0]}) < $signed({1'h0, sel_137694}) ? {add_137691, array_index_137466[2:0]} : sel_137694;
  assign concat_137779 = {1'h0, ($signed({1'h0, add_137630}) < $signed({1'h0, sel_137632}) ? add_137630 : sel_137632) == ($signed({1'h0, add_137634}) < $signed({1'h0, sel_137636}) ? add_137634 : sel_137636)};
  assign add_137794 = concat_137779 + 2'h1;
  assign add_137814 = array_index_137463[11:1] + 11'h79d;
  assign sel_137816 = $signed({1'h0, add_137752, array_index_137361[0]}) < $signed({1'h0, sel_137754}) ? {add_137752, array_index_137361[0]} : sel_137754;
  assign add_137818 = array_index_137466[11:1] + 11'h79d;
  assign sel_137820 = $signed({1'h0, add_137756, array_index_137364[0]}) < $signed({1'h0, sel_137758}) ? {add_137756, array_index_137364[0]} : sel_137758;
  assign add_137822 = array_index_137565[11:1] + 11'h347;
  assign sel_137824 = $signed({1'h0, add_137760, array_index_137463[0]}) < $signed({1'h0, sel_137762}) ? {add_137760, array_index_137463[0]} : sel_137762;
  assign add_137826 = array_index_137568[11:1] + 11'h347;
  assign sel_137828 = $signed({1'h0, add_137764, array_index_137466[0]}) < $signed({1'h0, sel_137766}) ? {add_137764, array_index_137466[0]} : sel_137766;
  assign concat_137831 = {1'h0, ($signed({1'h0, add_137696, array_index_137565[0]}) < $signed({1'h0, sel_137699}) ? {add_137696, array_index_137565[0]} : sel_137699) == ($signed({1'h0, add_137701, array_index_137568[0]}) < $signed({1'h0, sel_137704}) ? {add_137701, array_index_137568[0]} : sel_137704) ? add_137794 : concat_137779};
  assign add_137842 = concat_137831 + 3'h1;
  assign add_137856 = array_index_137565[11:1] + 11'h79d;
  assign sel_137858 = $signed({1'h0, add_137814, array_index_137463[0]}) < $signed({1'h0, sel_137816}) ? {add_137814, array_index_137463[0]} : sel_137816;
  assign add_137860 = array_index_137568[11:1] + 11'h79d;
  assign sel_137862 = $signed({1'h0, add_137818, array_index_137466[0]}) < $signed({1'h0, sel_137820}) ? {add_137818, array_index_137466[0]} : sel_137820;
  assign concat_137865 = {1'h0, ($signed({1'h0, add_137768, array_index_137565[2:0]}) < $signed({1'h0, sel_137771}) ? {add_137768, array_index_137565[2:0]} : sel_137771) == ($signed({1'h0, add_137773, array_index_137568[2:0]}) < $signed({1'h0, sel_137776}) ? {add_137773, array_index_137568[2:0]} : sel_137776) ? add_137842 : concat_137831};
  assign add_137872 = concat_137865 + 4'h1;
  assign concat_137881 = {1'h0, ($signed({1'h0, add_137822, array_index_137565[0]}) < $signed({1'h0, sel_137824}) ? {add_137822, array_index_137565[0]} : sel_137824) == ($signed({1'h0, add_137826, array_index_137568[0]}) < $signed({1'h0, sel_137828}) ? {add_137826, array_index_137568[0]} : sel_137828) ? add_137872 : concat_137865};
  assign add_137884 = concat_137881 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_137856, array_index_137565[0]}) < $signed({1'h0, sel_137858}) ? {add_137856, array_index_137565[0]} : sel_137858) == ($signed({1'h0, add_137860, array_index_137568[0]}) < $signed({1'h0, sel_137862}) ? {add_137860, array_index_137568[0]} : sel_137862) ? add_137884 : concat_137881}, {set1_unflattened[74], set1_unflattened[73], set1_unflattened[72], set1_unflattened[71], set1_unflattened[70], set1_unflattened[69], set1_unflattened[68], set1_unflattened[67], set1_unflattened[66], set1_unflattened[65], set1_unflattened[64], set1_unflattened[63], set1_unflattened[62], set1_unflattened[61], set1_unflattened[60], set1_unflattened[59], set1_unflattened[58], set1_unflattened[57], set1_unflattened[56], set1_unflattened[55], set1_unflattened[54], set1_unflattened[53], set1_unflattened[52], set1_unflattened[51], set1_unflattened[50], set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[74], set2_unflattened[73], set2_unflattened[72], set2_unflattened[71], set2_unflattened[70], set2_unflattened[69], set2_unflattened[68], set2_unflattened[67], set2_unflattened[66], set2_unflattened[65], set2_unflattened[64], set2_unflattened[63], set2_unflattened[62], set2_unflattened[61], set2_unflattened[60], set2_unflattened[59], set2_unflattened[58], set2_unflattened[57], set2_unflattened[56], set2_unflattened[55], set2_unflattened[54], set2_unflattened[53], set2_unflattened[52], set2_unflattened[51], set2_unflattened[50], set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
