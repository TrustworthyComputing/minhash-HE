module min_hash(
  input wire [479:0] set1,
  input wire [479:0] set2,
  output wire [975:0] out
);
  wire [15:0] set1_unflattened[30];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  wire [15:0] set2_unflattened[30];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  wire [15:0] array_index_257761;
  wire [15:0] array_index_257762;
  wire [11:0] add_257769;
  wire [11:0] add_257772;
  wire [15:0] array_index_257775;
  wire [15:0] array_index_257778;
  wire [11:0] add_257782;
  wire [11:0] add_257784;
  wire [11:0] add_257799;
  wire [11:0] sel_257801;
  wire [11:0] add_257804;
  wire [11:0] sel_257806;
  wire [15:0] array_index_257817;
  wire [15:0] array_index_257820;
  wire [9:0] add_257824;
  wire [9:0] add_257827;
  wire [11:0] add_257830;
  wire [11:0] sel_257832;
  wire [11:0] add_257834;
  wire [11:0] sel_257836;
  wire [11:0] add_257853;
  wire [11:0] sel_257855;
  wire [11:0] add_257858;
  wire [11:0] sel_257860;
  wire [15:0] array_index_257877;
  wire [15:0] array_index_257880;
  wire [9:0] add_257884;
  wire [9:0] add_257886;
  wire [9:0] add_257888;
  wire [11:0] sel_257891;
  wire [9:0] add_257893;
  wire [11:0] sel_257896;
  wire [11:0] add_257898;
  wire [11:0] sel_257900;
  wire [11:0] add_257902;
  wire [11:0] sel_257904;
  wire [11:0] add_257925;
  wire [11:0] sel_257927;
  wire [11:0] add_257930;
  wire [11:0] sel_257932;
  wire [15:0] array_index_257955;
  wire [15:0] array_index_257958;
  wire [11:0] add_257962;
  wire [11:0] add_257964;
  wire [9:0] add_257966;
  wire [11:0] sel_257968;
  wire [9:0] add_257970;
  wire [11:0] sel_257972;
  wire [9:0] add_257974;
  wire [11:0] sel_257977;
  wire [9:0] add_257979;
  wire [11:0] sel_257982;
  wire [11:0] add_257984;
  wire [11:0] sel_257986;
  wire [11:0] add_257988;
  wire [11:0] sel_257990;
  wire [11:0] add_258015;
  wire [11:0] sel_258017;
  wire [11:0] add_258020;
  wire [11:0] sel_258022;
  wire [15:0] array_index_258049;
  wire [15:0] array_index_258052;
  wire [11:0] add_258056;
  wire [11:0] add_258058;
  wire [11:0] add_258060;
  wire [11:0] sel_258062;
  wire [11:0] add_258064;
  wire [11:0] sel_258066;
  wire [9:0] add_258068;
  wire [11:0] sel_258070;
  wire [9:0] add_258072;
  wire [11:0] sel_258074;
  wire [9:0] add_258076;
  wire [11:0] sel_258079;
  wire [9:0] add_258081;
  wire [11:0] sel_258084;
  wire [11:0] add_258086;
  wire [11:0] sel_258088;
  wire [11:0] add_258090;
  wire [11:0] sel_258092;
  wire [11:0] add_258121;
  wire [11:0] sel_258123;
  wire [11:0] add_258126;
  wire [11:0] sel_258128;
  wire [15:0] array_index_258159;
  wire [15:0] array_index_258162;
  wire [11:0] add_258166;
  wire [11:0] add_258168;
  wire [11:0] add_258170;
  wire [11:0] sel_258172;
  wire [11:0] add_258174;
  wire [11:0] sel_258176;
  wire [11:0] add_258178;
  wire [11:0] sel_258180;
  wire [11:0] add_258182;
  wire [11:0] sel_258184;
  wire [9:0] add_258186;
  wire [11:0] sel_258188;
  wire [9:0] add_258190;
  wire [11:0] sel_258192;
  wire [9:0] add_258194;
  wire [11:0] sel_258197;
  wire [9:0] add_258199;
  wire [11:0] sel_258202;
  wire [11:0] add_258204;
  wire [11:0] sel_258206;
  wire [11:0] add_258208;
  wire [11:0] sel_258210;
  wire [11:0] add_258243;
  wire [11:0] sel_258245;
  wire [11:0] add_258248;
  wire [11:0] sel_258250;
  wire [15:0] array_index_258285;
  wire [15:0] array_index_258288;
  wire [11:0] add_258292;
  wire [11:0] add_258294;
  wire [11:0] add_258296;
  wire [11:0] sel_258298;
  wire [11:0] add_258300;
  wire [11:0] sel_258302;
  wire [11:0] add_258304;
  wire [11:0] sel_258306;
  wire [11:0] add_258308;
  wire [11:0] sel_258310;
  wire [11:0] add_258312;
  wire [11:0] sel_258314;
  wire [11:0] add_258316;
  wire [11:0] sel_258318;
  wire [9:0] add_258320;
  wire [11:0] sel_258322;
  wire [9:0] add_258324;
  wire [11:0] sel_258326;
  wire [9:0] add_258328;
  wire [11:0] sel_258331;
  wire [9:0] add_258333;
  wire [11:0] sel_258336;
  wire [11:0] add_258338;
  wire [11:0] sel_258340;
  wire [11:0] add_258342;
  wire [11:0] sel_258344;
  wire [11:0] add_258381;
  wire [11:0] sel_258383;
  wire [11:0] add_258386;
  wire [11:0] sel_258388;
  wire [15:0] array_index_258427;
  wire [15:0] array_index_258430;
  wire [11:0] add_258434;
  wire [11:0] add_258436;
  wire [11:0] add_258438;
  wire [11:0] sel_258440;
  wire [11:0] add_258442;
  wire [11:0] sel_258444;
  wire [11:0] add_258446;
  wire [11:0] sel_258448;
  wire [11:0] add_258450;
  wire [11:0] sel_258452;
  wire [11:0] add_258454;
  wire [11:0] sel_258456;
  wire [11:0] add_258458;
  wire [11:0] sel_258460;
  wire [11:0] add_258462;
  wire [11:0] sel_258464;
  wire [11:0] add_258466;
  wire [11:0] sel_258468;
  wire [9:0] add_258470;
  wire [11:0] sel_258472;
  wire [9:0] add_258474;
  wire [11:0] sel_258476;
  wire [9:0] add_258478;
  wire [11:0] sel_258481;
  wire [9:0] add_258483;
  wire [11:0] sel_258486;
  wire [11:0] add_258488;
  wire [11:0] sel_258490;
  wire [11:0] add_258492;
  wire [11:0] sel_258494;
  wire [11:0] add_258535;
  wire [11:0] sel_258537;
  wire [11:0] add_258540;
  wire [11:0] sel_258542;
  wire [15:0] array_index_258585;
  wire [15:0] array_index_258588;
  wire [11:0] add_258592;
  wire [11:0] add_258594;
  wire [11:0] add_258596;
  wire [11:0] sel_258598;
  wire [11:0] add_258600;
  wire [11:0] sel_258602;
  wire [11:0] add_258604;
  wire [11:0] sel_258606;
  wire [11:0] add_258608;
  wire [11:0] sel_258610;
  wire [11:0] add_258612;
  wire [11:0] sel_258614;
  wire [11:0] add_258616;
  wire [11:0] sel_258618;
  wire [11:0] add_258620;
  wire [11:0] sel_258622;
  wire [11:0] add_258624;
  wire [11:0] sel_258626;
  wire [11:0] add_258628;
  wire [11:0] sel_258630;
  wire [11:0] add_258632;
  wire [11:0] sel_258634;
  wire [9:0] add_258636;
  wire [11:0] sel_258638;
  wire [9:0] add_258640;
  wire [11:0] sel_258642;
  wire [9:0] add_258644;
  wire [11:0] sel_258647;
  wire [9:0] add_258649;
  wire [11:0] sel_258652;
  wire [11:0] add_258654;
  wire [11:0] sel_258656;
  wire [11:0] add_258658;
  wire [11:0] sel_258660;
  wire [11:0] add_258705;
  wire [11:0] sel_258707;
  wire [11:0] add_258710;
  wire [11:0] sel_258712;
  wire [15:0] array_index_258761;
  wire [15:0] array_index_258764;
  wire [10:0] add_258768;
  wire [10:0] add_258771;
  wire [11:0] add_258774;
  wire [11:0] sel_258776;
  wire [11:0] add_258778;
  wire [11:0] sel_258780;
  wire [11:0] add_258782;
  wire [11:0] sel_258784;
  wire [11:0] add_258786;
  wire [11:0] sel_258788;
  wire [11:0] add_258790;
  wire [11:0] sel_258792;
  wire [11:0] add_258794;
  wire [11:0] sel_258796;
  wire [11:0] add_258798;
  wire [11:0] sel_258800;
  wire [11:0] add_258802;
  wire [11:0] sel_258804;
  wire [11:0] add_258806;
  wire [11:0] sel_258808;
  wire [11:0] add_258810;
  wire [11:0] sel_258812;
  wire [11:0] add_258814;
  wire [11:0] sel_258816;
  wire [11:0] add_258818;
  wire [11:0] sel_258820;
  wire [9:0] add_258822;
  wire [11:0] sel_258824;
  wire [9:0] add_258826;
  wire [11:0] sel_258828;
  wire [9:0] add_258830;
  wire [11:0] sel_258833;
  wire [9:0] add_258835;
  wire [11:0] sel_258838;
  wire [11:0] add_258840;
  wire [11:0] sel_258842;
  wire [11:0] add_258844;
  wire [11:0] sel_258846;
  wire [11:0] add_258895;
  wire [11:0] sel_258897;
  wire [11:0] add_258900;
  wire [11:0] sel_258902;
  wire [15:0] array_index_258957;
  wire [15:0] array_index_258960;
  wire [10:0] add_258964;
  wire [10:0] add_258966;
  wire [10:0] add_258968;
  wire [11:0] sel_258971;
  wire [10:0] add_258973;
  wire [11:0] sel_258976;
  wire [11:0] add_258978;
  wire [11:0] sel_258980;
  wire [11:0] add_258982;
  wire [11:0] sel_258984;
  wire [11:0] add_258986;
  wire [11:0] sel_258988;
  wire [11:0] add_258990;
  wire [11:0] sel_258992;
  wire [11:0] add_258994;
  wire [11:0] sel_258996;
  wire [11:0] add_258998;
  wire [11:0] sel_259000;
  wire [11:0] add_259002;
  wire [11:0] sel_259004;
  wire [11:0] add_259006;
  wire [11:0] sel_259008;
  wire [11:0] add_259010;
  wire [11:0] sel_259012;
  wire [11:0] add_259014;
  wire [11:0] sel_259016;
  wire [11:0] add_259018;
  wire [11:0] sel_259020;
  wire [11:0] add_259022;
  wire [11:0] sel_259024;
  wire [9:0] add_259026;
  wire [11:0] sel_259028;
  wire [9:0] add_259030;
  wire [11:0] sel_259032;
  wire [9:0] add_259034;
  wire [11:0] sel_259037;
  wire [9:0] add_259039;
  wire [11:0] sel_259042;
  wire [11:0] add_259044;
  wire [11:0] sel_259046;
  wire [11:0] add_259048;
  wire [11:0] sel_259050;
  wire [11:0] add_259103;
  wire [11:0] sel_259105;
  wire [11:0] add_259108;
  wire [11:0] sel_259110;
  wire [15:0] array_index_259171;
  wire [15:0] array_index_259174;
  wire [11:0] add_259178;
  wire [11:0] add_259180;
  wire [10:0] add_259182;
  wire [11:0] sel_259184;
  wire [10:0] add_259186;
  wire [11:0] sel_259188;
  wire [10:0] add_259190;
  wire [11:0] sel_259193;
  wire [10:0] add_259195;
  wire [11:0] sel_259198;
  wire [11:0] add_259200;
  wire [11:0] sel_259202;
  wire [11:0] add_259204;
  wire [11:0] sel_259206;
  wire [11:0] add_259208;
  wire [11:0] sel_259210;
  wire [11:0] add_259212;
  wire [11:0] sel_259214;
  wire [11:0] add_259216;
  wire [11:0] sel_259218;
  wire [11:0] add_259220;
  wire [11:0] sel_259222;
  wire [11:0] add_259224;
  wire [11:0] sel_259226;
  wire [11:0] add_259228;
  wire [11:0] sel_259230;
  wire [11:0] add_259232;
  wire [11:0] sel_259234;
  wire [11:0] add_259236;
  wire [11:0] sel_259238;
  wire [11:0] add_259240;
  wire [11:0] sel_259242;
  wire [11:0] add_259244;
  wire [11:0] sel_259246;
  wire [9:0] add_259248;
  wire [11:0] sel_259250;
  wire [9:0] add_259252;
  wire [11:0] sel_259254;
  wire [9:0] add_259256;
  wire [11:0] sel_259259;
  wire [9:0] add_259261;
  wire [11:0] sel_259264;
  wire [11:0] add_259266;
  wire [11:0] sel_259268;
  wire [11:0] add_259270;
  wire [11:0] sel_259272;
  wire [11:0] add_259329;
  wire [11:0] sel_259331;
  wire [11:0] add_259334;
  wire [11:0] sel_259336;
  wire [15:0] array_index_259401;
  wire [15:0] array_index_259404;
  wire [11:0] add_259408;
  wire [11:0] add_259410;
  wire [11:0] add_259412;
  wire [11:0] sel_259414;
  wire [11:0] add_259416;
  wire [11:0] sel_259418;
  wire [10:0] add_259420;
  wire [11:0] sel_259422;
  wire [10:0] add_259424;
  wire [11:0] sel_259426;
  wire [10:0] add_259428;
  wire [11:0] sel_259431;
  wire [10:0] add_259433;
  wire [11:0] sel_259436;
  wire [11:0] add_259438;
  wire [11:0] sel_259440;
  wire [11:0] add_259442;
  wire [11:0] sel_259444;
  wire [11:0] add_259446;
  wire [11:0] sel_259448;
  wire [11:0] add_259450;
  wire [11:0] sel_259452;
  wire [11:0] add_259454;
  wire [11:0] sel_259456;
  wire [11:0] add_259458;
  wire [11:0] sel_259460;
  wire [11:0] add_259462;
  wire [11:0] sel_259464;
  wire [11:0] add_259466;
  wire [11:0] sel_259468;
  wire [11:0] add_259470;
  wire [11:0] sel_259472;
  wire [11:0] add_259474;
  wire [11:0] sel_259476;
  wire [11:0] add_259478;
  wire [11:0] sel_259480;
  wire [11:0] add_259482;
  wire [11:0] sel_259484;
  wire [9:0] add_259486;
  wire [11:0] sel_259488;
  wire [9:0] add_259490;
  wire [11:0] sel_259492;
  wire [9:0] add_259494;
  wire [11:0] sel_259497;
  wire [9:0] add_259499;
  wire [11:0] sel_259502;
  wire [11:0] add_259504;
  wire [11:0] sel_259506;
  wire [11:0] add_259508;
  wire [11:0] sel_259510;
  wire [11:0] add_259571;
  wire [11:0] sel_259573;
  wire [11:0] add_259576;
  wire [11:0] sel_259578;
  wire [15:0] array_index_259647;
  wire [15:0] array_index_259650;
  wire [10:0] add_259654;
  wire [10:0] add_259656;
  wire [11:0] add_259658;
  wire [11:0] sel_259660;
  wire [11:0] add_259662;
  wire [11:0] sel_259664;
  wire [11:0] add_259666;
  wire [11:0] sel_259668;
  wire [11:0] add_259670;
  wire [11:0] sel_259672;
  wire [10:0] add_259674;
  wire [11:0] sel_259676;
  wire [10:0] add_259678;
  wire [11:0] sel_259680;
  wire [10:0] add_259682;
  wire [11:0] sel_259685;
  wire [10:0] add_259687;
  wire [11:0] sel_259690;
  wire [11:0] add_259692;
  wire [11:0] sel_259694;
  wire [11:0] add_259696;
  wire [11:0] sel_259698;
  wire [11:0] add_259700;
  wire [11:0] sel_259702;
  wire [11:0] add_259704;
  wire [11:0] sel_259706;
  wire [11:0] add_259708;
  wire [11:0] sel_259710;
  wire [11:0] add_259712;
  wire [11:0] sel_259714;
  wire [11:0] add_259716;
  wire [11:0] sel_259718;
  wire [11:0] add_259720;
  wire [11:0] sel_259722;
  wire [11:0] add_259724;
  wire [11:0] sel_259726;
  wire [11:0] add_259728;
  wire [11:0] sel_259730;
  wire [11:0] add_259732;
  wire [11:0] sel_259734;
  wire [11:0] add_259736;
  wire [11:0] sel_259738;
  wire [9:0] add_259740;
  wire [11:0] sel_259742;
  wire [9:0] add_259744;
  wire [11:0] sel_259746;
  wire [9:0] add_259748;
  wire [11:0] sel_259751;
  wire [9:0] add_259753;
  wire [11:0] sel_259756;
  wire [11:0] add_259758;
  wire [11:0] sel_259760;
  wire [11:0] add_259762;
  wire [11:0] sel_259764;
  wire [11:0] add_259829;
  wire [11:0] sel_259831;
  wire [11:0] add_259834;
  wire [11:0] sel_259836;
  wire [15:0] array_index_259911;
  wire [15:0] array_index_259914;
  wire [11:0] add_259918;
  wire [11:0] add_259920;
  wire [10:0] add_259922;
  wire [11:0] sel_259924;
  wire [10:0] add_259926;
  wire [11:0] sel_259928;
  wire [11:0] add_259930;
  wire [11:0] sel_259932;
  wire [11:0] add_259934;
  wire [11:0] sel_259936;
  wire [11:0] add_259938;
  wire [11:0] sel_259940;
  wire [11:0] add_259942;
  wire [11:0] sel_259944;
  wire [10:0] add_259946;
  wire [11:0] sel_259948;
  wire [10:0] add_259950;
  wire [11:0] sel_259952;
  wire [10:0] add_259954;
  wire [11:0] sel_259957;
  wire [10:0] add_259959;
  wire [11:0] sel_259962;
  wire [11:0] add_259964;
  wire [11:0] sel_259966;
  wire [11:0] add_259968;
  wire [11:0] sel_259970;
  wire [11:0] add_259972;
  wire [11:0] sel_259974;
  wire [11:0] add_259976;
  wire [11:0] sel_259978;
  wire [11:0] add_259980;
  wire [11:0] sel_259982;
  wire [11:0] add_259984;
  wire [11:0] sel_259986;
  wire [11:0] add_259988;
  wire [11:0] sel_259990;
  wire [11:0] add_259992;
  wire [11:0] sel_259994;
  wire [11:0] add_259996;
  wire [11:0] sel_259998;
  wire [11:0] add_260000;
  wire [11:0] sel_260002;
  wire [11:0] add_260004;
  wire [11:0] sel_260006;
  wire [11:0] add_260008;
  wire [11:0] sel_260010;
  wire [9:0] add_260012;
  wire [11:0] sel_260014;
  wire [9:0] add_260016;
  wire [11:0] sel_260018;
  wire [9:0] add_260020;
  wire [11:0] sel_260023;
  wire [9:0] add_260025;
  wire [11:0] sel_260028;
  wire [11:0] add_260030;
  wire [11:0] sel_260032;
  wire [11:0] add_260034;
  wire [11:0] sel_260036;
  wire [11:0] add_260107;
  wire [11:0] sel_260109;
  wire [11:0] add_260112;
  wire [11:0] sel_260114;
  wire [10:0] add_260116;
  wire [10:0] add_260118;
  wire [15:0] array_index_260195;
  wire [15:0] array_index_260198;
  wire [11:0] add_260208;
  wire [11:0] sel_260210;
  wire [11:0] add_260212;
  wire [11:0] sel_260214;
  wire [10:0] add_260216;
  wire [11:0] sel_260218;
  wire [10:0] add_260220;
  wire [11:0] sel_260222;
  wire [11:0] add_260224;
  wire [11:0] sel_260226;
  wire [11:0] add_260228;
  wire [11:0] sel_260230;
  wire [11:0] add_260232;
  wire [11:0] sel_260234;
  wire [11:0] add_260236;
  wire [11:0] sel_260238;
  wire [10:0] add_260240;
  wire [11:0] sel_260242;
  wire [10:0] add_260244;
  wire [11:0] sel_260246;
  wire [10:0] add_260248;
  wire [11:0] sel_260251;
  wire [10:0] add_260253;
  wire [11:0] sel_260256;
  wire [11:0] add_260258;
  wire [11:0] sel_260260;
  wire [11:0] add_260262;
  wire [11:0] sel_260264;
  wire [11:0] add_260266;
  wire [11:0] sel_260268;
  wire [11:0] add_260270;
  wire [11:0] sel_260272;
  wire [11:0] add_260274;
  wire [11:0] sel_260276;
  wire [11:0] add_260278;
  wire [11:0] sel_260280;
  wire [11:0] add_260282;
  wire [11:0] sel_260284;
  wire [11:0] add_260286;
  wire [11:0] sel_260288;
  wire [11:0] add_260290;
  wire [11:0] sel_260292;
  wire [11:0] add_260294;
  wire [11:0] sel_260296;
  wire [11:0] add_260298;
  wire [11:0] sel_260300;
  wire [11:0] add_260302;
  wire [11:0] sel_260304;
  wire [9:0] add_260306;
  wire [11:0] sel_260308;
  wire [9:0] add_260310;
  wire [11:0] sel_260312;
  wire [9:0] add_260314;
  wire [11:0] sel_260317;
  wire [9:0] add_260319;
  wire [11:0] sel_260322;
  wire [11:0] add_260324;
  wire [11:0] sel_260326;
  wire [11:0] add_260328;
  wire [11:0] sel_260330;
  wire [11:0] add_260338;
  wire [11:0] add_260340;
  wire [11:0] add_260411;
  wire [11:0] sel_260413;
  wire [11:0] add_260416;
  wire [11:0] sel_260418;
  wire [10:0] add_260426;
  wire [11:0] sel_260428;
  wire [10:0] add_260430;
  wire [11:0] sel_260432;
  wire [15:0] array_index_260507;
  wire [15:0] array_index_260510;
  wire [10:0] add_260514;
  wire [10:0] add_260516;
  wire [11:0] add_260528;
  wire [11:0] sel_260530;
  wire [11:0] add_260532;
  wire [11:0] sel_260534;
  wire [10:0] add_260536;
  wire [11:0] sel_260538;
  wire [10:0] add_260540;
  wire [11:0] sel_260542;
  wire [11:0] add_260544;
  wire [11:0] sel_260546;
  wire [11:0] add_260548;
  wire [11:0] sel_260550;
  wire [11:0] add_260552;
  wire [11:0] sel_260554;
  wire [11:0] add_260556;
  wire [11:0] sel_260558;
  wire [10:0] add_260560;
  wire [11:0] sel_260562;
  wire [10:0] add_260564;
  wire [11:0] sel_260566;
  wire [10:0] add_260568;
  wire [11:0] sel_260571;
  wire [10:0] add_260573;
  wire [11:0] sel_260576;
  wire [11:0] add_260578;
  wire [11:0] sel_260580;
  wire [11:0] add_260582;
  wire [11:0] sel_260584;
  wire [11:0] add_260586;
  wire [11:0] sel_260588;
  wire [11:0] add_260590;
  wire [11:0] sel_260592;
  wire [11:0] add_260594;
  wire [11:0] sel_260596;
  wire [11:0] add_260598;
  wire [11:0] sel_260600;
  wire [11:0] add_260602;
  wire [11:0] sel_260604;
  wire [11:0] add_260606;
  wire [11:0] sel_260608;
  wire [11:0] add_260610;
  wire [11:0] sel_260612;
  wire [11:0] add_260614;
  wire [11:0] sel_260616;
  wire [11:0] add_260618;
  wire [11:0] sel_260620;
  wire [11:0] add_260622;
  wire [11:0] sel_260624;
  wire [9:0] add_260626;
  wire [11:0] sel_260628;
  wire [9:0] add_260630;
  wire [11:0] sel_260632;
  wire [9:0] add_260634;
  wire [11:0] sel_260637;
  wire [9:0] add_260639;
  wire [11:0] sel_260642;
  wire [11:0] add_260644;
  wire [11:0] sel_260646;
  wire [11:0] add_260648;
  wire [11:0] sel_260650;
  wire [11:0] add_260664;
  wire [11:0] sel_260666;
  wire [11:0] add_260668;
  wire [11:0] sel_260670;
  wire [11:0] add_260739;
  wire [11:0] sel_260741;
  wire [11:0] add_260744;
  wire [11:0] sel_260746;
  wire [11:0] add_260748;
  wire [11:0] add_260750;
  wire [10:0] add_260764;
  wire [11:0] sel_260766;
  wire [10:0] add_260768;
  wire [11:0] sel_260770;
  wire [15:0] array_index_260845;
  wire [15:0] array_index_260848;
  wire [10:0] add_260858;
  wire [11:0] sel_260860;
  wire [10:0] add_260862;
  wire [11:0] sel_260864;
  wire [11:0] add_260874;
  wire [11:0] sel_260876;
  wire [11:0] add_260878;
  wire [11:0] sel_260880;
  wire [10:0] add_260882;
  wire [11:0] sel_260884;
  wire [10:0] add_260886;
  wire [11:0] sel_260888;
  wire [11:0] add_260890;
  wire [11:0] sel_260892;
  wire [11:0] add_260894;
  wire [11:0] sel_260896;
  wire [11:0] add_260898;
  wire [11:0] sel_260900;
  wire [11:0] add_260902;
  wire [11:0] sel_260904;
  wire [10:0] add_260906;
  wire [11:0] sel_260908;
  wire [10:0] add_260910;
  wire [11:0] sel_260912;
  wire [10:0] add_260914;
  wire [11:0] sel_260917;
  wire [10:0] add_260919;
  wire [11:0] sel_260922;
  wire [11:0] add_260924;
  wire [11:0] sel_260926;
  wire [11:0] add_260928;
  wire [11:0] sel_260930;
  wire [11:0] add_260932;
  wire [11:0] sel_260934;
  wire [11:0] add_260936;
  wire [11:0] sel_260938;
  wire [11:0] add_260940;
  wire [11:0] sel_260942;
  wire [11:0] add_260944;
  wire [11:0] sel_260946;
  wire [11:0] add_260948;
  wire [11:0] sel_260950;
  wire [11:0] add_260952;
  wire [11:0] sel_260954;
  wire [11:0] add_260956;
  wire [11:0] sel_260958;
  wire [11:0] add_260960;
  wire [11:0] sel_260962;
  wire [11:0] add_260964;
  wire [11:0] sel_260966;
  wire [11:0] add_260968;
  wire [11:0] sel_260970;
  wire [9:0] add_260972;
  wire [11:0] sel_260974;
  wire [9:0] add_260976;
  wire [11:0] sel_260978;
  wire [9:0] add_260980;
  wire [11:0] sel_260983;
  wire [9:0] add_260985;
  wire [11:0] sel_260988;
  wire [11:0] add_260990;
  wire [11:0] sel_260992;
  wire [11:0] add_260994;
  wire [11:0] sel_260996;
  wire [11:0] add_261004;
  wire [11:0] add_261006;
  wire [11:0] add_261018;
  wire [11:0] sel_261020;
  wire [11:0] add_261022;
  wire [11:0] sel_261024;
  wire [11:0] add_261093;
  wire [11:0] sel_261095;
  wire [11:0] add_261098;
  wire [11:0] sel_261100;
  wire [11:0] add_261108;
  wire [11:0] sel_261110;
  wire [11:0] add_261112;
  wire [11:0] sel_261114;
  wire [10:0] add_261126;
  wire [11:0] sel_261128;
  wire [10:0] add_261130;
  wire [11:0] sel_261132;
  wire [15:0] array_index_261207;
  wire [15:0] array_index_261210;
  wire [9:0] add_261214;
  wire [9:0] add_261216;
  wire [10:0] add_261228;
  wire [11:0] sel_261230;
  wire [10:0] add_261232;
  wire [11:0] sel_261234;
  wire [11:0] add_261244;
  wire [11:0] sel_261246;
  wire [11:0] add_261248;
  wire [11:0] sel_261250;
  wire [10:0] add_261252;
  wire [11:0] sel_261254;
  wire [10:0] add_261256;
  wire [11:0] sel_261258;
  wire [11:0] add_261260;
  wire [11:0] sel_261262;
  wire [11:0] add_261264;
  wire [11:0] sel_261266;
  wire [11:0] add_261268;
  wire [11:0] sel_261270;
  wire [11:0] add_261272;
  wire [11:0] sel_261274;
  wire [10:0] add_261276;
  wire [11:0] sel_261278;
  wire [10:0] add_261280;
  wire [11:0] sel_261282;
  wire [10:0] add_261284;
  wire [11:0] sel_261287;
  wire [10:0] add_261289;
  wire [11:0] sel_261292;
  wire [11:0] add_261294;
  wire [11:0] sel_261296;
  wire [11:0] add_261298;
  wire [11:0] sel_261300;
  wire [11:0] add_261302;
  wire [11:0] sel_261304;
  wire [11:0] add_261306;
  wire [11:0] sel_261308;
  wire [11:0] add_261310;
  wire [11:0] sel_261312;
  wire [11:0] add_261314;
  wire [11:0] sel_261316;
  wire [11:0] add_261318;
  wire [11:0] sel_261320;
  wire [11:0] add_261322;
  wire [11:0] sel_261324;
  wire [11:0] add_261326;
  wire [11:0] sel_261328;
  wire [11:0] add_261330;
  wire [11:0] sel_261332;
  wire [11:0] add_261334;
  wire [11:0] sel_261336;
  wire [11:0] add_261338;
  wire [11:0] sel_261340;
  wire [9:0] add_261342;
  wire [11:0] sel_261344;
  wire [9:0] add_261346;
  wire [11:0] sel_261348;
  wire [9:0] add_261350;
  wire [11:0] sel_261353;
  wire [9:0] add_261355;
  wire [11:0] sel_261358;
  wire [11:0] add_261360;
  wire [11:0] sel_261362;
  wire [11:0] add_261364;
  wire [11:0] sel_261366;
  wire [11:0] add_261380;
  wire [11:0] sel_261382;
  wire [11:0] add_261384;
  wire [11:0] sel_261386;
  wire [11:0] add_261396;
  wire [11:0] sel_261398;
  wire [11:0] add_261400;
  wire [11:0] sel_261402;
  wire [11:0] add_261471;
  wire [11:0] sel_261473;
  wire [11:0] add_261476;
  wire [11:0] sel_261478;
  wire [11:0] add_261480;
  wire [11:0] add_261482;
  wire [11:0] add_261496;
  wire [11:0] sel_261498;
  wire [11:0] add_261500;
  wire [11:0] sel_261502;
  wire [10:0] add_261514;
  wire [11:0] sel_261516;
  wire [10:0] add_261518;
  wire [11:0] sel_261520;
  wire [15:0] array_index_261595;
  wire [15:0] array_index_261598;
  wire [9:0] add_261608;
  wire [11:0] sel_261610;
  wire [9:0] add_261612;
  wire [11:0] sel_261614;
  wire [10:0] add_261624;
  wire [11:0] sel_261626;
  wire [10:0] add_261628;
  wire [11:0] sel_261630;
  wire [11:0] add_261640;
  wire [11:0] sel_261642;
  wire [11:0] add_261644;
  wire [11:0] sel_261646;
  wire [10:0] add_261648;
  wire [11:0] sel_261650;
  wire [10:0] add_261652;
  wire [11:0] sel_261654;
  wire [11:0] add_261656;
  wire [11:0] sel_261658;
  wire [11:0] add_261660;
  wire [11:0] sel_261662;
  wire [11:0] add_261664;
  wire [11:0] sel_261666;
  wire [11:0] add_261668;
  wire [11:0] sel_261670;
  wire [10:0] add_261672;
  wire [11:0] sel_261674;
  wire [10:0] add_261676;
  wire [11:0] sel_261678;
  wire [10:0] add_261680;
  wire [11:0] sel_261683;
  wire [10:0] add_261685;
  wire [11:0] sel_261688;
  wire [11:0] add_261690;
  wire [11:0] sel_261692;
  wire [11:0] add_261694;
  wire [11:0] sel_261696;
  wire [11:0] add_261698;
  wire [11:0] sel_261700;
  wire [11:0] add_261702;
  wire [11:0] sel_261704;
  wire [11:0] add_261706;
  wire [11:0] sel_261708;
  wire [11:0] add_261710;
  wire [11:0] sel_261712;
  wire [11:0] add_261714;
  wire [11:0] sel_261716;
  wire [11:0] add_261718;
  wire [11:0] sel_261720;
  wire [11:0] add_261722;
  wire [11:0] sel_261724;
  wire [11:0] add_261726;
  wire [11:0] sel_261728;
  wire [11:0] add_261730;
  wire [11:0] sel_261732;
  wire [11:0] add_261734;
  wire [11:0] sel_261736;
  wire [9:0] add_261738;
  wire [11:0] sel_261740;
  wire [9:0] add_261742;
  wire [11:0] sel_261744;
  wire [9:0] add_261746;
  wire [11:0] sel_261749;
  wire [9:0] add_261751;
  wire [11:0] sel_261754;
  wire [11:0] add_261756;
  wire [11:0] sel_261758;
  wire [11:0] add_261760;
  wire [11:0] sel_261762;
  wire [9:0] add_261770;
  wire [9:0] add_261772;
  wire [11:0] add_261784;
  wire [11:0] sel_261786;
  wire [11:0] add_261788;
  wire [11:0] sel_261790;
  wire [11:0] add_261800;
  wire [11:0] sel_261802;
  wire [11:0] add_261804;
  wire [11:0] sel_261806;
  wire [11:0] add_261875;
  wire [11:0] sel_261877;
  wire [11:0] add_261880;
  wire [11:0] sel_261882;
  wire [11:0] add_261890;
  wire [11:0] sel_261892;
  wire [11:0] add_261894;
  wire [11:0] sel_261896;
  wire [11:0] add_261908;
  wire [11:0] sel_261910;
  wire [11:0] add_261912;
  wire [11:0] sel_261914;
  wire [10:0] add_261926;
  wire [11:0] sel_261928;
  wire [10:0] add_261930;
  wire [11:0] sel_261932;
  wire [15:0] array_index_262007;
  wire [15:0] array_index_262010;
  wire [11:0] add_262014;
  wire [11:0] add_262016;
  wire [9:0] add_262030;
  wire [11:0] sel_262032;
  wire [9:0] add_262034;
  wire [11:0] sel_262036;
  wire [10:0] add_262046;
  wire [11:0] sel_262048;
  wire [10:0] add_262050;
  wire [11:0] sel_262052;
  wire [11:0] add_262062;
  wire [11:0] sel_262064;
  wire [11:0] add_262066;
  wire [11:0] sel_262068;
  wire [10:0] add_262070;
  wire [11:0] sel_262072;
  wire [10:0] add_262074;
  wire [11:0] sel_262076;
  wire [11:0] add_262078;
  wire [11:0] sel_262080;
  wire [11:0] add_262082;
  wire [11:0] sel_262084;
  wire [11:0] add_262086;
  wire [11:0] sel_262088;
  wire [11:0] add_262090;
  wire [11:0] sel_262092;
  wire [10:0] add_262094;
  wire [11:0] sel_262096;
  wire [10:0] add_262098;
  wire [11:0] sel_262100;
  wire [10:0] add_262102;
  wire [11:0] sel_262105;
  wire [10:0] add_262107;
  wire [11:0] sel_262110;
  wire [11:0] add_262112;
  wire [11:0] sel_262114;
  wire [11:0] add_262116;
  wire [11:0] sel_262118;
  wire [11:0] add_262120;
  wire [11:0] sel_262122;
  wire [11:0] add_262124;
  wire [11:0] sel_262126;
  wire [11:0] add_262128;
  wire [11:0] sel_262130;
  wire [11:0] add_262132;
  wire [11:0] sel_262134;
  wire [11:0] add_262136;
  wire [11:0] sel_262138;
  wire [11:0] add_262140;
  wire [11:0] sel_262142;
  wire [11:0] add_262144;
  wire [11:0] sel_262146;
  wire [11:0] add_262148;
  wire [11:0] sel_262150;
  wire [11:0] add_262152;
  wire [11:0] sel_262154;
  wire [11:0] add_262156;
  wire [11:0] sel_262158;
  wire [9:0] add_262160;
  wire [11:0] sel_262162;
  wire [9:0] add_262164;
  wire [11:0] sel_262166;
  wire [9:0] add_262168;
  wire [11:0] sel_262171;
  wire [9:0] add_262173;
  wire [11:0] sel_262176;
  wire [11:0] add_262178;
  wire [11:0] sel_262180;
  wire [11:0] add_262182;
  wire [11:0] sel_262184;
  wire [9:0] add_262196;
  wire [11:0] sel_262198;
  wire [9:0] add_262200;
  wire [11:0] sel_262202;
  wire [11:0] add_262212;
  wire [11:0] sel_262214;
  wire [11:0] add_262216;
  wire [11:0] sel_262218;
  wire [11:0] add_262228;
  wire [11:0] sel_262230;
  wire [11:0] add_262232;
  wire [11:0] sel_262234;
  wire [11:0] add_262303;
  wire [11:0] sel_262305;
  wire [11:0] add_262308;
  wire [11:0] sel_262310;
  wire [11:0] add_262322;
  wire [11:0] sel_262324;
  wire [11:0] add_262326;
  wire [11:0] sel_262328;
  wire [11:0] add_262340;
  wire [11:0] sel_262342;
  wire [11:0] add_262344;
  wire [11:0] sel_262346;
  wire [10:0] add_262358;
  wire [11:0] sel_262360;
  wire [10:0] add_262362;
  wire [11:0] sel_262364;
  wire [15:0] array_index_262439;
  wire [15:0] array_index_262442;
  wire [11:0] add_262446;
  wire [11:0] sel_262448;
  wire [11:0] add_262450;
  wire [11:0] sel_262452;
  wire [9:0] add_262464;
  wire [11:0] sel_262466;
  wire [9:0] add_262468;
  wire [11:0] sel_262470;
  wire [10:0] add_262480;
  wire [11:0] sel_262482;
  wire [10:0] add_262484;
  wire [11:0] sel_262486;
  wire [11:0] add_262496;
  wire [11:0] sel_262498;
  wire [11:0] add_262500;
  wire [11:0] sel_262502;
  wire [10:0] add_262504;
  wire [11:0] sel_262506;
  wire [10:0] add_262508;
  wire [11:0] sel_262510;
  wire [11:0] add_262512;
  wire [11:0] sel_262514;
  wire [11:0] add_262516;
  wire [11:0] sel_262518;
  wire [11:0] add_262520;
  wire [11:0] sel_262522;
  wire [11:0] add_262524;
  wire [11:0] sel_262526;
  wire [10:0] add_262528;
  wire [11:0] sel_262530;
  wire [10:0] add_262532;
  wire [11:0] sel_262534;
  wire [10:0] add_262536;
  wire [11:0] sel_262539;
  wire [10:0] add_262541;
  wire [11:0] sel_262544;
  wire [11:0] add_262546;
  wire [11:0] sel_262548;
  wire [11:0] add_262550;
  wire [11:0] sel_262552;
  wire [11:0] add_262554;
  wire [11:0] sel_262556;
  wire [11:0] add_262558;
  wire [11:0] sel_262560;
  wire [11:0] add_262562;
  wire [11:0] sel_262564;
  wire [11:0] add_262566;
  wire [11:0] sel_262568;
  wire [11:0] add_262570;
  wire [11:0] sel_262572;
  wire [11:0] add_262574;
  wire [11:0] sel_262576;
  wire [11:0] add_262578;
  wire [11:0] sel_262580;
  wire [11:0] add_262582;
  wire [11:0] sel_262584;
  wire [11:0] add_262586;
  wire [11:0] sel_262588;
  wire [11:0] add_262590;
  wire [11:0] sel_262592;
  wire [9:0] add_262594;
  wire [11:0] sel_262596;
  wire [9:0] add_262598;
  wire [11:0] sel_262600;
  wire [9:0] add_262602;
  wire [11:0] sel_262605;
  wire [9:0] add_262607;
  wire [11:0] sel_262610;
  wire [11:0] add_262612;
  wire [11:0] sel_262614;
  wire [11:0] add_262616;
  wire [11:0] sel_262618;
  wire [9:0] add_262630;
  wire [11:0] sel_262632;
  wire [9:0] add_262634;
  wire [11:0] sel_262636;
  wire [11:0] add_262646;
  wire [11:0] sel_262648;
  wire [11:0] add_262650;
  wire [11:0] sel_262652;
  wire [11:0] add_262662;
  wire [11:0] sel_262664;
  wire [11:0] add_262666;
  wire [11:0] sel_262668;
  wire [11:0] add_262737;
  wire [11:0] sel_262739;
  wire [11:0] add_262742;
  wire [11:0] sel_262744;
  wire [11:0] add_262754;
  wire [11:0] sel_262756;
  wire [11:0] add_262758;
  wire [11:0] sel_262760;
  wire [11:0] add_262772;
  wire [11:0] sel_262774;
  wire [11:0] add_262776;
  wire [11:0] sel_262778;
  wire [10:0] add_262790;
  wire [11:0] sel_262792;
  wire [10:0] add_262794;
  wire [11:0] sel_262796;
  wire [15:0] array_index_262871;
  wire [15:0] array_index_262874;
  wire [11:0] add_262878;
  wire [11:0] sel_262880;
  wire [11:0] add_262882;
  wire [11:0] sel_262884;
  wire [9:0] add_262896;
  wire [11:0] sel_262898;
  wire [9:0] add_262900;
  wire [11:0] sel_262902;
  wire [10:0] add_262912;
  wire [11:0] sel_262914;
  wire [10:0] add_262916;
  wire [11:0] sel_262918;
  wire [11:0] add_262928;
  wire [11:0] sel_262930;
  wire [11:0] add_262932;
  wire [11:0] sel_262934;
  wire [10:0] add_262936;
  wire [11:0] sel_262938;
  wire [10:0] add_262940;
  wire [11:0] sel_262942;
  wire [11:0] add_262944;
  wire [11:0] sel_262946;
  wire [11:0] add_262948;
  wire [11:0] sel_262950;
  wire [11:0] add_262952;
  wire [11:0] sel_262954;
  wire [11:0] add_262956;
  wire [11:0] sel_262958;
  wire [10:0] add_262960;
  wire [11:0] sel_262962;
  wire [10:0] add_262964;
  wire [11:0] sel_262966;
  wire [10:0] add_262968;
  wire [11:0] sel_262971;
  wire [10:0] add_262973;
  wire [11:0] sel_262976;
  wire [11:0] add_262978;
  wire [11:0] sel_262980;
  wire [11:0] add_262982;
  wire [11:0] sel_262984;
  wire [11:0] add_262986;
  wire [11:0] sel_262988;
  wire [11:0] add_262990;
  wire [11:0] sel_262992;
  wire [11:0] add_262994;
  wire [11:0] sel_262996;
  wire [11:0] add_262998;
  wire [11:0] sel_263000;
  wire [11:0] add_263002;
  wire [11:0] sel_263004;
  wire [11:0] add_263006;
  wire [11:0] sel_263008;
  wire [11:0] add_263010;
  wire [11:0] sel_263012;
  wire [11:0] add_263014;
  wire [11:0] sel_263016;
  wire [11:0] add_263018;
  wire [11:0] sel_263020;
  wire [11:0] add_263022;
  wire [11:0] sel_263024;
  wire [9:0] add_263026;
  wire [11:0] sel_263028;
  wire [9:0] add_263030;
  wire [11:0] sel_263032;
  wire [9:0] add_263034;
  wire [11:0] sel_263037;
  wire [9:0] add_263039;
  wire [11:0] sel_263042;
  wire [11:0] add_263044;
  wire [11:0] sel_263046;
  wire [11:0] add_263048;
  wire [11:0] sel_263050;
  wire [9:0] add_263062;
  wire [11:0] sel_263064;
  wire [9:0] add_263066;
  wire [11:0] sel_263068;
  wire [11:0] add_263078;
  wire [11:0] sel_263080;
  wire [11:0] add_263082;
  wire [11:0] sel_263084;
  wire [11:0] add_263094;
  wire [11:0] sel_263096;
  wire [11:0] add_263098;
  wire [11:0] sel_263100;
  wire [11:0] add_263169;
  wire [11:0] sel_263171;
  wire [11:0] add_263174;
  wire [11:0] sel_263176;
  wire [11:0] add_263186;
  wire [11:0] sel_263188;
  wire [11:0] add_263190;
  wire [11:0] sel_263192;
  wire [11:0] add_263204;
  wire [11:0] sel_263206;
  wire [11:0] add_263208;
  wire [11:0] sel_263210;
  wire [10:0] add_263222;
  wire [11:0] sel_263224;
  wire [10:0] add_263226;
  wire [11:0] sel_263228;
  wire [15:0] array_index_263303;
  wire [15:0] array_index_263306;
  wire [11:0] add_263310;
  wire [11:0] sel_263312;
  wire [11:0] add_263314;
  wire [11:0] sel_263316;
  wire [9:0] add_263328;
  wire [11:0] sel_263330;
  wire [9:0] add_263332;
  wire [11:0] sel_263334;
  wire [10:0] add_263344;
  wire [11:0] sel_263346;
  wire [10:0] add_263348;
  wire [11:0] sel_263350;
  wire [11:0] add_263360;
  wire [11:0] sel_263362;
  wire [11:0] add_263364;
  wire [11:0] sel_263366;
  wire [10:0] add_263368;
  wire [11:0] sel_263370;
  wire [10:0] add_263372;
  wire [11:0] sel_263374;
  wire [11:0] add_263376;
  wire [11:0] sel_263378;
  wire [11:0] add_263380;
  wire [11:0] sel_263382;
  wire [11:0] add_263384;
  wire [11:0] sel_263386;
  wire [11:0] add_263388;
  wire [11:0] sel_263390;
  wire [10:0] add_263392;
  wire [11:0] sel_263394;
  wire [10:0] add_263396;
  wire [11:0] sel_263398;
  wire [10:0] add_263400;
  wire [11:0] sel_263403;
  wire [10:0] add_263405;
  wire [11:0] sel_263408;
  wire [11:0] add_263410;
  wire [11:0] sel_263412;
  wire [11:0] add_263414;
  wire [11:0] sel_263416;
  wire [11:0] add_263418;
  wire [11:0] sel_263420;
  wire [11:0] add_263422;
  wire [11:0] sel_263424;
  wire [11:0] add_263426;
  wire [11:0] sel_263428;
  wire [11:0] add_263430;
  wire [11:0] sel_263432;
  wire [11:0] add_263434;
  wire [11:0] sel_263436;
  wire [11:0] add_263438;
  wire [11:0] sel_263440;
  wire [11:0] add_263442;
  wire [11:0] sel_263444;
  wire [11:0] add_263446;
  wire [11:0] sel_263448;
  wire [11:0] add_263450;
  wire [11:0] sel_263452;
  wire [11:0] add_263454;
  wire [11:0] sel_263456;
  wire [9:0] add_263458;
  wire [11:0] sel_263460;
  wire [9:0] add_263462;
  wire [11:0] sel_263464;
  wire [9:0] add_263466;
  wire [11:0] sel_263469;
  wire [9:0] add_263471;
  wire [11:0] sel_263474;
  wire [11:0] add_263476;
  wire [11:0] sel_263478;
  wire [11:0] add_263480;
  wire [11:0] sel_263482;
  wire [9:0] add_263494;
  wire [11:0] sel_263496;
  wire [9:0] add_263498;
  wire [11:0] sel_263500;
  wire [11:0] add_263510;
  wire [11:0] sel_263512;
  wire [11:0] add_263514;
  wire [11:0] sel_263516;
  wire [11:0] add_263526;
  wire [11:0] sel_263528;
  wire [11:0] add_263530;
  wire [11:0] sel_263532;
  wire [11:0] add_263601;
  wire [11:0] sel_263603;
  wire [11:0] add_263606;
  wire [11:0] sel_263608;
  wire [11:0] add_263618;
  wire [11:0] sel_263620;
  wire [11:0] add_263622;
  wire [11:0] sel_263624;
  wire [11:0] add_263636;
  wire [11:0] sel_263638;
  wire [11:0] add_263640;
  wire [11:0] sel_263642;
  wire [10:0] add_263654;
  wire [11:0] sel_263656;
  wire [10:0] add_263658;
  wire [11:0] sel_263660;
  wire [15:0] array_index_263735;
  wire [15:0] array_index_263738;
  wire [11:0] add_263742;
  wire [11:0] sel_263744;
  wire [11:0] add_263746;
  wire [11:0] sel_263748;
  wire [9:0] add_263760;
  wire [11:0] sel_263762;
  wire [9:0] add_263764;
  wire [11:0] sel_263766;
  wire [10:0] add_263776;
  wire [11:0] sel_263778;
  wire [10:0] add_263780;
  wire [11:0] sel_263782;
  wire [11:0] add_263792;
  wire [11:0] sel_263794;
  wire [11:0] add_263796;
  wire [11:0] sel_263798;
  wire [10:0] add_263800;
  wire [11:0] sel_263802;
  wire [10:0] add_263804;
  wire [11:0] sel_263806;
  wire [11:0] add_263808;
  wire [11:0] sel_263810;
  wire [11:0] add_263812;
  wire [11:0] sel_263814;
  wire [11:0] add_263816;
  wire [11:0] sel_263818;
  wire [11:0] add_263820;
  wire [11:0] sel_263822;
  wire [10:0] add_263824;
  wire [11:0] sel_263826;
  wire [10:0] add_263828;
  wire [11:0] sel_263830;
  wire [10:0] add_263832;
  wire [11:0] sel_263835;
  wire [10:0] add_263837;
  wire [11:0] sel_263840;
  wire [11:0] add_263842;
  wire [11:0] sel_263844;
  wire [11:0] add_263846;
  wire [11:0] sel_263848;
  wire [11:0] add_263850;
  wire [11:0] sel_263852;
  wire [11:0] add_263854;
  wire [11:0] sel_263856;
  wire [11:0] add_263858;
  wire [11:0] sel_263860;
  wire [11:0] add_263862;
  wire [11:0] sel_263864;
  wire [11:0] add_263866;
  wire [11:0] sel_263868;
  wire [11:0] add_263870;
  wire [11:0] sel_263872;
  wire [11:0] add_263874;
  wire [11:0] sel_263876;
  wire [11:0] add_263878;
  wire [11:0] sel_263880;
  wire [11:0] add_263882;
  wire [11:0] sel_263884;
  wire [11:0] add_263886;
  wire [11:0] sel_263888;
  wire [9:0] add_263890;
  wire [11:0] sel_263892;
  wire [9:0] add_263894;
  wire [11:0] sel_263896;
  wire [9:0] add_263898;
  wire [11:0] sel_263901;
  wire [9:0] add_263903;
  wire [11:0] sel_263906;
  wire [11:0] add_263908;
  wire [11:0] sel_263910;
  wire [11:0] add_263912;
  wire [11:0] sel_263914;
  wire [9:0] add_263926;
  wire [11:0] sel_263928;
  wire [9:0] add_263930;
  wire [11:0] sel_263932;
  wire [11:0] add_263942;
  wire [11:0] sel_263944;
  wire [11:0] add_263946;
  wire [11:0] sel_263948;
  wire [11:0] add_263958;
  wire [11:0] sel_263960;
  wire [11:0] add_263962;
  wire [11:0] sel_263964;
  wire [11:0] add_264033;
  wire [11:0] sel_264035;
  wire [11:0] add_264038;
  wire [11:0] sel_264040;
  wire [11:0] add_264050;
  wire [11:0] sel_264052;
  wire [11:0] add_264054;
  wire [11:0] sel_264056;
  wire [11:0] add_264068;
  wire [11:0] sel_264070;
  wire [11:0] add_264072;
  wire [11:0] sel_264074;
  wire [10:0] add_264086;
  wire [11:0] sel_264088;
  wire [10:0] add_264090;
  wire [11:0] sel_264092;
  wire [15:0] array_index_264167;
  wire [15:0] array_index_264170;
  wire [11:0] add_264174;
  wire [11:0] sel_264176;
  wire [11:0] add_264178;
  wire [11:0] sel_264180;
  wire [9:0] add_264192;
  wire [11:0] sel_264194;
  wire [9:0] add_264196;
  wire [11:0] sel_264198;
  wire [10:0] add_264208;
  wire [11:0] sel_264210;
  wire [10:0] add_264212;
  wire [11:0] sel_264214;
  wire [11:0] add_264224;
  wire [11:0] sel_264226;
  wire [11:0] add_264228;
  wire [11:0] sel_264230;
  wire [10:0] add_264232;
  wire [11:0] sel_264234;
  wire [10:0] add_264236;
  wire [11:0] sel_264238;
  wire [11:0] add_264240;
  wire [11:0] sel_264242;
  wire [11:0] add_264244;
  wire [11:0] sel_264246;
  wire [11:0] add_264248;
  wire [11:0] sel_264250;
  wire [11:0] add_264252;
  wire [11:0] sel_264254;
  wire [10:0] add_264256;
  wire [11:0] sel_264258;
  wire [10:0] add_264260;
  wire [11:0] sel_264262;
  wire [10:0] add_264264;
  wire [11:0] sel_264267;
  wire [10:0] add_264269;
  wire [11:0] sel_264272;
  wire [11:0] add_264274;
  wire [11:0] sel_264276;
  wire [11:0] add_264278;
  wire [11:0] sel_264280;
  wire [11:0] add_264282;
  wire [11:0] sel_264284;
  wire [11:0] add_264286;
  wire [11:0] sel_264288;
  wire [11:0] add_264290;
  wire [11:0] sel_264292;
  wire [11:0] add_264294;
  wire [11:0] sel_264296;
  wire [11:0] add_264298;
  wire [11:0] sel_264300;
  wire [11:0] add_264302;
  wire [11:0] sel_264304;
  wire [11:0] add_264306;
  wire [11:0] sel_264308;
  wire [11:0] add_264310;
  wire [11:0] sel_264312;
  wire [11:0] add_264314;
  wire [11:0] sel_264316;
  wire [11:0] add_264318;
  wire [11:0] sel_264320;
  wire [9:0] add_264322;
  wire [11:0] sel_264324;
  wire [9:0] add_264326;
  wire [11:0] sel_264328;
  wire [9:0] add_264330;
  wire [11:0] sel_264333;
  wire [9:0] add_264335;
  wire [11:0] sel_264338;
  wire [11:0] add_264340;
  wire [11:0] sel_264342;
  wire [11:0] add_264344;
  wire [11:0] sel_264346;
  wire [9:0] add_264358;
  wire [11:0] sel_264360;
  wire [9:0] add_264362;
  wire [11:0] sel_264364;
  wire [11:0] add_264374;
  wire [11:0] sel_264376;
  wire [11:0] add_264378;
  wire [11:0] sel_264380;
  wire [11:0] add_264390;
  wire [11:0] sel_264392;
  wire [11:0] add_264394;
  wire [11:0] sel_264396;
  wire [11:0] add_264465;
  wire [11:0] sel_264467;
  wire [11:0] add_264470;
  wire [11:0] sel_264472;
  wire [11:0] add_264482;
  wire [11:0] sel_264484;
  wire [11:0] add_264486;
  wire [11:0] sel_264488;
  wire [11:0] add_264500;
  wire [11:0] sel_264502;
  wire [11:0] add_264504;
  wire [11:0] sel_264506;
  wire [10:0] add_264518;
  wire [11:0] sel_264520;
  wire [10:0] add_264522;
  wire [11:0] sel_264524;
  wire [15:0] array_index_264599;
  wire [15:0] array_index_264602;
  wire [11:0] add_264606;
  wire [11:0] sel_264608;
  wire [11:0] add_264610;
  wire [11:0] sel_264612;
  wire [9:0] add_264624;
  wire [11:0] sel_264626;
  wire [9:0] add_264628;
  wire [11:0] sel_264630;
  wire [10:0] add_264640;
  wire [11:0] sel_264642;
  wire [10:0] add_264644;
  wire [11:0] sel_264646;
  wire [11:0] add_264656;
  wire [11:0] sel_264658;
  wire [11:0] add_264660;
  wire [11:0] sel_264662;
  wire [10:0] add_264664;
  wire [11:0] sel_264666;
  wire [10:0] add_264668;
  wire [11:0] sel_264670;
  wire [11:0] add_264672;
  wire [11:0] sel_264674;
  wire [11:0] add_264676;
  wire [11:0] sel_264678;
  wire [11:0] add_264680;
  wire [11:0] sel_264682;
  wire [11:0] add_264684;
  wire [11:0] sel_264686;
  wire [10:0] add_264688;
  wire [11:0] sel_264690;
  wire [10:0] add_264692;
  wire [11:0] sel_264694;
  wire [10:0] add_264696;
  wire [11:0] sel_264699;
  wire [10:0] add_264701;
  wire [11:0] sel_264704;
  wire [11:0] add_264706;
  wire [11:0] sel_264708;
  wire [11:0] add_264710;
  wire [11:0] sel_264712;
  wire [11:0] add_264714;
  wire [11:0] sel_264716;
  wire [11:0] add_264718;
  wire [11:0] sel_264720;
  wire [11:0] add_264722;
  wire [11:0] sel_264724;
  wire [11:0] add_264726;
  wire [11:0] sel_264728;
  wire [11:0] add_264730;
  wire [11:0] sel_264732;
  wire [11:0] add_264734;
  wire [11:0] sel_264736;
  wire [11:0] add_264738;
  wire [11:0] sel_264740;
  wire [11:0] add_264742;
  wire [11:0] sel_264744;
  wire [11:0] add_264746;
  wire [11:0] sel_264748;
  wire [11:0] add_264750;
  wire [11:0] sel_264752;
  wire [9:0] add_264754;
  wire [11:0] sel_264756;
  wire [9:0] add_264758;
  wire [11:0] sel_264760;
  wire [9:0] add_264762;
  wire [11:0] sel_264765;
  wire [9:0] add_264767;
  wire [11:0] sel_264770;
  wire [11:0] add_264772;
  wire [11:0] sel_264774;
  wire [11:0] add_264776;
  wire [11:0] sel_264778;
  wire [9:0] add_264790;
  wire [11:0] sel_264792;
  wire [9:0] add_264794;
  wire [11:0] sel_264796;
  wire [11:0] add_264806;
  wire [11:0] sel_264808;
  wire [11:0] add_264810;
  wire [11:0] sel_264812;
  wire [11:0] add_264822;
  wire [11:0] sel_264824;
  wire [11:0] add_264826;
  wire [11:0] sel_264828;
  wire [11:0] add_264897;
  wire [11:0] sel_264899;
  wire [11:0] add_264902;
  wire [11:0] sel_264904;
  wire [11:0] add_264914;
  wire [11:0] sel_264916;
  wire [11:0] add_264918;
  wire [11:0] sel_264920;
  wire [11:0] add_264932;
  wire [11:0] sel_264934;
  wire [11:0] add_264936;
  wire [11:0] sel_264938;
  wire [10:0] add_264950;
  wire [11:0] sel_264952;
  wire [10:0] add_264954;
  wire [11:0] sel_264956;
  wire [15:0] array_index_265031;
  wire [15:0] array_index_265034;
  wire [11:0] add_265038;
  wire [11:0] sel_265040;
  wire [11:0] add_265042;
  wire [11:0] sel_265044;
  wire [9:0] add_265056;
  wire [11:0] sel_265058;
  wire [9:0] add_265060;
  wire [11:0] sel_265062;
  wire [10:0] add_265072;
  wire [11:0] sel_265074;
  wire [10:0] add_265076;
  wire [11:0] sel_265078;
  wire [11:0] add_265088;
  wire [11:0] sel_265090;
  wire [11:0] add_265092;
  wire [11:0] sel_265094;
  wire [10:0] add_265096;
  wire [11:0] sel_265098;
  wire [10:0] add_265100;
  wire [11:0] sel_265102;
  wire [11:0] add_265104;
  wire [11:0] sel_265106;
  wire [11:0] add_265108;
  wire [11:0] sel_265110;
  wire [11:0] add_265112;
  wire [11:0] sel_265114;
  wire [11:0] add_265116;
  wire [11:0] sel_265118;
  wire [10:0] add_265120;
  wire [11:0] sel_265122;
  wire [10:0] add_265124;
  wire [11:0] sel_265126;
  wire [10:0] add_265128;
  wire [11:0] sel_265131;
  wire [10:0] add_265133;
  wire [11:0] sel_265136;
  wire [11:0] add_265138;
  wire [11:0] sel_265140;
  wire [11:0] add_265142;
  wire [11:0] sel_265144;
  wire [11:0] add_265146;
  wire [11:0] sel_265148;
  wire [11:0] add_265150;
  wire [11:0] sel_265152;
  wire [11:0] add_265154;
  wire [11:0] sel_265156;
  wire [11:0] add_265158;
  wire [11:0] sel_265160;
  wire [11:0] add_265162;
  wire [11:0] sel_265164;
  wire [11:0] add_265166;
  wire [11:0] sel_265168;
  wire [11:0] add_265170;
  wire [11:0] sel_265172;
  wire [11:0] add_265174;
  wire [11:0] sel_265176;
  wire [11:0] add_265178;
  wire [11:0] sel_265180;
  wire [11:0] add_265182;
  wire [11:0] sel_265184;
  wire [9:0] add_265186;
  wire [11:0] sel_265188;
  wire [9:0] add_265190;
  wire [11:0] sel_265192;
  wire [9:0] add_265194;
  wire [11:0] sel_265197;
  wire [9:0] add_265199;
  wire [11:0] sel_265202;
  wire [11:0] add_265204;
  wire [11:0] sel_265206;
  wire [11:0] add_265208;
  wire [11:0] sel_265210;
  wire [9:0] add_265222;
  wire [11:0] sel_265224;
  wire [9:0] add_265226;
  wire [11:0] sel_265228;
  wire [11:0] add_265238;
  wire [11:0] sel_265240;
  wire [11:0] add_265242;
  wire [11:0] sel_265244;
  wire [11:0] add_265254;
  wire [11:0] sel_265256;
  wire [11:0] add_265258;
  wire [11:0] sel_265260;
  wire [11:0] add_265329;
  wire [11:0] sel_265331;
  wire [11:0] add_265334;
  wire [11:0] sel_265336;
  wire [11:0] add_265346;
  wire [11:0] sel_265348;
  wire [11:0] add_265350;
  wire [11:0] sel_265352;
  wire [11:0] add_265364;
  wire [11:0] sel_265366;
  wire [11:0] add_265368;
  wire [11:0] sel_265370;
  wire [10:0] add_265382;
  wire [11:0] sel_265384;
  wire [10:0] add_265386;
  wire [11:0] sel_265388;
  wire [15:0] array_index_265463;
  wire [15:0] array_index_265466;
  wire [11:0] add_265470;
  wire [11:0] sel_265472;
  wire [11:0] add_265474;
  wire [11:0] sel_265476;
  wire [9:0] add_265488;
  wire [11:0] sel_265490;
  wire [9:0] add_265492;
  wire [11:0] sel_265494;
  wire [10:0] add_265504;
  wire [11:0] sel_265506;
  wire [10:0] add_265508;
  wire [11:0] sel_265510;
  wire [11:0] add_265520;
  wire [11:0] sel_265522;
  wire [11:0] add_265524;
  wire [11:0] sel_265526;
  wire [10:0] add_265528;
  wire [11:0] sel_265530;
  wire [10:0] add_265532;
  wire [11:0] sel_265534;
  wire [11:0] add_265536;
  wire [11:0] sel_265538;
  wire [11:0] add_265540;
  wire [11:0] sel_265542;
  wire [11:0] add_265544;
  wire [11:0] sel_265546;
  wire [11:0] add_265548;
  wire [11:0] sel_265550;
  wire [10:0] add_265552;
  wire [11:0] sel_265554;
  wire [10:0] add_265556;
  wire [11:0] sel_265558;
  wire [10:0] add_265560;
  wire [11:0] sel_265563;
  wire [10:0] add_265565;
  wire [11:0] sel_265568;
  wire [11:0] add_265570;
  wire [11:0] sel_265572;
  wire [11:0] add_265574;
  wire [11:0] sel_265576;
  wire [11:0] add_265578;
  wire [11:0] sel_265580;
  wire [11:0] add_265582;
  wire [11:0] sel_265584;
  wire [11:0] add_265586;
  wire [11:0] sel_265588;
  wire [11:0] add_265590;
  wire [11:0] sel_265592;
  wire [11:0] add_265594;
  wire [11:0] sel_265596;
  wire [11:0] add_265598;
  wire [11:0] sel_265600;
  wire [11:0] add_265602;
  wire [11:0] sel_265604;
  wire [11:0] add_265606;
  wire [11:0] sel_265608;
  wire [11:0] add_265610;
  wire [11:0] sel_265612;
  wire [11:0] add_265614;
  wire [11:0] sel_265616;
  wire [9:0] add_265618;
  wire [11:0] sel_265620;
  wire [9:0] add_265622;
  wire [11:0] sel_265624;
  wire [9:0] add_265626;
  wire [11:0] sel_265629;
  wire [9:0] add_265631;
  wire [11:0] sel_265634;
  wire [11:0] add_265636;
  wire [11:0] sel_265638;
  wire [11:0] add_265640;
  wire [11:0] sel_265642;
  wire [9:0] add_265654;
  wire [11:0] sel_265656;
  wire [9:0] add_265658;
  wire [11:0] sel_265660;
  wire [11:0] add_265670;
  wire [11:0] sel_265672;
  wire [11:0] add_265674;
  wire [11:0] sel_265676;
  wire [11:0] add_265686;
  wire [11:0] sel_265688;
  wire [11:0] add_265690;
  wire [11:0] sel_265692;
  wire [11:0] add_265760;
  wire [11:0] sel_265762;
  wire [11:0] add_265764;
  wire [11:0] sel_265766;
  wire [11:0] add_265776;
  wire [11:0] sel_265778;
  wire [11:0] add_265780;
  wire [11:0] sel_265782;
  wire [11:0] add_265794;
  wire [11:0] sel_265796;
  wire [11:0] add_265798;
  wire [11:0] sel_265800;
  wire [10:0] add_265812;
  wire [11:0] sel_265814;
  wire [10:0] add_265816;
  wire [11:0] sel_265818;
  wire [11:0] add_265898;
  wire [11:0] sel_265900;
  wire [11:0] add_265902;
  wire [11:0] sel_265904;
  wire [9:0] add_265916;
  wire [11:0] sel_265918;
  wire [9:0] add_265920;
  wire [11:0] sel_265922;
  wire [10:0] add_265932;
  wire [11:0] sel_265934;
  wire [10:0] add_265936;
  wire [11:0] sel_265938;
  wire [11:0] add_265948;
  wire [11:0] sel_265950;
  wire [11:0] add_265952;
  wire [11:0] sel_265954;
  wire [10:0] add_265956;
  wire [11:0] sel_265958;
  wire [10:0] add_265960;
  wire [11:0] sel_265962;
  wire [11:0] add_265964;
  wire [11:0] sel_265966;
  wire [11:0] add_265968;
  wire [11:0] sel_265970;
  wire [11:0] add_265972;
  wire [11:0] sel_265974;
  wire [11:0] add_265976;
  wire [11:0] sel_265978;
  wire [10:0] add_265980;
  wire [11:0] sel_265982;
  wire [10:0] add_265984;
  wire [11:0] sel_265986;
  wire [10:0] add_265988;
  wire [11:0] sel_265991;
  wire [10:0] add_265993;
  wire [11:0] sel_265996;
  wire [11:0] add_265998;
  wire [11:0] sel_266000;
  wire [11:0] add_266002;
  wire [11:0] sel_266004;
  wire [11:0] add_266006;
  wire [11:0] sel_266008;
  wire [11:0] add_266010;
  wire [11:0] sel_266012;
  wire [11:0] add_266014;
  wire [11:0] sel_266016;
  wire [11:0] add_266018;
  wire [11:0] sel_266020;
  wire [11:0] add_266022;
  wire [11:0] sel_266024;
  wire [11:0] add_266026;
  wire [11:0] sel_266028;
  wire [11:0] add_266030;
  wire [11:0] sel_266032;
  wire [11:0] add_266034;
  wire [11:0] sel_266036;
  wire [11:0] add_266038;
  wire [11:0] sel_266040;
  wire [11:0] add_266042;
  wire [11:0] sel_266044;
  wire [9:0] add_266046;
  wire [11:0] sel_266048;
  wire [9:0] add_266050;
  wire [11:0] sel_266052;
  wire [9:0] add_266054;
  wire [11:0] sel_266057;
  wire [9:0] add_266059;
  wire [11:0] sel_266062;
  wire [11:0] add_266064;
  wire [11:0] sel_266066;
  wire [11:0] add_266068;
  wire [11:0] sel_266070;
  wire [9:0] add_266078;
  wire [11:0] sel_266080;
  wire [9:0] add_266082;
  wire [11:0] sel_266084;
  wire [11:0] add_266094;
  wire [11:0] sel_266096;
  wire [11:0] add_266098;
  wire [11:0] sel_266100;
  wire [11:0] add_266110;
  wire [11:0] sel_266112;
  wire [11:0] add_266114;
  wire [11:0] sel_266116;
  wire [11:0] add_266194;
  wire [11:0] sel_266196;
  wire [11:0] add_266198;
  wire [11:0] sel_266200;
  wire [11:0] add_266212;
  wire [11:0] sel_266214;
  wire [11:0] add_266216;
  wire [11:0] sel_266218;
  wire [10:0] add_266230;
  wire [11:0] sel_266232;
  wire [10:0] add_266234;
  wire [11:0] sel_266236;
  wire [11:0] add_266312;
  wire [11:0] sel_266314;
  wire [11:0] add_266316;
  wire [11:0] sel_266318;
  wire [9:0] add_266330;
  wire [11:0] sel_266332;
  wire [9:0] add_266334;
  wire [11:0] sel_266336;
  wire [10:0] add_266346;
  wire [11:0] sel_266348;
  wire [10:0] add_266350;
  wire [11:0] sel_266352;
  wire [11:0] add_266362;
  wire [11:0] sel_266364;
  wire [11:0] add_266366;
  wire [11:0] sel_266368;
  wire [10:0] add_266370;
  wire [11:0] sel_266372;
  wire [10:0] add_266374;
  wire [11:0] sel_266376;
  wire [11:0] add_266378;
  wire [11:0] sel_266380;
  wire [11:0] add_266382;
  wire [11:0] sel_266384;
  wire [11:0] add_266386;
  wire [11:0] sel_266388;
  wire [11:0] add_266390;
  wire [11:0] sel_266392;
  wire [10:0] add_266394;
  wire [11:0] sel_266396;
  wire [10:0] add_266398;
  wire [11:0] sel_266400;
  wire [10:0] add_266402;
  wire [11:0] sel_266405;
  wire [10:0] add_266407;
  wire [11:0] sel_266410;
  wire [11:0] add_266412;
  wire [11:0] sel_266414;
  wire [11:0] add_266416;
  wire [11:0] sel_266418;
  wire [11:0] add_266420;
  wire [11:0] sel_266422;
  wire [11:0] add_266424;
  wire [11:0] sel_266426;
  wire [11:0] add_266428;
  wire [11:0] sel_266430;
  wire [11:0] add_266432;
  wire [11:0] sel_266434;
  wire [11:0] add_266436;
  wire [11:0] sel_266438;
  wire [11:0] add_266440;
  wire [11:0] sel_266442;
  wire [11:0] add_266444;
  wire [11:0] sel_266446;
  wire [11:0] add_266448;
  wire [11:0] sel_266450;
  wire [11:0] add_266452;
  wire [11:0] sel_266454;
  wire [11:0] add_266456;
  wire [11:0] sel_266458;
  wire [9:0] add_266460;
  wire [11:0] sel_266462;
  wire [9:0] add_266464;
  wire [11:0] sel_266466;
  wire [9:0] add_266468;
  wire [11:0] sel_266471;
  wire [9:0] add_266473;
  wire [11:0] sel_266476;
  wire [1:0] concat_266479;
  wire [9:0] add_266486;
  wire [11:0] sel_266488;
  wire [9:0] add_266490;
  wire [11:0] sel_266492;
  wire [11:0] add_266502;
  wire [11:0] sel_266504;
  wire [11:0] add_266506;
  wire [11:0] sel_266508;
  wire [11:0] add_266518;
  wire [11:0] sel_266520;
  wire [11:0] add_266522;
  wire [11:0] sel_266524;
  wire [1:0] add_266588;
  wire [11:0] add_266598;
  wire [11:0] sel_266600;
  wire [11:0] add_266602;
  wire [11:0] sel_266604;
  wire [11:0] add_266616;
  wire [11:0] sel_266618;
  wire [11:0] add_266620;
  wire [11:0] sel_266622;
  wire [10:0] add_266634;
  wire [11:0] sel_266636;
  wire [10:0] add_266638;
  wire [11:0] sel_266640;
  wire [11:0] add_266710;
  wire [11:0] sel_266712;
  wire [11:0] add_266714;
  wire [11:0] sel_266716;
  wire [9:0] add_266728;
  wire [11:0] sel_266730;
  wire [9:0] add_266732;
  wire [11:0] sel_266734;
  wire [10:0] add_266744;
  wire [11:0] sel_266746;
  wire [10:0] add_266748;
  wire [11:0] sel_266750;
  wire [11:0] add_266760;
  wire [11:0] sel_266762;
  wire [11:0] add_266764;
  wire [11:0] sel_266766;
  wire [10:0] add_266768;
  wire [11:0] sel_266770;
  wire [10:0] add_266772;
  wire [11:0] sel_266774;
  wire [11:0] add_266776;
  wire [11:0] sel_266778;
  wire [11:0] add_266780;
  wire [11:0] sel_266782;
  wire [11:0] add_266784;
  wire [11:0] sel_266786;
  wire [11:0] add_266788;
  wire [11:0] sel_266790;
  wire [10:0] add_266792;
  wire [11:0] sel_266794;
  wire [10:0] add_266796;
  wire [11:0] sel_266798;
  wire [10:0] add_266800;
  wire [11:0] sel_266803;
  wire [10:0] add_266805;
  wire [11:0] sel_266808;
  wire [11:0] add_266810;
  wire [11:0] sel_266812;
  wire [11:0] add_266814;
  wire [11:0] sel_266816;
  wire [11:0] add_266818;
  wire [11:0] sel_266820;
  wire [11:0] add_266822;
  wire [11:0] sel_266824;
  wire [11:0] add_266826;
  wire [11:0] sel_266828;
  wire [11:0] add_266830;
  wire [11:0] sel_266832;
  wire [11:0] add_266834;
  wire [11:0] sel_266836;
  wire [11:0] add_266838;
  wire [11:0] sel_266840;
  wire [11:0] add_266842;
  wire [11:0] sel_266844;
  wire [11:0] add_266846;
  wire [11:0] sel_266848;
  wire [11:0] add_266850;
  wire [11:0] sel_266852;
  wire [11:0] add_266854;
  wire [11:0] sel_266856;
  wire [9:0] add_266858;
  wire [11:0] sel_266860;
  wire [9:0] add_266862;
  wire [11:0] sel_266864;
  wire [2:0] concat_266867;
  wire [9:0] add_266874;
  wire [11:0] sel_266876;
  wire [9:0] add_266878;
  wire [11:0] sel_266880;
  wire [11:0] add_266890;
  wire [11:0] sel_266892;
  wire [11:0] add_266894;
  wire [11:0] sel_266896;
  wire [11:0] add_266906;
  wire [11:0] sel_266908;
  wire [11:0] add_266910;
  wire [11:0] sel_266912;
  wire [2:0] add_266972;
  wire [11:0] add_266982;
  wire [11:0] sel_266984;
  wire [11:0] add_266986;
  wire [11:0] sel_266988;
  wire [11:0] add_267000;
  wire [11:0] sel_267002;
  wire [11:0] add_267004;
  wire [11:0] sel_267006;
  wire [10:0] add_267018;
  wire [11:0] sel_267020;
  wire [10:0] add_267022;
  wire [11:0] sel_267024;
  wire [11:0] add_267088;
  wire [11:0] sel_267090;
  wire [11:0] add_267092;
  wire [11:0] sel_267094;
  wire [9:0] add_267106;
  wire [11:0] sel_267108;
  wire [9:0] add_267110;
  wire [11:0] sel_267112;
  wire [10:0] add_267122;
  wire [11:0] sel_267124;
  wire [10:0] add_267126;
  wire [11:0] sel_267128;
  wire [11:0] add_267138;
  wire [11:0] sel_267140;
  wire [11:0] add_267142;
  wire [11:0] sel_267144;
  wire [10:0] add_267146;
  wire [11:0] sel_267148;
  wire [10:0] add_267150;
  wire [11:0] sel_267152;
  wire [11:0] add_267154;
  wire [11:0] sel_267156;
  wire [11:0] add_267158;
  wire [11:0] sel_267160;
  wire [11:0] add_267162;
  wire [11:0] sel_267164;
  wire [11:0] add_267166;
  wire [11:0] sel_267168;
  wire [10:0] add_267170;
  wire [11:0] sel_267172;
  wire [10:0] add_267174;
  wire [11:0] sel_267176;
  wire [10:0] add_267178;
  wire [11:0] sel_267181;
  wire [10:0] add_267183;
  wire [11:0] sel_267186;
  wire [11:0] add_267188;
  wire [11:0] sel_267190;
  wire [11:0] add_267192;
  wire [11:0] sel_267194;
  wire [11:0] add_267196;
  wire [11:0] sel_267198;
  wire [11:0] add_267200;
  wire [11:0] sel_267202;
  wire [11:0] add_267204;
  wire [11:0] sel_267206;
  wire [11:0] add_267208;
  wire [11:0] sel_267210;
  wire [11:0] add_267212;
  wire [11:0] sel_267214;
  wire [11:0] add_267216;
  wire [11:0] sel_267218;
  wire [11:0] add_267220;
  wire [11:0] sel_267222;
  wire [11:0] add_267224;
  wire [11:0] sel_267226;
  wire [11:0] add_267228;
  wire [11:0] sel_267230;
  wire [11:0] add_267232;
  wire [11:0] sel_267234;
  wire [3:0] concat_267237;
  wire [9:0] add_267244;
  wire [11:0] sel_267246;
  wire [9:0] add_267248;
  wire [11:0] sel_267250;
  wire [11:0] add_267260;
  wire [11:0] sel_267262;
  wire [11:0] add_267264;
  wire [11:0] sel_267266;
  wire [11:0] add_267276;
  wire [11:0] sel_267278;
  wire [11:0] add_267280;
  wire [11:0] sel_267282;
  wire [3:0] add_267338;
  wire [11:0] add_267348;
  wire [11:0] sel_267350;
  wire [11:0] add_267352;
  wire [11:0] sel_267354;
  wire [11:0] add_267366;
  wire [11:0] sel_267368;
  wire [11:0] add_267370;
  wire [11:0] sel_267372;
  wire [10:0] add_267384;
  wire [11:0] sel_267386;
  wire [10:0] add_267388;
  wire [11:0] sel_267390;
  wire [11:0] add_267448;
  wire [11:0] sel_267450;
  wire [11:0] add_267452;
  wire [11:0] sel_267454;
  wire [9:0] add_267466;
  wire [11:0] sel_267468;
  wire [9:0] add_267470;
  wire [11:0] sel_267472;
  wire [10:0] add_267482;
  wire [11:0] sel_267484;
  wire [10:0] add_267486;
  wire [11:0] sel_267488;
  wire [11:0] add_267498;
  wire [11:0] sel_267500;
  wire [11:0] add_267502;
  wire [11:0] sel_267504;
  wire [10:0] add_267506;
  wire [11:0] sel_267508;
  wire [10:0] add_267510;
  wire [11:0] sel_267512;
  wire [11:0] add_267514;
  wire [11:0] sel_267516;
  wire [11:0] add_267518;
  wire [11:0] sel_267520;
  wire [11:0] add_267522;
  wire [11:0] sel_267524;
  wire [11:0] add_267526;
  wire [11:0] sel_267528;
  wire [10:0] add_267530;
  wire [11:0] sel_267532;
  wire [10:0] add_267534;
  wire [11:0] sel_267536;
  wire [10:0] add_267538;
  wire [11:0] sel_267541;
  wire [10:0] add_267543;
  wire [11:0] sel_267546;
  wire [11:0] add_267548;
  wire [11:0] sel_267550;
  wire [11:0] add_267552;
  wire [11:0] sel_267554;
  wire [11:0] add_267556;
  wire [11:0] sel_267558;
  wire [11:0] add_267560;
  wire [11:0] sel_267562;
  wire [11:0] add_267564;
  wire [11:0] sel_267566;
  wire [11:0] add_267568;
  wire [11:0] sel_267570;
  wire [11:0] add_267572;
  wire [11:0] sel_267574;
  wire [11:0] add_267576;
  wire [11:0] sel_267578;
  wire [11:0] add_267580;
  wire [11:0] sel_267582;
  wire [11:0] add_267584;
  wire [11:0] sel_267586;
  wire [4:0] concat_267589;
  wire [9:0] add_267596;
  wire [11:0] sel_267598;
  wire [9:0] add_267600;
  wire [11:0] sel_267602;
  wire [11:0] add_267612;
  wire [11:0] sel_267614;
  wire [11:0] add_267616;
  wire [11:0] sel_267618;
  wire [11:0] add_267628;
  wire [11:0] sel_267630;
  wire [11:0] add_267632;
  wire [11:0] sel_267634;
  wire [4:0] add_267686;
  wire [11:0] add_267696;
  wire [11:0] sel_267698;
  wire [11:0] add_267700;
  wire [11:0] sel_267702;
  wire [11:0] add_267714;
  wire [11:0] sel_267716;
  wire [11:0] add_267718;
  wire [11:0] sel_267720;
  wire [10:0] add_267732;
  wire [11:0] sel_267734;
  wire [10:0] add_267736;
  wire [11:0] sel_267738;
  wire [11:0] add_267792;
  wire [11:0] sel_267794;
  wire [11:0] add_267796;
  wire [11:0] sel_267798;
  wire [9:0] add_267810;
  wire [11:0] sel_267812;
  wire [9:0] add_267814;
  wire [11:0] sel_267816;
  wire [10:0] add_267826;
  wire [11:0] sel_267828;
  wire [10:0] add_267830;
  wire [11:0] sel_267832;
  wire [11:0] add_267842;
  wire [11:0] sel_267844;
  wire [11:0] add_267846;
  wire [11:0] sel_267848;
  wire [10:0] add_267850;
  wire [11:0] sel_267852;
  wire [10:0] add_267854;
  wire [11:0] sel_267856;
  wire [11:0] add_267858;
  wire [11:0] sel_267860;
  wire [11:0] add_267862;
  wire [11:0] sel_267864;
  wire [11:0] add_267866;
  wire [11:0] sel_267868;
  wire [11:0] add_267870;
  wire [11:0] sel_267872;
  wire [10:0] add_267874;
  wire [11:0] sel_267876;
  wire [10:0] add_267878;
  wire [11:0] sel_267880;
  wire [10:0] add_267882;
  wire [11:0] sel_267885;
  wire [10:0] add_267887;
  wire [11:0] sel_267890;
  wire [11:0] add_267892;
  wire [11:0] sel_267894;
  wire [11:0] add_267896;
  wire [11:0] sel_267898;
  wire [11:0] add_267900;
  wire [11:0] sel_267902;
  wire [11:0] add_267904;
  wire [11:0] sel_267906;
  wire [11:0] add_267908;
  wire [11:0] sel_267910;
  wire [11:0] add_267912;
  wire [11:0] sel_267914;
  wire [11:0] add_267916;
  wire [11:0] sel_267918;
  wire [11:0] add_267920;
  wire [11:0] sel_267922;
  wire [5:0] concat_267925;
  wire [9:0] add_267932;
  wire [11:0] sel_267934;
  wire [9:0] add_267936;
  wire [11:0] sel_267938;
  wire [11:0] add_267948;
  wire [11:0] sel_267950;
  wire [11:0] add_267952;
  wire [11:0] sel_267954;
  wire [11:0] add_267964;
  wire [11:0] sel_267966;
  wire [11:0] add_267968;
  wire [11:0] sel_267970;
  wire [5:0] add_268018;
  wire [11:0] add_268028;
  wire [11:0] sel_268030;
  wire [11:0] add_268032;
  wire [11:0] sel_268034;
  wire [11:0] add_268046;
  wire [11:0] sel_268048;
  wire [11:0] add_268050;
  wire [11:0] sel_268052;
  wire [10:0] add_268064;
  wire [11:0] sel_268066;
  wire [10:0] add_268068;
  wire [11:0] sel_268070;
  wire [11:0] add_268120;
  wire [11:0] sel_268122;
  wire [11:0] add_268124;
  wire [11:0] sel_268126;
  wire [9:0] add_268138;
  wire [11:0] sel_268140;
  wire [9:0] add_268142;
  wire [11:0] sel_268144;
  wire [10:0] add_268154;
  wire [11:0] sel_268156;
  wire [10:0] add_268158;
  wire [11:0] sel_268160;
  wire [11:0] add_268170;
  wire [11:0] sel_268172;
  wire [11:0] add_268174;
  wire [11:0] sel_268176;
  wire [10:0] add_268178;
  wire [11:0] sel_268180;
  wire [10:0] add_268182;
  wire [11:0] sel_268184;
  wire [11:0] add_268186;
  wire [11:0] sel_268188;
  wire [11:0] add_268190;
  wire [11:0] sel_268192;
  wire [11:0] add_268194;
  wire [11:0] sel_268196;
  wire [11:0] add_268198;
  wire [11:0] sel_268200;
  wire [10:0] add_268202;
  wire [11:0] sel_268204;
  wire [10:0] add_268206;
  wire [11:0] sel_268208;
  wire [10:0] add_268210;
  wire [11:0] sel_268213;
  wire [10:0] add_268215;
  wire [11:0] sel_268218;
  wire [11:0] add_268220;
  wire [11:0] sel_268222;
  wire [11:0] add_268224;
  wire [11:0] sel_268226;
  wire [11:0] add_268228;
  wire [11:0] sel_268230;
  wire [11:0] add_268232;
  wire [11:0] sel_268234;
  wire [11:0] add_268236;
  wire [11:0] sel_268238;
  wire [11:0] add_268240;
  wire [11:0] sel_268242;
  wire [6:0] concat_268245;
  wire [9:0] add_268252;
  wire [11:0] sel_268254;
  wire [9:0] add_268256;
  wire [11:0] sel_268258;
  wire [11:0] add_268268;
  wire [11:0] sel_268270;
  wire [11:0] add_268272;
  wire [11:0] sel_268274;
  wire [11:0] add_268284;
  wire [11:0] sel_268286;
  wire [11:0] add_268288;
  wire [11:0] sel_268290;
  wire [6:0] add_268334;
  wire [11:0] add_268344;
  wire [11:0] sel_268346;
  wire [11:0] add_268348;
  wire [11:0] sel_268350;
  wire [11:0] add_268362;
  wire [11:0] sel_268364;
  wire [11:0] add_268366;
  wire [11:0] sel_268368;
  wire [10:0] add_268380;
  wire [11:0] sel_268382;
  wire [10:0] add_268384;
  wire [11:0] sel_268386;
  wire [11:0] add_268432;
  wire [11:0] sel_268434;
  wire [11:0] add_268436;
  wire [11:0] sel_268438;
  wire [9:0] add_268450;
  wire [11:0] sel_268452;
  wire [9:0] add_268454;
  wire [11:0] sel_268456;
  wire [10:0] add_268466;
  wire [11:0] sel_268468;
  wire [10:0] add_268470;
  wire [11:0] sel_268472;
  wire [11:0] add_268482;
  wire [11:0] sel_268484;
  wire [11:0] add_268486;
  wire [11:0] sel_268488;
  wire [10:0] add_268490;
  wire [11:0] sel_268492;
  wire [10:0] add_268494;
  wire [11:0] sel_268496;
  wire [11:0] add_268498;
  wire [11:0] sel_268500;
  wire [11:0] add_268502;
  wire [11:0] sel_268504;
  wire [11:0] add_268506;
  wire [11:0] sel_268508;
  wire [11:0] add_268510;
  wire [11:0] sel_268512;
  wire [10:0] add_268514;
  wire [11:0] sel_268516;
  wire [10:0] add_268518;
  wire [11:0] sel_268520;
  wire [10:0] add_268522;
  wire [11:0] sel_268525;
  wire [10:0] add_268527;
  wire [11:0] sel_268530;
  wire [11:0] add_268532;
  wire [11:0] sel_268534;
  wire [11:0] add_268536;
  wire [11:0] sel_268538;
  wire [11:0] add_268540;
  wire [11:0] sel_268542;
  wire [11:0] add_268544;
  wire [11:0] sel_268546;
  wire [7:0] concat_268549;
  wire [9:0] add_268556;
  wire [11:0] sel_268558;
  wire [9:0] add_268560;
  wire [11:0] sel_268562;
  wire [11:0] add_268572;
  wire [11:0] sel_268574;
  wire [11:0] add_268576;
  wire [11:0] sel_268578;
  wire [11:0] add_268588;
  wire [11:0] sel_268590;
  wire [11:0] add_268592;
  wire [11:0] sel_268594;
  wire [7:0] add_268634;
  wire [11:0] add_268644;
  wire [11:0] sel_268646;
  wire [11:0] add_268648;
  wire [11:0] sel_268650;
  wire [11:0] add_268662;
  wire [11:0] sel_268664;
  wire [11:0] add_268666;
  wire [11:0] sel_268668;
  wire [10:0] add_268680;
  wire [11:0] sel_268682;
  wire [10:0] add_268684;
  wire [11:0] sel_268686;
  wire [11:0] add_268728;
  wire [11:0] sel_268730;
  wire [11:0] add_268732;
  wire [11:0] sel_268734;
  wire [9:0] add_268746;
  wire [11:0] sel_268748;
  wire [9:0] add_268750;
  wire [11:0] sel_268752;
  wire [10:0] add_268762;
  wire [11:0] sel_268764;
  wire [10:0] add_268766;
  wire [11:0] sel_268768;
  wire [11:0] add_268778;
  wire [11:0] sel_268780;
  wire [11:0] add_268782;
  wire [11:0] sel_268784;
  wire [10:0] add_268786;
  wire [11:0] sel_268788;
  wire [10:0] add_268790;
  wire [11:0] sel_268792;
  wire [11:0] add_268794;
  wire [11:0] sel_268796;
  wire [11:0] add_268798;
  wire [11:0] sel_268800;
  wire [11:0] add_268802;
  wire [11:0] sel_268804;
  wire [11:0] add_268806;
  wire [11:0] sel_268808;
  wire [10:0] add_268810;
  wire [11:0] sel_268812;
  wire [10:0] add_268814;
  wire [11:0] sel_268816;
  wire [10:0] add_268818;
  wire [11:0] sel_268821;
  wire [10:0] add_268823;
  wire [11:0] sel_268826;
  wire [11:0] add_268828;
  wire [11:0] sel_268830;
  wire [11:0] add_268832;
  wire [11:0] sel_268834;
  wire [8:0] concat_268837;
  wire [9:0] add_268844;
  wire [11:0] sel_268846;
  wire [9:0] add_268848;
  wire [11:0] sel_268850;
  wire [11:0] add_268860;
  wire [11:0] sel_268862;
  wire [11:0] add_268864;
  wire [11:0] sel_268866;
  wire [11:0] add_268876;
  wire [11:0] sel_268878;
  wire [11:0] add_268880;
  wire [11:0] sel_268882;
  wire [8:0] add_268918;
  wire [11:0] add_268928;
  wire [11:0] sel_268930;
  wire [11:0] add_268932;
  wire [11:0] sel_268934;
  wire [11:0] add_268946;
  wire [11:0] sel_268948;
  wire [11:0] add_268950;
  wire [11:0] sel_268952;
  wire [10:0] add_268964;
  wire [11:0] sel_268966;
  wire [10:0] add_268968;
  wire [11:0] sel_268970;
  wire [11:0] add_269008;
  wire [11:0] sel_269010;
  wire [11:0] add_269012;
  wire [11:0] sel_269014;
  wire [9:0] add_269026;
  wire [11:0] sel_269028;
  wire [9:0] add_269030;
  wire [11:0] sel_269032;
  wire [10:0] add_269042;
  wire [11:0] sel_269044;
  wire [10:0] add_269046;
  wire [11:0] sel_269048;
  wire [11:0] add_269058;
  wire [11:0] sel_269060;
  wire [11:0] add_269062;
  wire [11:0] sel_269064;
  wire [10:0] add_269066;
  wire [11:0] sel_269068;
  wire [10:0] add_269070;
  wire [11:0] sel_269072;
  wire [11:0] add_269074;
  wire [11:0] sel_269076;
  wire [11:0] add_269078;
  wire [11:0] sel_269080;
  wire [11:0] add_269082;
  wire [11:0] sel_269084;
  wire [11:0] add_269086;
  wire [11:0] sel_269088;
  wire [10:0] add_269090;
  wire [11:0] sel_269092;
  wire [10:0] add_269094;
  wire [11:0] sel_269096;
  wire [10:0] add_269098;
  wire [11:0] sel_269101;
  wire [10:0] add_269103;
  wire [11:0] sel_269106;
  wire [9:0] concat_269109;
  wire [9:0] add_269116;
  wire [11:0] sel_269118;
  wire [9:0] add_269120;
  wire [11:0] sel_269122;
  wire [11:0] add_269132;
  wire [11:0] sel_269134;
  wire [11:0] add_269136;
  wire [11:0] sel_269138;
  wire [11:0] add_269148;
  wire [11:0] sel_269150;
  wire [11:0] add_269152;
  wire [11:0] sel_269154;
  wire [9:0] add_269186;
  wire [11:0] add_269196;
  wire [11:0] sel_269198;
  wire [11:0] add_269200;
  wire [11:0] sel_269202;
  wire [11:0] add_269214;
  wire [11:0] sel_269216;
  wire [11:0] add_269218;
  wire [11:0] sel_269220;
  wire [10:0] add_269232;
  wire [11:0] sel_269234;
  wire [10:0] add_269236;
  wire [11:0] sel_269238;
  wire [11:0] add_269270;
  wire [11:0] sel_269272;
  wire [11:0] add_269274;
  wire [11:0] sel_269276;
  wire [9:0] add_269288;
  wire [11:0] sel_269290;
  wire [9:0] add_269292;
  wire [11:0] sel_269294;
  wire [10:0] add_269304;
  wire [11:0] sel_269306;
  wire [10:0] add_269308;
  wire [11:0] sel_269310;
  wire [11:0] add_269320;
  wire [11:0] sel_269322;
  wire [11:0] add_269324;
  wire [11:0] sel_269326;
  wire [10:0] add_269328;
  wire [11:0] sel_269330;
  wire [10:0] add_269332;
  wire [11:0] sel_269334;
  wire [11:0] add_269336;
  wire [11:0] sel_269338;
  wire [11:0] add_269340;
  wire [11:0] sel_269342;
  wire [11:0] add_269344;
  wire [11:0] sel_269346;
  wire [11:0] add_269348;
  wire [11:0] sel_269350;
  wire [10:0] add_269352;
  wire [11:0] sel_269354;
  wire [10:0] add_269356;
  wire [11:0] sel_269358;
  wire [10:0] concat_269361;
  wire [9:0] add_269368;
  wire [11:0] sel_269370;
  wire [9:0] add_269372;
  wire [11:0] sel_269374;
  wire [11:0] add_269384;
  wire [11:0] sel_269386;
  wire [11:0] add_269388;
  wire [11:0] sel_269390;
  wire [11:0] add_269400;
  wire [11:0] sel_269402;
  wire [11:0] add_269404;
  wire [11:0] sel_269406;
  wire [10:0] add_269434;
  wire [11:0] add_269444;
  wire [11:0] sel_269446;
  wire [11:0] add_269448;
  wire [11:0] sel_269450;
  wire [11:0] add_269462;
  wire [11:0] sel_269464;
  wire [11:0] add_269466;
  wire [11:0] sel_269468;
  wire [10:0] add_269480;
  wire [11:0] sel_269482;
  wire [10:0] add_269484;
  wire [11:0] sel_269486;
  wire [11:0] add_269512;
  wire [11:0] sel_269514;
  wire [11:0] add_269516;
  wire [11:0] sel_269518;
  wire [9:0] add_269530;
  wire [11:0] sel_269532;
  wire [9:0] add_269534;
  wire [11:0] sel_269536;
  wire [10:0] add_269546;
  wire [11:0] sel_269548;
  wire [10:0] add_269550;
  wire [11:0] sel_269552;
  wire [11:0] add_269562;
  wire [11:0] sel_269564;
  wire [11:0] add_269566;
  wire [11:0] sel_269568;
  wire [10:0] add_269570;
  wire [11:0] sel_269572;
  wire [10:0] add_269574;
  wire [11:0] sel_269576;
  wire [11:0] add_269578;
  wire [11:0] sel_269580;
  wire [11:0] add_269582;
  wire [11:0] sel_269584;
  wire [11:0] add_269586;
  wire [11:0] sel_269588;
  wire [11:0] add_269590;
  wire [11:0] sel_269592;
  wire [11:0] concat_269595;
  wire [9:0] add_269602;
  wire [11:0] sel_269604;
  wire [9:0] add_269606;
  wire [11:0] sel_269608;
  wire [11:0] add_269618;
  wire [11:0] sel_269620;
  wire [11:0] add_269622;
  wire [11:0] sel_269624;
  wire [11:0] add_269634;
  wire [11:0] sel_269636;
  wire [11:0] add_269638;
  wire [11:0] sel_269640;
  wire [11:0] add_269664;
  wire [11:0] add_269674;
  wire [11:0] sel_269676;
  wire [11:0] add_269678;
  wire [11:0] sel_269680;
  wire [11:0] add_269692;
  wire [11:0] sel_269694;
  wire [11:0] add_269696;
  wire [11:0] sel_269698;
  wire [10:0] add_269710;
  wire [11:0] sel_269712;
  wire [10:0] add_269714;
  wire [11:0] sel_269716;
  wire [11:0] add_269736;
  wire [11:0] sel_269738;
  wire [11:0] add_269740;
  wire [11:0] sel_269742;
  wire [9:0] add_269754;
  wire [11:0] sel_269756;
  wire [9:0] add_269758;
  wire [11:0] sel_269760;
  wire [10:0] add_269770;
  wire [11:0] sel_269772;
  wire [10:0] add_269774;
  wire [11:0] sel_269776;
  wire [11:0] add_269786;
  wire [11:0] sel_269788;
  wire [11:0] add_269790;
  wire [11:0] sel_269792;
  wire [10:0] add_269794;
  wire [11:0] sel_269796;
  wire [10:0] add_269798;
  wire [11:0] sel_269800;
  wire [11:0] add_269802;
  wire [11:0] sel_269804;
  wire [11:0] add_269806;
  wire [11:0] sel_269808;
  wire [12:0] concat_269811;
  wire [9:0] add_269818;
  wire [11:0] sel_269820;
  wire [9:0] add_269822;
  wire [11:0] sel_269824;
  wire [11:0] add_269834;
  wire [11:0] sel_269836;
  wire [11:0] add_269838;
  wire [11:0] sel_269840;
  wire [11:0] add_269850;
  wire [11:0] sel_269852;
  wire [11:0] add_269854;
  wire [11:0] sel_269856;
  wire [12:0] add_269876;
  wire [11:0] add_269886;
  wire [11:0] sel_269888;
  wire [11:0] add_269890;
  wire [11:0] sel_269892;
  wire [11:0] add_269904;
  wire [11:0] sel_269906;
  wire [11:0] add_269908;
  wire [11:0] sel_269910;
  wire [10:0] add_269922;
  wire [11:0] sel_269924;
  wire [10:0] add_269926;
  wire [11:0] sel_269928;
  wire [11:0] add_269944;
  wire [11:0] sel_269946;
  wire [11:0] add_269948;
  wire [11:0] sel_269950;
  wire [9:0] add_269962;
  wire [11:0] sel_269964;
  wire [9:0] add_269966;
  wire [11:0] sel_269968;
  wire [10:0] add_269978;
  wire [11:0] sel_269980;
  wire [10:0] add_269982;
  wire [11:0] sel_269984;
  wire [11:0] add_269994;
  wire [11:0] sel_269996;
  wire [11:0] add_269998;
  wire [11:0] sel_270000;
  wire [10:0] add_270002;
  wire [11:0] sel_270004;
  wire [10:0] add_270006;
  wire [11:0] sel_270008;
  wire [13:0] concat_270011;
  wire [9:0] add_270018;
  wire [11:0] sel_270020;
  wire [9:0] add_270022;
  wire [11:0] sel_270024;
  wire [11:0] add_270034;
  wire [11:0] sel_270036;
  wire [11:0] add_270038;
  wire [11:0] sel_270040;
  wire [11:0] add_270050;
  wire [11:0] sel_270052;
  wire [11:0] add_270054;
  wire [11:0] sel_270056;
  wire [13:0] add_270072;
  wire [11:0] add_270082;
  wire [11:0] sel_270084;
  wire [11:0] add_270086;
  wire [11:0] sel_270088;
  wire [11:0] add_270100;
  wire [11:0] sel_270102;
  wire [11:0] add_270104;
  wire [11:0] sel_270106;
  wire [10:0] add_270118;
  wire [11:0] sel_270120;
  wire [10:0] add_270122;
  wire [11:0] sel_270124;
  wire [11:0] add_270136;
  wire [11:0] sel_270138;
  wire [11:0] add_270140;
  wire [11:0] sel_270142;
  wire [9:0] add_270154;
  wire [11:0] sel_270156;
  wire [9:0] add_270158;
  wire [11:0] sel_270160;
  wire [10:0] add_270170;
  wire [11:0] sel_270172;
  wire [10:0] add_270174;
  wire [11:0] sel_270176;
  wire [11:0] add_270186;
  wire [11:0] sel_270188;
  wire [11:0] add_270190;
  wire [11:0] sel_270192;
  wire [14:0] concat_270195;
  wire [9:0] add_270202;
  wire [11:0] sel_270204;
  wire [9:0] add_270206;
  wire [11:0] sel_270208;
  wire [11:0] add_270218;
  wire [11:0] sel_270220;
  wire [11:0] add_270222;
  wire [11:0] sel_270224;
  wire [11:0] add_270234;
  wire [11:0] sel_270236;
  wire [11:0] add_270238;
  wire [11:0] sel_270240;
  wire [14:0] add_270252;
  wire [11:0] add_270262;
  wire [11:0] sel_270264;
  wire [11:0] add_270266;
  wire [11:0] sel_270268;
  wire [11:0] add_270280;
  wire [11:0] sel_270282;
  wire [11:0] add_270284;
  wire [11:0] sel_270286;
  wire [10:0] add_270298;
  wire [11:0] sel_270300;
  wire [10:0] add_270302;
  wire [11:0] sel_270304;
  wire [11:0] add_270310;
  wire [11:0] sel_270312;
  wire [11:0] add_270314;
  wire [11:0] sel_270316;
  wire [9:0] add_270328;
  wire [11:0] sel_270330;
  wire [9:0] add_270332;
  wire [11:0] sel_270334;
  wire [10:0] add_270344;
  wire [11:0] sel_270346;
  wire [10:0] add_270348;
  wire [11:0] sel_270350;
  wire [15:0] concat_270361;
  wire [9:0] add_270368;
  wire [11:0] sel_270370;
  wire [9:0] add_270372;
  wire [11:0] sel_270374;
  wire [11:0] add_270384;
  wire [11:0] sel_270386;
  wire [11:0] add_270388;
  wire [11:0] sel_270390;
  wire [11:0] add_270400;
  wire [11:0] sel_270402;
  wire [11:0] add_270404;
  wire [11:0] sel_270406;
  wire [15:0] add_270412;
  wire [11:0] add_270422;
  wire [11:0] sel_270424;
  wire [11:0] add_270426;
  wire [11:0] sel_270428;
  wire [11:0] add_270440;
  wire [11:0] sel_270442;
  wire [11:0] add_270444;
  wire [11:0] sel_270446;
  wire [15:0] sel_270459;
  wire [11:0] add_270462;
  wire [11:0] sel_270464;
  wire [11:0] add_270466;
  wire [11:0] sel_270468;
  wire [9:0] add_270480;
  wire [11:0] sel_270482;
  wire [9:0] add_270484;
  wire [11:0] sel_270486;
  wire [10:0] add_270496;
  wire [11:0] sel_270498;
  wire [10:0] add_270500;
  wire [11:0] sel_270502;
  wire [15:0] add_270506;
  wire [9:0] add_270512;
  wire [11:0] sel_270514;
  wire [9:0] add_270516;
  wire [11:0] sel_270518;
  wire [11:0] add_270528;
  wire [11:0] sel_270530;
  wire [11:0] add_270532;
  wire [11:0] sel_270534;
  wire [15:0] sel_270545;
  wire [11:0] add_270556;
  wire [11:0] sel_270558;
  wire [11:0] add_270560;
  wire [11:0] sel_270562;
  wire [11:0] add_270574;
  wire [11:0] sel_270576;
  wire [11:0] add_270578;
  wire [11:0] sel_270580;
  wire [15:0] add_270586;
  wire [11:0] add_270588;
  wire [11:0] sel_270590;
  wire [11:0] add_270592;
  wire [11:0] sel_270594;
  wire [9:0] add_270606;
  wire [11:0] sel_270608;
  wire [9:0] add_270610;
  wire [11:0] sel_270612;
  wire [15:0] sel_270623;
  wire [9:0] add_270630;
  wire [11:0] sel_270632;
  wire [9:0] add_270634;
  wire [11:0] sel_270636;
  wire [11:0] add_270646;
  wire [11:0] sel_270648;
  wire [11:0] add_270650;
  wire [11:0] sel_270652;
  wire [15:0] add_270656;
  wire [11:0] add_270666;
  wire [11:0] sel_270668;
  wire [11:0] add_270670;
  wire [11:0] sel_270672;
  wire [15:0] sel_270685;
  wire [11:0] add_270688;
  wire [11:0] sel_270690;
  wire [11:0] add_270692;
  wire [11:0] sel_270694;
  wire [9:0] add_270706;
  wire [11:0] sel_270708;
  wire [9:0] add_270710;
  wire [11:0] sel_270712;
  wire [15:0] add_270716;
  wire [9:0] add_270722;
  wire [11:0] sel_270724;
  wire [9:0] add_270726;
  wire [11:0] sel_270728;
  wire [15:0] sel_270739;
  wire [11:0] add_270750;
  wire [11:0] sel_270752;
  wire [11:0] add_270754;
  wire [11:0] sel_270756;
  wire [15:0] add_270762;
  wire [11:0] add_270764;
  wire [11:0] sel_270766;
  wire [11:0] add_270768;
  wire [11:0] sel_270770;
  wire [15:0] sel_270783;
  wire [9:0] add_270790;
  wire [11:0] sel_270792;
  wire [9:0] add_270794;
  wire [11:0] sel_270796;
  wire [15:0] add_270800;
  wire [15:0] sel_270811;
  wire [11:0] add_270814;
  wire [11:0] sel_270816;
  wire [11:0] add_270818;
  wire [11:0] sel_270820;
  wire [15:0] add_270826;
  wire [15:0] sel_270833;
  wire [15:0] add_270838;
  wire [15:0] sel_270841;
  wire [15:0] add_270844;
  assign array_index_257761 = set1_unflattened[5'h00];
  assign array_index_257762 = set2_unflattened[5'h00];
  assign add_257769 = array_index_257761[11:0] + 12'h193;
  assign add_257772 = array_index_257762[11:0] + 12'h193;
  assign array_index_257775 = set1_unflattened[5'h01];
  assign array_index_257778 = set2_unflattened[5'h01];
  assign add_257782 = array_index_257761[11:0] + 12'hffb;
  assign add_257784 = array_index_257762[11:0] + 12'hffb;
  assign add_257799 = array_index_257775[11:0] + 12'h193;
  assign sel_257801 = $signed({1'h0, add_257769}) < $signed(13'h0fff) ? add_257769 : 12'hfff;
  assign add_257804 = array_index_257778[11:0] + 12'h193;
  assign sel_257806 = $signed({1'h0, add_257772}) < $signed(13'h0fff) ? add_257772 : 12'hfff;
  assign array_index_257817 = set1_unflattened[5'h02];
  assign array_index_257820 = set2_unflattened[5'h02];
  assign add_257824 = array_index_257761[11:2] + 10'h035;
  assign add_257827 = array_index_257762[11:2] + 10'h035;
  assign add_257830 = array_index_257775[11:0] + 12'hffb;
  assign sel_257832 = $signed({1'h0, add_257782}) < $signed(13'h0fff) ? add_257782 : 12'hfff;
  assign add_257834 = array_index_257778[11:0] + 12'hffb;
  assign sel_257836 = $signed({1'h0, add_257784}) < $signed(13'h0fff) ? add_257784 : 12'hfff;
  assign add_257853 = array_index_257817[11:0] + 12'h193;
  assign sel_257855 = $signed({1'h0, add_257799}) < $signed({1'h0, sel_257801}) ? add_257799 : sel_257801;
  assign add_257858 = array_index_257820[11:0] + 12'h193;
  assign sel_257860 = $signed({1'h0, add_257804}) < $signed({1'h0, sel_257806}) ? add_257804 : sel_257806;
  assign array_index_257877 = set1_unflattened[5'h03];
  assign array_index_257880 = set2_unflattened[5'h03];
  assign add_257884 = array_index_257761[11:2] + 10'h36b;
  assign add_257886 = array_index_257762[11:2] + 10'h36b;
  assign add_257888 = array_index_257775[11:2] + 10'h035;
  assign sel_257891 = $signed({1'h0, add_257824, array_index_257761[1:0]}) < $signed(13'h0fff) ? {add_257824, array_index_257761[1:0]} : 12'hfff;
  assign add_257893 = array_index_257778[11:2] + 10'h035;
  assign sel_257896 = $signed({1'h0, add_257827, array_index_257762[1:0]}) < $signed(13'h0fff) ? {add_257827, array_index_257762[1:0]} : 12'hfff;
  assign add_257898 = array_index_257817[11:0] + 12'hffb;
  assign sel_257900 = $signed({1'h0, add_257830}) < $signed({1'h0, sel_257832}) ? add_257830 : sel_257832;
  assign add_257902 = array_index_257820[11:0] + 12'hffb;
  assign sel_257904 = $signed({1'h0, add_257834}) < $signed({1'h0, sel_257836}) ? add_257834 : sel_257836;
  assign add_257925 = array_index_257877[11:0] + 12'h193;
  assign sel_257927 = $signed({1'h0, add_257853}) < $signed({1'h0, sel_257855}) ? add_257853 : sel_257855;
  assign add_257930 = array_index_257880[11:0] + 12'h193;
  assign sel_257932 = $signed({1'h0, add_257858}) < $signed({1'h0, sel_257860}) ? add_257858 : sel_257860;
  assign array_index_257955 = set1_unflattened[5'h04];
  assign array_index_257958 = set2_unflattened[5'h04];
  assign add_257962 = array_index_257761[11:0] + 12'h561;
  assign add_257964 = array_index_257762[11:0] + 12'h561;
  assign add_257966 = array_index_257775[11:2] + 10'h36b;
  assign sel_257968 = $signed({1'h0, add_257884, array_index_257761[1:0]}) < $signed(13'h0fff) ? {add_257884, array_index_257761[1:0]} : 12'hfff;
  assign add_257970 = array_index_257778[11:2] + 10'h36b;
  assign sel_257972 = $signed({1'h0, add_257886, array_index_257762[1:0]}) < $signed(13'h0fff) ? {add_257886, array_index_257762[1:0]} : 12'hfff;
  assign add_257974 = array_index_257817[11:2] + 10'h035;
  assign sel_257977 = $signed({1'h0, add_257888, array_index_257775[1:0]}) < $signed({1'h0, sel_257891}) ? {add_257888, array_index_257775[1:0]} : sel_257891;
  assign add_257979 = array_index_257820[11:2] + 10'h035;
  assign sel_257982 = $signed({1'h0, add_257893, array_index_257778[1:0]}) < $signed({1'h0, sel_257896}) ? {add_257893, array_index_257778[1:0]} : sel_257896;
  assign add_257984 = array_index_257877[11:0] + 12'hffb;
  assign sel_257986 = $signed({1'h0, add_257898}) < $signed({1'h0, sel_257900}) ? add_257898 : sel_257900;
  assign add_257988 = array_index_257880[11:0] + 12'hffb;
  assign sel_257990 = $signed({1'h0, add_257902}) < $signed({1'h0, sel_257904}) ? add_257902 : sel_257904;
  assign add_258015 = array_index_257955[11:0] + 12'h193;
  assign sel_258017 = $signed({1'h0, add_257925}) < $signed({1'h0, sel_257927}) ? add_257925 : sel_257927;
  assign add_258020 = array_index_257958[11:0] + 12'h193;
  assign sel_258022 = $signed({1'h0, add_257930}) < $signed({1'h0, sel_257932}) ? add_257930 : sel_257932;
  assign array_index_258049 = set1_unflattened[5'h05];
  assign array_index_258052 = set2_unflattened[5'h05];
  assign add_258056 = array_index_257761[11:0] + 12'h7b1;
  assign add_258058 = array_index_257762[11:0] + 12'h7b1;
  assign add_258060 = array_index_257775[11:0] + 12'h561;
  assign sel_258062 = $signed({1'h0, add_257962}) < $signed(13'h0fff) ? add_257962 : 12'hfff;
  assign add_258064 = array_index_257778[11:0] + 12'h561;
  assign sel_258066 = $signed({1'h0, add_257964}) < $signed(13'h0fff) ? add_257964 : 12'hfff;
  assign add_258068 = array_index_257817[11:2] + 10'h36b;
  assign sel_258070 = $signed({1'h0, add_257966, array_index_257775[1:0]}) < $signed({1'h0, sel_257968}) ? {add_257966, array_index_257775[1:0]} : sel_257968;
  assign add_258072 = array_index_257820[11:2] + 10'h36b;
  assign sel_258074 = $signed({1'h0, add_257970, array_index_257778[1:0]}) < $signed({1'h0, sel_257972}) ? {add_257970, array_index_257778[1:0]} : sel_257972;
  assign add_258076 = array_index_257877[11:2] + 10'h035;
  assign sel_258079 = $signed({1'h0, add_257974, array_index_257817[1:0]}) < $signed({1'h0, sel_257977}) ? {add_257974, array_index_257817[1:0]} : sel_257977;
  assign add_258081 = array_index_257880[11:2] + 10'h035;
  assign sel_258084 = $signed({1'h0, add_257979, array_index_257820[1:0]}) < $signed({1'h0, sel_257982}) ? {add_257979, array_index_257820[1:0]} : sel_257982;
  assign add_258086 = array_index_257955[11:0] + 12'hffb;
  assign sel_258088 = $signed({1'h0, add_257984}) < $signed({1'h0, sel_257986}) ? add_257984 : sel_257986;
  assign add_258090 = array_index_257958[11:0] + 12'hffb;
  assign sel_258092 = $signed({1'h0, add_257988}) < $signed({1'h0, sel_257990}) ? add_257988 : sel_257990;
  assign add_258121 = array_index_258049[11:0] + 12'h193;
  assign sel_258123 = $signed({1'h0, add_258015}) < $signed({1'h0, sel_258017}) ? add_258015 : sel_258017;
  assign add_258126 = array_index_258052[11:0] + 12'h193;
  assign sel_258128 = $signed({1'h0, add_258020}) < $signed({1'h0, sel_258022}) ? add_258020 : sel_258022;
  assign array_index_258159 = set1_unflattened[5'h06];
  assign array_index_258162 = set2_unflattened[5'h06];
  assign add_258166 = array_index_257761[11:0] + 12'hb01;
  assign add_258168 = array_index_257762[11:0] + 12'hb01;
  assign add_258170 = array_index_257775[11:0] + 12'h7b1;
  assign sel_258172 = $signed({1'h0, add_258056}) < $signed(13'h0fff) ? add_258056 : 12'hfff;
  assign add_258174 = array_index_257778[11:0] + 12'h7b1;
  assign sel_258176 = $signed({1'h0, add_258058}) < $signed(13'h0fff) ? add_258058 : 12'hfff;
  assign add_258178 = array_index_257817[11:0] + 12'h561;
  assign sel_258180 = $signed({1'h0, add_258060}) < $signed({1'h0, sel_258062}) ? add_258060 : sel_258062;
  assign add_258182 = array_index_257820[11:0] + 12'h561;
  assign sel_258184 = $signed({1'h0, add_258064}) < $signed({1'h0, sel_258066}) ? add_258064 : sel_258066;
  assign add_258186 = array_index_257877[11:2] + 10'h36b;
  assign sel_258188 = $signed({1'h0, add_258068, array_index_257817[1:0]}) < $signed({1'h0, sel_258070}) ? {add_258068, array_index_257817[1:0]} : sel_258070;
  assign add_258190 = array_index_257880[11:2] + 10'h36b;
  assign sel_258192 = $signed({1'h0, add_258072, array_index_257820[1:0]}) < $signed({1'h0, sel_258074}) ? {add_258072, array_index_257820[1:0]} : sel_258074;
  assign add_258194 = array_index_257955[11:2] + 10'h035;
  assign sel_258197 = $signed({1'h0, add_258076, array_index_257877[1:0]}) < $signed({1'h0, sel_258079}) ? {add_258076, array_index_257877[1:0]} : sel_258079;
  assign add_258199 = array_index_257958[11:2] + 10'h035;
  assign sel_258202 = $signed({1'h0, add_258081, array_index_257880[1:0]}) < $signed({1'h0, sel_258084}) ? {add_258081, array_index_257880[1:0]} : sel_258084;
  assign add_258204 = array_index_258049[11:0] + 12'hffb;
  assign sel_258206 = $signed({1'h0, add_258086}) < $signed({1'h0, sel_258088}) ? add_258086 : sel_258088;
  assign add_258208 = array_index_258052[11:0] + 12'hffb;
  assign sel_258210 = $signed({1'h0, add_258090}) < $signed({1'h0, sel_258092}) ? add_258090 : sel_258092;
  assign add_258243 = array_index_258159[11:0] + 12'h193;
  assign sel_258245 = $signed({1'h0, add_258121}) < $signed({1'h0, sel_258123}) ? add_258121 : sel_258123;
  assign add_258248 = array_index_258162[11:0] + 12'h193;
  assign sel_258250 = $signed({1'h0, add_258126}) < $signed({1'h0, sel_258128}) ? add_258126 : sel_258128;
  assign array_index_258285 = set1_unflattened[5'h07];
  assign array_index_258288 = set2_unflattened[5'h07];
  assign add_258292 = array_index_257761[11:0] + 12'h103;
  assign add_258294 = array_index_257762[11:0] + 12'h103;
  assign add_258296 = array_index_257775[11:0] + 12'hb01;
  assign sel_258298 = $signed({1'h0, add_258166}) < $signed(13'h0fff) ? add_258166 : 12'hfff;
  assign add_258300 = array_index_257778[11:0] + 12'hb01;
  assign sel_258302 = $signed({1'h0, add_258168}) < $signed(13'h0fff) ? add_258168 : 12'hfff;
  assign add_258304 = array_index_257817[11:0] + 12'h7b1;
  assign sel_258306 = $signed({1'h0, add_258170}) < $signed({1'h0, sel_258172}) ? add_258170 : sel_258172;
  assign add_258308 = array_index_257820[11:0] + 12'h7b1;
  assign sel_258310 = $signed({1'h0, add_258174}) < $signed({1'h0, sel_258176}) ? add_258174 : sel_258176;
  assign add_258312 = array_index_257877[11:0] + 12'h561;
  assign sel_258314 = $signed({1'h0, add_258178}) < $signed({1'h0, sel_258180}) ? add_258178 : sel_258180;
  assign add_258316 = array_index_257880[11:0] + 12'h561;
  assign sel_258318 = $signed({1'h0, add_258182}) < $signed({1'h0, sel_258184}) ? add_258182 : sel_258184;
  assign add_258320 = array_index_257955[11:2] + 10'h36b;
  assign sel_258322 = $signed({1'h0, add_258186, array_index_257877[1:0]}) < $signed({1'h0, sel_258188}) ? {add_258186, array_index_257877[1:0]} : sel_258188;
  assign add_258324 = array_index_257958[11:2] + 10'h36b;
  assign sel_258326 = $signed({1'h0, add_258190, array_index_257880[1:0]}) < $signed({1'h0, sel_258192}) ? {add_258190, array_index_257880[1:0]} : sel_258192;
  assign add_258328 = array_index_258049[11:2] + 10'h035;
  assign sel_258331 = $signed({1'h0, add_258194, array_index_257955[1:0]}) < $signed({1'h0, sel_258197}) ? {add_258194, array_index_257955[1:0]} : sel_258197;
  assign add_258333 = array_index_258052[11:2] + 10'h035;
  assign sel_258336 = $signed({1'h0, add_258199, array_index_257958[1:0]}) < $signed({1'h0, sel_258202}) ? {add_258199, array_index_257958[1:0]} : sel_258202;
  assign add_258338 = array_index_258159[11:0] + 12'hffb;
  assign sel_258340 = $signed({1'h0, add_258204}) < $signed({1'h0, sel_258206}) ? add_258204 : sel_258206;
  assign add_258342 = array_index_258162[11:0] + 12'hffb;
  assign sel_258344 = $signed({1'h0, add_258208}) < $signed({1'h0, sel_258210}) ? add_258208 : sel_258210;
  assign add_258381 = array_index_258285[11:0] + 12'h193;
  assign sel_258383 = $signed({1'h0, add_258243}) < $signed({1'h0, sel_258245}) ? add_258243 : sel_258245;
  assign add_258386 = array_index_258288[11:0] + 12'h193;
  assign sel_258388 = $signed({1'h0, add_258248}) < $signed({1'h0, sel_258250}) ? add_258248 : sel_258250;
  assign array_index_258427 = set1_unflattened[5'h08];
  assign array_index_258430 = set2_unflattened[5'h08];
  assign add_258434 = array_index_257761[11:0] + 12'hb55;
  assign add_258436 = array_index_257762[11:0] + 12'hb55;
  assign add_258438 = array_index_257775[11:0] + 12'h103;
  assign sel_258440 = $signed({1'h0, add_258292}) < $signed(13'h0fff) ? add_258292 : 12'hfff;
  assign add_258442 = array_index_257778[11:0] + 12'h103;
  assign sel_258444 = $signed({1'h0, add_258294}) < $signed(13'h0fff) ? add_258294 : 12'hfff;
  assign add_258446 = array_index_257817[11:0] + 12'hb01;
  assign sel_258448 = $signed({1'h0, add_258296}) < $signed({1'h0, sel_258298}) ? add_258296 : sel_258298;
  assign add_258450 = array_index_257820[11:0] + 12'hb01;
  assign sel_258452 = $signed({1'h0, add_258300}) < $signed({1'h0, sel_258302}) ? add_258300 : sel_258302;
  assign add_258454 = array_index_257877[11:0] + 12'h7b1;
  assign sel_258456 = $signed({1'h0, add_258304}) < $signed({1'h0, sel_258306}) ? add_258304 : sel_258306;
  assign add_258458 = array_index_257880[11:0] + 12'h7b1;
  assign sel_258460 = $signed({1'h0, add_258308}) < $signed({1'h0, sel_258310}) ? add_258308 : sel_258310;
  assign add_258462 = array_index_257955[11:0] + 12'h561;
  assign sel_258464 = $signed({1'h0, add_258312}) < $signed({1'h0, sel_258314}) ? add_258312 : sel_258314;
  assign add_258466 = array_index_257958[11:0] + 12'h561;
  assign sel_258468 = $signed({1'h0, add_258316}) < $signed({1'h0, sel_258318}) ? add_258316 : sel_258318;
  assign add_258470 = array_index_258049[11:2] + 10'h36b;
  assign sel_258472 = $signed({1'h0, add_258320, array_index_257955[1:0]}) < $signed({1'h0, sel_258322}) ? {add_258320, array_index_257955[1:0]} : sel_258322;
  assign add_258474 = array_index_258052[11:2] + 10'h36b;
  assign sel_258476 = $signed({1'h0, add_258324, array_index_257958[1:0]}) < $signed({1'h0, sel_258326}) ? {add_258324, array_index_257958[1:0]} : sel_258326;
  assign add_258478 = array_index_258159[11:2] + 10'h035;
  assign sel_258481 = $signed({1'h0, add_258328, array_index_258049[1:0]}) < $signed({1'h0, sel_258331}) ? {add_258328, array_index_258049[1:0]} : sel_258331;
  assign add_258483 = array_index_258162[11:2] + 10'h035;
  assign sel_258486 = $signed({1'h0, add_258333, array_index_258052[1:0]}) < $signed({1'h0, sel_258336}) ? {add_258333, array_index_258052[1:0]} : sel_258336;
  assign add_258488 = array_index_258285[11:0] + 12'hffb;
  assign sel_258490 = $signed({1'h0, add_258338}) < $signed({1'h0, sel_258340}) ? add_258338 : sel_258340;
  assign add_258492 = array_index_258288[11:0] + 12'hffb;
  assign sel_258494 = $signed({1'h0, add_258342}) < $signed({1'h0, sel_258344}) ? add_258342 : sel_258344;
  assign add_258535 = array_index_258427[11:0] + 12'h193;
  assign sel_258537 = $signed({1'h0, add_258381}) < $signed({1'h0, sel_258383}) ? add_258381 : sel_258383;
  assign add_258540 = array_index_258430[11:0] + 12'h193;
  assign sel_258542 = $signed({1'h0, add_258386}) < $signed({1'h0, sel_258388}) ? add_258386 : sel_258388;
  assign array_index_258585 = set1_unflattened[5'h09];
  assign array_index_258588 = set2_unflattened[5'h09];
  assign add_258592 = array_index_257761[11:0] + 12'h30f;
  assign add_258594 = array_index_257762[11:0] + 12'h30f;
  assign add_258596 = array_index_257775[11:0] + 12'hb55;
  assign sel_258598 = $signed({1'h0, add_258434}) < $signed(13'h0fff) ? add_258434 : 12'hfff;
  assign add_258600 = array_index_257778[11:0] + 12'hb55;
  assign sel_258602 = $signed({1'h0, add_258436}) < $signed(13'h0fff) ? add_258436 : 12'hfff;
  assign add_258604 = array_index_257817[11:0] + 12'h103;
  assign sel_258606 = $signed({1'h0, add_258438}) < $signed({1'h0, sel_258440}) ? add_258438 : sel_258440;
  assign add_258608 = array_index_257820[11:0] + 12'h103;
  assign sel_258610 = $signed({1'h0, add_258442}) < $signed({1'h0, sel_258444}) ? add_258442 : sel_258444;
  assign add_258612 = array_index_257877[11:0] + 12'hb01;
  assign sel_258614 = $signed({1'h0, add_258446}) < $signed({1'h0, sel_258448}) ? add_258446 : sel_258448;
  assign add_258616 = array_index_257880[11:0] + 12'hb01;
  assign sel_258618 = $signed({1'h0, add_258450}) < $signed({1'h0, sel_258452}) ? add_258450 : sel_258452;
  assign add_258620 = array_index_257955[11:0] + 12'h7b1;
  assign sel_258622 = $signed({1'h0, add_258454}) < $signed({1'h0, sel_258456}) ? add_258454 : sel_258456;
  assign add_258624 = array_index_257958[11:0] + 12'h7b1;
  assign sel_258626 = $signed({1'h0, add_258458}) < $signed({1'h0, sel_258460}) ? add_258458 : sel_258460;
  assign add_258628 = array_index_258049[11:0] + 12'h561;
  assign sel_258630 = $signed({1'h0, add_258462}) < $signed({1'h0, sel_258464}) ? add_258462 : sel_258464;
  assign add_258632 = array_index_258052[11:0] + 12'h561;
  assign sel_258634 = $signed({1'h0, add_258466}) < $signed({1'h0, sel_258468}) ? add_258466 : sel_258468;
  assign add_258636 = array_index_258159[11:2] + 10'h36b;
  assign sel_258638 = $signed({1'h0, add_258470, array_index_258049[1:0]}) < $signed({1'h0, sel_258472}) ? {add_258470, array_index_258049[1:0]} : sel_258472;
  assign add_258640 = array_index_258162[11:2] + 10'h36b;
  assign sel_258642 = $signed({1'h0, add_258474, array_index_258052[1:0]}) < $signed({1'h0, sel_258476}) ? {add_258474, array_index_258052[1:0]} : sel_258476;
  assign add_258644 = array_index_258285[11:2] + 10'h035;
  assign sel_258647 = $signed({1'h0, add_258478, array_index_258159[1:0]}) < $signed({1'h0, sel_258481}) ? {add_258478, array_index_258159[1:0]} : sel_258481;
  assign add_258649 = array_index_258288[11:2] + 10'h035;
  assign sel_258652 = $signed({1'h0, add_258483, array_index_258162[1:0]}) < $signed({1'h0, sel_258486}) ? {add_258483, array_index_258162[1:0]} : sel_258486;
  assign add_258654 = array_index_258427[11:0] + 12'hffb;
  assign sel_258656 = $signed({1'h0, add_258488}) < $signed({1'h0, sel_258490}) ? add_258488 : sel_258490;
  assign add_258658 = array_index_258430[11:0] + 12'hffb;
  assign sel_258660 = $signed({1'h0, add_258492}) < $signed({1'h0, sel_258494}) ? add_258492 : sel_258494;
  assign add_258705 = array_index_258585[11:0] + 12'h193;
  assign sel_258707 = $signed({1'h0, add_258535}) < $signed({1'h0, sel_258537}) ? add_258535 : sel_258537;
  assign add_258710 = array_index_258588[11:0] + 12'h193;
  assign sel_258712 = $signed({1'h0, add_258540}) < $signed({1'h0, sel_258542}) ? add_258540 : sel_258542;
  assign array_index_258761 = set1_unflattened[5'h0a];
  assign array_index_258764 = set2_unflattened[5'h0a];
  assign add_258768 = array_index_257761[11:1] + 11'h345;
  assign add_258771 = array_index_257762[11:1] + 11'h345;
  assign add_258774 = array_index_257775[11:0] + 12'h30f;
  assign sel_258776 = $signed({1'h0, add_258592}) < $signed(13'h0fff) ? add_258592 : 12'hfff;
  assign add_258778 = array_index_257778[11:0] + 12'h30f;
  assign sel_258780 = $signed({1'h0, add_258594}) < $signed(13'h0fff) ? add_258594 : 12'hfff;
  assign add_258782 = array_index_257817[11:0] + 12'hb55;
  assign sel_258784 = $signed({1'h0, add_258596}) < $signed({1'h0, sel_258598}) ? add_258596 : sel_258598;
  assign add_258786 = array_index_257820[11:0] + 12'hb55;
  assign sel_258788 = $signed({1'h0, add_258600}) < $signed({1'h0, sel_258602}) ? add_258600 : sel_258602;
  assign add_258790 = array_index_257877[11:0] + 12'h103;
  assign sel_258792 = $signed({1'h0, add_258604}) < $signed({1'h0, sel_258606}) ? add_258604 : sel_258606;
  assign add_258794 = array_index_257880[11:0] + 12'h103;
  assign sel_258796 = $signed({1'h0, add_258608}) < $signed({1'h0, sel_258610}) ? add_258608 : sel_258610;
  assign add_258798 = array_index_257955[11:0] + 12'hb01;
  assign sel_258800 = $signed({1'h0, add_258612}) < $signed({1'h0, sel_258614}) ? add_258612 : sel_258614;
  assign add_258802 = array_index_257958[11:0] + 12'hb01;
  assign sel_258804 = $signed({1'h0, add_258616}) < $signed({1'h0, sel_258618}) ? add_258616 : sel_258618;
  assign add_258806 = array_index_258049[11:0] + 12'h7b1;
  assign sel_258808 = $signed({1'h0, add_258620}) < $signed({1'h0, sel_258622}) ? add_258620 : sel_258622;
  assign add_258810 = array_index_258052[11:0] + 12'h7b1;
  assign sel_258812 = $signed({1'h0, add_258624}) < $signed({1'h0, sel_258626}) ? add_258624 : sel_258626;
  assign add_258814 = array_index_258159[11:0] + 12'h561;
  assign sel_258816 = $signed({1'h0, add_258628}) < $signed({1'h0, sel_258630}) ? add_258628 : sel_258630;
  assign add_258818 = array_index_258162[11:0] + 12'h561;
  assign sel_258820 = $signed({1'h0, add_258632}) < $signed({1'h0, sel_258634}) ? add_258632 : sel_258634;
  assign add_258822 = array_index_258285[11:2] + 10'h36b;
  assign sel_258824 = $signed({1'h0, add_258636, array_index_258159[1:0]}) < $signed({1'h0, sel_258638}) ? {add_258636, array_index_258159[1:0]} : sel_258638;
  assign add_258826 = array_index_258288[11:2] + 10'h36b;
  assign sel_258828 = $signed({1'h0, add_258640, array_index_258162[1:0]}) < $signed({1'h0, sel_258642}) ? {add_258640, array_index_258162[1:0]} : sel_258642;
  assign add_258830 = array_index_258427[11:2] + 10'h035;
  assign sel_258833 = $signed({1'h0, add_258644, array_index_258285[1:0]}) < $signed({1'h0, sel_258647}) ? {add_258644, array_index_258285[1:0]} : sel_258647;
  assign add_258835 = array_index_258430[11:2] + 10'h035;
  assign sel_258838 = $signed({1'h0, add_258649, array_index_258288[1:0]}) < $signed({1'h0, sel_258652}) ? {add_258649, array_index_258288[1:0]} : sel_258652;
  assign add_258840 = array_index_258585[11:0] + 12'hffb;
  assign sel_258842 = $signed({1'h0, add_258654}) < $signed({1'h0, sel_258656}) ? add_258654 : sel_258656;
  assign add_258844 = array_index_258588[11:0] + 12'hffb;
  assign sel_258846 = $signed({1'h0, add_258658}) < $signed({1'h0, sel_258660}) ? add_258658 : sel_258660;
  assign add_258895 = array_index_258761[11:0] + 12'h193;
  assign sel_258897 = $signed({1'h0, add_258705}) < $signed({1'h0, sel_258707}) ? add_258705 : sel_258707;
  assign add_258900 = array_index_258764[11:0] + 12'h193;
  assign sel_258902 = $signed({1'h0, add_258710}) < $signed({1'h0, sel_258712}) ? add_258710 : sel_258712;
  assign array_index_258957 = set1_unflattened[5'h0b];
  assign array_index_258960 = set2_unflattened[5'h0b];
  assign add_258964 = array_index_257761[11:1] + 11'h499;
  assign add_258966 = array_index_257762[11:1] + 11'h499;
  assign add_258968 = array_index_257775[11:1] + 11'h345;
  assign sel_258971 = $signed({1'h0, add_258768, array_index_257761[0]}) < $signed(13'h0fff) ? {add_258768, array_index_257761[0]} : 12'hfff;
  assign add_258973 = array_index_257778[11:1] + 11'h345;
  assign sel_258976 = $signed({1'h0, add_258771, array_index_257762[0]}) < $signed(13'h0fff) ? {add_258771, array_index_257762[0]} : 12'hfff;
  assign add_258978 = array_index_257817[11:0] + 12'h30f;
  assign sel_258980 = $signed({1'h0, add_258774}) < $signed({1'h0, sel_258776}) ? add_258774 : sel_258776;
  assign add_258982 = array_index_257820[11:0] + 12'h30f;
  assign sel_258984 = $signed({1'h0, add_258778}) < $signed({1'h0, sel_258780}) ? add_258778 : sel_258780;
  assign add_258986 = array_index_257877[11:0] + 12'hb55;
  assign sel_258988 = $signed({1'h0, add_258782}) < $signed({1'h0, sel_258784}) ? add_258782 : sel_258784;
  assign add_258990 = array_index_257880[11:0] + 12'hb55;
  assign sel_258992 = $signed({1'h0, add_258786}) < $signed({1'h0, sel_258788}) ? add_258786 : sel_258788;
  assign add_258994 = array_index_257955[11:0] + 12'h103;
  assign sel_258996 = $signed({1'h0, add_258790}) < $signed({1'h0, sel_258792}) ? add_258790 : sel_258792;
  assign add_258998 = array_index_257958[11:0] + 12'h103;
  assign sel_259000 = $signed({1'h0, add_258794}) < $signed({1'h0, sel_258796}) ? add_258794 : sel_258796;
  assign add_259002 = array_index_258049[11:0] + 12'hb01;
  assign sel_259004 = $signed({1'h0, add_258798}) < $signed({1'h0, sel_258800}) ? add_258798 : sel_258800;
  assign add_259006 = array_index_258052[11:0] + 12'hb01;
  assign sel_259008 = $signed({1'h0, add_258802}) < $signed({1'h0, sel_258804}) ? add_258802 : sel_258804;
  assign add_259010 = array_index_258159[11:0] + 12'h7b1;
  assign sel_259012 = $signed({1'h0, add_258806}) < $signed({1'h0, sel_258808}) ? add_258806 : sel_258808;
  assign add_259014 = array_index_258162[11:0] + 12'h7b1;
  assign sel_259016 = $signed({1'h0, add_258810}) < $signed({1'h0, sel_258812}) ? add_258810 : sel_258812;
  assign add_259018 = array_index_258285[11:0] + 12'h561;
  assign sel_259020 = $signed({1'h0, add_258814}) < $signed({1'h0, sel_258816}) ? add_258814 : sel_258816;
  assign add_259022 = array_index_258288[11:0] + 12'h561;
  assign sel_259024 = $signed({1'h0, add_258818}) < $signed({1'h0, sel_258820}) ? add_258818 : sel_258820;
  assign add_259026 = array_index_258427[11:2] + 10'h36b;
  assign sel_259028 = $signed({1'h0, add_258822, array_index_258285[1:0]}) < $signed({1'h0, sel_258824}) ? {add_258822, array_index_258285[1:0]} : sel_258824;
  assign add_259030 = array_index_258430[11:2] + 10'h36b;
  assign sel_259032 = $signed({1'h0, add_258826, array_index_258288[1:0]}) < $signed({1'h0, sel_258828}) ? {add_258826, array_index_258288[1:0]} : sel_258828;
  assign add_259034 = array_index_258585[11:2] + 10'h035;
  assign sel_259037 = $signed({1'h0, add_258830, array_index_258427[1:0]}) < $signed({1'h0, sel_258833}) ? {add_258830, array_index_258427[1:0]} : sel_258833;
  assign add_259039 = array_index_258588[11:2] + 10'h035;
  assign sel_259042 = $signed({1'h0, add_258835, array_index_258430[1:0]}) < $signed({1'h0, sel_258838}) ? {add_258835, array_index_258430[1:0]} : sel_258838;
  assign add_259044 = array_index_258761[11:0] + 12'hffb;
  assign sel_259046 = $signed({1'h0, add_258840}) < $signed({1'h0, sel_258842}) ? add_258840 : sel_258842;
  assign add_259048 = array_index_258764[11:0] + 12'hffb;
  assign sel_259050 = $signed({1'h0, add_258844}) < $signed({1'h0, sel_258846}) ? add_258844 : sel_258846;
  assign add_259103 = array_index_258957[11:0] + 12'h193;
  assign sel_259105 = $signed({1'h0, add_258895}) < $signed({1'h0, sel_258897}) ? add_258895 : sel_258897;
  assign add_259108 = array_index_258960[11:0] + 12'h193;
  assign sel_259110 = $signed({1'h0, add_258900}) < $signed({1'h0, sel_258902}) ? add_258900 : sel_258902;
  assign array_index_259171 = set1_unflattened[5'h0c];
  assign array_index_259174 = set2_unflattened[5'h0c];
  assign add_259178 = array_index_257761[11:0] + 12'ha6f;
  assign add_259180 = array_index_257762[11:0] + 12'ha6f;
  assign add_259182 = array_index_257775[11:1] + 11'h499;
  assign sel_259184 = $signed({1'h0, add_258964, array_index_257761[0]}) < $signed(13'h0fff) ? {add_258964, array_index_257761[0]} : 12'hfff;
  assign add_259186 = array_index_257778[11:1] + 11'h499;
  assign sel_259188 = $signed({1'h0, add_258966, array_index_257762[0]}) < $signed(13'h0fff) ? {add_258966, array_index_257762[0]} : 12'hfff;
  assign add_259190 = array_index_257817[11:1] + 11'h345;
  assign sel_259193 = $signed({1'h0, add_258968, array_index_257775[0]}) < $signed({1'h0, sel_258971}) ? {add_258968, array_index_257775[0]} : sel_258971;
  assign add_259195 = array_index_257820[11:1] + 11'h345;
  assign sel_259198 = $signed({1'h0, add_258973, array_index_257778[0]}) < $signed({1'h0, sel_258976}) ? {add_258973, array_index_257778[0]} : sel_258976;
  assign add_259200 = array_index_257877[11:0] + 12'h30f;
  assign sel_259202 = $signed({1'h0, add_258978}) < $signed({1'h0, sel_258980}) ? add_258978 : sel_258980;
  assign add_259204 = array_index_257880[11:0] + 12'h30f;
  assign sel_259206 = $signed({1'h0, add_258982}) < $signed({1'h0, sel_258984}) ? add_258982 : sel_258984;
  assign add_259208 = array_index_257955[11:0] + 12'hb55;
  assign sel_259210 = $signed({1'h0, add_258986}) < $signed({1'h0, sel_258988}) ? add_258986 : sel_258988;
  assign add_259212 = array_index_257958[11:0] + 12'hb55;
  assign sel_259214 = $signed({1'h0, add_258990}) < $signed({1'h0, sel_258992}) ? add_258990 : sel_258992;
  assign add_259216 = array_index_258049[11:0] + 12'h103;
  assign sel_259218 = $signed({1'h0, add_258994}) < $signed({1'h0, sel_258996}) ? add_258994 : sel_258996;
  assign add_259220 = array_index_258052[11:0] + 12'h103;
  assign sel_259222 = $signed({1'h0, add_258998}) < $signed({1'h0, sel_259000}) ? add_258998 : sel_259000;
  assign add_259224 = array_index_258159[11:0] + 12'hb01;
  assign sel_259226 = $signed({1'h0, add_259002}) < $signed({1'h0, sel_259004}) ? add_259002 : sel_259004;
  assign add_259228 = array_index_258162[11:0] + 12'hb01;
  assign sel_259230 = $signed({1'h0, add_259006}) < $signed({1'h0, sel_259008}) ? add_259006 : sel_259008;
  assign add_259232 = array_index_258285[11:0] + 12'h7b1;
  assign sel_259234 = $signed({1'h0, add_259010}) < $signed({1'h0, sel_259012}) ? add_259010 : sel_259012;
  assign add_259236 = array_index_258288[11:0] + 12'h7b1;
  assign sel_259238 = $signed({1'h0, add_259014}) < $signed({1'h0, sel_259016}) ? add_259014 : sel_259016;
  assign add_259240 = array_index_258427[11:0] + 12'h561;
  assign sel_259242 = $signed({1'h0, add_259018}) < $signed({1'h0, sel_259020}) ? add_259018 : sel_259020;
  assign add_259244 = array_index_258430[11:0] + 12'h561;
  assign sel_259246 = $signed({1'h0, add_259022}) < $signed({1'h0, sel_259024}) ? add_259022 : sel_259024;
  assign add_259248 = array_index_258585[11:2] + 10'h36b;
  assign sel_259250 = $signed({1'h0, add_259026, array_index_258427[1:0]}) < $signed({1'h0, sel_259028}) ? {add_259026, array_index_258427[1:0]} : sel_259028;
  assign add_259252 = array_index_258588[11:2] + 10'h36b;
  assign sel_259254 = $signed({1'h0, add_259030, array_index_258430[1:0]}) < $signed({1'h0, sel_259032}) ? {add_259030, array_index_258430[1:0]} : sel_259032;
  assign add_259256 = array_index_258761[11:2] + 10'h035;
  assign sel_259259 = $signed({1'h0, add_259034, array_index_258585[1:0]}) < $signed({1'h0, sel_259037}) ? {add_259034, array_index_258585[1:0]} : sel_259037;
  assign add_259261 = array_index_258764[11:2] + 10'h035;
  assign sel_259264 = $signed({1'h0, add_259039, array_index_258588[1:0]}) < $signed({1'h0, sel_259042}) ? {add_259039, array_index_258588[1:0]} : sel_259042;
  assign add_259266 = array_index_258957[11:0] + 12'hffb;
  assign sel_259268 = $signed({1'h0, add_259044}) < $signed({1'h0, sel_259046}) ? add_259044 : sel_259046;
  assign add_259270 = array_index_258960[11:0] + 12'hffb;
  assign sel_259272 = $signed({1'h0, add_259048}) < $signed({1'h0, sel_259050}) ? add_259048 : sel_259050;
  assign add_259329 = array_index_259171[11:0] + 12'h193;
  assign sel_259331 = $signed({1'h0, add_259103}) < $signed({1'h0, sel_259105}) ? add_259103 : sel_259105;
  assign add_259334 = array_index_259174[11:0] + 12'h193;
  assign sel_259336 = $signed({1'h0, add_259108}) < $signed({1'h0, sel_259110}) ? add_259108 : sel_259110;
  assign array_index_259401 = set1_unflattened[5'h0d];
  assign array_index_259404 = set2_unflattened[5'h0d];
  assign add_259408 = array_index_257761[11:0] + 12'h59d;
  assign add_259410 = array_index_257762[11:0] + 12'h59d;
  assign add_259412 = array_index_257775[11:0] + 12'ha6f;
  assign sel_259414 = $signed({1'h0, add_259178}) < $signed(13'h0fff) ? add_259178 : 12'hfff;
  assign add_259416 = array_index_257778[11:0] + 12'ha6f;
  assign sel_259418 = $signed({1'h0, add_259180}) < $signed(13'h0fff) ? add_259180 : 12'hfff;
  assign add_259420 = array_index_257817[11:1] + 11'h499;
  assign sel_259422 = $signed({1'h0, add_259182, array_index_257775[0]}) < $signed({1'h0, sel_259184}) ? {add_259182, array_index_257775[0]} : sel_259184;
  assign add_259424 = array_index_257820[11:1] + 11'h499;
  assign sel_259426 = $signed({1'h0, add_259186, array_index_257778[0]}) < $signed({1'h0, sel_259188}) ? {add_259186, array_index_257778[0]} : sel_259188;
  assign add_259428 = array_index_257877[11:1] + 11'h345;
  assign sel_259431 = $signed({1'h0, add_259190, array_index_257817[0]}) < $signed({1'h0, sel_259193}) ? {add_259190, array_index_257817[0]} : sel_259193;
  assign add_259433 = array_index_257880[11:1] + 11'h345;
  assign sel_259436 = $signed({1'h0, add_259195, array_index_257820[0]}) < $signed({1'h0, sel_259198}) ? {add_259195, array_index_257820[0]} : sel_259198;
  assign add_259438 = array_index_257955[11:0] + 12'h30f;
  assign sel_259440 = $signed({1'h0, add_259200}) < $signed({1'h0, sel_259202}) ? add_259200 : sel_259202;
  assign add_259442 = array_index_257958[11:0] + 12'h30f;
  assign sel_259444 = $signed({1'h0, add_259204}) < $signed({1'h0, sel_259206}) ? add_259204 : sel_259206;
  assign add_259446 = array_index_258049[11:0] + 12'hb55;
  assign sel_259448 = $signed({1'h0, add_259208}) < $signed({1'h0, sel_259210}) ? add_259208 : sel_259210;
  assign add_259450 = array_index_258052[11:0] + 12'hb55;
  assign sel_259452 = $signed({1'h0, add_259212}) < $signed({1'h0, sel_259214}) ? add_259212 : sel_259214;
  assign add_259454 = array_index_258159[11:0] + 12'h103;
  assign sel_259456 = $signed({1'h0, add_259216}) < $signed({1'h0, sel_259218}) ? add_259216 : sel_259218;
  assign add_259458 = array_index_258162[11:0] + 12'h103;
  assign sel_259460 = $signed({1'h0, add_259220}) < $signed({1'h0, sel_259222}) ? add_259220 : sel_259222;
  assign add_259462 = array_index_258285[11:0] + 12'hb01;
  assign sel_259464 = $signed({1'h0, add_259224}) < $signed({1'h0, sel_259226}) ? add_259224 : sel_259226;
  assign add_259466 = array_index_258288[11:0] + 12'hb01;
  assign sel_259468 = $signed({1'h0, add_259228}) < $signed({1'h0, sel_259230}) ? add_259228 : sel_259230;
  assign add_259470 = array_index_258427[11:0] + 12'h7b1;
  assign sel_259472 = $signed({1'h0, add_259232}) < $signed({1'h0, sel_259234}) ? add_259232 : sel_259234;
  assign add_259474 = array_index_258430[11:0] + 12'h7b1;
  assign sel_259476 = $signed({1'h0, add_259236}) < $signed({1'h0, sel_259238}) ? add_259236 : sel_259238;
  assign add_259478 = array_index_258585[11:0] + 12'h561;
  assign sel_259480 = $signed({1'h0, add_259240}) < $signed({1'h0, sel_259242}) ? add_259240 : sel_259242;
  assign add_259482 = array_index_258588[11:0] + 12'h561;
  assign sel_259484 = $signed({1'h0, add_259244}) < $signed({1'h0, sel_259246}) ? add_259244 : sel_259246;
  assign add_259486 = array_index_258761[11:2] + 10'h36b;
  assign sel_259488 = $signed({1'h0, add_259248, array_index_258585[1:0]}) < $signed({1'h0, sel_259250}) ? {add_259248, array_index_258585[1:0]} : sel_259250;
  assign add_259490 = array_index_258764[11:2] + 10'h36b;
  assign sel_259492 = $signed({1'h0, add_259252, array_index_258588[1:0]}) < $signed({1'h0, sel_259254}) ? {add_259252, array_index_258588[1:0]} : sel_259254;
  assign add_259494 = array_index_258957[11:2] + 10'h035;
  assign sel_259497 = $signed({1'h0, add_259256, array_index_258761[1:0]}) < $signed({1'h0, sel_259259}) ? {add_259256, array_index_258761[1:0]} : sel_259259;
  assign add_259499 = array_index_258960[11:2] + 10'h035;
  assign sel_259502 = $signed({1'h0, add_259261, array_index_258764[1:0]}) < $signed({1'h0, sel_259264}) ? {add_259261, array_index_258764[1:0]} : sel_259264;
  assign add_259504 = array_index_259171[11:0] + 12'hffb;
  assign sel_259506 = $signed({1'h0, add_259266}) < $signed({1'h0, sel_259268}) ? add_259266 : sel_259268;
  assign add_259508 = array_index_259174[11:0] + 12'hffb;
  assign sel_259510 = $signed({1'h0, add_259270}) < $signed({1'h0, sel_259272}) ? add_259270 : sel_259272;
  assign add_259571 = array_index_259401[11:0] + 12'h193;
  assign sel_259573 = $signed({1'h0, add_259329}) < $signed({1'h0, sel_259331}) ? add_259329 : sel_259331;
  assign add_259576 = array_index_259404[11:0] + 12'h193;
  assign sel_259578 = $signed({1'h0, add_259334}) < $signed({1'h0, sel_259336}) ? add_259334 : sel_259336;
  assign array_index_259647 = set1_unflattened[5'h0e];
  assign array_index_259650 = set2_unflattened[5'h0e];
  assign add_259654 = array_index_257761[11:1] + 11'h079;
  assign add_259656 = array_index_257762[11:1] + 11'h079;
  assign add_259658 = array_index_257775[11:0] + 12'h59d;
  assign sel_259660 = $signed({1'h0, add_259408}) < $signed(13'h0fff) ? add_259408 : 12'hfff;
  assign add_259662 = array_index_257778[11:0] + 12'h59d;
  assign sel_259664 = $signed({1'h0, add_259410}) < $signed(13'h0fff) ? add_259410 : 12'hfff;
  assign add_259666 = array_index_257817[11:0] + 12'ha6f;
  assign sel_259668 = $signed({1'h0, add_259412}) < $signed({1'h0, sel_259414}) ? add_259412 : sel_259414;
  assign add_259670 = array_index_257820[11:0] + 12'ha6f;
  assign sel_259672 = $signed({1'h0, add_259416}) < $signed({1'h0, sel_259418}) ? add_259416 : sel_259418;
  assign add_259674 = array_index_257877[11:1] + 11'h499;
  assign sel_259676 = $signed({1'h0, add_259420, array_index_257817[0]}) < $signed({1'h0, sel_259422}) ? {add_259420, array_index_257817[0]} : sel_259422;
  assign add_259678 = array_index_257880[11:1] + 11'h499;
  assign sel_259680 = $signed({1'h0, add_259424, array_index_257820[0]}) < $signed({1'h0, sel_259426}) ? {add_259424, array_index_257820[0]} : sel_259426;
  assign add_259682 = array_index_257955[11:1] + 11'h345;
  assign sel_259685 = $signed({1'h0, add_259428, array_index_257877[0]}) < $signed({1'h0, sel_259431}) ? {add_259428, array_index_257877[0]} : sel_259431;
  assign add_259687 = array_index_257958[11:1] + 11'h345;
  assign sel_259690 = $signed({1'h0, add_259433, array_index_257880[0]}) < $signed({1'h0, sel_259436}) ? {add_259433, array_index_257880[0]} : sel_259436;
  assign add_259692 = array_index_258049[11:0] + 12'h30f;
  assign sel_259694 = $signed({1'h0, add_259438}) < $signed({1'h0, sel_259440}) ? add_259438 : sel_259440;
  assign add_259696 = array_index_258052[11:0] + 12'h30f;
  assign sel_259698 = $signed({1'h0, add_259442}) < $signed({1'h0, sel_259444}) ? add_259442 : sel_259444;
  assign add_259700 = array_index_258159[11:0] + 12'hb55;
  assign sel_259702 = $signed({1'h0, add_259446}) < $signed({1'h0, sel_259448}) ? add_259446 : sel_259448;
  assign add_259704 = array_index_258162[11:0] + 12'hb55;
  assign sel_259706 = $signed({1'h0, add_259450}) < $signed({1'h0, sel_259452}) ? add_259450 : sel_259452;
  assign add_259708 = array_index_258285[11:0] + 12'h103;
  assign sel_259710 = $signed({1'h0, add_259454}) < $signed({1'h0, sel_259456}) ? add_259454 : sel_259456;
  assign add_259712 = array_index_258288[11:0] + 12'h103;
  assign sel_259714 = $signed({1'h0, add_259458}) < $signed({1'h0, sel_259460}) ? add_259458 : sel_259460;
  assign add_259716 = array_index_258427[11:0] + 12'hb01;
  assign sel_259718 = $signed({1'h0, add_259462}) < $signed({1'h0, sel_259464}) ? add_259462 : sel_259464;
  assign add_259720 = array_index_258430[11:0] + 12'hb01;
  assign sel_259722 = $signed({1'h0, add_259466}) < $signed({1'h0, sel_259468}) ? add_259466 : sel_259468;
  assign add_259724 = array_index_258585[11:0] + 12'h7b1;
  assign sel_259726 = $signed({1'h0, add_259470}) < $signed({1'h0, sel_259472}) ? add_259470 : sel_259472;
  assign add_259728 = array_index_258588[11:0] + 12'h7b1;
  assign sel_259730 = $signed({1'h0, add_259474}) < $signed({1'h0, sel_259476}) ? add_259474 : sel_259476;
  assign add_259732 = array_index_258761[11:0] + 12'h561;
  assign sel_259734 = $signed({1'h0, add_259478}) < $signed({1'h0, sel_259480}) ? add_259478 : sel_259480;
  assign add_259736 = array_index_258764[11:0] + 12'h561;
  assign sel_259738 = $signed({1'h0, add_259482}) < $signed({1'h0, sel_259484}) ? add_259482 : sel_259484;
  assign add_259740 = array_index_258957[11:2] + 10'h36b;
  assign sel_259742 = $signed({1'h0, add_259486, array_index_258761[1:0]}) < $signed({1'h0, sel_259488}) ? {add_259486, array_index_258761[1:0]} : sel_259488;
  assign add_259744 = array_index_258960[11:2] + 10'h36b;
  assign sel_259746 = $signed({1'h0, add_259490, array_index_258764[1:0]}) < $signed({1'h0, sel_259492}) ? {add_259490, array_index_258764[1:0]} : sel_259492;
  assign add_259748 = array_index_259171[11:2] + 10'h035;
  assign sel_259751 = $signed({1'h0, add_259494, array_index_258957[1:0]}) < $signed({1'h0, sel_259497}) ? {add_259494, array_index_258957[1:0]} : sel_259497;
  assign add_259753 = array_index_259174[11:2] + 10'h035;
  assign sel_259756 = $signed({1'h0, add_259499, array_index_258960[1:0]}) < $signed({1'h0, sel_259502}) ? {add_259499, array_index_258960[1:0]} : sel_259502;
  assign add_259758 = array_index_259401[11:0] + 12'hffb;
  assign sel_259760 = $signed({1'h0, add_259504}) < $signed({1'h0, sel_259506}) ? add_259504 : sel_259506;
  assign add_259762 = array_index_259404[11:0] + 12'hffb;
  assign sel_259764 = $signed({1'h0, add_259508}) < $signed({1'h0, sel_259510}) ? add_259508 : sel_259510;
  assign add_259829 = array_index_259647[11:0] + 12'h193;
  assign sel_259831 = $signed({1'h0, add_259571}) < $signed({1'h0, sel_259573}) ? add_259571 : sel_259573;
  assign add_259834 = array_index_259650[11:0] + 12'h193;
  assign sel_259836 = $signed({1'h0, add_259576}) < $signed({1'h0, sel_259578}) ? add_259576 : sel_259578;
  assign array_index_259911 = set1_unflattened[5'h0f];
  assign array_index_259914 = set2_unflattened[5'h0f];
  assign add_259918 = array_index_257761[11:0] + 12'h141;
  assign add_259920 = array_index_257762[11:0] + 12'h141;
  assign add_259922 = array_index_257775[11:1] + 11'h079;
  assign sel_259924 = $signed({1'h0, add_259654, array_index_257761[0]}) < $signed(13'h0fff) ? {add_259654, array_index_257761[0]} : 12'hfff;
  assign add_259926 = array_index_257778[11:1] + 11'h079;
  assign sel_259928 = $signed({1'h0, add_259656, array_index_257762[0]}) < $signed(13'h0fff) ? {add_259656, array_index_257762[0]} : 12'hfff;
  assign add_259930 = array_index_257817[11:0] + 12'h59d;
  assign sel_259932 = $signed({1'h0, add_259658}) < $signed({1'h0, sel_259660}) ? add_259658 : sel_259660;
  assign add_259934 = array_index_257820[11:0] + 12'h59d;
  assign sel_259936 = $signed({1'h0, add_259662}) < $signed({1'h0, sel_259664}) ? add_259662 : sel_259664;
  assign add_259938 = array_index_257877[11:0] + 12'ha6f;
  assign sel_259940 = $signed({1'h0, add_259666}) < $signed({1'h0, sel_259668}) ? add_259666 : sel_259668;
  assign add_259942 = array_index_257880[11:0] + 12'ha6f;
  assign sel_259944 = $signed({1'h0, add_259670}) < $signed({1'h0, sel_259672}) ? add_259670 : sel_259672;
  assign add_259946 = array_index_257955[11:1] + 11'h499;
  assign sel_259948 = $signed({1'h0, add_259674, array_index_257877[0]}) < $signed({1'h0, sel_259676}) ? {add_259674, array_index_257877[0]} : sel_259676;
  assign add_259950 = array_index_257958[11:1] + 11'h499;
  assign sel_259952 = $signed({1'h0, add_259678, array_index_257880[0]}) < $signed({1'h0, sel_259680}) ? {add_259678, array_index_257880[0]} : sel_259680;
  assign add_259954 = array_index_258049[11:1] + 11'h345;
  assign sel_259957 = $signed({1'h0, add_259682, array_index_257955[0]}) < $signed({1'h0, sel_259685}) ? {add_259682, array_index_257955[0]} : sel_259685;
  assign add_259959 = array_index_258052[11:1] + 11'h345;
  assign sel_259962 = $signed({1'h0, add_259687, array_index_257958[0]}) < $signed({1'h0, sel_259690}) ? {add_259687, array_index_257958[0]} : sel_259690;
  assign add_259964 = array_index_258159[11:0] + 12'h30f;
  assign sel_259966 = $signed({1'h0, add_259692}) < $signed({1'h0, sel_259694}) ? add_259692 : sel_259694;
  assign add_259968 = array_index_258162[11:0] + 12'h30f;
  assign sel_259970 = $signed({1'h0, add_259696}) < $signed({1'h0, sel_259698}) ? add_259696 : sel_259698;
  assign add_259972 = array_index_258285[11:0] + 12'hb55;
  assign sel_259974 = $signed({1'h0, add_259700}) < $signed({1'h0, sel_259702}) ? add_259700 : sel_259702;
  assign add_259976 = array_index_258288[11:0] + 12'hb55;
  assign sel_259978 = $signed({1'h0, add_259704}) < $signed({1'h0, sel_259706}) ? add_259704 : sel_259706;
  assign add_259980 = array_index_258427[11:0] + 12'h103;
  assign sel_259982 = $signed({1'h0, add_259708}) < $signed({1'h0, sel_259710}) ? add_259708 : sel_259710;
  assign add_259984 = array_index_258430[11:0] + 12'h103;
  assign sel_259986 = $signed({1'h0, add_259712}) < $signed({1'h0, sel_259714}) ? add_259712 : sel_259714;
  assign add_259988 = array_index_258585[11:0] + 12'hb01;
  assign sel_259990 = $signed({1'h0, add_259716}) < $signed({1'h0, sel_259718}) ? add_259716 : sel_259718;
  assign add_259992 = array_index_258588[11:0] + 12'hb01;
  assign sel_259994 = $signed({1'h0, add_259720}) < $signed({1'h0, sel_259722}) ? add_259720 : sel_259722;
  assign add_259996 = array_index_258761[11:0] + 12'h7b1;
  assign sel_259998 = $signed({1'h0, add_259724}) < $signed({1'h0, sel_259726}) ? add_259724 : sel_259726;
  assign add_260000 = array_index_258764[11:0] + 12'h7b1;
  assign sel_260002 = $signed({1'h0, add_259728}) < $signed({1'h0, sel_259730}) ? add_259728 : sel_259730;
  assign add_260004 = array_index_258957[11:0] + 12'h561;
  assign sel_260006 = $signed({1'h0, add_259732}) < $signed({1'h0, sel_259734}) ? add_259732 : sel_259734;
  assign add_260008 = array_index_258960[11:0] + 12'h561;
  assign sel_260010 = $signed({1'h0, add_259736}) < $signed({1'h0, sel_259738}) ? add_259736 : sel_259738;
  assign add_260012 = array_index_259171[11:2] + 10'h36b;
  assign sel_260014 = $signed({1'h0, add_259740, array_index_258957[1:0]}) < $signed({1'h0, sel_259742}) ? {add_259740, array_index_258957[1:0]} : sel_259742;
  assign add_260016 = array_index_259174[11:2] + 10'h36b;
  assign sel_260018 = $signed({1'h0, add_259744, array_index_258960[1:0]}) < $signed({1'h0, sel_259746}) ? {add_259744, array_index_258960[1:0]} : sel_259746;
  assign add_260020 = array_index_259401[11:2] + 10'h035;
  assign sel_260023 = $signed({1'h0, add_259748, array_index_259171[1:0]}) < $signed({1'h0, sel_259751}) ? {add_259748, array_index_259171[1:0]} : sel_259751;
  assign add_260025 = array_index_259404[11:2] + 10'h035;
  assign sel_260028 = $signed({1'h0, add_259753, array_index_259174[1:0]}) < $signed({1'h0, sel_259756}) ? {add_259753, array_index_259174[1:0]} : sel_259756;
  assign add_260030 = array_index_259647[11:0] + 12'hffb;
  assign sel_260032 = $signed({1'h0, add_259758}) < $signed({1'h0, sel_259760}) ? add_259758 : sel_259760;
  assign add_260034 = array_index_259650[11:0] + 12'hffb;
  assign sel_260036 = $signed({1'h0, add_259762}) < $signed({1'h0, sel_259764}) ? add_259762 : sel_259764;
  assign add_260107 = array_index_259911[11:0] + 12'h193;
  assign sel_260109 = $signed({1'h0, add_259829}) < $signed({1'h0, sel_259831}) ? add_259829 : sel_259831;
  assign add_260112 = array_index_259914[11:0] + 12'h193;
  assign sel_260114 = $signed({1'h0, add_259834}) < $signed({1'h0, sel_259836}) ? add_259834 : sel_259836;
  assign add_260116 = array_index_257761[11:1] + 11'h7b5;
  assign add_260118 = array_index_257762[11:1] + 11'h7b5;
  assign array_index_260195 = set1_unflattened[5'h10];
  assign array_index_260198 = set2_unflattened[5'h10];
  assign add_260208 = array_index_257775[11:0] + 12'h141;
  assign sel_260210 = $signed({1'h0, add_259918}) < $signed(13'h0fff) ? add_259918 : 12'hfff;
  assign add_260212 = array_index_257778[11:0] + 12'h141;
  assign sel_260214 = $signed({1'h0, add_259920}) < $signed(13'h0fff) ? add_259920 : 12'hfff;
  assign add_260216 = array_index_257817[11:1] + 11'h079;
  assign sel_260218 = $signed({1'h0, add_259922, array_index_257775[0]}) < $signed({1'h0, sel_259924}) ? {add_259922, array_index_257775[0]} : sel_259924;
  assign add_260220 = array_index_257820[11:1] + 11'h079;
  assign sel_260222 = $signed({1'h0, add_259926, array_index_257778[0]}) < $signed({1'h0, sel_259928}) ? {add_259926, array_index_257778[0]} : sel_259928;
  assign add_260224 = array_index_257877[11:0] + 12'h59d;
  assign sel_260226 = $signed({1'h0, add_259930}) < $signed({1'h0, sel_259932}) ? add_259930 : sel_259932;
  assign add_260228 = array_index_257880[11:0] + 12'h59d;
  assign sel_260230 = $signed({1'h0, add_259934}) < $signed({1'h0, sel_259936}) ? add_259934 : sel_259936;
  assign add_260232 = array_index_257955[11:0] + 12'ha6f;
  assign sel_260234 = $signed({1'h0, add_259938}) < $signed({1'h0, sel_259940}) ? add_259938 : sel_259940;
  assign add_260236 = array_index_257958[11:0] + 12'ha6f;
  assign sel_260238 = $signed({1'h0, add_259942}) < $signed({1'h0, sel_259944}) ? add_259942 : sel_259944;
  assign add_260240 = array_index_258049[11:1] + 11'h499;
  assign sel_260242 = $signed({1'h0, add_259946, array_index_257955[0]}) < $signed({1'h0, sel_259948}) ? {add_259946, array_index_257955[0]} : sel_259948;
  assign add_260244 = array_index_258052[11:1] + 11'h499;
  assign sel_260246 = $signed({1'h0, add_259950, array_index_257958[0]}) < $signed({1'h0, sel_259952}) ? {add_259950, array_index_257958[0]} : sel_259952;
  assign add_260248 = array_index_258159[11:1] + 11'h345;
  assign sel_260251 = $signed({1'h0, add_259954, array_index_258049[0]}) < $signed({1'h0, sel_259957}) ? {add_259954, array_index_258049[0]} : sel_259957;
  assign add_260253 = array_index_258162[11:1] + 11'h345;
  assign sel_260256 = $signed({1'h0, add_259959, array_index_258052[0]}) < $signed({1'h0, sel_259962}) ? {add_259959, array_index_258052[0]} : sel_259962;
  assign add_260258 = array_index_258285[11:0] + 12'h30f;
  assign sel_260260 = $signed({1'h0, add_259964}) < $signed({1'h0, sel_259966}) ? add_259964 : sel_259966;
  assign add_260262 = array_index_258288[11:0] + 12'h30f;
  assign sel_260264 = $signed({1'h0, add_259968}) < $signed({1'h0, sel_259970}) ? add_259968 : sel_259970;
  assign add_260266 = array_index_258427[11:0] + 12'hb55;
  assign sel_260268 = $signed({1'h0, add_259972}) < $signed({1'h0, sel_259974}) ? add_259972 : sel_259974;
  assign add_260270 = array_index_258430[11:0] + 12'hb55;
  assign sel_260272 = $signed({1'h0, add_259976}) < $signed({1'h0, sel_259978}) ? add_259976 : sel_259978;
  assign add_260274 = array_index_258585[11:0] + 12'h103;
  assign sel_260276 = $signed({1'h0, add_259980}) < $signed({1'h0, sel_259982}) ? add_259980 : sel_259982;
  assign add_260278 = array_index_258588[11:0] + 12'h103;
  assign sel_260280 = $signed({1'h0, add_259984}) < $signed({1'h0, sel_259986}) ? add_259984 : sel_259986;
  assign add_260282 = array_index_258761[11:0] + 12'hb01;
  assign sel_260284 = $signed({1'h0, add_259988}) < $signed({1'h0, sel_259990}) ? add_259988 : sel_259990;
  assign add_260286 = array_index_258764[11:0] + 12'hb01;
  assign sel_260288 = $signed({1'h0, add_259992}) < $signed({1'h0, sel_259994}) ? add_259992 : sel_259994;
  assign add_260290 = array_index_258957[11:0] + 12'h7b1;
  assign sel_260292 = $signed({1'h0, add_259996}) < $signed({1'h0, sel_259998}) ? add_259996 : sel_259998;
  assign add_260294 = array_index_258960[11:0] + 12'h7b1;
  assign sel_260296 = $signed({1'h0, add_260000}) < $signed({1'h0, sel_260002}) ? add_260000 : sel_260002;
  assign add_260298 = array_index_259171[11:0] + 12'h561;
  assign sel_260300 = $signed({1'h0, add_260004}) < $signed({1'h0, sel_260006}) ? add_260004 : sel_260006;
  assign add_260302 = array_index_259174[11:0] + 12'h561;
  assign sel_260304 = $signed({1'h0, add_260008}) < $signed({1'h0, sel_260010}) ? add_260008 : sel_260010;
  assign add_260306 = array_index_259401[11:2] + 10'h36b;
  assign sel_260308 = $signed({1'h0, add_260012, array_index_259171[1:0]}) < $signed({1'h0, sel_260014}) ? {add_260012, array_index_259171[1:0]} : sel_260014;
  assign add_260310 = array_index_259404[11:2] + 10'h36b;
  assign sel_260312 = $signed({1'h0, add_260016, array_index_259174[1:0]}) < $signed({1'h0, sel_260018}) ? {add_260016, array_index_259174[1:0]} : sel_260018;
  assign add_260314 = array_index_259647[11:2] + 10'h035;
  assign sel_260317 = $signed({1'h0, add_260020, array_index_259401[1:0]}) < $signed({1'h0, sel_260023}) ? {add_260020, array_index_259401[1:0]} : sel_260023;
  assign add_260319 = array_index_259650[11:2] + 10'h035;
  assign sel_260322 = $signed({1'h0, add_260025, array_index_259404[1:0]}) < $signed({1'h0, sel_260028}) ? {add_260025, array_index_259404[1:0]} : sel_260028;
  assign add_260324 = array_index_259911[11:0] + 12'hffb;
  assign sel_260326 = $signed({1'h0, add_260030}) < $signed({1'h0, sel_260032}) ? add_260030 : sel_260032;
  assign add_260328 = array_index_259914[11:0] + 12'hffb;
  assign sel_260330 = $signed({1'h0, add_260034}) < $signed({1'h0, sel_260036}) ? add_260034 : sel_260036;
  assign add_260338 = array_index_257761[11:0] + 12'h30b;
  assign add_260340 = array_index_257762[11:0] + 12'h30b;
  assign add_260411 = array_index_260195[11:0] + 12'h193;
  assign sel_260413 = $signed({1'h0, add_260107}) < $signed({1'h0, sel_260109}) ? add_260107 : sel_260109;
  assign add_260416 = array_index_260198[11:0] + 12'h193;
  assign sel_260418 = $signed({1'h0, add_260112}) < $signed({1'h0, sel_260114}) ? add_260112 : sel_260114;
  assign add_260426 = array_index_257775[11:1] + 11'h7b5;
  assign sel_260428 = $signed({1'h0, add_260116, array_index_257761[0]}) < $signed(13'h0fff) ? {add_260116, array_index_257761[0]} : 12'hfff;
  assign add_260430 = array_index_257778[11:1] + 11'h7b5;
  assign sel_260432 = $signed({1'h0, add_260118, array_index_257762[0]}) < $signed(13'h0fff) ? {add_260118, array_index_257762[0]} : 12'hfff;
  assign array_index_260507 = set1_unflattened[5'h11];
  assign array_index_260510 = set2_unflattened[5'h11];
  assign add_260514 = array_index_257761[11:1] + 11'h1e7;
  assign add_260516 = array_index_257762[11:1] + 11'h1e7;
  assign add_260528 = array_index_257817[11:0] + 12'h141;
  assign sel_260530 = $signed({1'h0, add_260208}) < $signed({1'h0, sel_260210}) ? add_260208 : sel_260210;
  assign add_260532 = array_index_257820[11:0] + 12'h141;
  assign sel_260534 = $signed({1'h0, add_260212}) < $signed({1'h0, sel_260214}) ? add_260212 : sel_260214;
  assign add_260536 = array_index_257877[11:1] + 11'h079;
  assign sel_260538 = $signed({1'h0, add_260216, array_index_257817[0]}) < $signed({1'h0, sel_260218}) ? {add_260216, array_index_257817[0]} : sel_260218;
  assign add_260540 = array_index_257880[11:1] + 11'h079;
  assign sel_260542 = $signed({1'h0, add_260220, array_index_257820[0]}) < $signed({1'h0, sel_260222}) ? {add_260220, array_index_257820[0]} : sel_260222;
  assign add_260544 = array_index_257955[11:0] + 12'h59d;
  assign sel_260546 = $signed({1'h0, add_260224}) < $signed({1'h0, sel_260226}) ? add_260224 : sel_260226;
  assign add_260548 = array_index_257958[11:0] + 12'h59d;
  assign sel_260550 = $signed({1'h0, add_260228}) < $signed({1'h0, sel_260230}) ? add_260228 : sel_260230;
  assign add_260552 = array_index_258049[11:0] + 12'ha6f;
  assign sel_260554 = $signed({1'h0, add_260232}) < $signed({1'h0, sel_260234}) ? add_260232 : sel_260234;
  assign add_260556 = array_index_258052[11:0] + 12'ha6f;
  assign sel_260558 = $signed({1'h0, add_260236}) < $signed({1'h0, sel_260238}) ? add_260236 : sel_260238;
  assign add_260560 = array_index_258159[11:1] + 11'h499;
  assign sel_260562 = $signed({1'h0, add_260240, array_index_258049[0]}) < $signed({1'h0, sel_260242}) ? {add_260240, array_index_258049[0]} : sel_260242;
  assign add_260564 = array_index_258162[11:1] + 11'h499;
  assign sel_260566 = $signed({1'h0, add_260244, array_index_258052[0]}) < $signed({1'h0, sel_260246}) ? {add_260244, array_index_258052[0]} : sel_260246;
  assign add_260568 = array_index_258285[11:1] + 11'h345;
  assign sel_260571 = $signed({1'h0, add_260248, array_index_258159[0]}) < $signed({1'h0, sel_260251}) ? {add_260248, array_index_258159[0]} : sel_260251;
  assign add_260573 = array_index_258288[11:1] + 11'h345;
  assign sel_260576 = $signed({1'h0, add_260253, array_index_258162[0]}) < $signed({1'h0, sel_260256}) ? {add_260253, array_index_258162[0]} : sel_260256;
  assign add_260578 = array_index_258427[11:0] + 12'h30f;
  assign sel_260580 = $signed({1'h0, add_260258}) < $signed({1'h0, sel_260260}) ? add_260258 : sel_260260;
  assign add_260582 = array_index_258430[11:0] + 12'h30f;
  assign sel_260584 = $signed({1'h0, add_260262}) < $signed({1'h0, sel_260264}) ? add_260262 : sel_260264;
  assign add_260586 = array_index_258585[11:0] + 12'hb55;
  assign sel_260588 = $signed({1'h0, add_260266}) < $signed({1'h0, sel_260268}) ? add_260266 : sel_260268;
  assign add_260590 = array_index_258588[11:0] + 12'hb55;
  assign sel_260592 = $signed({1'h0, add_260270}) < $signed({1'h0, sel_260272}) ? add_260270 : sel_260272;
  assign add_260594 = array_index_258761[11:0] + 12'h103;
  assign sel_260596 = $signed({1'h0, add_260274}) < $signed({1'h0, sel_260276}) ? add_260274 : sel_260276;
  assign add_260598 = array_index_258764[11:0] + 12'h103;
  assign sel_260600 = $signed({1'h0, add_260278}) < $signed({1'h0, sel_260280}) ? add_260278 : sel_260280;
  assign add_260602 = array_index_258957[11:0] + 12'hb01;
  assign sel_260604 = $signed({1'h0, add_260282}) < $signed({1'h0, sel_260284}) ? add_260282 : sel_260284;
  assign add_260606 = array_index_258960[11:0] + 12'hb01;
  assign sel_260608 = $signed({1'h0, add_260286}) < $signed({1'h0, sel_260288}) ? add_260286 : sel_260288;
  assign add_260610 = array_index_259171[11:0] + 12'h7b1;
  assign sel_260612 = $signed({1'h0, add_260290}) < $signed({1'h0, sel_260292}) ? add_260290 : sel_260292;
  assign add_260614 = array_index_259174[11:0] + 12'h7b1;
  assign sel_260616 = $signed({1'h0, add_260294}) < $signed({1'h0, sel_260296}) ? add_260294 : sel_260296;
  assign add_260618 = array_index_259401[11:0] + 12'h561;
  assign sel_260620 = $signed({1'h0, add_260298}) < $signed({1'h0, sel_260300}) ? add_260298 : sel_260300;
  assign add_260622 = array_index_259404[11:0] + 12'h561;
  assign sel_260624 = $signed({1'h0, add_260302}) < $signed({1'h0, sel_260304}) ? add_260302 : sel_260304;
  assign add_260626 = array_index_259647[11:2] + 10'h36b;
  assign sel_260628 = $signed({1'h0, add_260306, array_index_259401[1:0]}) < $signed({1'h0, sel_260308}) ? {add_260306, array_index_259401[1:0]} : sel_260308;
  assign add_260630 = array_index_259650[11:2] + 10'h36b;
  assign sel_260632 = $signed({1'h0, add_260310, array_index_259404[1:0]}) < $signed({1'h0, sel_260312}) ? {add_260310, array_index_259404[1:0]} : sel_260312;
  assign add_260634 = array_index_259911[11:2] + 10'h035;
  assign sel_260637 = $signed({1'h0, add_260314, array_index_259647[1:0]}) < $signed({1'h0, sel_260317}) ? {add_260314, array_index_259647[1:0]} : sel_260317;
  assign add_260639 = array_index_259914[11:2] + 10'h035;
  assign sel_260642 = $signed({1'h0, add_260319, array_index_259650[1:0]}) < $signed({1'h0, sel_260322}) ? {add_260319, array_index_259650[1:0]} : sel_260322;
  assign add_260644 = array_index_260195[11:0] + 12'hffb;
  assign sel_260646 = $signed({1'h0, add_260324}) < $signed({1'h0, sel_260326}) ? add_260324 : sel_260326;
  assign add_260648 = array_index_260198[11:0] + 12'hffb;
  assign sel_260650 = $signed({1'h0, add_260328}) < $signed({1'h0, sel_260330}) ? add_260328 : sel_260330;
  assign add_260664 = array_index_257775[11:0] + 12'h30b;
  assign sel_260666 = $signed({1'h0, add_260338}) < $signed(13'h0fff) ? add_260338 : 12'hfff;
  assign add_260668 = array_index_257778[11:0] + 12'h30b;
  assign sel_260670 = $signed({1'h0, add_260340}) < $signed(13'h0fff) ? add_260340 : 12'hfff;
  assign add_260739 = array_index_260507[11:0] + 12'h193;
  assign sel_260741 = $signed({1'h0, add_260411}) < $signed({1'h0, sel_260413}) ? add_260411 : sel_260413;
  assign add_260744 = array_index_260510[11:0] + 12'h193;
  assign sel_260746 = $signed({1'h0, add_260416}) < $signed({1'h0, sel_260418}) ? add_260416 : sel_260418;
  assign add_260748 = array_index_257761[11:0] + 12'h83f;
  assign add_260750 = array_index_257762[11:0] + 12'h83f;
  assign add_260764 = array_index_257817[11:1] + 11'h7b5;
  assign sel_260766 = $signed({1'h0, add_260426, array_index_257775[0]}) < $signed({1'h0, sel_260428}) ? {add_260426, array_index_257775[0]} : sel_260428;
  assign add_260768 = array_index_257820[11:1] + 11'h7b5;
  assign sel_260770 = $signed({1'h0, add_260430, array_index_257778[0]}) < $signed({1'h0, sel_260432}) ? {add_260430, array_index_257778[0]} : sel_260432;
  assign array_index_260845 = set1_unflattened[5'h12];
  assign array_index_260848 = set2_unflattened[5'h12];
  assign add_260858 = array_index_257775[11:1] + 11'h1e7;
  assign sel_260860 = $signed({1'h0, add_260514, array_index_257761[0]}) < $signed(13'h0fff) ? {add_260514, array_index_257761[0]} : 12'hfff;
  assign add_260862 = array_index_257778[11:1] + 11'h1e7;
  assign sel_260864 = $signed({1'h0, add_260516, array_index_257762[0]}) < $signed(13'h0fff) ? {add_260516, array_index_257762[0]} : 12'hfff;
  assign add_260874 = array_index_257877[11:0] + 12'h141;
  assign sel_260876 = $signed({1'h0, add_260528}) < $signed({1'h0, sel_260530}) ? add_260528 : sel_260530;
  assign add_260878 = array_index_257880[11:0] + 12'h141;
  assign sel_260880 = $signed({1'h0, add_260532}) < $signed({1'h0, sel_260534}) ? add_260532 : sel_260534;
  assign add_260882 = array_index_257955[11:1] + 11'h079;
  assign sel_260884 = $signed({1'h0, add_260536, array_index_257877[0]}) < $signed({1'h0, sel_260538}) ? {add_260536, array_index_257877[0]} : sel_260538;
  assign add_260886 = array_index_257958[11:1] + 11'h079;
  assign sel_260888 = $signed({1'h0, add_260540, array_index_257880[0]}) < $signed({1'h0, sel_260542}) ? {add_260540, array_index_257880[0]} : sel_260542;
  assign add_260890 = array_index_258049[11:0] + 12'h59d;
  assign sel_260892 = $signed({1'h0, add_260544}) < $signed({1'h0, sel_260546}) ? add_260544 : sel_260546;
  assign add_260894 = array_index_258052[11:0] + 12'h59d;
  assign sel_260896 = $signed({1'h0, add_260548}) < $signed({1'h0, sel_260550}) ? add_260548 : sel_260550;
  assign add_260898 = array_index_258159[11:0] + 12'ha6f;
  assign sel_260900 = $signed({1'h0, add_260552}) < $signed({1'h0, sel_260554}) ? add_260552 : sel_260554;
  assign add_260902 = array_index_258162[11:0] + 12'ha6f;
  assign sel_260904 = $signed({1'h0, add_260556}) < $signed({1'h0, sel_260558}) ? add_260556 : sel_260558;
  assign add_260906 = array_index_258285[11:1] + 11'h499;
  assign sel_260908 = $signed({1'h0, add_260560, array_index_258159[0]}) < $signed({1'h0, sel_260562}) ? {add_260560, array_index_258159[0]} : sel_260562;
  assign add_260910 = array_index_258288[11:1] + 11'h499;
  assign sel_260912 = $signed({1'h0, add_260564, array_index_258162[0]}) < $signed({1'h0, sel_260566}) ? {add_260564, array_index_258162[0]} : sel_260566;
  assign add_260914 = array_index_258427[11:1] + 11'h345;
  assign sel_260917 = $signed({1'h0, add_260568, array_index_258285[0]}) < $signed({1'h0, sel_260571}) ? {add_260568, array_index_258285[0]} : sel_260571;
  assign add_260919 = array_index_258430[11:1] + 11'h345;
  assign sel_260922 = $signed({1'h0, add_260573, array_index_258288[0]}) < $signed({1'h0, sel_260576}) ? {add_260573, array_index_258288[0]} : sel_260576;
  assign add_260924 = array_index_258585[11:0] + 12'h30f;
  assign sel_260926 = $signed({1'h0, add_260578}) < $signed({1'h0, sel_260580}) ? add_260578 : sel_260580;
  assign add_260928 = array_index_258588[11:0] + 12'h30f;
  assign sel_260930 = $signed({1'h0, add_260582}) < $signed({1'h0, sel_260584}) ? add_260582 : sel_260584;
  assign add_260932 = array_index_258761[11:0] + 12'hb55;
  assign sel_260934 = $signed({1'h0, add_260586}) < $signed({1'h0, sel_260588}) ? add_260586 : sel_260588;
  assign add_260936 = array_index_258764[11:0] + 12'hb55;
  assign sel_260938 = $signed({1'h0, add_260590}) < $signed({1'h0, sel_260592}) ? add_260590 : sel_260592;
  assign add_260940 = array_index_258957[11:0] + 12'h103;
  assign sel_260942 = $signed({1'h0, add_260594}) < $signed({1'h0, sel_260596}) ? add_260594 : sel_260596;
  assign add_260944 = array_index_258960[11:0] + 12'h103;
  assign sel_260946 = $signed({1'h0, add_260598}) < $signed({1'h0, sel_260600}) ? add_260598 : sel_260600;
  assign add_260948 = array_index_259171[11:0] + 12'hb01;
  assign sel_260950 = $signed({1'h0, add_260602}) < $signed({1'h0, sel_260604}) ? add_260602 : sel_260604;
  assign add_260952 = array_index_259174[11:0] + 12'hb01;
  assign sel_260954 = $signed({1'h0, add_260606}) < $signed({1'h0, sel_260608}) ? add_260606 : sel_260608;
  assign add_260956 = array_index_259401[11:0] + 12'h7b1;
  assign sel_260958 = $signed({1'h0, add_260610}) < $signed({1'h0, sel_260612}) ? add_260610 : sel_260612;
  assign add_260960 = array_index_259404[11:0] + 12'h7b1;
  assign sel_260962 = $signed({1'h0, add_260614}) < $signed({1'h0, sel_260616}) ? add_260614 : sel_260616;
  assign add_260964 = array_index_259647[11:0] + 12'h561;
  assign sel_260966 = $signed({1'h0, add_260618}) < $signed({1'h0, sel_260620}) ? add_260618 : sel_260620;
  assign add_260968 = array_index_259650[11:0] + 12'h561;
  assign sel_260970 = $signed({1'h0, add_260622}) < $signed({1'h0, sel_260624}) ? add_260622 : sel_260624;
  assign add_260972 = array_index_259911[11:2] + 10'h36b;
  assign sel_260974 = $signed({1'h0, add_260626, array_index_259647[1:0]}) < $signed({1'h0, sel_260628}) ? {add_260626, array_index_259647[1:0]} : sel_260628;
  assign add_260976 = array_index_259914[11:2] + 10'h36b;
  assign sel_260978 = $signed({1'h0, add_260630, array_index_259650[1:0]}) < $signed({1'h0, sel_260632}) ? {add_260630, array_index_259650[1:0]} : sel_260632;
  assign add_260980 = array_index_260195[11:2] + 10'h035;
  assign sel_260983 = $signed({1'h0, add_260634, array_index_259911[1:0]}) < $signed({1'h0, sel_260637}) ? {add_260634, array_index_259911[1:0]} : sel_260637;
  assign add_260985 = array_index_260198[11:2] + 10'h035;
  assign sel_260988 = $signed({1'h0, add_260639, array_index_259914[1:0]}) < $signed({1'h0, sel_260642}) ? {add_260639, array_index_259914[1:0]} : sel_260642;
  assign add_260990 = array_index_260507[11:0] + 12'hffb;
  assign sel_260992 = $signed({1'h0, add_260644}) < $signed({1'h0, sel_260646}) ? add_260644 : sel_260646;
  assign add_260994 = array_index_260510[11:0] + 12'hffb;
  assign sel_260996 = $signed({1'h0, add_260648}) < $signed({1'h0, sel_260650}) ? add_260648 : sel_260650;
  assign add_261004 = array_index_257761[11:0] + 12'h9cf;
  assign add_261006 = array_index_257762[11:0] + 12'h9cf;
  assign add_261018 = array_index_257817[11:0] + 12'h30b;
  assign sel_261020 = $signed({1'h0, add_260664}) < $signed({1'h0, sel_260666}) ? add_260664 : sel_260666;
  assign add_261022 = array_index_257820[11:0] + 12'h30b;
  assign sel_261024 = $signed({1'h0, add_260668}) < $signed({1'h0, sel_260670}) ? add_260668 : sel_260670;
  assign add_261093 = array_index_260845[11:0] + 12'h193;
  assign sel_261095 = $signed({1'h0, add_260739}) < $signed({1'h0, sel_260741}) ? add_260739 : sel_260741;
  assign add_261098 = array_index_260848[11:0] + 12'h193;
  assign sel_261100 = $signed({1'h0, add_260744}) < $signed({1'h0, sel_260746}) ? add_260744 : sel_260746;
  assign add_261108 = array_index_257775[11:0] + 12'h83f;
  assign sel_261110 = $signed({1'h0, add_260748}) < $signed(13'h0fff) ? add_260748 : 12'hfff;
  assign add_261112 = array_index_257778[11:0] + 12'h83f;
  assign sel_261114 = $signed({1'h0, add_260750}) < $signed(13'h0fff) ? add_260750 : 12'hfff;
  assign add_261126 = array_index_257877[11:1] + 11'h7b5;
  assign sel_261128 = $signed({1'h0, add_260764, array_index_257817[0]}) < $signed({1'h0, sel_260766}) ? {add_260764, array_index_257817[0]} : sel_260766;
  assign add_261130 = array_index_257880[11:1] + 11'h7b5;
  assign sel_261132 = $signed({1'h0, add_260768, array_index_257820[0]}) < $signed({1'h0, sel_260770}) ? {add_260768, array_index_257820[0]} : sel_260770;
  assign array_index_261207 = set1_unflattened[5'h13];
  assign array_index_261210 = set2_unflattened[5'h13];
  assign add_261214 = array_index_257761[11:2] + 10'h2b3;
  assign add_261216 = array_index_257762[11:2] + 10'h2b3;
  assign add_261228 = array_index_257817[11:1] + 11'h1e7;
  assign sel_261230 = $signed({1'h0, add_260858, array_index_257775[0]}) < $signed({1'h0, sel_260860}) ? {add_260858, array_index_257775[0]} : sel_260860;
  assign add_261232 = array_index_257820[11:1] + 11'h1e7;
  assign sel_261234 = $signed({1'h0, add_260862, array_index_257778[0]}) < $signed({1'h0, sel_260864}) ? {add_260862, array_index_257778[0]} : sel_260864;
  assign add_261244 = array_index_257955[11:0] + 12'h141;
  assign sel_261246 = $signed({1'h0, add_260874}) < $signed({1'h0, sel_260876}) ? add_260874 : sel_260876;
  assign add_261248 = array_index_257958[11:0] + 12'h141;
  assign sel_261250 = $signed({1'h0, add_260878}) < $signed({1'h0, sel_260880}) ? add_260878 : sel_260880;
  assign add_261252 = array_index_258049[11:1] + 11'h079;
  assign sel_261254 = $signed({1'h0, add_260882, array_index_257955[0]}) < $signed({1'h0, sel_260884}) ? {add_260882, array_index_257955[0]} : sel_260884;
  assign add_261256 = array_index_258052[11:1] + 11'h079;
  assign sel_261258 = $signed({1'h0, add_260886, array_index_257958[0]}) < $signed({1'h0, sel_260888}) ? {add_260886, array_index_257958[0]} : sel_260888;
  assign add_261260 = array_index_258159[11:0] + 12'h59d;
  assign sel_261262 = $signed({1'h0, add_260890}) < $signed({1'h0, sel_260892}) ? add_260890 : sel_260892;
  assign add_261264 = array_index_258162[11:0] + 12'h59d;
  assign sel_261266 = $signed({1'h0, add_260894}) < $signed({1'h0, sel_260896}) ? add_260894 : sel_260896;
  assign add_261268 = array_index_258285[11:0] + 12'ha6f;
  assign sel_261270 = $signed({1'h0, add_260898}) < $signed({1'h0, sel_260900}) ? add_260898 : sel_260900;
  assign add_261272 = array_index_258288[11:0] + 12'ha6f;
  assign sel_261274 = $signed({1'h0, add_260902}) < $signed({1'h0, sel_260904}) ? add_260902 : sel_260904;
  assign add_261276 = array_index_258427[11:1] + 11'h499;
  assign sel_261278 = $signed({1'h0, add_260906, array_index_258285[0]}) < $signed({1'h0, sel_260908}) ? {add_260906, array_index_258285[0]} : sel_260908;
  assign add_261280 = array_index_258430[11:1] + 11'h499;
  assign sel_261282 = $signed({1'h0, add_260910, array_index_258288[0]}) < $signed({1'h0, sel_260912}) ? {add_260910, array_index_258288[0]} : sel_260912;
  assign add_261284 = array_index_258585[11:1] + 11'h345;
  assign sel_261287 = $signed({1'h0, add_260914, array_index_258427[0]}) < $signed({1'h0, sel_260917}) ? {add_260914, array_index_258427[0]} : sel_260917;
  assign add_261289 = array_index_258588[11:1] + 11'h345;
  assign sel_261292 = $signed({1'h0, add_260919, array_index_258430[0]}) < $signed({1'h0, sel_260922}) ? {add_260919, array_index_258430[0]} : sel_260922;
  assign add_261294 = array_index_258761[11:0] + 12'h30f;
  assign sel_261296 = $signed({1'h0, add_260924}) < $signed({1'h0, sel_260926}) ? add_260924 : sel_260926;
  assign add_261298 = array_index_258764[11:0] + 12'h30f;
  assign sel_261300 = $signed({1'h0, add_260928}) < $signed({1'h0, sel_260930}) ? add_260928 : sel_260930;
  assign add_261302 = array_index_258957[11:0] + 12'hb55;
  assign sel_261304 = $signed({1'h0, add_260932}) < $signed({1'h0, sel_260934}) ? add_260932 : sel_260934;
  assign add_261306 = array_index_258960[11:0] + 12'hb55;
  assign sel_261308 = $signed({1'h0, add_260936}) < $signed({1'h0, sel_260938}) ? add_260936 : sel_260938;
  assign add_261310 = array_index_259171[11:0] + 12'h103;
  assign sel_261312 = $signed({1'h0, add_260940}) < $signed({1'h0, sel_260942}) ? add_260940 : sel_260942;
  assign add_261314 = array_index_259174[11:0] + 12'h103;
  assign sel_261316 = $signed({1'h0, add_260944}) < $signed({1'h0, sel_260946}) ? add_260944 : sel_260946;
  assign add_261318 = array_index_259401[11:0] + 12'hb01;
  assign sel_261320 = $signed({1'h0, add_260948}) < $signed({1'h0, sel_260950}) ? add_260948 : sel_260950;
  assign add_261322 = array_index_259404[11:0] + 12'hb01;
  assign sel_261324 = $signed({1'h0, add_260952}) < $signed({1'h0, sel_260954}) ? add_260952 : sel_260954;
  assign add_261326 = array_index_259647[11:0] + 12'h7b1;
  assign sel_261328 = $signed({1'h0, add_260956}) < $signed({1'h0, sel_260958}) ? add_260956 : sel_260958;
  assign add_261330 = array_index_259650[11:0] + 12'h7b1;
  assign sel_261332 = $signed({1'h0, add_260960}) < $signed({1'h0, sel_260962}) ? add_260960 : sel_260962;
  assign add_261334 = array_index_259911[11:0] + 12'h561;
  assign sel_261336 = $signed({1'h0, add_260964}) < $signed({1'h0, sel_260966}) ? add_260964 : sel_260966;
  assign add_261338 = array_index_259914[11:0] + 12'h561;
  assign sel_261340 = $signed({1'h0, add_260968}) < $signed({1'h0, sel_260970}) ? add_260968 : sel_260970;
  assign add_261342 = array_index_260195[11:2] + 10'h36b;
  assign sel_261344 = $signed({1'h0, add_260972, array_index_259911[1:0]}) < $signed({1'h0, sel_260974}) ? {add_260972, array_index_259911[1:0]} : sel_260974;
  assign add_261346 = array_index_260198[11:2] + 10'h36b;
  assign sel_261348 = $signed({1'h0, add_260976, array_index_259914[1:0]}) < $signed({1'h0, sel_260978}) ? {add_260976, array_index_259914[1:0]} : sel_260978;
  assign add_261350 = array_index_260507[11:2] + 10'h035;
  assign sel_261353 = $signed({1'h0, add_260980, array_index_260195[1:0]}) < $signed({1'h0, sel_260983}) ? {add_260980, array_index_260195[1:0]} : sel_260983;
  assign add_261355 = array_index_260510[11:2] + 10'h035;
  assign sel_261358 = $signed({1'h0, add_260985, array_index_260198[1:0]}) < $signed({1'h0, sel_260988}) ? {add_260985, array_index_260198[1:0]} : sel_260988;
  assign add_261360 = array_index_260845[11:0] + 12'hffb;
  assign sel_261362 = $signed({1'h0, add_260990}) < $signed({1'h0, sel_260992}) ? add_260990 : sel_260992;
  assign add_261364 = array_index_260848[11:0] + 12'hffb;
  assign sel_261366 = $signed({1'h0, add_260994}) < $signed({1'h0, sel_260996}) ? add_260994 : sel_260996;
  assign add_261380 = array_index_257775[11:0] + 12'h9cf;
  assign sel_261382 = $signed({1'h0, add_261004}) < $signed(13'h0fff) ? add_261004 : 12'hfff;
  assign add_261384 = array_index_257778[11:0] + 12'h9cf;
  assign sel_261386 = $signed({1'h0, add_261006}) < $signed(13'h0fff) ? add_261006 : 12'hfff;
  assign add_261396 = array_index_257877[11:0] + 12'h30b;
  assign sel_261398 = $signed({1'h0, add_261018}) < $signed({1'h0, sel_261020}) ? add_261018 : sel_261020;
  assign add_261400 = array_index_257880[11:0] + 12'h30b;
  assign sel_261402 = $signed({1'h0, add_261022}) < $signed({1'h0, sel_261024}) ? add_261022 : sel_261024;
  assign add_261471 = array_index_261207[11:0] + 12'h193;
  assign sel_261473 = $signed({1'h0, add_261093}) < $signed({1'h0, sel_261095}) ? add_261093 : sel_261095;
  assign add_261476 = array_index_261210[11:0] + 12'h193;
  assign sel_261478 = $signed({1'h0, add_261098}) < $signed({1'h0, sel_261100}) ? add_261098 : sel_261100;
  assign add_261480 = array_index_257761[11:0] + 12'hc05;
  assign add_261482 = array_index_257762[11:0] + 12'hc05;
  assign add_261496 = array_index_257817[11:0] + 12'h83f;
  assign sel_261498 = $signed({1'h0, add_261108}) < $signed({1'h0, sel_261110}) ? add_261108 : sel_261110;
  assign add_261500 = array_index_257820[11:0] + 12'h83f;
  assign sel_261502 = $signed({1'h0, add_261112}) < $signed({1'h0, sel_261114}) ? add_261112 : sel_261114;
  assign add_261514 = array_index_257955[11:1] + 11'h7b5;
  assign sel_261516 = $signed({1'h0, add_261126, array_index_257877[0]}) < $signed({1'h0, sel_261128}) ? {add_261126, array_index_257877[0]} : sel_261128;
  assign add_261518 = array_index_257958[11:1] + 11'h7b5;
  assign sel_261520 = $signed({1'h0, add_261130, array_index_257880[0]}) < $signed({1'h0, sel_261132}) ? {add_261130, array_index_257880[0]} : sel_261132;
  assign array_index_261595 = set1_unflattened[5'h14];
  assign array_index_261598 = set2_unflattened[5'h14];
  assign add_261608 = array_index_257775[11:2] + 10'h2b3;
  assign sel_261610 = $signed({1'h0, add_261214, array_index_257761[1:0]}) < $signed(13'h0fff) ? {add_261214, array_index_257761[1:0]} : 12'hfff;
  assign add_261612 = array_index_257778[11:2] + 10'h2b3;
  assign sel_261614 = $signed({1'h0, add_261216, array_index_257762[1:0]}) < $signed(13'h0fff) ? {add_261216, array_index_257762[1:0]} : 12'hfff;
  assign add_261624 = array_index_257877[11:1] + 11'h1e7;
  assign sel_261626 = $signed({1'h0, add_261228, array_index_257817[0]}) < $signed({1'h0, sel_261230}) ? {add_261228, array_index_257817[0]} : sel_261230;
  assign add_261628 = array_index_257880[11:1] + 11'h1e7;
  assign sel_261630 = $signed({1'h0, add_261232, array_index_257820[0]}) < $signed({1'h0, sel_261234}) ? {add_261232, array_index_257820[0]} : sel_261234;
  assign add_261640 = array_index_258049[11:0] + 12'h141;
  assign sel_261642 = $signed({1'h0, add_261244}) < $signed({1'h0, sel_261246}) ? add_261244 : sel_261246;
  assign add_261644 = array_index_258052[11:0] + 12'h141;
  assign sel_261646 = $signed({1'h0, add_261248}) < $signed({1'h0, sel_261250}) ? add_261248 : sel_261250;
  assign add_261648 = array_index_258159[11:1] + 11'h079;
  assign sel_261650 = $signed({1'h0, add_261252, array_index_258049[0]}) < $signed({1'h0, sel_261254}) ? {add_261252, array_index_258049[0]} : sel_261254;
  assign add_261652 = array_index_258162[11:1] + 11'h079;
  assign sel_261654 = $signed({1'h0, add_261256, array_index_258052[0]}) < $signed({1'h0, sel_261258}) ? {add_261256, array_index_258052[0]} : sel_261258;
  assign add_261656 = array_index_258285[11:0] + 12'h59d;
  assign sel_261658 = $signed({1'h0, add_261260}) < $signed({1'h0, sel_261262}) ? add_261260 : sel_261262;
  assign add_261660 = array_index_258288[11:0] + 12'h59d;
  assign sel_261662 = $signed({1'h0, add_261264}) < $signed({1'h0, sel_261266}) ? add_261264 : sel_261266;
  assign add_261664 = array_index_258427[11:0] + 12'ha6f;
  assign sel_261666 = $signed({1'h0, add_261268}) < $signed({1'h0, sel_261270}) ? add_261268 : sel_261270;
  assign add_261668 = array_index_258430[11:0] + 12'ha6f;
  assign sel_261670 = $signed({1'h0, add_261272}) < $signed({1'h0, sel_261274}) ? add_261272 : sel_261274;
  assign add_261672 = array_index_258585[11:1] + 11'h499;
  assign sel_261674 = $signed({1'h0, add_261276, array_index_258427[0]}) < $signed({1'h0, sel_261278}) ? {add_261276, array_index_258427[0]} : sel_261278;
  assign add_261676 = array_index_258588[11:1] + 11'h499;
  assign sel_261678 = $signed({1'h0, add_261280, array_index_258430[0]}) < $signed({1'h0, sel_261282}) ? {add_261280, array_index_258430[0]} : sel_261282;
  assign add_261680 = array_index_258761[11:1] + 11'h345;
  assign sel_261683 = $signed({1'h0, add_261284, array_index_258585[0]}) < $signed({1'h0, sel_261287}) ? {add_261284, array_index_258585[0]} : sel_261287;
  assign add_261685 = array_index_258764[11:1] + 11'h345;
  assign sel_261688 = $signed({1'h0, add_261289, array_index_258588[0]}) < $signed({1'h0, sel_261292}) ? {add_261289, array_index_258588[0]} : sel_261292;
  assign add_261690 = array_index_258957[11:0] + 12'h30f;
  assign sel_261692 = $signed({1'h0, add_261294}) < $signed({1'h0, sel_261296}) ? add_261294 : sel_261296;
  assign add_261694 = array_index_258960[11:0] + 12'h30f;
  assign sel_261696 = $signed({1'h0, add_261298}) < $signed({1'h0, sel_261300}) ? add_261298 : sel_261300;
  assign add_261698 = array_index_259171[11:0] + 12'hb55;
  assign sel_261700 = $signed({1'h0, add_261302}) < $signed({1'h0, sel_261304}) ? add_261302 : sel_261304;
  assign add_261702 = array_index_259174[11:0] + 12'hb55;
  assign sel_261704 = $signed({1'h0, add_261306}) < $signed({1'h0, sel_261308}) ? add_261306 : sel_261308;
  assign add_261706 = array_index_259401[11:0] + 12'h103;
  assign sel_261708 = $signed({1'h0, add_261310}) < $signed({1'h0, sel_261312}) ? add_261310 : sel_261312;
  assign add_261710 = array_index_259404[11:0] + 12'h103;
  assign sel_261712 = $signed({1'h0, add_261314}) < $signed({1'h0, sel_261316}) ? add_261314 : sel_261316;
  assign add_261714 = array_index_259647[11:0] + 12'hb01;
  assign sel_261716 = $signed({1'h0, add_261318}) < $signed({1'h0, sel_261320}) ? add_261318 : sel_261320;
  assign add_261718 = array_index_259650[11:0] + 12'hb01;
  assign sel_261720 = $signed({1'h0, add_261322}) < $signed({1'h0, sel_261324}) ? add_261322 : sel_261324;
  assign add_261722 = array_index_259911[11:0] + 12'h7b1;
  assign sel_261724 = $signed({1'h0, add_261326}) < $signed({1'h0, sel_261328}) ? add_261326 : sel_261328;
  assign add_261726 = array_index_259914[11:0] + 12'h7b1;
  assign sel_261728 = $signed({1'h0, add_261330}) < $signed({1'h0, sel_261332}) ? add_261330 : sel_261332;
  assign add_261730 = array_index_260195[11:0] + 12'h561;
  assign sel_261732 = $signed({1'h0, add_261334}) < $signed({1'h0, sel_261336}) ? add_261334 : sel_261336;
  assign add_261734 = array_index_260198[11:0] + 12'h561;
  assign sel_261736 = $signed({1'h0, add_261338}) < $signed({1'h0, sel_261340}) ? add_261338 : sel_261340;
  assign add_261738 = array_index_260507[11:2] + 10'h36b;
  assign sel_261740 = $signed({1'h0, add_261342, array_index_260195[1:0]}) < $signed({1'h0, sel_261344}) ? {add_261342, array_index_260195[1:0]} : sel_261344;
  assign add_261742 = array_index_260510[11:2] + 10'h36b;
  assign sel_261744 = $signed({1'h0, add_261346, array_index_260198[1:0]}) < $signed({1'h0, sel_261348}) ? {add_261346, array_index_260198[1:0]} : sel_261348;
  assign add_261746 = array_index_260845[11:2] + 10'h035;
  assign sel_261749 = $signed({1'h0, add_261350, array_index_260507[1:0]}) < $signed({1'h0, sel_261353}) ? {add_261350, array_index_260507[1:0]} : sel_261353;
  assign add_261751 = array_index_260848[11:2] + 10'h035;
  assign sel_261754 = $signed({1'h0, add_261355, array_index_260510[1:0]}) < $signed({1'h0, sel_261358}) ? {add_261355, array_index_260510[1:0]} : sel_261358;
  assign add_261756 = array_index_261207[11:0] + 12'hffb;
  assign sel_261758 = $signed({1'h0, add_261360}) < $signed({1'h0, sel_261362}) ? add_261360 : sel_261362;
  assign add_261760 = array_index_261210[11:0] + 12'hffb;
  assign sel_261762 = $signed({1'h0, add_261364}) < $signed({1'h0, sel_261366}) ? add_261364 : sel_261366;
  assign add_261770 = array_index_257761[11:2] + 10'h29b;
  assign add_261772 = array_index_257762[11:2] + 10'h29b;
  assign add_261784 = array_index_257817[11:0] + 12'h9cf;
  assign sel_261786 = $signed({1'h0, add_261380}) < $signed({1'h0, sel_261382}) ? add_261380 : sel_261382;
  assign add_261788 = array_index_257820[11:0] + 12'h9cf;
  assign sel_261790 = $signed({1'h0, add_261384}) < $signed({1'h0, sel_261386}) ? add_261384 : sel_261386;
  assign add_261800 = array_index_257955[11:0] + 12'h30b;
  assign sel_261802 = $signed({1'h0, add_261396}) < $signed({1'h0, sel_261398}) ? add_261396 : sel_261398;
  assign add_261804 = array_index_257958[11:0] + 12'h30b;
  assign sel_261806 = $signed({1'h0, add_261400}) < $signed({1'h0, sel_261402}) ? add_261400 : sel_261402;
  assign add_261875 = array_index_261595[11:0] + 12'h193;
  assign sel_261877 = $signed({1'h0, add_261471}) < $signed({1'h0, sel_261473}) ? add_261471 : sel_261473;
  assign add_261880 = array_index_261598[11:0] + 12'h193;
  assign sel_261882 = $signed({1'h0, add_261476}) < $signed({1'h0, sel_261478}) ? add_261476 : sel_261478;
  assign add_261890 = array_index_257775[11:0] + 12'hc05;
  assign sel_261892 = $signed({1'h0, add_261480}) < $signed(13'h0fff) ? add_261480 : 12'hfff;
  assign add_261894 = array_index_257778[11:0] + 12'hc05;
  assign sel_261896 = $signed({1'h0, add_261482}) < $signed(13'h0fff) ? add_261482 : 12'hfff;
  assign add_261908 = array_index_257877[11:0] + 12'h83f;
  assign sel_261910 = $signed({1'h0, add_261496}) < $signed({1'h0, sel_261498}) ? add_261496 : sel_261498;
  assign add_261912 = array_index_257880[11:0] + 12'h83f;
  assign sel_261914 = $signed({1'h0, add_261500}) < $signed({1'h0, sel_261502}) ? add_261500 : sel_261502;
  assign add_261926 = array_index_258049[11:1] + 11'h7b5;
  assign sel_261928 = $signed({1'h0, add_261514, array_index_257955[0]}) < $signed({1'h0, sel_261516}) ? {add_261514, array_index_257955[0]} : sel_261516;
  assign add_261930 = array_index_258052[11:1] + 11'h7b5;
  assign sel_261932 = $signed({1'h0, add_261518, array_index_257958[0]}) < $signed({1'h0, sel_261520}) ? {add_261518, array_index_257958[0]} : sel_261520;
  assign array_index_262007 = set1_unflattened[5'h15];
  assign array_index_262010 = set2_unflattened[5'h15];
  assign add_262014 = array_index_257761[11:0] + 12'hdab;
  assign add_262016 = array_index_257762[11:0] + 12'hdab;
  assign add_262030 = array_index_257817[11:2] + 10'h2b3;
  assign sel_262032 = $signed({1'h0, add_261608, array_index_257775[1:0]}) < $signed({1'h0, sel_261610}) ? {add_261608, array_index_257775[1:0]} : sel_261610;
  assign add_262034 = array_index_257820[11:2] + 10'h2b3;
  assign sel_262036 = $signed({1'h0, add_261612, array_index_257778[1:0]}) < $signed({1'h0, sel_261614}) ? {add_261612, array_index_257778[1:0]} : sel_261614;
  assign add_262046 = array_index_257955[11:1] + 11'h1e7;
  assign sel_262048 = $signed({1'h0, add_261624, array_index_257877[0]}) < $signed({1'h0, sel_261626}) ? {add_261624, array_index_257877[0]} : sel_261626;
  assign add_262050 = array_index_257958[11:1] + 11'h1e7;
  assign sel_262052 = $signed({1'h0, add_261628, array_index_257880[0]}) < $signed({1'h0, sel_261630}) ? {add_261628, array_index_257880[0]} : sel_261630;
  assign add_262062 = array_index_258159[11:0] + 12'h141;
  assign sel_262064 = $signed({1'h0, add_261640}) < $signed({1'h0, sel_261642}) ? add_261640 : sel_261642;
  assign add_262066 = array_index_258162[11:0] + 12'h141;
  assign sel_262068 = $signed({1'h0, add_261644}) < $signed({1'h0, sel_261646}) ? add_261644 : sel_261646;
  assign add_262070 = array_index_258285[11:1] + 11'h079;
  assign sel_262072 = $signed({1'h0, add_261648, array_index_258159[0]}) < $signed({1'h0, sel_261650}) ? {add_261648, array_index_258159[0]} : sel_261650;
  assign add_262074 = array_index_258288[11:1] + 11'h079;
  assign sel_262076 = $signed({1'h0, add_261652, array_index_258162[0]}) < $signed({1'h0, sel_261654}) ? {add_261652, array_index_258162[0]} : sel_261654;
  assign add_262078 = array_index_258427[11:0] + 12'h59d;
  assign sel_262080 = $signed({1'h0, add_261656}) < $signed({1'h0, sel_261658}) ? add_261656 : sel_261658;
  assign add_262082 = array_index_258430[11:0] + 12'h59d;
  assign sel_262084 = $signed({1'h0, add_261660}) < $signed({1'h0, sel_261662}) ? add_261660 : sel_261662;
  assign add_262086 = array_index_258585[11:0] + 12'ha6f;
  assign sel_262088 = $signed({1'h0, add_261664}) < $signed({1'h0, sel_261666}) ? add_261664 : sel_261666;
  assign add_262090 = array_index_258588[11:0] + 12'ha6f;
  assign sel_262092 = $signed({1'h0, add_261668}) < $signed({1'h0, sel_261670}) ? add_261668 : sel_261670;
  assign add_262094 = array_index_258761[11:1] + 11'h499;
  assign sel_262096 = $signed({1'h0, add_261672, array_index_258585[0]}) < $signed({1'h0, sel_261674}) ? {add_261672, array_index_258585[0]} : sel_261674;
  assign add_262098 = array_index_258764[11:1] + 11'h499;
  assign sel_262100 = $signed({1'h0, add_261676, array_index_258588[0]}) < $signed({1'h0, sel_261678}) ? {add_261676, array_index_258588[0]} : sel_261678;
  assign add_262102 = array_index_258957[11:1] + 11'h345;
  assign sel_262105 = $signed({1'h0, add_261680, array_index_258761[0]}) < $signed({1'h0, sel_261683}) ? {add_261680, array_index_258761[0]} : sel_261683;
  assign add_262107 = array_index_258960[11:1] + 11'h345;
  assign sel_262110 = $signed({1'h0, add_261685, array_index_258764[0]}) < $signed({1'h0, sel_261688}) ? {add_261685, array_index_258764[0]} : sel_261688;
  assign add_262112 = array_index_259171[11:0] + 12'h30f;
  assign sel_262114 = $signed({1'h0, add_261690}) < $signed({1'h0, sel_261692}) ? add_261690 : sel_261692;
  assign add_262116 = array_index_259174[11:0] + 12'h30f;
  assign sel_262118 = $signed({1'h0, add_261694}) < $signed({1'h0, sel_261696}) ? add_261694 : sel_261696;
  assign add_262120 = array_index_259401[11:0] + 12'hb55;
  assign sel_262122 = $signed({1'h0, add_261698}) < $signed({1'h0, sel_261700}) ? add_261698 : sel_261700;
  assign add_262124 = array_index_259404[11:0] + 12'hb55;
  assign sel_262126 = $signed({1'h0, add_261702}) < $signed({1'h0, sel_261704}) ? add_261702 : sel_261704;
  assign add_262128 = array_index_259647[11:0] + 12'h103;
  assign sel_262130 = $signed({1'h0, add_261706}) < $signed({1'h0, sel_261708}) ? add_261706 : sel_261708;
  assign add_262132 = array_index_259650[11:0] + 12'h103;
  assign sel_262134 = $signed({1'h0, add_261710}) < $signed({1'h0, sel_261712}) ? add_261710 : sel_261712;
  assign add_262136 = array_index_259911[11:0] + 12'hb01;
  assign sel_262138 = $signed({1'h0, add_261714}) < $signed({1'h0, sel_261716}) ? add_261714 : sel_261716;
  assign add_262140 = array_index_259914[11:0] + 12'hb01;
  assign sel_262142 = $signed({1'h0, add_261718}) < $signed({1'h0, sel_261720}) ? add_261718 : sel_261720;
  assign add_262144 = array_index_260195[11:0] + 12'h7b1;
  assign sel_262146 = $signed({1'h0, add_261722}) < $signed({1'h0, sel_261724}) ? add_261722 : sel_261724;
  assign add_262148 = array_index_260198[11:0] + 12'h7b1;
  assign sel_262150 = $signed({1'h0, add_261726}) < $signed({1'h0, sel_261728}) ? add_261726 : sel_261728;
  assign add_262152 = array_index_260507[11:0] + 12'h561;
  assign sel_262154 = $signed({1'h0, add_261730}) < $signed({1'h0, sel_261732}) ? add_261730 : sel_261732;
  assign add_262156 = array_index_260510[11:0] + 12'h561;
  assign sel_262158 = $signed({1'h0, add_261734}) < $signed({1'h0, sel_261736}) ? add_261734 : sel_261736;
  assign add_262160 = array_index_260845[11:2] + 10'h36b;
  assign sel_262162 = $signed({1'h0, add_261738, array_index_260507[1:0]}) < $signed({1'h0, sel_261740}) ? {add_261738, array_index_260507[1:0]} : sel_261740;
  assign add_262164 = array_index_260848[11:2] + 10'h36b;
  assign sel_262166 = $signed({1'h0, add_261742, array_index_260510[1:0]}) < $signed({1'h0, sel_261744}) ? {add_261742, array_index_260510[1:0]} : sel_261744;
  assign add_262168 = array_index_261207[11:2] + 10'h035;
  assign sel_262171 = $signed({1'h0, add_261746, array_index_260845[1:0]}) < $signed({1'h0, sel_261749}) ? {add_261746, array_index_260845[1:0]} : sel_261749;
  assign add_262173 = array_index_261210[11:2] + 10'h035;
  assign sel_262176 = $signed({1'h0, add_261751, array_index_260848[1:0]}) < $signed({1'h0, sel_261754}) ? {add_261751, array_index_260848[1:0]} : sel_261754;
  assign add_262178 = array_index_261595[11:0] + 12'hffb;
  assign sel_262180 = $signed({1'h0, add_261756}) < $signed({1'h0, sel_261758}) ? add_261756 : sel_261758;
  assign add_262182 = array_index_261598[11:0] + 12'hffb;
  assign sel_262184 = $signed({1'h0, add_261760}) < $signed({1'h0, sel_261762}) ? add_261760 : sel_261762;
  assign add_262196 = array_index_257775[11:2] + 10'h29b;
  assign sel_262198 = $signed({1'h0, add_261770, array_index_257761[1:0]}) < $signed(13'h0fff) ? {add_261770, array_index_257761[1:0]} : 12'hfff;
  assign add_262200 = array_index_257778[11:2] + 10'h29b;
  assign sel_262202 = $signed({1'h0, add_261772, array_index_257762[1:0]}) < $signed(13'h0fff) ? {add_261772, array_index_257762[1:0]} : 12'hfff;
  assign add_262212 = array_index_257877[11:0] + 12'h9cf;
  assign sel_262214 = $signed({1'h0, add_261784}) < $signed({1'h0, sel_261786}) ? add_261784 : sel_261786;
  assign add_262216 = array_index_257880[11:0] + 12'h9cf;
  assign sel_262218 = $signed({1'h0, add_261788}) < $signed({1'h0, sel_261790}) ? add_261788 : sel_261790;
  assign add_262228 = array_index_258049[11:0] + 12'h30b;
  assign sel_262230 = $signed({1'h0, add_261800}) < $signed({1'h0, sel_261802}) ? add_261800 : sel_261802;
  assign add_262232 = array_index_258052[11:0] + 12'h30b;
  assign sel_262234 = $signed({1'h0, add_261804}) < $signed({1'h0, sel_261806}) ? add_261804 : sel_261806;
  assign add_262303 = array_index_262007[11:0] + 12'h193;
  assign sel_262305 = $signed({1'h0, add_261875}) < $signed({1'h0, sel_261877}) ? add_261875 : sel_261877;
  assign add_262308 = array_index_262010[11:0] + 12'h193;
  assign sel_262310 = $signed({1'h0, add_261880}) < $signed({1'h0, sel_261882}) ? add_261880 : sel_261882;
  assign add_262322 = array_index_257817[11:0] + 12'hc05;
  assign sel_262324 = $signed({1'h0, add_261890}) < $signed({1'h0, sel_261892}) ? add_261890 : sel_261892;
  assign add_262326 = array_index_257820[11:0] + 12'hc05;
  assign sel_262328 = $signed({1'h0, add_261894}) < $signed({1'h0, sel_261896}) ? add_261894 : sel_261896;
  assign add_262340 = array_index_257955[11:0] + 12'h83f;
  assign sel_262342 = $signed({1'h0, add_261908}) < $signed({1'h0, sel_261910}) ? add_261908 : sel_261910;
  assign add_262344 = array_index_257958[11:0] + 12'h83f;
  assign sel_262346 = $signed({1'h0, add_261912}) < $signed({1'h0, sel_261914}) ? add_261912 : sel_261914;
  assign add_262358 = array_index_258159[11:1] + 11'h7b5;
  assign sel_262360 = $signed({1'h0, add_261926, array_index_258049[0]}) < $signed({1'h0, sel_261928}) ? {add_261926, array_index_258049[0]} : sel_261928;
  assign add_262362 = array_index_258162[11:1] + 11'h7b5;
  assign sel_262364 = $signed({1'h0, add_261930, array_index_258052[0]}) < $signed({1'h0, sel_261932}) ? {add_261930, array_index_258052[0]} : sel_261932;
  assign array_index_262439 = set1_unflattened[5'h16];
  assign array_index_262442 = set2_unflattened[5'h16];
  assign add_262446 = array_index_257775[11:0] + 12'hdab;
  assign sel_262448 = $signed({1'h0, add_262014}) < $signed(13'h0fff) ? add_262014 : 12'hfff;
  assign add_262450 = array_index_257778[11:0] + 12'hdab;
  assign sel_262452 = $signed({1'h0, add_262016}) < $signed(13'h0fff) ? add_262016 : 12'hfff;
  assign add_262464 = array_index_257877[11:2] + 10'h2b3;
  assign sel_262466 = $signed({1'h0, add_262030, array_index_257817[1:0]}) < $signed({1'h0, sel_262032}) ? {add_262030, array_index_257817[1:0]} : sel_262032;
  assign add_262468 = array_index_257880[11:2] + 10'h2b3;
  assign sel_262470 = $signed({1'h0, add_262034, array_index_257820[1:0]}) < $signed({1'h0, sel_262036}) ? {add_262034, array_index_257820[1:0]} : sel_262036;
  assign add_262480 = array_index_258049[11:1] + 11'h1e7;
  assign sel_262482 = $signed({1'h0, add_262046, array_index_257955[0]}) < $signed({1'h0, sel_262048}) ? {add_262046, array_index_257955[0]} : sel_262048;
  assign add_262484 = array_index_258052[11:1] + 11'h1e7;
  assign sel_262486 = $signed({1'h0, add_262050, array_index_257958[0]}) < $signed({1'h0, sel_262052}) ? {add_262050, array_index_257958[0]} : sel_262052;
  assign add_262496 = array_index_258285[11:0] + 12'h141;
  assign sel_262498 = $signed({1'h0, add_262062}) < $signed({1'h0, sel_262064}) ? add_262062 : sel_262064;
  assign add_262500 = array_index_258288[11:0] + 12'h141;
  assign sel_262502 = $signed({1'h0, add_262066}) < $signed({1'h0, sel_262068}) ? add_262066 : sel_262068;
  assign add_262504 = array_index_258427[11:1] + 11'h079;
  assign sel_262506 = $signed({1'h0, add_262070, array_index_258285[0]}) < $signed({1'h0, sel_262072}) ? {add_262070, array_index_258285[0]} : sel_262072;
  assign add_262508 = array_index_258430[11:1] + 11'h079;
  assign sel_262510 = $signed({1'h0, add_262074, array_index_258288[0]}) < $signed({1'h0, sel_262076}) ? {add_262074, array_index_258288[0]} : sel_262076;
  assign add_262512 = array_index_258585[11:0] + 12'h59d;
  assign sel_262514 = $signed({1'h0, add_262078}) < $signed({1'h0, sel_262080}) ? add_262078 : sel_262080;
  assign add_262516 = array_index_258588[11:0] + 12'h59d;
  assign sel_262518 = $signed({1'h0, add_262082}) < $signed({1'h0, sel_262084}) ? add_262082 : sel_262084;
  assign add_262520 = array_index_258761[11:0] + 12'ha6f;
  assign sel_262522 = $signed({1'h0, add_262086}) < $signed({1'h0, sel_262088}) ? add_262086 : sel_262088;
  assign add_262524 = array_index_258764[11:0] + 12'ha6f;
  assign sel_262526 = $signed({1'h0, add_262090}) < $signed({1'h0, sel_262092}) ? add_262090 : sel_262092;
  assign add_262528 = array_index_258957[11:1] + 11'h499;
  assign sel_262530 = $signed({1'h0, add_262094, array_index_258761[0]}) < $signed({1'h0, sel_262096}) ? {add_262094, array_index_258761[0]} : sel_262096;
  assign add_262532 = array_index_258960[11:1] + 11'h499;
  assign sel_262534 = $signed({1'h0, add_262098, array_index_258764[0]}) < $signed({1'h0, sel_262100}) ? {add_262098, array_index_258764[0]} : sel_262100;
  assign add_262536 = array_index_259171[11:1] + 11'h345;
  assign sel_262539 = $signed({1'h0, add_262102, array_index_258957[0]}) < $signed({1'h0, sel_262105}) ? {add_262102, array_index_258957[0]} : sel_262105;
  assign add_262541 = array_index_259174[11:1] + 11'h345;
  assign sel_262544 = $signed({1'h0, add_262107, array_index_258960[0]}) < $signed({1'h0, sel_262110}) ? {add_262107, array_index_258960[0]} : sel_262110;
  assign add_262546 = array_index_259401[11:0] + 12'h30f;
  assign sel_262548 = $signed({1'h0, add_262112}) < $signed({1'h0, sel_262114}) ? add_262112 : sel_262114;
  assign add_262550 = array_index_259404[11:0] + 12'h30f;
  assign sel_262552 = $signed({1'h0, add_262116}) < $signed({1'h0, sel_262118}) ? add_262116 : sel_262118;
  assign add_262554 = array_index_259647[11:0] + 12'hb55;
  assign sel_262556 = $signed({1'h0, add_262120}) < $signed({1'h0, sel_262122}) ? add_262120 : sel_262122;
  assign add_262558 = array_index_259650[11:0] + 12'hb55;
  assign sel_262560 = $signed({1'h0, add_262124}) < $signed({1'h0, sel_262126}) ? add_262124 : sel_262126;
  assign add_262562 = array_index_259911[11:0] + 12'h103;
  assign sel_262564 = $signed({1'h0, add_262128}) < $signed({1'h0, sel_262130}) ? add_262128 : sel_262130;
  assign add_262566 = array_index_259914[11:0] + 12'h103;
  assign sel_262568 = $signed({1'h0, add_262132}) < $signed({1'h0, sel_262134}) ? add_262132 : sel_262134;
  assign add_262570 = array_index_260195[11:0] + 12'hb01;
  assign sel_262572 = $signed({1'h0, add_262136}) < $signed({1'h0, sel_262138}) ? add_262136 : sel_262138;
  assign add_262574 = array_index_260198[11:0] + 12'hb01;
  assign sel_262576 = $signed({1'h0, add_262140}) < $signed({1'h0, sel_262142}) ? add_262140 : sel_262142;
  assign add_262578 = array_index_260507[11:0] + 12'h7b1;
  assign sel_262580 = $signed({1'h0, add_262144}) < $signed({1'h0, sel_262146}) ? add_262144 : sel_262146;
  assign add_262582 = array_index_260510[11:0] + 12'h7b1;
  assign sel_262584 = $signed({1'h0, add_262148}) < $signed({1'h0, sel_262150}) ? add_262148 : sel_262150;
  assign add_262586 = array_index_260845[11:0] + 12'h561;
  assign sel_262588 = $signed({1'h0, add_262152}) < $signed({1'h0, sel_262154}) ? add_262152 : sel_262154;
  assign add_262590 = array_index_260848[11:0] + 12'h561;
  assign sel_262592 = $signed({1'h0, add_262156}) < $signed({1'h0, sel_262158}) ? add_262156 : sel_262158;
  assign add_262594 = array_index_261207[11:2] + 10'h36b;
  assign sel_262596 = $signed({1'h0, add_262160, array_index_260845[1:0]}) < $signed({1'h0, sel_262162}) ? {add_262160, array_index_260845[1:0]} : sel_262162;
  assign add_262598 = array_index_261210[11:2] + 10'h36b;
  assign sel_262600 = $signed({1'h0, add_262164, array_index_260848[1:0]}) < $signed({1'h0, sel_262166}) ? {add_262164, array_index_260848[1:0]} : sel_262166;
  assign add_262602 = array_index_261595[11:2] + 10'h035;
  assign sel_262605 = $signed({1'h0, add_262168, array_index_261207[1:0]}) < $signed({1'h0, sel_262171}) ? {add_262168, array_index_261207[1:0]} : sel_262171;
  assign add_262607 = array_index_261598[11:2] + 10'h035;
  assign sel_262610 = $signed({1'h0, add_262173, array_index_261210[1:0]}) < $signed({1'h0, sel_262176}) ? {add_262173, array_index_261210[1:0]} : sel_262176;
  assign add_262612 = array_index_262007[11:0] + 12'hffb;
  assign sel_262614 = $signed({1'h0, add_262178}) < $signed({1'h0, sel_262180}) ? add_262178 : sel_262180;
  assign add_262616 = array_index_262010[11:0] + 12'hffb;
  assign sel_262618 = $signed({1'h0, add_262182}) < $signed({1'h0, sel_262184}) ? add_262182 : sel_262184;
  assign add_262630 = array_index_257817[11:2] + 10'h29b;
  assign sel_262632 = $signed({1'h0, add_262196, array_index_257775[1:0]}) < $signed({1'h0, sel_262198}) ? {add_262196, array_index_257775[1:0]} : sel_262198;
  assign add_262634 = array_index_257820[11:2] + 10'h29b;
  assign sel_262636 = $signed({1'h0, add_262200, array_index_257778[1:0]}) < $signed({1'h0, sel_262202}) ? {add_262200, array_index_257778[1:0]} : sel_262202;
  assign add_262646 = array_index_257955[11:0] + 12'h9cf;
  assign sel_262648 = $signed({1'h0, add_262212}) < $signed({1'h0, sel_262214}) ? add_262212 : sel_262214;
  assign add_262650 = array_index_257958[11:0] + 12'h9cf;
  assign sel_262652 = $signed({1'h0, add_262216}) < $signed({1'h0, sel_262218}) ? add_262216 : sel_262218;
  assign add_262662 = array_index_258159[11:0] + 12'h30b;
  assign sel_262664 = $signed({1'h0, add_262228}) < $signed({1'h0, sel_262230}) ? add_262228 : sel_262230;
  assign add_262666 = array_index_258162[11:0] + 12'h30b;
  assign sel_262668 = $signed({1'h0, add_262232}) < $signed({1'h0, sel_262234}) ? add_262232 : sel_262234;
  assign add_262737 = array_index_262439[11:0] + 12'h193;
  assign sel_262739 = $signed({1'h0, add_262303}) < $signed({1'h0, sel_262305}) ? add_262303 : sel_262305;
  assign add_262742 = array_index_262442[11:0] + 12'h193;
  assign sel_262744 = $signed({1'h0, add_262308}) < $signed({1'h0, sel_262310}) ? add_262308 : sel_262310;
  assign add_262754 = array_index_257877[11:0] + 12'hc05;
  assign sel_262756 = $signed({1'h0, add_262322}) < $signed({1'h0, sel_262324}) ? add_262322 : sel_262324;
  assign add_262758 = array_index_257880[11:0] + 12'hc05;
  assign sel_262760 = $signed({1'h0, add_262326}) < $signed({1'h0, sel_262328}) ? add_262326 : sel_262328;
  assign add_262772 = array_index_258049[11:0] + 12'h83f;
  assign sel_262774 = $signed({1'h0, add_262340}) < $signed({1'h0, sel_262342}) ? add_262340 : sel_262342;
  assign add_262776 = array_index_258052[11:0] + 12'h83f;
  assign sel_262778 = $signed({1'h0, add_262344}) < $signed({1'h0, sel_262346}) ? add_262344 : sel_262346;
  assign add_262790 = array_index_258285[11:1] + 11'h7b5;
  assign sel_262792 = $signed({1'h0, add_262358, array_index_258159[0]}) < $signed({1'h0, sel_262360}) ? {add_262358, array_index_258159[0]} : sel_262360;
  assign add_262794 = array_index_258288[11:1] + 11'h7b5;
  assign sel_262796 = $signed({1'h0, add_262362, array_index_258162[0]}) < $signed({1'h0, sel_262364}) ? {add_262362, array_index_258162[0]} : sel_262364;
  assign array_index_262871 = set1_unflattened[5'h17];
  assign array_index_262874 = set2_unflattened[5'h17];
  assign add_262878 = array_index_257817[11:0] + 12'hdab;
  assign sel_262880 = $signed({1'h0, add_262446}) < $signed({1'h0, sel_262448}) ? add_262446 : sel_262448;
  assign add_262882 = array_index_257820[11:0] + 12'hdab;
  assign sel_262884 = $signed({1'h0, add_262450}) < $signed({1'h0, sel_262452}) ? add_262450 : sel_262452;
  assign add_262896 = array_index_257955[11:2] + 10'h2b3;
  assign sel_262898 = $signed({1'h0, add_262464, array_index_257877[1:0]}) < $signed({1'h0, sel_262466}) ? {add_262464, array_index_257877[1:0]} : sel_262466;
  assign add_262900 = array_index_257958[11:2] + 10'h2b3;
  assign sel_262902 = $signed({1'h0, add_262468, array_index_257880[1:0]}) < $signed({1'h0, sel_262470}) ? {add_262468, array_index_257880[1:0]} : sel_262470;
  assign add_262912 = array_index_258159[11:1] + 11'h1e7;
  assign sel_262914 = $signed({1'h0, add_262480, array_index_258049[0]}) < $signed({1'h0, sel_262482}) ? {add_262480, array_index_258049[0]} : sel_262482;
  assign add_262916 = array_index_258162[11:1] + 11'h1e7;
  assign sel_262918 = $signed({1'h0, add_262484, array_index_258052[0]}) < $signed({1'h0, sel_262486}) ? {add_262484, array_index_258052[0]} : sel_262486;
  assign add_262928 = array_index_258427[11:0] + 12'h141;
  assign sel_262930 = $signed({1'h0, add_262496}) < $signed({1'h0, sel_262498}) ? add_262496 : sel_262498;
  assign add_262932 = array_index_258430[11:0] + 12'h141;
  assign sel_262934 = $signed({1'h0, add_262500}) < $signed({1'h0, sel_262502}) ? add_262500 : sel_262502;
  assign add_262936 = array_index_258585[11:1] + 11'h079;
  assign sel_262938 = $signed({1'h0, add_262504, array_index_258427[0]}) < $signed({1'h0, sel_262506}) ? {add_262504, array_index_258427[0]} : sel_262506;
  assign add_262940 = array_index_258588[11:1] + 11'h079;
  assign sel_262942 = $signed({1'h0, add_262508, array_index_258430[0]}) < $signed({1'h0, sel_262510}) ? {add_262508, array_index_258430[0]} : sel_262510;
  assign add_262944 = array_index_258761[11:0] + 12'h59d;
  assign sel_262946 = $signed({1'h0, add_262512}) < $signed({1'h0, sel_262514}) ? add_262512 : sel_262514;
  assign add_262948 = array_index_258764[11:0] + 12'h59d;
  assign sel_262950 = $signed({1'h0, add_262516}) < $signed({1'h0, sel_262518}) ? add_262516 : sel_262518;
  assign add_262952 = array_index_258957[11:0] + 12'ha6f;
  assign sel_262954 = $signed({1'h0, add_262520}) < $signed({1'h0, sel_262522}) ? add_262520 : sel_262522;
  assign add_262956 = array_index_258960[11:0] + 12'ha6f;
  assign sel_262958 = $signed({1'h0, add_262524}) < $signed({1'h0, sel_262526}) ? add_262524 : sel_262526;
  assign add_262960 = array_index_259171[11:1] + 11'h499;
  assign sel_262962 = $signed({1'h0, add_262528, array_index_258957[0]}) < $signed({1'h0, sel_262530}) ? {add_262528, array_index_258957[0]} : sel_262530;
  assign add_262964 = array_index_259174[11:1] + 11'h499;
  assign sel_262966 = $signed({1'h0, add_262532, array_index_258960[0]}) < $signed({1'h0, sel_262534}) ? {add_262532, array_index_258960[0]} : sel_262534;
  assign add_262968 = array_index_259401[11:1] + 11'h345;
  assign sel_262971 = $signed({1'h0, add_262536, array_index_259171[0]}) < $signed({1'h0, sel_262539}) ? {add_262536, array_index_259171[0]} : sel_262539;
  assign add_262973 = array_index_259404[11:1] + 11'h345;
  assign sel_262976 = $signed({1'h0, add_262541, array_index_259174[0]}) < $signed({1'h0, sel_262544}) ? {add_262541, array_index_259174[0]} : sel_262544;
  assign add_262978 = array_index_259647[11:0] + 12'h30f;
  assign sel_262980 = $signed({1'h0, add_262546}) < $signed({1'h0, sel_262548}) ? add_262546 : sel_262548;
  assign add_262982 = array_index_259650[11:0] + 12'h30f;
  assign sel_262984 = $signed({1'h0, add_262550}) < $signed({1'h0, sel_262552}) ? add_262550 : sel_262552;
  assign add_262986 = array_index_259911[11:0] + 12'hb55;
  assign sel_262988 = $signed({1'h0, add_262554}) < $signed({1'h0, sel_262556}) ? add_262554 : sel_262556;
  assign add_262990 = array_index_259914[11:0] + 12'hb55;
  assign sel_262992 = $signed({1'h0, add_262558}) < $signed({1'h0, sel_262560}) ? add_262558 : sel_262560;
  assign add_262994 = array_index_260195[11:0] + 12'h103;
  assign sel_262996 = $signed({1'h0, add_262562}) < $signed({1'h0, sel_262564}) ? add_262562 : sel_262564;
  assign add_262998 = array_index_260198[11:0] + 12'h103;
  assign sel_263000 = $signed({1'h0, add_262566}) < $signed({1'h0, sel_262568}) ? add_262566 : sel_262568;
  assign add_263002 = array_index_260507[11:0] + 12'hb01;
  assign sel_263004 = $signed({1'h0, add_262570}) < $signed({1'h0, sel_262572}) ? add_262570 : sel_262572;
  assign add_263006 = array_index_260510[11:0] + 12'hb01;
  assign sel_263008 = $signed({1'h0, add_262574}) < $signed({1'h0, sel_262576}) ? add_262574 : sel_262576;
  assign add_263010 = array_index_260845[11:0] + 12'h7b1;
  assign sel_263012 = $signed({1'h0, add_262578}) < $signed({1'h0, sel_262580}) ? add_262578 : sel_262580;
  assign add_263014 = array_index_260848[11:0] + 12'h7b1;
  assign sel_263016 = $signed({1'h0, add_262582}) < $signed({1'h0, sel_262584}) ? add_262582 : sel_262584;
  assign add_263018 = array_index_261207[11:0] + 12'h561;
  assign sel_263020 = $signed({1'h0, add_262586}) < $signed({1'h0, sel_262588}) ? add_262586 : sel_262588;
  assign add_263022 = array_index_261210[11:0] + 12'h561;
  assign sel_263024 = $signed({1'h0, add_262590}) < $signed({1'h0, sel_262592}) ? add_262590 : sel_262592;
  assign add_263026 = array_index_261595[11:2] + 10'h36b;
  assign sel_263028 = $signed({1'h0, add_262594, array_index_261207[1:0]}) < $signed({1'h0, sel_262596}) ? {add_262594, array_index_261207[1:0]} : sel_262596;
  assign add_263030 = array_index_261598[11:2] + 10'h36b;
  assign sel_263032 = $signed({1'h0, add_262598, array_index_261210[1:0]}) < $signed({1'h0, sel_262600}) ? {add_262598, array_index_261210[1:0]} : sel_262600;
  assign add_263034 = array_index_262007[11:2] + 10'h035;
  assign sel_263037 = $signed({1'h0, add_262602, array_index_261595[1:0]}) < $signed({1'h0, sel_262605}) ? {add_262602, array_index_261595[1:0]} : sel_262605;
  assign add_263039 = array_index_262010[11:2] + 10'h035;
  assign sel_263042 = $signed({1'h0, add_262607, array_index_261598[1:0]}) < $signed({1'h0, sel_262610}) ? {add_262607, array_index_261598[1:0]} : sel_262610;
  assign add_263044 = array_index_262439[11:0] + 12'hffb;
  assign sel_263046 = $signed({1'h0, add_262612}) < $signed({1'h0, sel_262614}) ? add_262612 : sel_262614;
  assign add_263048 = array_index_262442[11:0] + 12'hffb;
  assign sel_263050 = $signed({1'h0, add_262616}) < $signed({1'h0, sel_262618}) ? add_262616 : sel_262618;
  assign add_263062 = array_index_257877[11:2] + 10'h29b;
  assign sel_263064 = $signed({1'h0, add_262630, array_index_257817[1:0]}) < $signed({1'h0, sel_262632}) ? {add_262630, array_index_257817[1:0]} : sel_262632;
  assign add_263066 = array_index_257880[11:2] + 10'h29b;
  assign sel_263068 = $signed({1'h0, add_262634, array_index_257820[1:0]}) < $signed({1'h0, sel_262636}) ? {add_262634, array_index_257820[1:0]} : sel_262636;
  assign add_263078 = array_index_258049[11:0] + 12'h9cf;
  assign sel_263080 = $signed({1'h0, add_262646}) < $signed({1'h0, sel_262648}) ? add_262646 : sel_262648;
  assign add_263082 = array_index_258052[11:0] + 12'h9cf;
  assign sel_263084 = $signed({1'h0, add_262650}) < $signed({1'h0, sel_262652}) ? add_262650 : sel_262652;
  assign add_263094 = array_index_258285[11:0] + 12'h30b;
  assign sel_263096 = $signed({1'h0, add_262662}) < $signed({1'h0, sel_262664}) ? add_262662 : sel_262664;
  assign add_263098 = array_index_258288[11:0] + 12'h30b;
  assign sel_263100 = $signed({1'h0, add_262666}) < $signed({1'h0, sel_262668}) ? add_262666 : sel_262668;
  assign add_263169 = array_index_262871[11:0] + 12'h193;
  assign sel_263171 = $signed({1'h0, add_262737}) < $signed({1'h0, sel_262739}) ? add_262737 : sel_262739;
  assign add_263174 = array_index_262874[11:0] + 12'h193;
  assign sel_263176 = $signed({1'h0, add_262742}) < $signed({1'h0, sel_262744}) ? add_262742 : sel_262744;
  assign add_263186 = array_index_257955[11:0] + 12'hc05;
  assign sel_263188 = $signed({1'h0, add_262754}) < $signed({1'h0, sel_262756}) ? add_262754 : sel_262756;
  assign add_263190 = array_index_257958[11:0] + 12'hc05;
  assign sel_263192 = $signed({1'h0, add_262758}) < $signed({1'h0, sel_262760}) ? add_262758 : sel_262760;
  assign add_263204 = array_index_258159[11:0] + 12'h83f;
  assign sel_263206 = $signed({1'h0, add_262772}) < $signed({1'h0, sel_262774}) ? add_262772 : sel_262774;
  assign add_263208 = array_index_258162[11:0] + 12'h83f;
  assign sel_263210 = $signed({1'h0, add_262776}) < $signed({1'h0, sel_262778}) ? add_262776 : sel_262778;
  assign add_263222 = array_index_258427[11:1] + 11'h7b5;
  assign sel_263224 = $signed({1'h0, add_262790, array_index_258285[0]}) < $signed({1'h0, sel_262792}) ? {add_262790, array_index_258285[0]} : sel_262792;
  assign add_263226 = array_index_258430[11:1] + 11'h7b5;
  assign sel_263228 = $signed({1'h0, add_262794, array_index_258288[0]}) < $signed({1'h0, sel_262796}) ? {add_262794, array_index_258288[0]} : sel_262796;
  assign array_index_263303 = set1_unflattened[5'h18];
  assign array_index_263306 = set2_unflattened[5'h18];
  assign add_263310 = array_index_257877[11:0] + 12'hdab;
  assign sel_263312 = $signed({1'h0, add_262878}) < $signed({1'h0, sel_262880}) ? add_262878 : sel_262880;
  assign add_263314 = array_index_257880[11:0] + 12'hdab;
  assign sel_263316 = $signed({1'h0, add_262882}) < $signed({1'h0, sel_262884}) ? add_262882 : sel_262884;
  assign add_263328 = array_index_258049[11:2] + 10'h2b3;
  assign sel_263330 = $signed({1'h0, add_262896, array_index_257955[1:0]}) < $signed({1'h0, sel_262898}) ? {add_262896, array_index_257955[1:0]} : sel_262898;
  assign add_263332 = array_index_258052[11:2] + 10'h2b3;
  assign sel_263334 = $signed({1'h0, add_262900, array_index_257958[1:0]}) < $signed({1'h0, sel_262902}) ? {add_262900, array_index_257958[1:0]} : sel_262902;
  assign add_263344 = array_index_258285[11:1] + 11'h1e7;
  assign sel_263346 = $signed({1'h0, add_262912, array_index_258159[0]}) < $signed({1'h0, sel_262914}) ? {add_262912, array_index_258159[0]} : sel_262914;
  assign add_263348 = array_index_258288[11:1] + 11'h1e7;
  assign sel_263350 = $signed({1'h0, add_262916, array_index_258162[0]}) < $signed({1'h0, sel_262918}) ? {add_262916, array_index_258162[0]} : sel_262918;
  assign add_263360 = array_index_258585[11:0] + 12'h141;
  assign sel_263362 = $signed({1'h0, add_262928}) < $signed({1'h0, sel_262930}) ? add_262928 : sel_262930;
  assign add_263364 = array_index_258588[11:0] + 12'h141;
  assign sel_263366 = $signed({1'h0, add_262932}) < $signed({1'h0, sel_262934}) ? add_262932 : sel_262934;
  assign add_263368 = array_index_258761[11:1] + 11'h079;
  assign sel_263370 = $signed({1'h0, add_262936, array_index_258585[0]}) < $signed({1'h0, sel_262938}) ? {add_262936, array_index_258585[0]} : sel_262938;
  assign add_263372 = array_index_258764[11:1] + 11'h079;
  assign sel_263374 = $signed({1'h0, add_262940, array_index_258588[0]}) < $signed({1'h0, sel_262942}) ? {add_262940, array_index_258588[0]} : sel_262942;
  assign add_263376 = array_index_258957[11:0] + 12'h59d;
  assign sel_263378 = $signed({1'h0, add_262944}) < $signed({1'h0, sel_262946}) ? add_262944 : sel_262946;
  assign add_263380 = array_index_258960[11:0] + 12'h59d;
  assign sel_263382 = $signed({1'h0, add_262948}) < $signed({1'h0, sel_262950}) ? add_262948 : sel_262950;
  assign add_263384 = array_index_259171[11:0] + 12'ha6f;
  assign sel_263386 = $signed({1'h0, add_262952}) < $signed({1'h0, sel_262954}) ? add_262952 : sel_262954;
  assign add_263388 = array_index_259174[11:0] + 12'ha6f;
  assign sel_263390 = $signed({1'h0, add_262956}) < $signed({1'h0, sel_262958}) ? add_262956 : sel_262958;
  assign add_263392 = array_index_259401[11:1] + 11'h499;
  assign sel_263394 = $signed({1'h0, add_262960, array_index_259171[0]}) < $signed({1'h0, sel_262962}) ? {add_262960, array_index_259171[0]} : sel_262962;
  assign add_263396 = array_index_259404[11:1] + 11'h499;
  assign sel_263398 = $signed({1'h0, add_262964, array_index_259174[0]}) < $signed({1'h0, sel_262966}) ? {add_262964, array_index_259174[0]} : sel_262966;
  assign add_263400 = array_index_259647[11:1] + 11'h345;
  assign sel_263403 = $signed({1'h0, add_262968, array_index_259401[0]}) < $signed({1'h0, sel_262971}) ? {add_262968, array_index_259401[0]} : sel_262971;
  assign add_263405 = array_index_259650[11:1] + 11'h345;
  assign sel_263408 = $signed({1'h0, add_262973, array_index_259404[0]}) < $signed({1'h0, sel_262976}) ? {add_262973, array_index_259404[0]} : sel_262976;
  assign add_263410 = array_index_259911[11:0] + 12'h30f;
  assign sel_263412 = $signed({1'h0, add_262978}) < $signed({1'h0, sel_262980}) ? add_262978 : sel_262980;
  assign add_263414 = array_index_259914[11:0] + 12'h30f;
  assign sel_263416 = $signed({1'h0, add_262982}) < $signed({1'h0, sel_262984}) ? add_262982 : sel_262984;
  assign add_263418 = array_index_260195[11:0] + 12'hb55;
  assign sel_263420 = $signed({1'h0, add_262986}) < $signed({1'h0, sel_262988}) ? add_262986 : sel_262988;
  assign add_263422 = array_index_260198[11:0] + 12'hb55;
  assign sel_263424 = $signed({1'h0, add_262990}) < $signed({1'h0, sel_262992}) ? add_262990 : sel_262992;
  assign add_263426 = array_index_260507[11:0] + 12'h103;
  assign sel_263428 = $signed({1'h0, add_262994}) < $signed({1'h0, sel_262996}) ? add_262994 : sel_262996;
  assign add_263430 = array_index_260510[11:0] + 12'h103;
  assign sel_263432 = $signed({1'h0, add_262998}) < $signed({1'h0, sel_263000}) ? add_262998 : sel_263000;
  assign add_263434 = array_index_260845[11:0] + 12'hb01;
  assign sel_263436 = $signed({1'h0, add_263002}) < $signed({1'h0, sel_263004}) ? add_263002 : sel_263004;
  assign add_263438 = array_index_260848[11:0] + 12'hb01;
  assign sel_263440 = $signed({1'h0, add_263006}) < $signed({1'h0, sel_263008}) ? add_263006 : sel_263008;
  assign add_263442 = array_index_261207[11:0] + 12'h7b1;
  assign sel_263444 = $signed({1'h0, add_263010}) < $signed({1'h0, sel_263012}) ? add_263010 : sel_263012;
  assign add_263446 = array_index_261210[11:0] + 12'h7b1;
  assign sel_263448 = $signed({1'h0, add_263014}) < $signed({1'h0, sel_263016}) ? add_263014 : sel_263016;
  assign add_263450 = array_index_261595[11:0] + 12'h561;
  assign sel_263452 = $signed({1'h0, add_263018}) < $signed({1'h0, sel_263020}) ? add_263018 : sel_263020;
  assign add_263454 = array_index_261598[11:0] + 12'h561;
  assign sel_263456 = $signed({1'h0, add_263022}) < $signed({1'h0, sel_263024}) ? add_263022 : sel_263024;
  assign add_263458 = array_index_262007[11:2] + 10'h36b;
  assign sel_263460 = $signed({1'h0, add_263026, array_index_261595[1:0]}) < $signed({1'h0, sel_263028}) ? {add_263026, array_index_261595[1:0]} : sel_263028;
  assign add_263462 = array_index_262010[11:2] + 10'h36b;
  assign sel_263464 = $signed({1'h0, add_263030, array_index_261598[1:0]}) < $signed({1'h0, sel_263032}) ? {add_263030, array_index_261598[1:0]} : sel_263032;
  assign add_263466 = array_index_262439[11:2] + 10'h035;
  assign sel_263469 = $signed({1'h0, add_263034, array_index_262007[1:0]}) < $signed({1'h0, sel_263037}) ? {add_263034, array_index_262007[1:0]} : sel_263037;
  assign add_263471 = array_index_262442[11:2] + 10'h035;
  assign sel_263474 = $signed({1'h0, add_263039, array_index_262010[1:0]}) < $signed({1'h0, sel_263042}) ? {add_263039, array_index_262010[1:0]} : sel_263042;
  assign add_263476 = array_index_262871[11:0] + 12'hffb;
  assign sel_263478 = $signed({1'h0, add_263044}) < $signed({1'h0, sel_263046}) ? add_263044 : sel_263046;
  assign add_263480 = array_index_262874[11:0] + 12'hffb;
  assign sel_263482 = $signed({1'h0, add_263048}) < $signed({1'h0, sel_263050}) ? add_263048 : sel_263050;
  assign add_263494 = array_index_257955[11:2] + 10'h29b;
  assign sel_263496 = $signed({1'h0, add_263062, array_index_257877[1:0]}) < $signed({1'h0, sel_263064}) ? {add_263062, array_index_257877[1:0]} : sel_263064;
  assign add_263498 = array_index_257958[11:2] + 10'h29b;
  assign sel_263500 = $signed({1'h0, add_263066, array_index_257880[1:0]}) < $signed({1'h0, sel_263068}) ? {add_263066, array_index_257880[1:0]} : sel_263068;
  assign add_263510 = array_index_258159[11:0] + 12'h9cf;
  assign sel_263512 = $signed({1'h0, add_263078}) < $signed({1'h0, sel_263080}) ? add_263078 : sel_263080;
  assign add_263514 = array_index_258162[11:0] + 12'h9cf;
  assign sel_263516 = $signed({1'h0, add_263082}) < $signed({1'h0, sel_263084}) ? add_263082 : sel_263084;
  assign add_263526 = array_index_258427[11:0] + 12'h30b;
  assign sel_263528 = $signed({1'h0, add_263094}) < $signed({1'h0, sel_263096}) ? add_263094 : sel_263096;
  assign add_263530 = array_index_258430[11:0] + 12'h30b;
  assign sel_263532 = $signed({1'h0, add_263098}) < $signed({1'h0, sel_263100}) ? add_263098 : sel_263100;
  assign add_263601 = array_index_263303[11:0] + 12'h193;
  assign sel_263603 = $signed({1'h0, add_263169}) < $signed({1'h0, sel_263171}) ? add_263169 : sel_263171;
  assign add_263606 = array_index_263306[11:0] + 12'h193;
  assign sel_263608 = $signed({1'h0, add_263174}) < $signed({1'h0, sel_263176}) ? add_263174 : sel_263176;
  assign add_263618 = array_index_258049[11:0] + 12'hc05;
  assign sel_263620 = $signed({1'h0, add_263186}) < $signed({1'h0, sel_263188}) ? add_263186 : sel_263188;
  assign add_263622 = array_index_258052[11:0] + 12'hc05;
  assign sel_263624 = $signed({1'h0, add_263190}) < $signed({1'h0, sel_263192}) ? add_263190 : sel_263192;
  assign add_263636 = array_index_258285[11:0] + 12'h83f;
  assign sel_263638 = $signed({1'h0, add_263204}) < $signed({1'h0, sel_263206}) ? add_263204 : sel_263206;
  assign add_263640 = array_index_258288[11:0] + 12'h83f;
  assign sel_263642 = $signed({1'h0, add_263208}) < $signed({1'h0, sel_263210}) ? add_263208 : sel_263210;
  assign add_263654 = array_index_258585[11:1] + 11'h7b5;
  assign sel_263656 = $signed({1'h0, add_263222, array_index_258427[0]}) < $signed({1'h0, sel_263224}) ? {add_263222, array_index_258427[0]} : sel_263224;
  assign add_263658 = array_index_258588[11:1] + 11'h7b5;
  assign sel_263660 = $signed({1'h0, add_263226, array_index_258430[0]}) < $signed({1'h0, sel_263228}) ? {add_263226, array_index_258430[0]} : sel_263228;
  assign array_index_263735 = set1_unflattened[5'h19];
  assign array_index_263738 = set2_unflattened[5'h19];
  assign add_263742 = array_index_257955[11:0] + 12'hdab;
  assign sel_263744 = $signed({1'h0, add_263310}) < $signed({1'h0, sel_263312}) ? add_263310 : sel_263312;
  assign add_263746 = array_index_257958[11:0] + 12'hdab;
  assign sel_263748 = $signed({1'h0, add_263314}) < $signed({1'h0, sel_263316}) ? add_263314 : sel_263316;
  assign add_263760 = array_index_258159[11:2] + 10'h2b3;
  assign sel_263762 = $signed({1'h0, add_263328, array_index_258049[1:0]}) < $signed({1'h0, sel_263330}) ? {add_263328, array_index_258049[1:0]} : sel_263330;
  assign add_263764 = array_index_258162[11:2] + 10'h2b3;
  assign sel_263766 = $signed({1'h0, add_263332, array_index_258052[1:0]}) < $signed({1'h0, sel_263334}) ? {add_263332, array_index_258052[1:0]} : sel_263334;
  assign add_263776 = array_index_258427[11:1] + 11'h1e7;
  assign sel_263778 = $signed({1'h0, add_263344, array_index_258285[0]}) < $signed({1'h0, sel_263346}) ? {add_263344, array_index_258285[0]} : sel_263346;
  assign add_263780 = array_index_258430[11:1] + 11'h1e7;
  assign sel_263782 = $signed({1'h0, add_263348, array_index_258288[0]}) < $signed({1'h0, sel_263350}) ? {add_263348, array_index_258288[0]} : sel_263350;
  assign add_263792 = array_index_258761[11:0] + 12'h141;
  assign sel_263794 = $signed({1'h0, add_263360}) < $signed({1'h0, sel_263362}) ? add_263360 : sel_263362;
  assign add_263796 = array_index_258764[11:0] + 12'h141;
  assign sel_263798 = $signed({1'h0, add_263364}) < $signed({1'h0, sel_263366}) ? add_263364 : sel_263366;
  assign add_263800 = array_index_258957[11:1] + 11'h079;
  assign sel_263802 = $signed({1'h0, add_263368, array_index_258761[0]}) < $signed({1'h0, sel_263370}) ? {add_263368, array_index_258761[0]} : sel_263370;
  assign add_263804 = array_index_258960[11:1] + 11'h079;
  assign sel_263806 = $signed({1'h0, add_263372, array_index_258764[0]}) < $signed({1'h0, sel_263374}) ? {add_263372, array_index_258764[0]} : sel_263374;
  assign add_263808 = array_index_259171[11:0] + 12'h59d;
  assign sel_263810 = $signed({1'h0, add_263376}) < $signed({1'h0, sel_263378}) ? add_263376 : sel_263378;
  assign add_263812 = array_index_259174[11:0] + 12'h59d;
  assign sel_263814 = $signed({1'h0, add_263380}) < $signed({1'h0, sel_263382}) ? add_263380 : sel_263382;
  assign add_263816 = array_index_259401[11:0] + 12'ha6f;
  assign sel_263818 = $signed({1'h0, add_263384}) < $signed({1'h0, sel_263386}) ? add_263384 : sel_263386;
  assign add_263820 = array_index_259404[11:0] + 12'ha6f;
  assign sel_263822 = $signed({1'h0, add_263388}) < $signed({1'h0, sel_263390}) ? add_263388 : sel_263390;
  assign add_263824 = array_index_259647[11:1] + 11'h499;
  assign sel_263826 = $signed({1'h0, add_263392, array_index_259401[0]}) < $signed({1'h0, sel_263394}) ? {add_263392, array_index_259401[0]} : sel_263394;
  assign add_263828 = array_index_259650[11:1] + 11'h499;
  assign sel_263830 = $signed({1'h0, add_263396, array_index_259404[0]}) < $signed({1'h0, sel_263398}) ? {add_263396, array_index_259404[0]} : sel_263398;
  assign add_263832 = array_index_259911[11:1] + 11'h345;
  assign sel_263835 = $signed({1'h0, add_263400, array_index_259647[0]}) < $signed({1'h0, sel_263403}) ? {add_263400, array_index_259647[0]} : sel_263403;
  assign add_263837 = array_index_259914[11:1] + 11'h345;
  assign sel_263840 = $signed({1'h0, add_263405, array_index_259650[0]}) < $signed({1'h0, sel_263408}) ? {add_263405, array_index_259650[0]} : sel_263408;
  assign add_263842 = array_index_260195[11:0] + 12'h30f;
  assign sel_263844 = $signed({1'h0, add_263410}) < $signed({1'h0, sel_263412}) ? add_263410 : sel_263412;
  assign add_263846 = array_index_260198[11:0] + 12'h30f;
  assign sel_263848 = $signed({1'h0, add_263414}) < $signed({1'h0, sel_263416}) ? add_263414 : sel_263416;
  assign add_263850 = array_index_260507[11:0] + 12'hb55;
  assign sel_263852 = $signed({1'h0, add_263418}) < $signed({1'h0, sel_263420}) ? add_263418 : sel_263420;
  assign add_263854 = array_index_260510[11:0] + 12'hb55;
  assign sel_263856 = $signed({1'h0, add_263422}) < $signed({1'h0, sel_263424}) ? add_263422 : sel_263424;
  assign add_263858 = array_index_260845[11:0] + 12'h103;
  assign sel_263860 = $signed({1'h0, add_263426}) < $signed({1'h0, sel_263428}) ? add_263426 : sel_263428;
  assign add_263862 = array_index_260848[11:0] + 12'h103;
  assign sel_263864 = $signed({1'h0, add_263430}) < $signed({1'h0, sel_263432}) ? add_263430 : sel_263432;
  assign add_263866 = array_index_261207[11:0] + 12'hb01;
  assign sel_263868 = $signed({1'h0, add_263434}) < $signed({1'h0, sel_263436}) ? add_263434 : sel_263436;
  assign add_263870 = array_index_261210[11:0] + 12'hb01;
  assign sel_263872 = $signed({1'h0, add_263438}) < $signed({1'h0, sel_263440}) ? add_263438 : sel_263440;
  assign add_263874 = array_index_261595[11:0] + 12'h7b1;
  assign sel_263876 = $signed({1'h0, add_263442}) < $signed({1'h0, sel_263444}) ? add_263442 : sel_263444;
  assign add_263878 = array_index_261598[11:0] + 12'h7b1;
  assign sel_263880 = $signed({1'h0, add_263446}) < $signed({1'h0, sel_263448}) ? add_263446 : sel_263448;
  assign add_263882 = array_index_262007[11:0] + 12'h561;
  assign sel_263884 = $signed({1'h0, add_263450}) < $signed({1'h0, sel_263452}) ? add_263450 : sel_263452;
  assign add_263886 = array_index_262010[11:0] + 12'h561;
  assign sel_263888 = $signed({1'h0, add_263454}) < $signed({1'h0, sel_263456}) ? add_263454 : sel_263456;
  assign add_263890 = array_index_262439[11:2] + 10'h36b;
  assign sel_263892 = $signed({1'h0, add_263458, array_index_262007[1:0]}) < $signed({1'h0, sel_263460}) ? {add_263458, array_index_262007[1:0]} : sel_263460;
  assign add_263894 = array_index_262442[11:2] + 10'h36b;
  assign sel_263896 = $signed({1'h0, add_263462, array_index_262010[1:0]}) < $signed({1'h0, sel_263464}) ? {add_263462, array_index_262010[1:0]} : sel_263464;
  assign add_263898 = array_index_262871[11:2] + 10'h035;
  assign sel_263901 = $signed({1'h0, add_263466, array_index_262439[1:0]}) < $signed({1'h0, sel_263469}) ? {add_263466, array_index_262439[1:0]} : sel_263469;
  assign add_263903 = array_index_262874[11:2] + 10'h035;
  assign sel_263906 = $signed({1'h0, add_263471, array_index_262442[1:0]}) < $signed({1'h0, sel_263474}) ? {add_263471, array_index_262442[1:0]} : sel_263474;
  assign add_263908 = array_index_263303[11:0] + 12'hffb;
  assign sel_263910 = $signed({1'h0, add_263476}) < $signed({1'h0, sel_263478}) ? add_263476 : sel_263478;
  assign add_263912 = array_index_263306[11:0] + 12'hffb;
  assign sel_263914 = $signed({1'h0, add_263480}) < $signed({1'h0, sel_263482}) ? add_263480 : sel_263482;
  assign add_263926 = array_index_258049[11:2] + 10'h29b;
  assign sel_263928 = $signed({1'h0, add_263494, array_index_257955[1:0]}) < $signed({1'h0, sel_263496}) ? {add_263494, array_index_257955[1:0]} : sel_263496;
  assign add_263930 = array_index_258052[11:2] + 10'h29b;
  assign sel_263932 = $signed({1'h0, add_263498, array_index_257958[1:0]}) < $signed({1'h0, sel_263500}) ? {add_263498, array_index_257958[1:0]} : sel_263500;
  assign add_263942 = array_index_258285[11:0] + 12'h9cf;
  assign sel_263944 = $signed({1'h0, add_263510}) < $signed({1'h0, sel_263512}) ? add_263510 : sel_263512;
  assign add_263946 = array_index_258288[11:0] + 12'h9cf;
  assign sel_263948 = $signed({1'h0, add_263514}) < $signed({1'h0, sel_263516}) ? add_263514 : sel_263516;
  assign add_263958 = array_index_258585[11:0] + 12'h30b;
  assign sel_263960 = $signed({1'h0, add_263526}) < $signed({1'h0, sel_263528}) ? add_263526 : sel_263528;
  assign add_263962 = array_index_258588[11:0] + 12'h30b;
  assign sel_263964 = $signed({1'h0, add_263530}) < $signed({1'h0, sel_263532}) ? add_263530 : sel_263532;
  assign add_264033 = array_index_263735[11:0] + 12'h193;
  assign sel_264035 = $signed({1'h0, add_263601}) < $signed({1'h0, sel_263603}) ? add_263601 : sel_263603;
  assign add_264038 = array_index_263738[11:0] + 12'h193;
  assign sel_264040 = $signed({1'h0, add_263606}) < $signed({1'h0, sel_263608}) ? add_263606 : sel_263608;
  assign add_264050 = array_index_258159[11:0] + 12'hc05;
  assign sel_264052 = $signed({1'h0, add_263618}) < $signed({1'h0, sel_263620}) ? add_263618 : sel_263620;
  assign add_264054 = array_index_258162[11:0] + 12'hc05;
  assign sel_264056 = $signed({1'h0, add_263622}) < $signed({1'h0, sel_263624}) ? add_263622 : sel_263624;
  assign add_264068 = array_index_258427[11:0] + 12'h83f;
  assign sel_264070 = $signed({1'h0, add_263636}) < $signed({1'h0, sel_263638}) ? add_263636 : sel_263638;
  assign add_264072 = array_index_258430[11:0] + 12'h83f;
  assign sel_264074 = $signed({1'h0, add_263640}) < $signed({1'h0, sel_263642}) ? add_263640 : sel_263642;
  assign add_264086 = array_index_258761[11:1] + 11'h7b5;
  assign sel_264088 = $signed({1'h0, add_263654, array_index_258585[0]}) < $signed({1'h0, sel_263656}) ? {add_263654, array_index_258585[0]} : sel_263656;
  assign add_264090 = array_index_258764[11:1] + 11'h7b5;
  assign sel_264092 = $signed({1'h0, add_263658, array_index_258588[0]}) < $signed({1'h0, sel_263660}) ? {add_263658, array_index_258588[0]} : sel_263660;
  assign array_index_264167 = set1_unflattened[5'h1a];
  assign array_index_264170 = set2_unflattened[5'h1a];
  assign add_264174 = array_index_258049[11:0] + 12'hdab;
  assign sel_264176 = $signed({1'h0, add_263742}) < $signed({1'h0, sel_263744}) ? add_263742 : sel_263744;
  assign add_264178 = array_index_258052[11:0] + 12'hdab;
  assign sel_264180 = $signed({1'h0, add_263746}) < $signed({1'h0, sel_263748}) ? add_263746 : sel_263748;
  assign add_264192 = array_index_258285[11:2] + 10'h2b3;
  assign sel_264194 = $signed({1'h0, add_263760, array_index_258159[1:0]}) < $signed({1'h0, sel_263762}) ? {add_263760, array_index_258159[1:0]} : sel_263762;
  assign add_264196 = array_index_258288[11:2] + 10'h2b3;
  assign sel_264198 = $signed({1'h0, add_263764, array_index_258162[1:0]}) < $signed({1'h0, sel_263766}) ? {add_263764, array_index_258162[1:0]} : sel_263766;
  assign add_264208 = array_index_258585[11:1] + 11'h1e7;
  assign sel_264210 = $signed({1'h0, add_263776, array_index_258427[0]}) < $signed({1'h0, sel_263778}) ? {add_263776, array_index_258427[0]} : sel_263778;
  assign add_264212 = array_index_258588[11:1] + 11'h1e7;
  assign sel_264214 = $signed({1'h0, add_263780, array_index_258430[0]}) < $signed({1'h0, sel_263782}) ? {add_263780, array_index_258430[0]} : sel_263782;
  assign add_264224 = array_index_258957[11:0] + 12'h141;
  assign sel_264226 = $signed({1'h0, add_263792}) < $signed({1'h0, sel_263794}) ? add_263792 : sel_263794;
  assign add_264228 = array_index_258960[11:0] + 12'h141;
  assign sel_264230 = $signed({1'h0, add_263796}) < $signed({1'h0, sel_263798}) ? add_263796 : sel_263798;
  assign add_264232 = array_index_259171[11:1] + 11'h079;
  assign sel_264234 = $signed({1'h0, add_263800, array_index_258957[0]}) < $signed({1'h0, sel_263802}) ? {add_263800, array_index_258957[0]} : sel_263802;
  assign add_264236 = array_index_259174[11:1] + 11'h079;
  assign sel_264238 = $signed({1'h0, add_263804, array_index_258960[0]}) < $signed({1'h0, sel_263806}) ? {add_263804, array_index_258960[0]} : sel_263806;
  assign add_264240 = array_index_259401[11:0] + 12'h59d;
  assign sel_264242 = $signed({1'h0, add_263808}) < $signed({1'h0, sel_263810}) ? add_263808 : sel_263810;
  assign add_264244 = array_index_259404[11:0] + 12'h59d;
  assign sel_264246 = $signed({1'h0, add_263812}) < $signed({1'h0, sel_263814}) ? add_263812 : sel_263814;
  assign add_264248 = array_index_259647[11:0] + 12'ha6f;
  assign sel_264250 = $signed({1'h0, add_263816}) < $signed({1'h0, sel_263818}) ? add_263816 : sel_263818;
  assign add_264252 = array_index_259650[11:0] + 12'ha6f;
  assign sel_264254 = $signed({1'h0, add_263820}) < $signed({1'h0, sel_263822}) ? add_263820 : sel_263822;
  assign add_264256 = array_index_259911[11:1] + 11'h499;
  assign sel_264258 = $signed({1'h0, add_263824, array_index_259647[0]}) < $signed({1'h0, sel_263826}) ? {add_263824, array_index_259647[0]} : sel_263826;
  assign add_264260 = array_index_259914[11:1] + 11'h499;
  assign sel_264262 = $signed({1'h0, add_263828, array_index_259650[0]}) < $signed({1'h0, sel_263830}) ? {add_263828, array_index_259650[0]} : sel_263830;
  assign add_264264 = array_index_260195[11:1] + 11'h345;
  assign sel_264267 = $signed({1'h0, add_263832, array_index_259911[0]}) < $signed({1'h0, sel_263835}) ? {add_263832, array_index_259911[0]} : sel_263835;
  assign add_264269 = array_index_260198[11:1] + 11'h345;
  assign sel_264272 = $signed({1'h0, add_263837, array_index_259914[0]}) < $signed({1'h0, sel_263840}) ? {add_263837, array_index_259914[0]} : sel_263840;
  assign add_264274 = array_index_260507[11:0] + 12'h30f;
  assign sel_264276 = $signed({1'h0, add_263842}) < $signed({1'h0, sel_263844}) ? add_263842 : sel_263844;
  assign add_264278 = array_index_260510[11:0] + 12'h30f;
  assign sel_264280 = $signed({1'h0, add_263846}) < $signed({1'h0, sel_263848}) ? add_263846 : sel_263848;
  assign add_264282 = array_index_260845[11:0] + 12'hb55;
  assign sel_264284 = $signed({1'h0, add_263850}) < $signed({1'h0, sel_263852}) ? add_263850 : sel_263852;
  assign add_264286 = array_index_260848[11:0] + 12'hb55;
  assign sel_264288 = $signed({1'h0, add_263854}) < $signed({1'h0, sel_263856}) ? add_263854 : sel_263856;
  assign add_264290 = array_index_261207[11:0] + 12'h103;
  assign sel_264292 = $signed({1'h0, add_263858}) < $signed({1'h0, sel_263860}) ? add_263858 : sel_263860;
  assign add_264294 = array_index_261210[11:0] + 12'h103;
  assign sel_264296 = $signed({1'h0, add_263862}) < $signed({1'h0, sel_263864}) ? add_263862 : sel_263864;
  assign add_264298 = array_index_261595[11:0] + 12'hb01;
  assign sel_264300 = $signed({1'h0, add_263866}) < $signed({1'h0, sel_263868}) ? add_263866 : sel_263868;
  assign add_264302 = array_index_261598[11:0] + 12'hb01;
  assign sel_264304 = $signed({1'h0, add_263870}) < $signed({1'h0, sel_263872}) ? add_263870 : sel_263872;
  assign add_264306 = array_index_262007[11:0] + 12'h7b1;
  assign sel_264308 = $signed({1'h0, add_263874}) < $signed({1'h0, sel_263876}) ? add_263874 : sel_263876;
  assign add_264310 = array_index_262010[11:0] + 12'h7b1;
  assign sel_264312 = $signed({1'h0, add_263878}) < $signed({1'h0, sel_263880}) ? add_263878 : sel_263880;
  assign add_264314 = array_index_262439[11:0] + 12'h561;
  assign sel_264316 = $signed({1'h0, add_263882}) < $signed({1'h0, sel_263884}) ? add_263882 : sel_263884;
  assign add_264318 = array_index_262442[11:0] + 12'h561;
  assign sel_264320 = $signed({1'h0, add_263886}) < $signed({1'h0, sel_263888}) ? add_263886 : sel_263888;
  assign add_264322 = array_index_262871[11:2] + 10'h36b;
  assign sel_264324 = $signed({1'h0, add_263890, array_index_262439[1:0]}) < $signed({1'h0, sel_263892}) ? {add_263890, array_index_262439[1:0]} : sel_263892;
  assign add_264326 = array_index_262874[11:2] + 10'h36b;
  assign sel_264328 = $signed({1'h0, add_263894, array_index_262442[1:0]}) < $signed({1'h0, sel_263896}) ? {add_263894, array_index_262442[1:0]} : sel_263896;
  assign add_264330 = array_index_263303[11:2] + 10'h035;
  assign sel_264333 = $signed({1'h0, add_263898, array_index_262871[1:0]}) < $signed({1'h0, sel_263901}) ? {add_263898, array_index_262871[1:0]} : sel_263901;
  assign add_264335 = array_index_263306[11:2] + 10'h035;
  assign sel_264338 = $signed({1'h0, add_263903, array_index_262874[1:0]}) < $signed({1'h0, sel_263906}) ? {add_263903, array_index_262874[1:0]} : sel_263906;
  assign add_264340 = array_index_263735[11:0] + 12'hffb;
  assign sel_264342 = $signed({1'h0, add_263908}) < $signed({1'h0, sel_263910}) ? add_263908 : sel_263910;
  assign add_264344 = array_index_263738[11:0] + 12'hffb;
  assign sel_264346 = $signed({1'h0, add_263912}) < $signed({1'h0, sel_263914}) ? add_263912 : sel_263914;
  assign add_264358 = array_index_258159[11:2] + 10'h29b;
  assign sel_264360 = $signed({1'h0, add_263926, array_index_258049[1:0]}) < $signed({1'h0, sel_263928}) ? {add_263926, array_index_258049[1:0]} : sel_263928;
  assign add_264362 = array_index_258162[11:2] + 10'h29b;
  assign sel_264364 = $signed({1'h0, add_263930, array_index_258052[1:0]}) < $signed({1'h0, sel_263932}) ? {add_263930, array_index_258052[1:0]} : sel_263932;
  assign add_264374 = array_index_258427[11:0] + 12'h9cf;
  assign sel_264376 = $signed({1'h0, add_263942}) < $signed({1'h0, sel_263944}) ? add_263942 : sel_263944;
  assign add_264378 = array_index_258430[11:0] + 12'h9cf;
  assign sel_264380 = $signed({1'h0, add_263946}) < $signed({1'h0, sel_263948}) ? add_263946 : sel_263948;
  assign add_264390 = array_index_258761[11:0] + 12'h30b;
  assign sel_264392 = $signed({1'h0, add_263958}) < $signed({1'h0, sel_263960}) ? add_263958 : sel_263960;
  assign add_264394 = array_index_258764[11:0] + 12'h30b;
  assign sel_264396 = $signed({1'h0, add_263962}) < $signed({1'h0, sel_263964}) ? add_263962 : sel_263964;
  assign add_264465 = array_index_264167[11:0] + 12'h193;
  assign sel_264467 = $signed({1'h0, add_264033}) < $signed({1'h0, sel_264035}) ? add_264033 : sel_264035;
  assign add_264470 = array_index_264170[11:0] + 12'h193;
  assign sel_264472 = $signed({1'h0, add_264038}) < $signed({1'h0, sel_264040}) ? add_264038 : sel_264040;
  assign add_264482 = array_index_258285[11:0] + 12'hc05;
  assign sel_264484 = $signed({1'h0, add_264050}) < $signed({1'h0, sel_264052}) ? add_264050 : sel_264052;
  assign add_264486 = array_index_258288[11:0] + 12'hc05;
  assign sel_264488 = $signed({1'h0, add_264054}) < $signed({1'h0, sel_264056}) ? add_264054 : sel_264056;
  assign add_264500 = array_index_258585[11:0] + 12'h83f;
  assign sel_264502 = $signed({1'h0, add_264068}) < $signed({1'h0, sel_264070}) ? add_264068 : sel_264070;
  assign add_264504 = array_index_258588[11:0] + 12'h83f;
  assign sel_264506 = $signed({1'h0, add_264072}) < $signed({1'h0, sel_264074}) ? add_264072 : sel_264074;
  assign add_264518 = array_index_258957[11:1] + 11'h7b5;
  assign sel_264520 = $signed({1'h0, add_264086, array_index_258761[0]}) < $signed({1'h0, sel_264088}) ? {add_264086, array_index_258761[0]} : sel_264088;
  assign add_264522 = array_index_258960[11:1] + 11'h7b5;
  assign sel_264524 = $signed({1'h0, add_264090, array_index_258764[0]}) < $signed({1'h0, sel_264092}) ? {add_264090, array_index_258764[0]} : sel_264092;
  assign array_index_264599 = set1_unflattened[5'h1b];
  assign array_index_264602 = set2_unflattened[5'h1b];
  assign add_264606 = array_index_258159[11:0] + 12'hdab;
  assign sel_264608 = $signed({1'h0, add_264174}) < $signed({1'h0, sel_264176}) ? add_264174 : sel_264176;
  assign add_264610 = array_index_258162[11:0] + 12'hdab;
  assign sel_264612 = $signed({1'h0, add_264178}) < $signed({1'h0, sel_264180}) ? add_264178 : sel_264180;
  assign add_264624 = array_index_258427[11:2] + 10'h2b3;
  assign sel_264626 = $signed({1'h0, add_264192, array_index_258285[1:0]}) < $signed({1'h0, sel_264194}) ? {add_264192, array_index_258285[1:0]} : sel_264194;
  assign add_264628 = array_index_258430[11:2] + 10'h2b3;
  assign sel_264630 = $signed({1'h0, add_264196, array_index_258288[1:0]}) < $signed({1'h0, sel_264198}) ? {add_264196, array_index_258288[1:0]} : sel_264198;
  assign add_264640 = array_index_258761[11:1] + 11'h1e7;
  assign sel_264642 = $signed({1'h0, add_264208, array_index_258585[0]}) < $signed({1'h0, sel_264210}) ? {add_264208, array_index_258585[0]} : sel_264210;
  assign add_264644 = array_index_258764[11:1] + 11'h1e7;
  assign sel_264646 = $signed({1'h0, add_264212, array_index_258588[0]}) < $signed({1'h0, sel_264214}) ? {add_264212, array_index_258588[0]} : sel_264214;
  assign add_264656 = array_index_259171[11:0] + 12'h141;
  assign sel_264658 = $signed({1'h0, add_264224}) < $signed({1'h0, sel_264226}) ? add_264224 : sel_264226;
  assign add_264660 = array_index_259174[11:0] + 12'h141;
  assign sel_264662 = $signed({1'h0, add_264228}) < $signed({1'h0, sel_264230}) ? add_264228 : sel_264230;
  assign add_264664 = array_index_259401[11:1] + 11'h079;
  assign sel_264666 = $signed({1'h0, add_264232, array_index_259171[0]}) < $signed({1'h0, sel_264234}) ? {add_264232, array_index_259171[0]} : sel_264234;
  assign add_264668 = array_index_259404[11:1] + 11'h079;
  assign sel_264670 = $signed({1'h0, add_264236, array_index_259174[0]}) < $signed({1'h0, sel_264238}) ? {add_264236, array_index_259174[0]} : sel_264238;
  assign add_264672 = array_index_259647[11:0] + 12'h59d;
  assign sel_264674 = $signed({1'h0, add_264240}) < $signed({1'h0, sel_264242}) ? add_264240 : sel_264242;
  assign add_264676 = array_index_259650[11:0] + 12'h59d;
  assign sel_264678 = $signed({1'h0, add_264244}) < $signed({1'h0, sel_264246}) ? add_264244 : sel_264246;
  assign add_264680 = array_index_259911[11:0] + 12'ha6f;
  assign sel_264682 = $signed({1'h0, add_264248}) < $signed({1'h0, sel_264250}) ? add_264248 : sel_264250;
  assign add_264684 = array_index_259914[11:0] + 12'ha6f;
  assign sel_264686 = $signed({1'h0, add_264252}) < $signed({1'h0, sel_264254}) ? add_264252 : sel_264254;
  assign add_264688 = array_index_260195[11:1] + 11'h499;
  assign sel_264690 = $signed({1'h0, add_264256, array_index_259911[0]}) < $signed({1'h0, sel_264258}) ? {add_264256, array_index_259911[0]} : sel_264258;
  assign add_264692 = array_index_260198[11:1] + 11'h499;
  assign sel_264694 = $signed({1'h0, add_264260, array_index_259914[0]}) < $signed({1'h0, sel_264262}) ? {add_264260, array_index_259914[0]} : sel_264262;
  assign add_264696 = array_index_260507[11:1] + 11'h345;
  assign sel_264699 = $signed({1'h0, add_264264, array_index_260195[0]}) < $signed({1'h0, sel_264267}) ? {add_264264, array_index_260195[0]} : sel_264267;
  assign add_264701 = array_index_260510[11:1] + 11'h345;
  assign sel_264704 = $signed({1'h0, add_264269, array_index_260198[0]}) < $signed({1'h0, sel_264272}) ? {add_264269, array_index_260198[0]} : sel_264272;
  assign add_264706 = array_index_260845[11:0] + 12'h30f;
  assign sel_264708 = $signed({1'h0, add_264274}) < $signed({1'h0, sel_264276}) ? add_264274 : sel_264276;
  assign add_264710 = array_index_260848[11:0] + 12'h30f;
  assign sel_264712 = $signed({1'h0, add_264278}) < $signed({1'h0, sel_264280}) ? add_264278 : sel_264280;
  assign add_264714 = array_index_261207[11:0] + 12'hb55;
  assign sel_264716 = $signed({1'h0, add_264282}) < $signed({1'h0, sel_264284}) ? add_264282 : sel_264284;
  assign add_264718 = array_index_261210[11:0] + 12'hb55;
  assign sel_264720 = $signed({1'h0, add_264286}) < $signed({1'h0, sel_264288}) ? add_264286 : sel_264288;
  assign add_264722 = array_index_261595[11:0] + 12'h103;
  assign sel_264724 = $signed({1'h0, add_264290}) < $signed({1'h0, sel_264292}) ? add_264290 : sel_264292;
  assign add_264726 = array_index_261598[11:0] + 12'h103;
  assign sel_264728 = $signed({1'h0, add_264294}) < $signed({1'h0, sel_264296}) ? add_264294 : sel_264296;
  assign add_264730 = array_index_262007[11:0] + 12'hb01;
  assign sel_264732 = $signed({1'h0, add_264298}) < $signed({1'h0, sel_264300}) ? add_264298 : sel_264300;
  assign add_264734 = array_index_262010[11:0] + 12'hb01;
  assign sel_264736 = $signed({1'h0, add_264302}) < $signed({1'h0, sel_264304}) ? add_264302 : sel_264304;
  assign add_264738 = array_index_262439[11:0] + 12'h7b1;
  assign sel_264740 = $signed({1'h0, add_264306}) < $signed({1'h0, sel_264308}) ? add_264306 : sel_264308;
  assign add_264742 = array_index_262442[11:0] + 12'h7b1;
  assign sel_264744 = $signed({1'h0, add_264310}) < $signed({1'h0, sel_264312}) ? add_264310 : sel_264312;
  assign add_264746 = array_index_262871[11:0] + 12'h561;
  assign sel_264748 = $signed({1'h0, add_264314}) < $signed({1'h0, sel_264316}) ? add_264314 : sel_264316;
  assign add_264750 = array_index_262874[11:0] + 12'h561;
  assign sel_264752 = $signed({1'h0, add_264318}) < $signed({1'h0, sel_264320}) ? add_264318 : sel_264320;
  assign add_264754 = array_index_263303[11:2] + 10'h36b;
  assign sel_264756 = $signed({1'h0, add_264322, array_index_262871[1:0]}) < $signed({1'h0, sel_264324}) ? {add_264322, array_index_262871[1:0]} : sel_264324;
  assign add_264758 = array_index_263306[11:2] + 10'h36b;
  assign sel_264760 = $signed({1'h0, add_264326, array_index_262874[1:0]}) < $signed({1'h0, sel_264328}) ? {add_264326, array_index_262874[1:0]} : sel_264328;
  assign add_264762 = array_index_263735[11:2] + 10'h035;
  assign sel_264765 = $signed({1'h0, add_264330, array_index_263303[1:0]}) < $signed({1'h0, sel_264333}) ? {add_264330, array_index_263303[1:0]} : sel_264333;
  assign add_264767 = array_index_263738[11:2] + 10'h035;
  assign sel_264770 = $signed({1'h0, add_264335, array_index_263306[1:0]}) < $signed({1'h0, sel_264338}) ? {add_264335, array_index_263306[1:0]} : sel_264338;
  assign add_264772 = array_index_264167[11:0] + 12'hffb;
  assign sel_264774 = $signed({1'h0, add_264340}) < $signed({1'h0, sel_264342}) ? add_264340 : sel_264342;
  assign add_264776 = array_index_264170[11:0] + 12'hffb;
  assign sel_264778 = $signed({1'h0, add_264344}) < $signed({1'h0, sel_264346}) ? add_264344 : sel_264346;
  assign add_264790 = array_index_258285[11:2] + 10'h29b;
  assign sel_264792 = $signed({1'h0, add_264358, array_index_258159[1:0]}) < $signed({1'h0, sel_264360}) ? {add_264358, array_index_258159[1:0]} : sel_264360;
  assign add_264794 = array_index_258288[11:2] + 10'h29b;
  assign sel_264796 = $signed({1'h0, add_264362, array_index_258162[1:0]}) < $signed({1'h0, sel_264364}) ? {add_264362, array_index_258162[1:0]} : sel_264364;
  assign add_264806 = array_index_258585[11:0] + 12'h9cf;
  assign sel_264808 = $signed({1'h0, add_264374}) < $signed({1'h0, sel_264376}) ? add_264374 : sel_264376;
  assign add_264810 = array_index_258588[11:0] + 12'h9cf;
  assign sel_264812 = $signed({1'h0, add_264378}) < $signed({1'h0, sel_264380}) ? add_264378 : sel_264380;
  assign add_264822 = array_index_258957[11:0] + 12'h30b;
  assign sel_264824 = $signed({1'h0, add_264390}) < $signed({1'h0, sel_264392}) ? add_264390 : sel_264392;
  assign add_264826 = array_index_258960[11:0] + 12'h30b;
  assign sel_264828 = $signed({1'h0, add_264394}) < $signed({1'h0, sel_264396}) ? add_264394 : sel_264396;
  assign add_264897 = array_index_264599[11:0] + 12'h193;
  assign sel_264899 = $signed({1'h0, add_264465}) < $signed({1'h0, sel_264467}) ? add_264465 : sel_264467;
  assign add_264902 = array_index_264602[11:0] + 12'h193;
  assign sel_264904 = $signed({1'h0, add_264470}) < $signed({1'h0, sel_264472}) ? add_264470 : sel_264472;
  assign add_264914 = array_index_258427[11:0] + 12'hc05;
  assign sel_264916 = $signed({1'h0, add_264482}) < $signed({1'h0, sel_264484}) ? add_264482 : sel_264484;
  assign add_264918 = array_index_258430[11:0] + 12'hc05;
  assign sel_264920 = $signed({1'h0, add_264486}) < $signed({1'h0, sel_264488}) ? add_264486 : sel_264488;
  assign add_264932 = array_index_258761[11:0] + 12'h83f;
  assign sel_264934 = $signed({1'h0, add_264500}) < $signed({1'h0, sel_264502}) ? add_264500 : sel_264502;
  assign add_264936 = array_index_258764[11:0] + 12'h83f;
  assign sel_264938 = $signed({1'h0, add_264504}) < $signed({1'h0, sel_264506}) ? add_264504 : sel_264506;
  assign add_264950 = array_index_259171[11:1] + 11'h7b5;
  assign sel_264952 = $signed({1'h0, add_264518, array_index_258957[0]}) < $signed({1'h0, sel_264520}) ? {add_264518, array_index_258957[0]} : sel_264520;
  assign add_264954 = array_index_259174[11:1] + 11'h7b5;
  assign sel_264956 = $signed({1'h0, add_264522, array_index_258960[0]}) < $signed({1'h0, sel_264524}) ? {add_264522, array_index_258960[0]} : sel_264524;
  assign array_index_265031 = set1_unflattened[5'h1c];
  assign array_index_265034 = set2_unflattened[5'h1c];
  assign add_265038 = array_index_258285[11:0] + 12'hdab;
  assign sel_265040 = $signed({1'h0, add_264606}) < $signed({1'h0, sel_264608}) ? add_264606 : sel_264608;
  assign add_265042 = array_index_258288[11:0] + 12'hdab;
  assign sel_265044 = $signed({1'h0, add_264610}) < $signed({1'h0, sel_264612}) ? add_264610 : sel_264612;
  assign add_265056 = array_index_258585[11:2] + 10'h2b3;
  assign sel_265058 = $signed({1'h0, add_264624, array_index_258427[1:0]}) < $signed({1'h0, sel_264626}) ? {add_264624, array_index_258427[1:0]} : sel_264626;
  assign add_265060 = array_index_258588[11:2] + 10'h2b3;
  assign sel_265062 = $signed({1'h0, add_264628, array_index_258430[1:0]}) < $signed({1'h0, sel_264630}) ? {add_264628, array_index_258430[1:0]} : sel_264630;
  assign add_265072 = array_index_258957[11:1] + 11'h1e7;
  assign sel_265074 = $signed({1'h0, add_264640, array_index_258761[0]}) < $signed({1'h0, sel_264642}) ? {add_264640, array_index_258761[0]} : sel_264642;
  assign add_265076 = array_index_258960[11:1] + 11'h1e7;
  assign sel_265078 = $signed({1'h0, add_264644, array_index_258764[0]}) < $signed({1'h0, sel_264646}) ? {add_264644, array_index_258764[0]} : sel_264646;
  assign add_265088 = array_index_259401[11:0] + 12'h141;
  assign sel_265090 = $signed({1'h0, add_264656}) < $signed({1'h0, sel_264658}) ? add_264656 : sel_264658;
  assign add_265092 = array_index_259404[11:0] + 12'h141;
  assign sel_265094 = $signed({1'h0, add_264660}) < $signed({1'h0, sel_264662}) ? add_264660 : sel_264662;
  assign add_265096 = array_index_259647[11:1] + 11'h079;
  assign sel_265098 = $signed({1'h0, add_264664, array_index_259401[0]}) < $signed({1'h0, sel_264666}) ? {add_264664, array_index_259401[0]} : sel_264666;
  assign add_265100 = array_index_259650[11:1] + 11'h079;
  assign sel_265102 = $signed({1'h0, add_264668, array_index_259404[0]}) < $signed({1'h0, sel_264670}) ? {add_264668, array_index_259404[0]} : sel_264670;
  assign add_265104 = array_index_259911[11:0] + 12'h59d;
  assign sel_265106 = $signed({1'h0, add_264672}) < $signed({1'h0, sel_264674}) ? add_264672 : sel_264674;
  assign add_265108 = array_index_259914[11:0] + 12'h59d;
  assign sel_265110 = $signed({1'h0, add_264676}) < $signed({1'h0, sel_264678}) ? add_264676 : sel_264678;
  assign add_265112 = array_index_260195[11:0] + 12'ha6f;
  assign sel_265114 = $signed({1'h0, add_264680}) < $signed({1'h0, sel_264682}) ? add_264680 : sel_264682;
  assign add_265116 = array_index_260198[11:0] + 12'ha6f;
  assign sel_265118 = $signed({1'h0, add_264684}) < $signed({1'h0, sel_264686}) ? add_264684 : sel_264686;
  assign add_265120 = array_index_260507[11:1] + 11'h499;
  assign sel_265122 = $signed({1'h0, add_264688, array_index_260195[0]}) < $signed({1'h0, sel_264690}) ? {add_264688, array_index_260195[0]} : sel_264690;
  assign add_265124 = array_index_260510[11:1] + 11'h499;
  assign sel_265126 = $signed({1'h0, add_264692, array_index_260198[0]}) < $signed({1'h0, sel_264694}) ? {add_264692, array_index_260198[0]} : sel_264694;
  assign add_265128 = array_index_260845[11:1] + 11'h345;
  assign sel_265131 = $signed({1'h0, add_264696, array_index_260507[0]}) < $signed({1'h0, sel_264699}) ? {add_264696, array_index_260507[0]} : sel_264699;
  assign add_265133 = array_index_260848[11:1] + 11'h345;
  assign sel_265136 = $signed({1'h0, add_264701, array_index_260510[0]}) < $signed({1'h0, sel_264704}) ? {add_264701, array_index_260510[0]} : sel_264704;
  assign add_265138 = array_index_261207[11:0] + 12'h30f;
  assign sel_265140 = $signed({1'h0, add_264706}) < $signed({1'h0, sel_264708}) ? add_264706 : sel_264708;
  assign add_265142 = array_index_261210[11:0] + 12'h30f;
  assign sel_265144 = $signed({1'h0, add_264710}) < $signed({1'h0, sel_264712}) ? add_264710 : sel_264712;
  assign add_265146 = array_index_261595[11:0] + 12'hb55;
  assign sel_265148 = $signed({1'h0, add_264714}) < $signed({1'h0, sel_264716}) ? add_264714 : sel_264716;
  assign add_265150 = array_index_261598[11:0] + 12'hb55;
  assign sel_265152 = $signed({1'h0, add_264718}) < $signed({1'h0, sel_264720}) ? add_264718 : sel_264720;
  assign add_265154 = array_index_262007[11:0] + 12'h103;
  assign sel_265156 = $signed({1'h0, add_264722}) < $signed({1'h0, sel_264724}) ? add_264722 : sel_264724;
  assign add_265158 = array_index_262010[11:0] + 12'h103;
  assign sel_265160 = $signed({1'h0, add_264726}) < $signed({1'h0, sel_264728}) ? add_264726 : sel_264728;
  assign add_265162 = array_index_262439[11:0] + 12'hb01;
  assign sel_265164 = $signed({1'h0, add_264730}) < $signed({1'h0, sel_264732}) ? add_264730 : sel_264732;
  assign add_265166 = array_index_262442[11:0] + 12'hb01;
  assign sel_265168 = $signed({1'h0, add_264734}) < $signed({1'h0, sel_264736}) ? add_264734 : sel_264736;
  assign add_265170 = array_index_262871[11:0] + 12'h7b1;
  assign sel_265172 = $signed({1'h0, add_264738}) < $signed({1'h0, sel_264740}) ? add_264738 : sel_264740;
  assign add_265174 = array_index_262874[11:0] + 12'h7b1;
  assign sel_265176 = $signed({1'h0, add_264742}) < $signed({1'h0, sel_264744}) ? add_264742 : sel_264744;
  assign add_265178 = array_index_263303[11:0] + 12'h561;
  assign sel_265180 = $signed({1'h0, add_264746}) < $signed({1'h0, sel_264748}) ? add_264746 : sel_264748;
  assign add_265182 = array_index_263306[11:0] + 12'h561;
  assign sel_265184 = $signed({1'h0, add_264750}) < $signed({1'h0, sel_264752}) ? add_264750 : sel_264752;
  assign add_265186 = array_index_263735[11:2] + 10'h36b;
  assign sel_265188 = $signed({1'h0, add_264754, array_index_263303[1:0]}) < $signed({1'h0, sel_264756}) ? {add_264754, array_index_263303[1:0]} : sel_264756;
  assign add_265190 = array_index_263738[11:2] + 10'h36b;
  assign sel_265192 = $signed({1'h0, add_264758, array_index_263306[1:0]}) < $signed({1'h0, sel_264760}) ? {add_264758, array_index_263306[1:0]} : sel_264760;
  assign add_265194 = array_index_264167[11:2] + 10'h035;
  assign sel_265197 = $signed({1'h0, add_264762, array_index_263735[1:0]}) < $signed({1'h0, sel_264765}) ? {add_264762, array_index_263735[1:0]} : sel_264765;
  assign add_265199 = array_index_264170[11:2] + 10'h035;
  assign sel_265202 = $signed({1'h0, add_264767, array_index_263738[1:0]}) < $signed({1'h0, sel_264770}) ? {add_264767, array_index_263738[1:0]} : sel_264770;
  assign add_265204 = array_index_264599[11:0] + 12'hffb;
  assign sel_265206 = $signed({1'h0, add_264772}) < $signed({1'h0, sel_264774}) ? add_264772 : sel_264774;
  assign add_265208 = array_index_264602[11:0] + 12'hffb;
  assign sel_265210 = $signed({1'h0, add_264776}) < $signed({1'h0, sel_264778}) ? add_264776 : sel_264778;
  assign add_265222 = array_index_258427[11:2] + 10'h29b;
  assign sel_265224 = $signed({1'h0, add_264790, array_index_258285[1:0]}) < $signed({1'h0, sel_264792}) ? {add_264790, array_index_258285[1:0]} : sel_264792;
  assign add_265226 = array_index_258430[11:2] + 10'h29b;
  assign sel_265228 = $signed({1'h0, add_264794, array_index_258288[1:0]}) < $signed({1'h0, sel_264796}) ? {add_264794, array_index_258288[1:0]} : sel_264796;
  assign add_265238 = array_index_258761[11:0] + 12'h9cf;
  assign sel_265240 = $signed({1'h0, add_264806}) < $signed({1'h0, sel_264808}) ? add_264806 : sel_264808;
  assign add_265242 = array_index_258764[11:0] + 12'h9cf;
  assign sel_265244 = $signed({1'h0, add_264810}) < $signed({1'h0, sel_264812}) ? add_264810 : sel_264812;
  assign add_265254 = array_index_259171[11:0] + 12'h30b;
  assign sel_265256 = $signed({1'h0, add_264822}) < $signed({1'h0, sel_264824}) ? add_264822 : sel_264824;
  assign add_265258 = array_index_259174[11:0] + 12'h30b;
  assign sel_265260 = $signed({1'h0, add_264826}) < $signed({1'h0, sel_264828}) ? add_264826 : sel_264828;
  assign add_265329 = array_index_265031[11:0] + 12'h193;
  assign sel_265331 = $signed({1'h0, add_264897}) < $signed({1'h0, sel_264899}) ? add_264897 : sel_264899;
  assign add_265334 = array_index_265034[11:0] + 12'h193;
  assign sel_265336 = $signed({1'h0, add_264902}) < $signed({1'h0, sel_264904}) ? add_264902 : sel_264904;
  assign add_265346 = array_index_258585[11:0] + 12'hc05;
  assign sel_265348 = $signed({1'h0, add_264914}) < $signed({1'h0, sel_264916}) ? add_264914 : sel_264916;
  assign add_265350 = array_index_258588[11:0] + 12'hc05;
  assign sel_265352 = $signed({1'h0, add_264918}) < $signed({1'h0, sel_264920}) ? add_264918 : sel_264920;
  assign add_265364 = array_index_258957[11:0] + 12'h83f;
  assign sel_265366 = $signed({1'h0, add_264932}) < $signed({1'h0, sel_264934}) ? add_264932 : sel_264934;
  assign add_265368 = array_index_258960[11:0] + 12'h83f;
  assign sel_265370 = $signed({1'h0, add_264936}) < $signed({1'h0, sel_264938}) ? add_264936 : sel_264938;
  assign add_265382 = array_index_259401[11:1] + 11'h7b5;
  assign sel_265384 = $signed({1'h0, add_264950, array_index_259171[0]}) < $signed({1'h0, sel_264952}) ? {add_264950, array_index_259171[0]} : sel_264952;
  assign add_265386 = array_index_259404[11:1] + 11'h7b5;
  assign sel_265388 = $signed({1'h0, add_264954, array_index_259174[0]}) < $signed({1'h0, sel_264956}) ? {add_264954, array_index_259174[0]} : sel_264956;
  assign array_index_265463 = set1_unflattened[5'h1d];
  assign array_index_265466 = set2_unflattened[5'h1d];
  assign add_265470 = array_index_258427[11:0] + 12'hdab;
  assign sel_265472 = $signed({1'h0, add_265038}) < $signed({1'h0, sel_265040}) ? add_265038 : sel_265040;
  assign add_265474 = array_index_258430[11:0] + 12'hdab;
  assign sel_265476 = $signed({1'h0, add_265042}) < $signed({1'h0, sel_265044}) ? add_265042 : sel_265044;
  assign add_265488 = array_index_258761[11:2] + 10'h2b3;
  assign sel_265490 = $signed({1'h0, add_265056, array_index_258585[1:0]}) < $signed({1'h0, sel_265058}) ? {add_265056, array_index_258585[1:0]} : sel_265058;
  assign add_265492 = array_index_258764[11:2] + 10'h2b3;
  assign sel_265494 = $signed({1'h0, add_265060, array_index_258588[1:0]}) < $signed({1'h0, sel_265062}) ? {add_265060, array_index_258588[1:0]} : sel_265062;
  assign add_265504 = array_index_259171[11:1] + 11'h1e7;
  assign sel_265506 = $signed({1'h0, add_265072, array_index_258957[0]}) < $signed({1'h0, sel_265074}) ? {add_265072, array_index_258957[0]} : sel_265074;
  assign add_265508 = array_index_259174[11:1] + 11'h1e7;
  assign sel_265510 = $signed({1'h0, add_265076, array_index_258960[0]}) < $signed({1'h0, sel_265078}) ? {add_265076, array_index_258960[0]} : sel_265078;
  assign add_265520 = array_index_259647[11:0] + 12'h141;
  assign sel_265522 = $signed({1'h0, add_265088}) < $signed({1'h0, sel_265090}) ? add_265088 : sel_265090;
  assign add_265524 = array_index_259650[11:0] + 12'h141;
  assign sel_265526 = $signed({1'h0, add_265092}) < $signed({1'h0, sel_265094}) ? add_265092 : sel_265094;
  assign add_265528 = array_index_259911[11:1] + 11'h079;
  assign sel_265530 = $signed({1'h0, add_265096, array_index_259647[0]}) < $signed({1'h0, sel_265098}) ? {add_265096, array_index_259647[0]} : sel_265098;
  assign add_265532 = array_index_259914[11:1] + 11'h079;
  assign sel_265534 = $signed({1'h0, add_265100, array_index_259650[0]}) < $signed({1'h0, sel_265102}) ? {add_265100, array_index_259650[0]} : sel_265102;
  assign add_265536 = array_index_260195[11:0] + 12'h59d;
  assign sel_265538 = $signed({1'h0, add_265104}) < $signed({1'h0, sel_265106}) ? add_265104 : sel_265106;
  assign add_265540 = array_index_260198[11:0] + 12'h59d;
  assign sel_265542 = $signed({1'h0, add_265108}) < $signed({1'h0, sel_265110}) ? add_265108 : sel_265110;
  assign add_265544 = array_index_260507[11:0] + 12'ha6f;
  assign sel_265546 = $signed({1'h0, add_265112}) < $signed({1'h0, sel_265114}) ? add_265112 : sel_265114;
  assign add_265548 = array_index_260510[11:0] + 12'ha6f;
  assign sel_265550 = $signed({1'h0, add_265116}) < $signed({1'h0, sel_265118}) ? add_265116 : sel_265118;
  assign add_265552 = array_index_260845[11:1] + 11'h499;
  assign sel_265554 = $signed({1'h0, add_265120, array_index_260507[0]}) < $signed({1'h0, sel_265122}) ? {add_265120, array_index_260507[0]} : sel_265122;
  assign add_265556 = array_index_260848[11:1] + 11'h499;
  assign sel_265558 = $signed({1'h0, add_265124, array_index_260510[0]}) < $signed({1'h0, sel_265126}) ? {add_265124, array_index_260510[0]} : sel_265126;
  assign add_265560 = array_index_261207[11:1] + 11'h345;
  assign sel_265563 = $signed({1'h0, add_265128, array_index_260845[0]}) < $signed({1'h0, sel_265131}) ? {add_265128, array_index_260845[0]} : sel_265131;
  assign add_265565 = array_index_261210[11:1] + 11'h345;
  assign sel_265568 = $signed({1'h0, add_265133, array_index_260848[0]}) < $signed({1'h0, sel_265136}) ? {add_265133, array_index_260848[0]} : sel_265136;
  assign add_265570 = array_index_261595[11:0] + 12'h30f;
  assign sel_265572 = $signed({1'h0, add_265138}) < $signed({1'h0, sel_265140}) ? add_265138 : sel_265140;
  assign add_265574 = array_index_261598[11:0] + 12'h30f;
  assign sel_265576 = $signed({1'h0, add_265142}) < $signed({1'h0, sel_265144}) ? add_265142 : sel_265144;
  assign add_265578 = array_index_262007[11:0] + 12'hb55;
  assign sel_265580 = $signed({1'h0, add_265146}) < $signed({1'h0, sel_265148}) ? add_265146 : sel_265148;
  assign add_265582 = array_index_262010[11:0] + 12'hb55;
  assign sel_265584 = $signed({1'h0, add_265150}) < $signed({1'h0, sel_265152}) ? add_265150 : sel_265152;
  assign add_265586 = array_index_262439[11:0] + 12'h103;
  assign sel_265588 = $signed({1'h0, add_265154}) < $signed({1'h0, sel_265156}) ? add_265154 : sel_265156;
  assign add_265590 = array_index_262442[11:0] + 12'h103;
  assign sel_265592 = $signed({1'h0, add_265158}) < $signed({1'h0, sel_265160}) ? add_265158 : sel_265160;
  assign add_265594 = array_index_262871[11:0] + 12'hb01;
  assign sel_265596 = $signed({1'h0, add_265162}) < $signed({1'h0, sel_265164}) ? add_265162 : sel_265164;
  assign add_265598 = array_index_262874[11:0] + 12'hb01;
  assign sel_265600 = $signed({1'h0, add_265166}) < $signed({1'h0, sel_265168}) ? add_265166 : sel_265168;
  assign add_265602 = array_index_263303[11:0] + 12'h7b1;
  assign sel_265604 = $signed({1'h0, add_265170}) < $signed({1'h0, sel_265172}) ? add_265170 : sel_265172;
  assign add_265606 = array_index_263306[11:0] + 12'h7b1;
  assign sel_265608 = $signed({1'h0, add_265174}) < $signed({1'h0, sel_265176}) ? add_265174 : sel_265176;
  assign add_265610 = array_index_263735[11:0] + 12'h561;
  assign sel_265612 = $signed({1'h0, add_265178}) < $signed({1'h0, sel_265180}) ? add_265178 : sel_265180;
  assign add_265614 = array_index_263738[11:0] + 12'h561;
  assign sel_265616 = $signed({1'h0, add_265182}) < $signed({1'h0, sel_265184}) ? add_265182 : sel_265184;
  assign add_265618 = array_index_264167[11:2] + 10'h36b;
  assign sel_265620 = $signed({1'h0, add_265186, array_index_263735[1:0]}) < $signed({1'h0, sel_265188}) ? {add_265186, array_index_263735[1:0]} : sel_265188;
  assign add_265622 = array_index_264170[11:2] + 10'h36b;
  assign sel_265624 = $signed({1'h0, add_265190, array_index_263738[1:0]}) < $signed({1'h0, sel_265192}) ? {add_265190, array_index_263738[1:0]} : sel_265192;
  assign add_265626 = array_index_264599[11:2] + 10'h035;
  assign sel_265629 = $signed({1'h0, add_265194, array_index_264167[1:0]}) < $signed({1'h0, sel_265197}) ? {add_265194, array_index_264167[1:0]} : sel_265197;
  assign add_265631 = array_index_264602[11:2] + 10'h035;
  assign sel_265634 = $signed({1'h0, add_265199, array_index_264170[1:0]}) < $signed({1'h0, sel_265202}) ? {add_265199, array_index_264170[1:0]} : sel_265202;
  assign add_265636 = array_index_265031[11:0] + 12'hffb;
  assign sel_265638 = $signed({1'h0, add_265204}) < $signed({1'h0, sel_265206}) ? add_265204 : sel_265206;
  assign add_265640 = array_index_265034[11:0] + 12'hffb;
  assign sel_265642 = $signed({1'h0, add_265208}) < $signed({1'h0, sel_265210}) ? add_265208 : sel_265210;
  assign add_265654 = array_index_258585[11:2] + 10'h29b;
  assign sel_265656 = $signed({1'h0, add_265222, array_index_258427[1:0]}) < $signed({1'h0, sel_265224}) ? {add_265222, array_index_258427[1:0]} : sel_265224;
  assign add_265658 = array_index_258588[11:2] + 10'h29b;
  assign sel_265660 = $signed({1'h0, add_265226, array_index_258430[1:0]}) < $signed({1'h0, sel_265228}) ? {add_265226, array_index_258430[1:0]} : sel_265228;
  assign add_265670 = array_index_258957[11:0] + 12'h9cf;
  assign sel_265672 = $signed({1'h0, add_265238}) < $signed({1'h0, sel_265240}) ? add_265238 : sel_265240;
  assign add_265674 = array_index_258960[11:0] + 12'h9cf;
  assign sel_265676 = $signed({1'h0, add_265242}) < $signed({1'h0, sel_265244}) ? add_265242 : sel_265244;
  assign add_265686 = array_index_259401[11:0] + 12'h30b;
  assign sel_265688 = $signed({1'h0, add_265254}) < $signed({1'h0, sel_265256}) ? add_265254 : sel_265256;
  assign add_265690 = array_index_259404[11:0] + 12'h30b;
  assign sel_265692 = $signed({1'h0, add_265258}) < $signed({1'h0, sel_265260}) ? add_265258 : sel_265260;
  assign add_265760 = array_index_265463[11:0] + 12'h193;
  assign sel_265762 = $signed({1'h0, add_265329}) < $signed({1'h0, sel_265331}) ? add_265329 : sel_265331;
  assign add_265764 = array_index_265466[11:0] + 12'h193;
  assign sel_265766 = $signed({1'h0, add_265334}) < $signed({1'h0, sel_265336}) ? add_265334 : sel_265336;
  assign add_265776 = array_index_258761[11:0] + 12'hc05;
  assign sel_265778 = $signed({1'h0, add_265346}) < $signed({1'h0, sel_265348}) ? add_265346 : sel_265348;
  assign add_265780 = array_index_258764[11:0] + 12'hc05;
  assign sel_265782 = $signed({1'h0, add_265350}) < $signed({1'h0, sel_265352}) ? add_265350 : sel_265352;
  assign add_265794 = array_index_259171[11:0] + 12'h83f;
  assign sel_265796 = $signed({1'h0, add_265364}) < $signed({1'h0, sel_265366}) ? add_265364 : sel_265366;
  assign add_265798 = array_index_259174[11:0] + 12'h83f;
  assign sel_265800 = $signed({1'h0, add_265368}) < $signed({1'h0, sel_265370}) ? add_265368 : sel_265370;
  assign add_265812 = array_index_259647[11:1] + 11'h7b5;
  assign sel_265814 = $signed({1'h0, add_265382, array_index_259401[0]}) < $signed({1'h0, sel_265384}) ? {add_265382, array_index_259401[0]} : sel_265384;
  assign add_265816 = array_index_259650[11:1] + 11'h7b5;
  assign sel_265818 = $signed({1'h0, add_265386, array_index_259404[0]}) < $signed({1'h0, sel_265388}) ? {add_265386, array_index_259404[0]} : sel_265388;
  assign add_265898 = array_index_258585[11:0] + 12'hdab;
  assign sel_265900 = $signed({1'h0, add_265470}) < $signed({1'h0, sel_265472}) ? add_265470 : sel_265472;
  assign add_265902 = array_index_258588[11:0] + 12'hdab;
  assign sel_265904 = $signed({1'h0, add_265474}) < $signed({1'h0, sel_265476}) ? add_265474 : sel_265476;
  assign add_265916 = array_index_258957[11:2] + 10'h2b3;
  assign sel_265918 = $signed({1'h0, add_265488, array_index_258761[1:0]}) < $signed({1'h0, sel_265490}) ? {add_265488, array_index_258761[1:0]} : sel_265490;
  assign add_265920 = array_index_258960[11:2] + 10'h2b3;
  assign sel_265922 = $signed({1'h0, add_265492, array_index_258764[1:0]}) < $signed({1'h0, sel_265494}) ? {add_265492, array_index_258764[1:0]} : sel_265494;
  assign add_265932 = array_index_259401[11:1] + 11'h1e7;
  assign sel_265934 = $signed({1'h0, add_265504, array_index_259171[0]}) < $signed({1'h0, sel_265506}) ? {add_265504, array_index_259171[0]} : sel_265506;
  assign add_265936 = array_index_259404[11:1] + 11'h1e7;
  assign sel_265938 = $signed({1'h0, add_265508, array_index_259174[0]}) < $signed({1'h0, sel_265510}) ? {add_265508, array_index_259174[0]} : sel_265510;
  assign add_265948 = array_index_259911[11:0] + 12'h141;
  assign sel_265950 = $signed({1'h0, add_265520}) < $signed({1'h0, sel_265522}) ? add_265520 : sel_265522;
  assign add_265952 = array_index_259914[11:0] + 12'h141;
  assign sel_265954 = $signed({1'h0, add_265524}) < $signed({1'h0, sel_265526}) ? add_265524 : sel_265526;
  assign add_265956 = array_index_260195[11:1] + 11'h079;
  assign sel_265958 = $signed({1'h0, add_265528, array_index_259911[0]}) < $signed({1'h0, sel_265530}) ? {add_265528, array_index_259911[0]} : sel_265530;
  assign add_265960 = array_index_260198[11:1] + 11'h079;
  assign sel_265962 = $signed({1'h0, add_265532, array_index_259914[0]}) < $signed({1'h0, sel_265534}) ? {add_265532, array_index_259914[0]} : sel_265534;
  assign add_265964 = array_index_260507[11:0] + 12'h59d;
  assign sel_265966 = $signed({1'h0, add_265536}) < $signed({1'h0, sel_265538}) ? add_265536 : sel_265538;
  assign add_265968 = array_index_260510[11:0] + 12'h59d;
  assign sel_265970 = $signed({1'h0, add_265540}) < $signed({1'h0, sel_265542}) ? add_265540 : sel_265542;
  assign add_265972 = array_index_260845[11:0] + 12'ha6f;
  assign sel_265974 = $signed({1'h0, add_265544}) < $signed({1'h0, sel_265546}) ? add_265544 : sel_265546;
  assign add_265976 = array_index_260848[11:0] + 12'ha6f;
  assign sel_265978 = $signed({1'h0, add_265548}) < $signed({1'h0, sel_265550}) ? add_265548 : sel_265550;
  assign add_265980 = array_index_261207[11:1] + 11'h499;
  assign sel_265982 = $signed({1'h0, add_265552, array_index_260845[0]}) < $signed({1'h0, sel_265554}) ? {add_265552, array_index_260845[0]} : sel_265554;
  assign add_265984 = array_index_261210[11:1] + 11'h499;
  assign sel_265986 = $signed({1'h0, add_265556, array_index_260848[0]}) < $signed({1'h0, sel_265558}) ? {add_265556, array_index_260848[0]} : sel_265558;
  assign add_265988 = array_index_261595[11:1] + 11'h345;
  assign sel_265991 = $signed({1'h0, add_265560, array_index_261207[0]}) < $signed({1'h0, sel_265563}) ? {add_265560, array_index_261207[0]} : sel_265563;
  assign add_265993 = array_index_261598[11:1] + 11'h345;
  assign sel_265996 = $signed({1'h0, add_265565, array_index_261210[0]}) < $signed({1'h0, sel_265568}) ? {add_265565, array_index_261210[0]} : sel_265568;
  assign add_265998 = array_index_262007[11:0] + 12'h30f;
  assign sel_266000 = $signed({1'h0, add_265570}) < $signed({1'h0, sel_265572}) ? add_265570 : sel_265572;
  assign add_266002 = array_index_262010[11:0] + 12'h30f;
  assign sel_266004 = $signed({1'h0, add_265574}) < $signed({1'h0, sel_265576}) ? add_265574 : sel_265576;
  assign add_266006 = array_index_262439[11:0] + 12'hb55;
  assign sel_266008 = $signed({1'h0, add_265578}) < $signed({1'h0, sel_265580}) ? add_265578 : sel_265580;
  assign add_266010 = array_index_262442[11:0] + 12'hb55;
  assign sel_266012 = $signed({1'h0, add_265582}) < $signed({1'h0, sel_265584}) ? add_265582 : sel_265584;
  assign add_266014 = array_index_262871[11:0] + 12'h103;
  assign sel_266016 = $signed({1'h0, add_265586}) < $signed({1'h0, sel_265588}) ? add_265586 : sel_265588;
  assign add_266018 = array_index_262874[11:0] + 12'h103;
  assign sel_266020 = $signed({1'h0, add_265590}) < $signed({1'h0, sel_265592}) ? add_265590 : sel_265592;
  assign add_266022 = array_index_263303[11:0] + 12'hb01;
  assign sel_266024 = $signed({1'h0, add_265594}) < $signed({1'h0, sel_265596}) ? add_265594 : sel_265596;
  assign add_266026 = array_index_263306[11:0] + 12'hb01;
  assign sel_266028 = $signed({1'h0, add_265598}) < $signed({1'h0, sel_265600}) ? add_265598 : sel_265600;
  assign add_266030 = array_index_263735[11:0] + 12'h7b1;
  assign sel_266032 = $signed({1'h0, add_265602}) < $signed({1'h0, sel_265604}) ? add_265602 : sel_265604;
  assign add_266034 = array_index_263738[11:0] + 12'h7b1;
  assign sel_266036 = $signed({1'h0, add_265606}) < $signed({1'h0, sel_265608}) ? add_265606 : sel_265608;
  assign add_266038 = array_index_264167[11:0] + 12'h561;
  assign sel_266040 = $signed({1'h0, add_265610}) < $signed({1'h0, sel_265612}) ? add_265610 : sel_265612;
  assign add_266042 = array_index_264170[11:0] + 12'h561;
  assign sel_266044 = $signed({1'h0, add_265614}) < $signed({1'h0, sel_265616}) ? add_265614 : sel_265616;
  assign add_266046 = array_index_264599[11:2] + 10'h36b;
  assign sel_266048 = $signed({1'h0, add_265618, array_index_264167[1:0]}) < $signed({1'h0, sel_265620}) ? {add_265618, array_index_264167[1:0]} : sel_265620;
  assign add_266050 = array_index_264602[11:2] + 10'h36b;
  assign sel_266052 = $signed({1'h0, add_265622, array_index_264170[1:0]}) < $signed({1'h0, sel_265624}) ? {add_265622, array_index_264170[1:0]} : sel_265624;
  assign add_266054 = array_index_265031[11:2] + 10'h035;
  assign sel_266057 = $signed({1'h0, add_265626, array_index_264599[1:0]}) < $signed({1'h0, sel_265629}) ? {add_265626, array_index_264599[1:0]} : sel_265629;
  assign add_266059 = array_index_265034[11:2] + 10'h035;
  assign sel_266062 = $signed({1'h0, add_265631, array_index_264602[1:0]}) < $signed({1'h0, sel_265634}) ? {add_265631, array_index_264602[1:0]} : sel_265634;
  assign add_266064 = array_index_265463[11:0] + 12'hffb;
  assign sel_266066 = $signed({1'h0, add_265636}) < $signed({1'h0, sel_265638}) ? add_265636 : sel_265638;
  assign add_266068 = array_index_265466[11:0] + 12'hffb;
  assign sel_266070 = $signed({1'h0, add_265640}) < $signed({1'h0, sel_265642}) ? add_265640 : sel_265642;
  assign add_266078 = array_index_258761[11:2] + 10'h29b;
  assign sel_266080 = $signed({1'h0, add_265654, array_index_258585[1:0]}) < $signed({1'h0, sel_265656}) ? {add_265654, array_index_258585[1:0]} : sel_265656;
  assign add_266082 = array_index_258764[11:2] + 10'h29b;
  assign sel_266084 = $signed({1'h0, add_265658, array_index_258588[1:0]}) < $signed({1'h0, sel_265660}) ? {add_265658, array_index_258588[1:0]} : sel_265660;
  assign add_266094 = array_index_259171[11:0] + 12'h9cf;
  assign sel_266096 = $signed({1'h0, add_265670}) < $signed({1'h0, sel_265672}) ? add_265670 : sel_265672;
  assign add_266098 = array_index_259174[11:0] + 12'h9cf;
  assign sel_266100 = $signed({1'h0, add_265674}) < $signed({1'h0, sel_265676}) ? add_265674 : sel_265676;
  assign add_266110 = array_index_259647[11:0] + 12'h30b;
  assign sel_266112 = $signed({1'h0, add_265686}) < $signed({1'h0, sel_265688}) ? add_265686 : sel_265688;
  assign add_266114 = array_index_259650[11:0] + 12'h30b;
  assign sel_266116 = $signed({1'h0, add_265690}) < $signed({1'h0, sel_265692}) ? add_265690 : sel_265692;
  assign add_266194 = array_index_258957[11:0] + 12'hc05;
  assign sel_266196 = $signed({1'h0, add_265776}) < $signed({1'h0, sel_265778}) ? add_265776 : sel_265778;
  assign add_266198 = array_index_258960[11:0] + 12'hc05;
  assign sel_266200 = $signed({1'h0, add_265780}) < $signed({1'h0, sel_265782}) ? add_265780 : sel_265782;
  assign add_266212 = array_index_259401[11:0] + 12'h83f;
  assign sel_266214 = $signed({1'h0, add_265794}) < $signed({1'h0, sel_265796}) ? add_265794 : sel_265796;
  assign add_266216 = array_index_259404[11:0] + 12'h83f;
  assign sel_266218 = $signed({1'h0, add_265798}) < $signed({1'h0, sel_265800}) ? add_265798 : sel_265800;
  assign add_266230 = array_index_259911[11:1] + 11'h7b5;
  assign sel_266232 = $signed({1'h0, add_265812, array_index_259647[0]}) < $signed({1'h0, sel_265814}) ? {add_265812, array_index_259647[0]} : sel_265814;
  assign add_266234 = array_index_259914[11:1] + 11'h7b5;
  assign sel_266236 = $signed({1'h0, add_265816, array_index_259650[0]}) < $signed({1'h0, sel_265818}) ? {add_265816, array_index_259650[0]} : sel_265818;
  assign add_266312 = array_index_258761[11:0] + 12'hdab;
  assign sel_266314 = $signed({1'h0, add_265898}) < $signed({1'h0, sel_265900}) ? add_265898 : sel_265900;
  assign add_266316 = array_index_258764[11:0] + 12'hdab;
  assign sel_266318 = $signed({1'h0, add_265902}) < $signed({1'h0, sel_265904}) ? add_265902 : sel_265904;
  assign add_266330 = array_index_259171[11:2] + 10'h2b3;
  assign sel_266332 = $signed({1'h0, add_265916, array_index_258957[1:0]}) < $signed({1'h0, sel_265918}) ? {add_265916, array_index_258957[1:0]} : sel_265918;
  assign add_266334 = array_index_259174[11:2] + 10'h2b3;
  assign sel_266336 = $signed({1'h0, add_265920, array_index_258960[1:0]}) < $signed({1'h0, sel_265922}) ? {add_265920, array_index_258960[1:0]} : sel_265922;
  assign add_266346 = array_index_259647[11:1] + 11'h1e7;
  assign sel_266348 = $signed({1'h0, add_265932, array_index_259401[0]}) < $signed({1'h0, sel_265934}) ? {add_265932, array_index_259401[0]} : sel_265934;
  assign add_266350 = array_index_259650[11:1] + 11'h1e7;
  assign sel_266352 = $signed({1'h0, add_265936, array_index_259404[0]}) < $signed({1'h0, sel_265938}) ? {add_265936, array_index_259404[0]} : sel_265938;
  assign add_266362 = array_index_260195[11:0] + 12'h141;
  assign sel_266364 = $signed({1'h0, add_265948}) < $signed({1'h0, sel_265950}) ? add_265948 : sel_265950;
  assign add_266366 = array_index_260198[11:0] + 12'h141;
  assign sel_266368 = $signed({1'h0, add_265952}) < $signed({1'h0, sel_265954}) ? add_265952 : sel_265954;
  assign add_266370 = array_index_260507[11:1] + 11'h079;
  assign sel_266372 = $signed({1'h0, add_265956, array_index_260195[0]}) < $signed({1'h0, sel_265958}) ? {add_265956, array_index_260195[0]} : sel_265958;
  assign add_266374 = array_index_260510[11:1] + 11'h079;
  assign sel_266376 = $signed({1'h0, add_265960, array_index_260198[0]}) < $signed({1'h0, sel_265962}) ? {add_265960, array_index_260198[0]} : sel_265962;
  assign add_266378 = array_index_260845[11:0] + 12'h59d;
  assign sel_266380 = $signed({1'h0, add_265964}) < $signed({1'h0, sel_265966}) ? add_265964 : sel_265966;
  assign add_266382 = array_index_260848[11:0] + 12'h59d;
  assign sel_266384 = $signed({1'h0, add_265968}) < $signed({1'h0, sel_265970}) ? add_265968 : sel_265970;
  assign add_266386 = array_index_261207[11:0] + 12'ha6f;
  assign sel_266388 = $signed({1'h0, add_265972}) < $signed({1'h0, sel_265974}) ? add_265972 : sel_265974;
  assign add_266390 = array_index_261210[11:0] + 12'ha6f;
  assign sel_266392 = $signed({1'h0, add_265976}) < $signed({1'h0, sel_265978}) ? add_265976 : sel_265978;
  assign add_266394 = array_index_261595[11:1] + 11'h499;
  assign sel_266396 = $signed({1'h0, add_265980, array_index_261207[0]}) < $signed({1'h0, sel_265982}) ? {add_265980, array_index_261207[0]} : sel_265982;
  assign add_266398 = array_index_261598[11:1] + 11'h499;
  assign sel_266400 = $signed({1'h0, add_265984, array_index_261210[0]}) < $signed({1'h0, sel_265986}) ? {add_265984, array_index_261210[0]} : sel_265986;
  assign add_266402 = array_index_262007[11:1] + 11'h345;
  assign sel_266405 = $signed({1'h0, add_265988, array_index_261595[0]}) < $signed({1'h0, sel_265991}) ? {add_265988, array_index_261595[0]} : sel_265991;
  assign add_266407 = array_index_262010[11:1] + 11'h345;
  assign sel_266410 = $signed({1'h0, add_265993, array_index_261598[0]}) < $signed({1'h0, sel_265996}) ? {add_265993, array_index_261598[0]} : sel_265996;
  assign add_266412 = array_index_262439[11:0] + 12'h30f;
  assign sel_266414 = $signed({1'h0, add_265998}) < $signed({1'h0, sel_266000}) ? add_265998 : sel_266000;
  assign add_266416 = array_index_262442[11:0] + 12'h30f;
  assign sel_266418 = $signed({1'h0, add_266002}) < $signed({1'h0, sel_266004}) ? add_266002 : sel_266004;
  assign add_266420 = array_index_262871[11:0] + 12'hb55;
  assign sel_266422 = $signed({1'h0, add_266006}) < $signed({1'h0, sel_266008}) ? add_266006 : sel_266008;
  assign add_266424 = array_index_262874[11:0] + 12'hb55;
  assign sel_266426 = $signed({1'h0, add_266010}) < $signed({1'h0, sel_266012}) ? add_266010 : sel_266012;
  assign add_266428 = array_index_263303[11:0] + 12'h103;
  assign sel_266430 = $signed({1'h0, add_266014}) < $signed({1'h0, sel_266016}) ? add_266014 : sel_266016;
  assign add_266432 = array_index_263306[11:0] + 12'h103;
  assign sel_266434 = $signed({1'h0, add_266018}) < $signed({1'h0, sel_266020}) ? add_266018 : sel_266020;
  assign add_266436 = array_index_263735[11:0] + 12'hb01;
  assign sel_266438 = $signed({1'h0, add_266022}) < $signed({1'h0, sel_266024}) ? add_266022 : sel_266024;
  assign add_266440 = array_index_263738[11:0] + 12'hb01;
  assign sel_266442 = $signed({1'h0, add_266026}) < $signed({1'h0, sel_266028}) ? add_266026 : sel_266028;
  assign add_266444 = array_index_264167[11:0] + 12'h7b1;
  assign sel_266446 = $signed({1'h0, add_266030}) < $signed({1'h0, sel_266032}) ? add_266030 : sel_266032;
  assign add_266448 = array_index_264170[11:0] + 12'h7b1;
  assign sel_266450 = $signed({1'h0, add_266034}) < $signed({1'h0, sel_266036}) ? add_266034 : sel_266036;
  assign add_266452 = array_index_264599[11:0] + 12'h561;
  assign sel_266454 = $signed({1'h0, add_266038}) < $signed({1'h0, sel_266040}) ? add_266038 : sel_266040;
  assign add_266456 = array_index_264602[11:0] + 12'h561;
  assign sel_266458 = $signed({1'h0, add_266042}) < $signed({1'h0, sel_266044}) ? add_266042 : sel_266044;
  assign add_266460 = array_index_265031[11:2] + 10'h36b;
  assign sel_266462 = $signed({1'h0, add_266046, array_index_264599[1:0]}) < $signed({1'h0, sel_266048}) ? {add_266046, array_index_264599[1:0]} : sel_266048;
  assign add_266464 = array_index_265034[11:2] + 10'h36b;
  assign sel_266466 = $signed({1'h0, add_266050, array_index_264602[1:0]}) < $signed({1'h0, sel_266052}) ? {add_266050, array_index_264602[1:0]} : sel_266052;
  assign add_266468 = array_index_265463[11:2] + 10'h035;
  assign sel_266471 = $signed({1'h0, add_266054, array_index_265031[1:0]}) < $signed({1'h0, sel_266057}) ? {add_266054, array_index_265031[1:0]} : sel_266057;
  assign add_266473 = array_index_265466[11:2] + 10'h035;
  assign sel_266476 = $signed({1'h0, add_266059, array_index_265034[1:0]}) < $signed({1'h0, sel_266062}) ? {add_266059, array_index_265034[1:0]} : sel_266062;
  assign concat_266479 = {1'h0, ($signed({1'h0, add_265760}) < $signed({1'h0, sel_265762}) ? add_265760 : sel_265762) == ($signed({1'h0, add_265764}) < $signed({1'h0, sel_265766}) ? add_265764 : sel_265766)};
  assign add_266486 = array_index_258957[11:2] + 10'h29b;
  assign sel_266488 = $signed({1'h0, add_266078, array_index_258761[1:0]}) < $signed({1'h0, sel_266080}) ? {add_266078, array_index_258761[1:0]} : sel_266080;
  assign add_266490 = array_index_258960[11:2] + 10'h29b;
  assign sel_266492 = $signed({1'h0, add_266082, array_index_258764[1:0]}) < $signed({1'h0, sel_266084}) ? {add_266082, array_index_258764[1:0]} : sel_266084;
  assign add_266502 = array_index_259401[11:0] + 12'h9cf;
  assign sel_266504 = $signed({1'h0, add_266094}) < $signed({1'h0, sel_266096}) ? add_266094 : sel_266096;
  assign add_266506 = array_index_259404[11:0] + 12'h9cf;
  assign sel_266508 = $signed({1'h0, add_266098}) < $signed({1'h0, sel_266100}) ? add_266098 : sel_266100;
  assign add_266518 = array_index_259911[11:0] + 12'h30b;
  assign sel_266520 = $signed({1'h0, add_266110}) < $signed({1'h0, sel_266112}) ? add_266110 : sel_266112;
  assign add_266522 = array_index_259914[11:0] + 12'h30b;
  assign sel_266524 = $signed({1'h0, add_266114}) < $signed({1'h0, sel_266116}) ? add_266114 : sel_266116;
  assign add_266588 = concat_266479 + 2'h1;
  assign add_266598 = array_index_259171[11:0] + 12'hc05;
  assign sel_266600 = $signed({1'h0, add_266194}) < $signed({1'h0, sel_266196}) ? add_266194 : sel_266196;
  assign add_266602 = array_index_259174[11:0] + 12'hc05;
  assign sel_266604 = $signed({1'h0, add_266198}) < $signed({1'h0, sel_266200}) ? add_266198 : sel_266200;
  assign add_266616 = array_index_259647[11:0] + 12'h83f;
  assign sel_266618 = $signed({1'h0, add_266212}) < $signed({1'h0, sel_266214}) ? add_266212 : sel_266214;
  assign add_266620 = array_index_259650[11:0] + 12'h83f;
  assign sel_266622 = $signed({1'h0, add_266216}) < $signed({1'h0, sel_266218}) ? add_266216 : sel_266218;
  assign add_266634 = array_index_260195[11:1] + 11'h7b5;
  assign sel_266636 = $signed({1'h0, add_266230, array_index_259911[0]}) < $signed({1'h0, sel_266232}) ? {add_266230, array_index_259911[0]} : sel_266232;
  assign add_266638 = array_index_260198[11:1] + 11'h7b5;
  assign sel_266640 = $signed({1'h0, add_266234, array_index_259914[0]}) < $signed({1'h0, sel_266236}) ? {add_266234, array_index_259914[0]} : sel_266236;
  assign add_266710 = array_index_258957[11:0] + 12'hdab;
  assign sel_266712 = $signed({1'h0, add_266312}) < $signed({1'h0, sel_266314}) ? add_266312 : sel_266314;
  assign add_266714 = array_index_258960[11:0] + 12'hdab;
  assign sel_266716 = $signed({1'h0, add_266316}) < $signed({1'h0, sel_266318}) ? add_266316 : sel_266318;
  assign add_266728 = array_index_259401[11:2] + 10'h2b3;
  assign sel_266730 = $signed({1'h0, add_266330, array_index_259171[1:0]}) < $signed({1'h0, sel_266332}) ? {add_266330, array_index_259171[1:0]} : sel_266332;
  assign add_266732 = array_index_259404[11:2] + 10'h2b3;
  assign sel_266734 = $signed({1'h0, add_266334, array_index_259174[1:0]}) < $signed({1'h0, sel_266336}) ? {add_266334, array_index_259174[1:0]} : sel_266336;
  assign add_266744 = array_index_259911[11:1] + 11'h1e7;
  assign sel_266746 = $signed({1'h0, add_266346, array_index_259647[0]}) < $signed({1'h0, sel_266348}) ? {add_266346, array_index_259647[0]} : sel_266348;
  assign add_266748 = array_index_259914[11:1] + 11'h1e7;
  assign sel_266750 = $signed({1'h0, add_266350, array_index_259650[0]}) < $signed({1'h0, sel_266352}) ? {add_266350, array_index_259650[0]} : sel_266352;
  assign add_266760 = array_index_260507[11:0] + 12'h141;
  assign sel_266762 = $signed({1'h0, add_266362}) < $signed({1'h0, sel_266364}) ? add_266362 : sel_266364;
  assign add_266764 = array_index_260510[11:0] + 12'h141;
  assign sel_266766 = $signed({1'h0, add_266366}) < $signed({1'h0, sel_266368}) ? add_266366 : sel_266368;
  assign add_266768 = array_index_260845[11:1] + 11'h079;
  assign sel_266770 = $signed({1'h0, add_266370, array_index_260507[0]}) < $signed({1'h0, sel_266372}) ? {add_266370, array_index_260507[0]} : sel_266372;
  assign add_266772 = array_index_260848[11:1] + 11'h079;
  assign sel_266774 = $signed({1'h0, add_266374, array_index_260510[0]}) < $signed({1'h0, sel_266376}) ? {add_266374, array_index_260510[0]} : sel_266376;
  assign add_266776 = array_index_261207[11:0] + 12'h59d;
  assign sel_266778 = $signed({1'h0, add_266378}) < $signed({1'h0, sel_266380}) ? add_266378 : sel_266380;
  assign add_266780 = array_index_261210[11:0] + 12'h59d;
  assign sel_266782 = $signed({1'h0, add_266382}) < $signed({1'h0, sel_266384}) ? add_266382 : sel_266384;
  assign add_266784 = array_index_261595[11:0] + 12'ha6f;
  assign sel_266786 = $signed({1'h0, add_266386}) < $signed({1'h0, sel_266388}) ? add_266386 : sel_266388;
  assign add_266788 = array_index_261598[11:0] + 12'ha6f;
  assign sel_266790 = $signed({1'h0, add_266390}) < $signed({1'h0, sel_266392}) ? add_266390 : sel_266392;
  assign add_266792 = array_index_262007[11:1] + 11'h499;
  assign sel_266794 = $signed({1'h0, add_266394, array_index_261595[0]}) < $signed({1'h0, sel_266396}) ? {add_266394, array_index_261595[0]} : sel_266396;
  assign add_266796 = array_index_262010[11:1] + 11'h499;
  assign sel_266798 = $signed({1'h0, add_266398, array_index_261598[0]}) < $signed({1'h0, sel_266400}) ? {add_266398, array_index_261598[0]} : sel_266400;
  assign add_266800 = array_index_262439[11:1] + 11'h345;
  assign sel_266803 = $signed({1'h0, add_266402, array_index_262007[0]}) < $signed({1'h0, sel_266405}) ? {add_266402, array_index_262007[0]} : sel_266405;
  assign add_266805 = array_index_262442[11:1] + 11'h345;
  assign sel_266808 = $signed({1'h0, add_266407, array_index_262010[0]}) < $signed({1'h0, sel_266410}) ? {add_266407, array_index_262010[0]} : sel_266410;
  assign add_266810 = array_index_262871[11:0] + 12'h30f;
  assign sel_266812 = $signed({1'h0, add_266412}) < $signed({1'h0, sel_266414}) ? add_266412 : sel_266414;
  assign add_266814 = array_index_262874[11:0] + 12'h30f;
  assign sel_266816 = $signed({1'h0, add_266416}) < $signed({1'h0, sel_266418}) ? add_266416 : sel_266418;
  assign add_266818 = array_index_263303[11:0] + 12'hb55;
  assign sel_266820 = $signed({1'h0, add_266420}) < $signed({1'h0, sel_266422}) ? add_266420 : sel_266422;
  assign add_266822 = array_index_263306[11:0] + 12'hb55;
  assign sel_266824 = $signed({1'h0, add_266424}) < $signed({1'h0, sel_266426}) ? add_266424 : sel_266426;
  assign add_266826 = array_index_263735[11:0] + 12'h103;
  assign sel_266828 = $signed({1'h0, add_266428}) < $signed({1'h0, sel_266430}) ? add_266428 : sel_266430;
  assign add_266830 = array_index_263738[11:0] + 12'h103;
  assign sel_266832 = $signed({1'h0, add_266432}) < $signed({1'h0, sel_266434}) ? add_266432 : sel_266434;
  assign add_266834 = array_index_264167[11:0] + 12'hb01;
  assign sel_266836 = $signed({1'h0, add_266436}) < $signed({1'h0, sel_266438}) ? add_266436 : sel_266438;
  assign add_266838 = array_index_264170[11:0] + 12'hb01;
  assign sel_266840 = $signed({1'h0, add_266440}) < $signed({1'h0, sel_266442}) ? add_266440 : sel_266442;
  assign add_266842 = array_index_264599[11:0] + 12'h7b1;
  assign sel_266844 = $signed({1'h0, add_266444}) < $signed({1'h0, sel_266446}) ? add_266444 : sel_266446;
  assign add_266846 = array_index_264602[11:0] + 12'h7b1;
  assign sel_266848 = $signed({1'h0, add_266448}) < $signed({1'h0, sel_266450}) ? add_266448 : sel_266450;
  assign add_266850 = array_index_265031[11:0] + 12'h561;
  assign sel_266852 = $signed({1'h0, add_266452}) < $signed({1'h0, sel_266454}) ? add_266452 : sel_266454;
  assign add_266854 = array_index_265034[11:0] + 12'h561;
  assign sel_266856 = $signed({1'h0, add_266456}) < $signed({1'h0, sel_266458}) ? add_266456 : sel_266458;
  assign add_266858 = array_index_265463[11:2] + 10'h36b;
  assign sel_266860 = $signed({1'h0, add_266460, array_index_265031[1:0]}) < $signed({1'h0, sel_266462}) ? {add_266460, array_index_265031[1:0]} : sel_266462;
  assign add_266862 = array_index_265466[11:2] + 10'h36b;
  assign sel_266864 = $signed({1'h0, add_266464, array_index_265034[1:0]}) < $signed({1'h0, sel_266466}) ? {add_266464, array_index_265034[1:0]} : sel_266466;
  assign concat_266867 = {1'h0, ($signed({1'h0, add_266064}) < $signed({1'h0, sel_266066}) ? add_266064 : sel_266066) == ($signed({1'h0, add_266068}) < $signed({1'h0, sel_266070}) ? add_266068 : sel_266070) ? add_266588 : concat_266479};
  assign add_266874 = array_index_259171[11:2] + 10'h29b;
  assign sel_266876 = $signed({1'h0, add_266486, array_index_258957[1:0]}) < $signed({1'h0, sel_266488}) ? {add_266486, array_index_258957[1:0]} : sel_266488;
  assign add_266878 = array_index_259174[11:2] + 10'h29b;
  assign sel_266880 = $signed({1'h0, add_266490, array_index_258960[1:0]}) < $signed({1'h0, sel_266492}) ? {add_266490, array_index_258960[1:0]} : sel_266492;
  assign add_266890 = array_index_259647[11:0] + 12'h9cf;
  assign sel_266892 = $signed({1'h0, add_266502}) < $signed({1'h0, sel_266504}) ? add_266502 : sel_266504;
  assign add_266894 = array_index_259650[11:0] + 12'h9cf;
  assign sel_266896 = $signed({1'h0, add_266506}) < $signed({1'h0, sel_266508}) ? add_266506 : sel_266508;
  assign add_266906 = array_index_260195[11:0] + 12'h30b;
  assign sel_266908 = $signed({1'h0, add_266518}) < $signed({1'h0, sel_266520}) ? add_266518 : sel_266520;
  assign add_266910 = array_index_260198[11:0] + 12'h30b;
  assign sel_266912 = $signed({1'h0, add_266522}) < $signed({1'h0, sel_266524}) ? add_266522 : sel_266524;
  assign add_266972 = concat_266867 + 3'h1;
  assign add_266982 = array_index_259401[11:0] + 12'hc05;
  assign sel_266984 = $signed({1'h0, add_266598}) < $signed({1'h0, sel_266600}) ? add_266598 : sel_266600;
  assign add_266986 = array_index_259404[11:0] + 12'hc05;
  assign sel_266988 = $signed({1'h0, add_266602}) < $signed({1'h0, sel_266604}) ? add_266602 : sel_266604;
  assign add_267000 = array_index_259911[11:0] + 12'h83f;
  assign sel_267002 = $signed({1'h0, add_266616}) < $signed({1'h0, sel_266618}) ? add_266616 : sel_266618;
  assign add_267004 = array_index_259914[11:0] + 12'h83f;
  assign sel_267006 = $signed({1'h0, add_266620}) < $signed({1'h0, sel_266622}) ? add_266620 : sel_266622;
  assign add_267018 = array_index_260507[11:1] + 11'h7b5;
  assign sel_267020 = $signed({1'h0, add_266634, array_index_260195[0]}) < $signed({1'h0, sel_266636}) ? {add_266634, array_index_260195[0]} : sel_266636;
  assign add_267022 = array_index_260510[11:1] + 11'h7b5;
  assign sel_267024 = $signed({1'h0, add_266638, array_index_260198[0]}) < $signed({1'h0, sel_266640}) ? {add_266638, array_index_260198[0]} : sel_266640;
  assign add_267088 = array_index_259171[11:0] + 12'hdab;
  assign sel_267090 = $signed({1'h0, add_266710}) < $signed({1'h0, sel_266712}) ? add_266710 : sel_266712;
  assign add_267092 = array_index_259174[11:0] + 12'hdab;
  assign sel_267094 = $signed({1'h0, add_266714}) < $signed({1'h0, sel_266716}) ? add_266714 : sel_266716;
  assign add_267106 = array_index_259647[11:2] + 10'h2b3;
  assign sel_267108 = $signed({1'h0, add_266728, array_index_259401[1:0]}) < $signed({1'h0, sel_266730}) ? {add_266728, array_index_259401[1:0]} : sel_266730;
  assign add_267110 = array_index_259650[11:2] + 10'h2b3;
  assign sel_267112 = $signed({1'h0, add_266732, array_index_259404[1:0]}) < $signed({1'h0, sel_266734}) ? {add_266732, array_index_259404[1:0]} : sel_266734;
  assign add_267122 = array_index_260195[11:1] + 11'h1e7;
  assign sel_267124 = $signed({1'h0, add_266744, array_index_259911[0]}) < $signed({1'h0, sel_266746}) ? {add_266744, array_index_259911[0]} : sel_266746;
  assign add_267126 = array_index_260198[11:1] + 11'h1e7;
  assign sel_267128 = $signed({1'h0, add_266748, array_index_259914[0]}) < $signed({1'h0, sel_266750}) ? {add_266748, array_index_259914[0]} : sel_266750;
  assign add_267138 = array_index_260845[11:0] + 12'h141;
  assign sel_267140 = $signed({1'h0, add_266760}) < $signed({1'h0, sel_266762}) ? add_266760 : sel_266762;
  assign add_267142 = array_index_260848[11:0] + 12'h141;
  assign sel_267144 = $signed({1'h0, add_266764}) < $signed({1'h0, sel_266766}) ? add_266764 : sel_266766;
  assign add_267146 = array_index_261207[11:1] + 11'h079;
  assign sel_267148 = $signed({1'h0, add_266768, array_index_260845[0]}) < $signed({1'h0, sel_266770}) ? {add_266768, array_index_260845[0]} : sel_266770;
  assign add_267150 = array_index_261210[11:1] + 11'h079;
  assign sel_267152 = $signed({1'h0, add_266772, array_index_260848[0]}) < $signed({1'h0, sel_266774}) ? {add_266772, array_index_260848[0]} : sel_266774;
  assign add_267154 = array_index_261595[11:0] + 12'h59d;
  assign sel_267156 = $signed({1'h0, add_266776}) < $signed({1'h0, sel_266778}) ? add_266776 : sel_266778;
  assign add_267158 = array_index_261598[11:0] + 12'h59d;
  assign sel_267160 = $signed({1'h0, add_266780}) < $signed({1'h0, sel_266782}) ? add_266780 : sel_266782;
  assign add_267162 = array_index_262007[11:0] + 12'ha6f;
  assign sel_267164 = $signed({1'h0, add_266784}) < $signed({1'h0, sel_266786}) ? add_266784 : sel_266786;
  assign add_267166 = array_index_262010[11:0] + 12'ha6f;
  assign sel_267168 = $signed({1'h0, add_266788}) < $signed({1'h0, sel_266790}) ? add_266788 : sel_266790;
  assign add_267170 = array_index_262439[11:1] + 11'h499;
  assign sel_267172 = $signed({1'h0, add_266792, array_index_262007[0]}) < $signed({1'h0, sel_266794}) ? {add_266792, array_index_262007[0]} : sel_266794;
  assign add_267174 = array_index_262442[11:1] + 11'h499;
  assign sel_267176 = $signed({1'h0, add_266796, array_index_262010[0]}) < $signed({1'h0, sel_266798}) ? {add_266796, array_index_262010[0]} : sel_266798;
  assign add_267178 = array_index_262871[11:1] + 11'h345;
  assign sel_267181 = $signed({1'h0, add_266800, array_index_262439[0]}) < $signed({1'h0, sel_266803}) ? {add_266800, array_index_262439[0]} : sel_266803;
  assign add_267183 = array_index_262874[11:1] + 11'h345;
  assign sel_267186 = $signed({1'h0, add_266805, array_index_262442[0]}) < $signed({1'h0, sel_266808}) ? {add_266805, array_index_262442[0]} : sel_266808;
  assign add_267188 = array_index_263303[11:0] + 12'h30f;
  assign sel_267190 = $signed({1'h0, add_266810}) < $signed({1'h0, sel_266812}) ? add_266810 : sel_266812;
  assign add_267192 = array_index_263306[11:0] + 12'h30f;
  assign sel_267194 = $signed({1'h0, add_266814}) < $signed({1'h0, sel_266816}) ? add_266814 : sel_266816;
  assign add_267196 = array_index_263735[11:0] + 12'hb55;
  assign sel_267198 = $signed({1'h0, add_266818}) < $signed({1'h0, sel_266820}) ? add_266818 : sel_266820;
  assign add_267200 = array_index_263738[11:0] + 12'hb55;
  assign sel_267202 = $signed({1'h0, add_266822}) < $signed({1'h0, sel_266824}) ? add_266822 : sel_266824;
  assign add_267204 = array_index_264167[11:0] + 12'h103;
  assign sel_267206 = $signed({1'h0, add_266826}) < $signed({1'h0, sel_266828}) ? add_266826 : sel_266828;
  assign add_267208 = array_index_264170[11:0] + 12'h103;
  assign sel_267210 = $signed({1'h0, add_266830}) < $signed({1'h0, sel_266832}) ? add_266830 : sel_266832;
  assign add_267212 = array_index_264599[11:0] + 12'hb01;
  assign sel_267214 = $signed({1'h0, add_266834}) < $signed({1'h0, sel_266836}) ? add_266834 : sel_266836;
  assign add_267216 = array_index_264602[11:0] + 12'hb01;
  assign sel_267218 = $signed({1'h0, add_266838}) < $signed({1'h0, sel_266840}) ? add_266838 : sel_266840;
  assign add_267220 = array_index_265031[11:0] + 12'h7b1;
  assign sel_267222 = $signed({1'h0, add_266842}) < $signed({1'h0, sel_266844}) ? add_266842 : sel_266844;
  assign add_267224 = array_index_265034[11:0] + 12'h7b1;
  assign sel_267226 = $signed({1'h0, add_266846}) < $signed({1'h0, sel_266848}) ? add_266846 : sel_266848;
  assign add_267228 = array_index_265463[11:0] + 12'h561;
  assign sel_267230 = $signed({1'h0, add_266850}) < $signed({1'h0, sel_266852}) ? add_266850 : sel_266852;
  assign add_267232 = array_index_265466[11:0] + 12'h561;
  assign sel_267234 = $signed({1'h0, add_266854}) < $signed({1'h0, sel_266856}) ? add_266854 : sel_266856;
  assign concat_267237 = {1'h0, ($signed({1'h0, add_266468, array_index_265463[1:0]}) < $signed({1'h0, sel_266471}) ? {add_266468, array_index_265463[1:0]} : sel_266471) == ($signed({1'h0, add_266473, array_index_265466[1:0]}) < $signed({1'h0, sel_266476}) ? {add_266473, array_index_265466[1:0]} : sel_266476) ? add_266972 : concat_266867};
  assign add_267244 = array_index_259401[11:2] + 10'h29b;
  assign sel_267246 = $signed({1'h0, add_266874, array_index_259171[1:0]}) < $signed({1'h0, sel_266876}) ? {add_266874, array_index_259171[1:0]} : sel_266876;
  assign add_267248 = array_index_259404[11:2] + 10'h29b;
  assign sel_267250 = $signed({1'h0, add_266878, array_index_259174[1:0]}) < $signed({1'h0, sel_266880}) ? {add_266878, array_index_259174[1:0]} : sel_266880;
  assign add_267260 = array_index_259911[11:0] + 12'h9cf;
  assign sel_267262 = $signed({1'h0, add_266890}) < $signed({1'h0, sel_266892}) ? add_266890 : sel_266892;
  assign add_267264 = array_index_259914[11:0] + 12'h9cf;
  assign sel_267266 = $signed({1'h0, add_266894}) < $signed({1'h0, sel_266896}) ? add_266894 : sel_266896;
  assign add_267276 = array_index_260507[11:0] + 12'h30b;
  assign sel_267278 = $signed({1'h0, add_266906}) < $signed({1'h0, sel_266908}) ? add_266906 : sel_266908;
  assign add_267280 = array_index_260510[11:0] + 12'h30b;
  assign sel_267282 = $signed({1'h0, add_266910}) < $signed({1'h0, sel_266912}) ? add_266910 : sel_266912;
  assign add_267338 = concat_267237 + 4'h1;
  assign add_267348 = array_index_259647[11:0] + 12'hc05;
  assign sel_267350 = $signed({1'h0, add_266982}) < $signed({1'h0, sel_266984}) ? add_266982 : sel_266984;
  assign add_267352 = array_index_259650[11:0] + 12'hc05;
  assign sel_267354 = $signed({1'h0, add_266986}) < $signed({1'h0, sel_266988}) ? add_266986 : sel_266988;
  assign add_267366 = array_index_260195[11:0] + 12'h83f;
  assign sel_267368 = $signed({1'h0, add_267000}) < $signed({1'h0, sel_267002}) ? add_267000 : sel_267002;
  assign add_267370 = array_index_260198[11:0] + 12'h83f;
  assign sel_267372 = $signed({1'h0, add_267004}) < $signed({1'h0, sel_267006}) ? add_267004 : sel_267006;
  assign add_267384 = array_index_260845[11:1] + 11'h7b5;
  assign sel_267386 = $signed({1'h0, add_267018, array_index_260507[0]}) < $signed({1'h0, sel_267020}) ? {add_267018, array_index_260507[0]} : sel_267020;
  assign add_267388 = array_index_260848[11:1] + 11'h7b5;
  assign sel_267390 = $signed({1'h0, add_267022, array_index_260510[0]}) < $signed({1'h0, sel_267024}) ? {add_267022, array_index_260510[0]} : sel_267024;
  assign add_267448 = array_index_259401[11:0] + 12'hdab;
  assign sel_267450 = $signed({1'h0, add_267088}) < $signed({1'h0, sel_267090}) ? add_267088 : sel_267090;
  assign add_267452 = array_index_259404[11:0] + 12'hdab;
  assign sel_267454 = $signed({1'h0, add_267092}) < $signed({1'h0, sel_267094}) ? add_267092 : sel_267094;
  assign add_267466 = array_index_259911[11:2] + 10'h2b3;
  assign sel_267468 = $signed({1'h0, add_267106, array_index_259647[1:0]}) < $signed({1'h0, sel_267108}) ? {add_267106, array_index_259647[1:0]} : sel_267108;
  assign add_267470 = array_index_259914[11:2] + 10'h2b3;
  assign sel_267472 = $signed({1'h0, add_267110, array_index_259650[1:0]}) < $signed({1'h0, sel_267112}) ? {add_267110, array_index_259650[1:0]} : sel_267112;
  assign add_267482 = array_index_260507[11:1] + 11'h1e7;
  assign sel_267484 = $signed({1'h0, add_267122, array_index_260195[0]}) < $signed({1'h0, sel_267124}) ? {add_267122, array_index_260195[0]} : sel_267124;
  assign add_267486 = array_index_260510[11:1] + 11'h1e7;
  assign sel_267488 = $signed({1'h0, add_267126, array_index_260198[0]}) < $signed({1'h0, sel_267128}) ? {add_267126, array_index_260198[0]} : sel_267128;
  assign add_267498 = array_index_261207[11:0] + 12'h141;
  assign sel_267500 = $signed({1'h0, add_267138}) < $signed({1'h0, sel_267140}) ? add_267138 : sel_267140;
  assign add_267502 = array_index_261210[11:0] + 12'h141;
  assign sel_267504 = $signed({1'h0, add_267142}) < $signed({1'h0, sel_267144}) ? add_267142 : sel_267144;
  assign add_267506 = array_index_261595[11:1] + 11'h079;
  assign sel_267508 = $signed({1'h0, add_267146, array_index_261207[0]}) < $signed({1'h0, sel_267148}) ? {add_267146, array_index_261207[0]} : sel_267148;
  assign add_267510 = array_index_261598[11:1] + 11'h079;
  assign sel_267512 = $signed({1'h0, add_267150, array_index_261210[0]}) < $signed({1'h0, sel_267152}) ? {add_267150, array_index_261210[0]} : sel_267152;
  assign add_267514 = array_index_262007[11:0] + 12'h59d;
  assign sel_267516 = $signed({1'h0, add_267154}) < $signed({1'h0, sel_267156}) ? add_267154 : sel_267156;
  assign add_267518 = array_index_262010[11:0] + 12'h59d;
  assign sel_267520 = $signed({1'h0, add_267158}) < $signed({1'h0, sel_267160}) ? add_267158 : sel_267160;
  assign add_267522 = array_index_262439[11:0] + 12'ha6f;
  assign sel_267524 = $signed({1'h0, add_267162}) < $signed({1'h0, sel_267164}) ? add_267162 : sel_267164;
  assign add_267526 = array_index_262442[11:0] + 12'ha6f;
  assign sel_267528 = $signed({1'h0, add_267166}) < $signed({1'h0, sel_267168}) ? add_267166 : sel_267168;
  assign add_267530 = array_index_262871[11:1] + 11'h499;
  assign sel_267532 = $signed({1'h0, add_267170, array_index_262439[0]}) < $signed({1'h0, sel_267172}) ? {add_267170, array_index_262439[0]} : sel_267172;
  assign add_267534 = array_index_262874[11:1] + 11'h499;
  assign sel_267536 = $signed({1'h0, add_267174, array_index_262442[0]}) < $signed({1'h0, sel_267176}) ? {add_267174, array_index_262442[0]} : sel_267176;
  assign add_267538 = array_index_263303[11:1] + 11'h345;
  assign sel_267541 = $signed({1'h0, add_267178, array_index_262871[0]}) < $signed({1'h0, sel_267181}) ? {add_267178, array_index_262871[0]} : sel_267181;
  assign add_267543 = array_index_263306[11:1] + 11'h345;
  assign sel_267546 = $signed({1'h0, add_267183, array_index_262874[0]}) < $signed({1'h0, sel_267186}) ? {add_267183, array_index_262874[0]} : sel_267186;
  assign add_267548 = array_index_263735[11:0] + 12'h30f;
  assign sel_267550 = $signed({1'h0, add_267188}) < $signed({1'h0, sel_267190}) ? add_267188 : sel_267190;
  assign add_267552 = array_index_263738[11:0] + 12'h30f;
  assign sel_267554 = $signed({1'h0, add_267192}) < $signed({1'h0, sel_267194}) ? add_267192 : sel_267194;
  assign add_267556 = array_index_264167[11:0] + 12'hb55;
  assign sel_267558 = $signed({1'h0, add_267196}) < $signed({1'h0, sel_267198}) ? add_267196 : sel_267198;
  assign add_267560 = array_index_264170[11:0] + 12'hb55;
  assign sel_267562 = $signed({1'h0, add_267200}) < $signed({1'h0, sel_267202}) ? add_267200 : sel_267202;
  assign add_267564 = array_index_264599[11:0] + 12'h103;
  assign sel_267566 = $signed({1'h0, add_267204}) < $signed({1'h0, sel_267206}) ? add_267204 : sel_267206;
  assign add_267568 = array_index_264602[11:0] + 12'h103;
  assign sel_267570 = $signed({1'h0, add_267208}) < $signed({1'h0, sel_267210}) ? add_267208 : sel_267210;
  assign add_267572 = array_index_265031[11:0] + 12'hb01;
  assign sel_267574 = $signed({1'h0, add_267212}) < $signed({1'h0, sel_267214}) ? add_267212 : sel_267214;
  assign add_267576 = array_index_265034[11:0] + 12'hb01;
  assign sel_267578 = $signed({1'h0, add_267216}) < $signed({1'h0, sel_267218}) ? add_267216 : sel_267218;
  assign add_267580 = array_index_265463[11:0] + 12'h7b1;
  assign sel_267582 = $signed({1'h0, add_267220}) < $signed({1'h0, sel_267222}) ? add_267220 : sel_267222;
  assign add_267584 = array_index_265466[11:0] + 12'h7b1;
  assign sel_267586 = $signed({1'h0, add_267224}) < $signed({1'h0, sel_267226}) ? add_267224 : sel_267226;
  assign concat_267589 = {1'h0, ($signed({1'h0, add_266858, array_index_265463[1:0]}) < $signed({1'h0, sel_266860}) ? {add_266858, array_index_265463[1:0]} : sel_266860) == ($signed({1'h0, add_266862, array_index_265466[1:0]}) < $signed({1'h0, sel_266864}) ? {add_266862, array_index_265466[1:0]} : sel_266864) ? add_267338 : concat_267237};
  assign add_267596 = array_index_259647[11:2] + 10'h29b;
  assign sel_267598 = $signed({1'h0, add_267244, array_index_259401[1:0]}) < $signed({1'h0, sel_267246}) ? {add_267244, array_index_259401[1:0]} : sel_267246;
  assign add_267600 = array_index_259650[11:2] + 10'h29b;
  assign sel_267602 = $signed({1'h0, add_267248, array_index_259404[1:0]}) < $signed({1'h0, sel_267250}) ? {add_267248, array_index_259404[1:0]} : sel_267250;
  assign add_267612 = array_index_260195[11:0] + 12'h9cf;
  assign sel_267614 = $signed({1'h0, add_267260}) < $signed({1'h0, sel_267262}) ? add_267260 : sel_267262;
  assign add_267616 = array_index_260198[11:0] + 12'h9cf;
  assign sel_267618 = $signed({1'h0, add_267264}) < $signed({1'h0, sel_267266}) ? add_267264 : sel_267266;
  assign add_267628 = array_index_260845[11:0] + 12'h30b;
  assign sel_267630 = $signed({1'h0, add_267276}) < $signed({1'h0, sel_267278}) ? add_267276 : sel_267278;
  assign add_267632 = array_index_260848[11:0] + 12'h30b;
  assign sel_267634 = $signed({1'h0, add_267280}) < $signed({1'h0, sel_267282}) ? add_267280 : sel_267282;
  assign add_267686 = concat_267589 + 5'h01;
  assign add_267696 = array_index_259911[11:0] + 12'hc05;
  assign sel_267698 = $signed({1'h0, add_267348}) < $signed({1'h0, sel_267350}) ? add_267348 : sel_267350;
  assign add_267700 = array_index_259914[11:0] + 12'hc05;
  assign sel_267702 = $signed({1'h0, add_267352}) < $signed({1'h0, sel_267354}) ? add_267352 : sel_267354;
  assign add_267714 = array_index_260507[11:0] + 12'h83f;
  assign sel_267716 = $signed({1'h0, add_267366}) < $signed({1'h0, sel_267368}) ? add_267366 : sel_267368;
  assign add_267718 = array_index_260510[11:0] + 12'h83f;
  assign sel_267720 = $signed({1'h0, add_267370}) < $signed({1'h0, sel_267372}) ? add_267370 : sel_267372;
  assign add_267732 = array_index_261207[11:1] + 11'h7b5;
  assign sel_267734 = $signed({1'h0, add_267384, array_index_260845[0]}) < $signed({1'h0, sel_267386}) ? {add_267384, array_index_260845[0]} : sel_267386;
  assign add_267736 = array_index_261210[11:1] + 11'h7b5;
  assign sel_267738 = $signed({1'h0, add_267388, array_index_260848[0]}) < $signed({1'h0, sel_267390}) ? {add_267388, array_index_260848[0]} : sel_267390;
  assign add_267792 = array_index_259647[11:0] + 12'hdab;
  assign sel_267794 = $signed({1'h0, add_267448}) < $signed({1'h0, sel_267450}) ? add_267448 : sel_267450;
  assign add_267796 = array_index_259650[11:0] + 12'hdab;
  assign sel_267798 = $signed({1'h0, add_267452}) < $signed({1'h0, sel_267454}) ? add_267452 : sel_267454;
  assign add_267810 = array_index_260195[11:2] + 10'h2b3;
  assign sel_267812 = $signed({1'h0, add_267466, array_index_259911[1:0]}) < $signed({1'h0, sel_267468}) ? {add_267466, array_index_259911[1:0]} : sel_267468;
  assign add_267814 = array_index_260198[11:2] + 10'h2b3;
  assign sel_267816 = $signed({1'h0, add_267470, array_index_259914[1:0]}) < $signed({1'h0, sel_267472}) ? {add_267470, array_index_259914[1:0]} : sel_267472;
  assign add_267826 = array_index_260845[11:1] + 11'h1e7;
  assign sel_267828 = $signed({1'h0, add_267482, array_index_260507[0]}) < $signed({1'h0, sel_267484}) ? {add_267482, array_index_260507[0]} : sel_267484;
  assign add_267830 = array_index_260848[11:1] + 11'h1e7;
  assign sel_267832 = $signed({1'h0, add_267486, array_index_260510[0]}) < $signed({1'h0, sel_267488}) ? {add_267486, array_index_260510[0]} : sel_267488;
  assign add_267842 = array_index_261595[11:0] + 12'h141;
  assign sel_267844 = $signed({1'h0, add_267498}) < $signed({1'h0, sel_267500}) ? add_267498 : sel_267500;
  assign add_267846 = array_index_261598[11:0] + 12'h141;
  assign sel_267848 = $signed({1'h0, add_267502}) < $signed({1'h0, sel_267504}) ? add_267502 : sel_267504;
  assign add_267850 = array_index_262007[11:1] + 11'h079;
  assign sel_267852 = $signed({1'h0, add_267506, array_index_261595[0]}) < $signed({1'h0, sel_267508}) ? {add_267506, array_index_261595[0]} : sel_267508;
  assign add_267854 = array_index_262010[11:1] + 11'h079;
  assign sel_267856 = $signed({1'h0, add_267510, array_index_261598[0]}) < $signed({1'h0, sel_267512}) ? {add_267510, array_index_261598[0]} : sel_267512;
  assign add_267858 = array_index_262439[11:0] + 12'h59d;
  assign sel_267860 = $signed({1'h0, add_267514}) < $signed({1'h0, sel_267516}) ? add_267514 : sel_267516;
  assign add_267862 = array_index_262442[11:0] + 12'h59d;
  assign sel_267864 = $signed({1'h0, add_267518}) < $signed({1'h0, sel_267520}) ? add_267518 : sel_267520;
  assign add_267866 = array_index_262871[11:0] + 12'ha6f;
  assign sel_267868 = $signed({1'h0, add_267522}) < $signed({1'h0, sel_267524}) ? add_267522 : sel_267524;
  assign add_267870 = array_index_262874[11:0] + 12'ha6f;
  assign sel_267872 = $signed({1'h0, add_267526}) < $signed({1'h0, sel_267528}) ? add_267526 : sel_267528;
  assign add_267874 = array_index_263303[11:1] + 11'h499;
  assign sel_267876 = $signed({1'h0, add_267530, array_index_262871[0]}) < $signed({1'h0, sel_267532}) ? {add_267530, array_index_262871[0]} : sel_267532;
  assign add_267878 = array_index_263306[11:1] + 11'h499;
  assign sel_267880 = $signed({1'h0, add_267534, array_index_262874[0]}) < $signed({1'h0, sel_267536}) ? {add_267534, array_index_262874[0]} : sel_267536;
  assign add_267882 = array_index_263735[11:1] + 11'h345;
  assign sel_267885 = $signed({1'h0, add_267538, array_index_263303[0]}) < $signed({1'h0, sel_267541}) ? {add_267538, array_index_263303[0]} : sel_267541;
  assign add_267887 = array_index_263738[11:1] + 11'h345;
  assign sel_267890 = $signed({1'h0, add_267543, array_index_263306[0]}) < $signed({1'h0, sel_267546}) ? {add_267543, array_index_263306[0]} : sel_267546;
  assign add_267892 = array_index_264167[11:0] + 12'h30f;
  assign sel_267894 = $signed({1'h0, add_267548}) < $signed({1'h0, sel_267550}) ? add_267548 : sel_267550;
  assign add_267896 = array_index_264170[11:0] + 12'h30f;
  assign sel_267898 = $signed({1'h0, add_267552}) < $signed({1'h0, sel_267554}) ? add_267552 : sel_267554;
  assign add_267900 = array_index_264599[11:0] + 12'hb55;
  assign sel_267902 = $signed({1'h0, add_267556}) < $signed({1'h0, sel_267558}) ? add_267556 : sel_267558;
  assign add_267904 = array_index_264602[11:0] + 12'hb55;
  assign sel_267906 = $signed({1'h0, add_267560}) < $signed({1'h0, sel_267562}) ? add_267560 : sel_267562;
  assign add_267908 = array_index_265031[11:0] + 12'h103;
  assign sel_267910 = $signed({1'h0, add_267564}) < $signed({1'h0, sel_267566}) ? add_267564 : sel_267566;
  assign add_267912 = array_index_265034[11:0] + 12'h103;
  assign sel_267914 = $signed({1'h0, add_267568}) < $signed({1'h0, sel_267570}) ? add_267568 : sel_267570;
  assign add_267916 = array_index_265463[11:0] + 12'hb01;
  assign sel_267918 = $signed({1'h0, add_267572}) < $signed({1'h0, sel_267574}) ? add_267572 : sel_267574;
  assign add_267920 = array_index_265466[11:0] + 12'hb01;
  assign sel_267922 = $signed({1'h0, add_267576}) < $signed({1'h0, sel_267578}) ? add_267576 : sel_267578;
  assign concat_267925 = {1'h0, ($signed({1'h0, add_267228}) < $signed({1'h0, sel_267230}) ? add_267228 : sel_267230) == ($signed({1'h0, add_267232}) < $signed({1'h0, sel_267234}) ? add_267232 : sel_267234) ? add_267686 : concat_267589};
  assign add_267932 = array_index_259911[11:2] + 10'h29b;
  assign sel_267934 = $signed({1'h0, add_267596, array_index_259647[1:0]}) < $signed({1'h0, sel_267598}) ? {add_267596, array_index_259647[1:0]} : sel_267598;
  assign add_267936 = array_index_259914[11:2] + 10'h29b;
  assign sel_267938 = $signed({1'h0, add_267600, array_index_259650[1:0]}) < $signed({1'h0, sel_267602}) ? {add_267600, array_index_259650[1:0]} : sel_267602;
  assign add_267948 = array_index_260507[11:0] + 12'h9cf;
  assign sel_267950 = $signed({1'h0, add_267612}) < $signed({1'h0, sel_267614}) ? add_267612 : sel_267614;
  assign add_267952 = array_index_260510[11:0] + 12'h9cf;
  assign sel_267954 = $signed({1'h0, add_267616}) < $signed({1'h0, sel_267618}) ? add_267616 : sel_267618;
  assign add_267964 = array_index_261207[11:0] + 12'h30b;
  assign sel_267966 = $signed({1'h0, add_267628}) < $signed({1'h0, sel_267630}) ? add_267628 : sel_267630;
  assign add_267968 = array_index_261210[11:0] + 12'h30b;
  assign sel_267970 = $signed({1'h0, add_267632}) < $signed({1'h0, sel_267634}) ? add_267632 : sel_267634;
  assign add_268018 = concat_267925 + 6'h01;
  assign add_268028 = array_index_260195[11:0] + 12'hc05;
  assign sel_268030 = $signed({1'h0, add_267696}) < $signed({1'h0, sel_267698}) ? add_267696 : sel_267698;
  assign add_268032 = array_index_260198[11:0] + 12'hc05;
  assign sel_268034 = $signed({1'h0, add_267700}) < $signed({1'h0, sel_267702}) ? add_267700 : sel_267702;
  assign add_268046 = array_index_260845[11:0] + 12'h83f;
  assign sel_268048 = $signed({1'h0, add_267714}) < $signed({1'h0, sel_267716}) ? add_267714 : sel_267716;
  assign add_268050 = array_index_260848[11:0] + 12'h83f;
  assign sel_268052 = $signed({1'h0, add_267718}) < $signed({1'h0, sel_267720}) ? add_267718 : sel_267720;
  assign add_268064 = array_index_261595[11:1] + 11'h7b5;
  assign sel_268066 = $signed({1'h0, add_267732, array_index_261207[0]}) < $signed({1'h0, sel_267734}) ? {add_267732, array_index_261207[0]} : sel_267734;
  assign add_268068 = array_index_261598[11:1] + 11'h7b5;
  assign sel_268070 = $signed({1'h0, add_267736, array_index_261210[0]}) < $signed({1'h0, sel_267738}) ? {add_267736, array_index_261210[0]} : sel_267738;
  assign add_268120 = array_index_259911[11:0] + 12'hdab;
  assign sel_268122 = $signed({1'h0, add_267792}) < $signed({1'h0, sel_267794}) ? add_267792 : sel_267794;
  assign add_268124 = array_index_259914[11:0] + 12'hdab;
  assign sel_268126 = $signed({1'h0, add_267796}) < $signed({1'h0, sel_267798}) ? add_267796 : sel_267798;
  assign add_268138 = array_index_260507[11:2] + 10'h2b3;
  assign sel_268140 = $signed({1'h0, add_267810, array_index_260195[1:0]}) < $signed({1'h0, sel_267812}) ? {add_267810, array_index_260195[1:0]} : sel_267812;
  assign add_268142 = array_index_260510[11:2] + 10'h2b3;
  assign sel_268144 = $signed({1'h0, add_267814, array_index_260198[1:0]}) < $signed({1'h0, sel_267816}) ? {add_267814, array_index_260198[1:0]} : sel_267816;
  assign add_268154 = array_index_261207[11:1] + 11'h1e7;
  assign sel_268156 = $signed({1'h0, add_267826, array_index_260845[0]}) < $signed({1'h0, sel_267828}) ? {add_267826, array_index_260845[0]} : sel_267828;
  assign add_268158 = array_index_261210[11:1] + 11'h1e7;
  assign sel_268160 = $signed({1'h0, add_267830, array_index_260848[0]}) < $signed({1'h0, sel_267832}) ? {add_267830, array_index_260848[0]} : sel_267832;
  assign add_268170 = array_index_262007[11:0] + 12'h141;
  assign sel_268172 = $signed({1'h0, add_267842}) < $signed({1'h0, sel_267844}) ? add_267842 : sel_267844;
  assign add_268174 = array_index_262010[11:0] + 12'h141;
  assign sel_268176 = $signed({1'h0, add_267846}) < $signed({1'h0, sel_267848}) ? add_267846 : sel_267848;
  assign add_268178 = array_index_262439[11:1] + 11'h079;
  assign sel_268180 = $signed({1'h0, add_267850, array_index_262007[0]}) < $signed({1'h0, sel_267852}) ? {add_267850, array_index_262007[0]} : sel_267852;
  assign add_268182 = array_index_262442[11:1] + 11'h079;
  assign sel_268184 = $signed({1'h0, add_267854, array_index_262010[0]}) < $signed({1'h0, sel_267856}) ? {add_267854, array_index_262010[0]} : sel_267856;
  assign add_268186 = array_index_262871[11:0] + 12'h59d;
  assign sel_268188 = $signed({1'h0, add_267858}) < $signed({1'h0, sel_267860}) ? add_267858 : sel_267860;
  assign add_268190 = array_index_262874[11:0] + 12'h59d;
  assign sel_268192 = $signed({1'h0, add_267862}) < $signed({1'h0, sel_267864}) ? add_267862 : sel_267864;
  assign add_268194 = array_index_263303[11:0] + 12'ha6f;
  assign sel_268196 = $signed({1'h0, add_267866}) < $signed({1'h0, sel_267868}) ? add_267866 : sel_267868;
  assign add_268198 = array_index_263306[11:0] + 12'ha6f;
  assign sel_268200 = $signed({1'h0, add_267870}) < $signed({1'h0, sel_267872}) ? add_267870 : sel_267872;
  assign add_268202 = array_index_263735[11:1] + 11'h499;
  assign sel_268204 = $signed({1'h0, add_267874, array_index_263303[0]}) < $signed({1'h0, sel_267876}) ? {add_267874, array_index_263303[0]} : sel_267876;
  assign add_268206 = array_index_263738[11:1] + 11'h499;
  assign sel_268208 = $signed({1'h0, add_267878, array_index_263306[0]}) < $signed({1'h0, sel_267880}) ? {add_267878, array_index_263306[0]} : sel_267880;
  assign add_268210 = array_index_264167[11:1] + 11'h345;
  assign sel_268213 = $signed({1'h0, add_267882, array_index_263735[0]}) < $signed({1'h0, sel_267885}) ? {add_267882, array_index_263735[0]} : sel_267885;
  assign add_268215 = array_index_264170[11:1] + 11'h345;
  assign sel_268218 = $signed({1'h0, add_267887, array_index_263738[0]}) < $signed({1'h0, sel_267890}) ? {add_267887, array_index_263738[0]} : sel_267890;
  assign add_268220 = array_index_264599[11:0] + 12'h30f;
  assign sel_268222 = $signed({1'h0, add_267892}) < $signed({1'h0, sel_267894}) ? add_267892 : sel_267894;
  assign add_268224 = array_index_264602[11:0] + 12'h30f;
  assign sel_268226 = $signed({1'h0, add_267896}) < $signed({1'h0, sel_267898}) ? add_267896 : sel_267898;
  assign add_268228 = array_index_265031[11:0] + 12'hb55;
  assign sel_268230 = $signed({1'h0, add_267900}) < $signed({1'h0, sel_267902}) ? add_267900 : sel_267902;
  assign add_268232 = array_index_265034[11:0] + 12'hb55;
  assign sel_268234 = $signed({1'h0, add_267904}) < $signed({1'h0, sel_267906}) ? add_267904 : sel_267906;
  assign add_268236 = array_index_265463[11:0] + 12'h103;
  assign sel_268238 = $signed({1'h0, add_267908}) < $signed({1'h0, sel_267910}) ? add_267908 : sel_267910;
  assign add_268240 = array_index_265466[11:0] + 12'h103;
  assign sel_268242 = $signed({1'h0, add_267912}) < $signed({1'h0, sel_267914}) ? add_267912 : sel_267914;
  assign concat_268245 = {1'h0, ($signed({1'h0, add_267580}) < $signed({1'h0, sel_267582}) ? add_267580 : sel_267582) == ($signed({1'h0, add_267584}) < $signed({1'h0, sel_267586}) ? add_267584 : sel_267586) ? add_268018 : concat_267925};
  assign add_268252 = array_index_260195[11:2] + 10'h29b;
  assign sel_268254 = $signed({1'h0, add_267932, array_index_259911[1:0]}) < $signed({1'h0, sel_267934}) ? {add_267932, array_index_259911[1:0]} : sel_267934;
  assign add_268256 = array_index_260198[11:2] + 10'h29b;
  assign sel_268258 = $signed({1'h0, add_267936, array_index_259914[1:0]}) < $signed({1'h0, sel_267938}) ? {add_267936, array_index_259914[1:0]} : sel_267938;
  assign add_268268 = array_index_260845[11:0] + 12'h9cf;
  assign sel_268270 = $signed({1'h0, add_267948}) < $signed({1'h0, sel_267950}) ? add_267948 : sel_267950;
  assign add_268272 = array_index_260848[11:0] + 12'h9cf;
  assign sel_268274 = $signed({1'h0, add_267952}) < $signed({1'h0, sel_267954}) ? add_267952 : sel_267954;
  assign add_268284 = array_index_261595[11:0] + 12'h30b;
  assign sel_268286 = $signed({1'h0, add_267964}) < $signed({1'h0, sel_267966}) ? add_267964 : sel_267966;
  assign add_268288 = array_index_261598[11:0] + 12'h30b;
  assign sel_268290 = $signed({1'h0, add_267968}) < $signed({1'h0, sel_267970}) ? add_267968 : sel_267970;
  assign add_268334 = concat_268245 + 7'h01;
  assign add_268344 = array_index_260507[11:0] + 12'hc05;
  assign sel_268346 = $signed({1'h0, add_268028}) < $signed({1'h0, sel_268030}) ? add_268028 : sel_268030;
  assign add_268348 = array_index_260510[11:0] + 12'hc05;
  assign sel_268350 = $signed({1'h0, add_268032}) < $signed({1'h0, sel_268034}) ? add_268032 : sel_268034;
  assign add_268362 = array_index_261207[11:0] + 12'h83f;
  assign sel_268364 = $signed({1'h0, add_268046}) < $signed({1'h0, sel_268048}) ? add_268046 : sel_268048;
  assign add_268366 = array_index_261210[11:0] + 12'h83f;
  assign sel_268368 = $signed({1'h0, add_268050}) < $signed({1'h0, sel_268052}) ? add_268050 : sel_268052;
  assign add_268380 = array_index_262007[11:1] + 11'h7b5;
  assign sel_268382 = $signed({1'h0, add_268064, array_index_261595[0]}) < $signed({1'h0, sel_268066}) ? {add_268064, array_index_261595[0]} : sel_268066;
  assign add_268384 = array_index_262010[11:1] + 11'h7b5;
  assign sel_268386 = $signed({1'h0, add_268068, array_index_261598[0]}) < $signed({1'h0, sel_268070}) ? {add_268068, array_index_261598[0]} : sel_268070;
  assign add_268432 = array_index_260195[11:0] + 12'hdab;
  assign sel_268434 = $signed({1'h0, add_268120}) < $signed({1'h0, sel_268122}) ? add_268120 : sel_268122;
  assign add_268436 = array_index_260198[11:0] + 12'hdab;
  assign sel_268438 = $signed({1'h0, add_268124}) < $signed({1'h0, sel_268126}) ? add_268124 : sel_268126;
  assign add_268450 = array_index_260845[11:2] + 10'h2b3;
  assign sel_268452 = $signed({1'h0, add_268138, array_index_260507[1:0]}) < $signed({1'h0, sel_268140}) ? {add_268138, array_index_260507[1:0]} : sel_268140;
  assign add_268454 = array_index_260848[11:2] + 10'h2b3;
  assign sel_268456 = $signed({1'h0, add_268142, array_index_260510[1:0]}) < $signed({1'h0, sel_268144}) ? {add_268142, array_index_260510[1:0]} : sel_268144;
  assign add_268466 = array_index_261595[11:1] + 11'h1e7;
  assign sel_268468 = $signed({1'h0, add_268154, array_index_261207[0]}) < $signed({1'h0, sel_268156}) ? {add_268154, array_index_261207[0]} : sel_268156;
  assign add_268470 = array_index_261598[11:1] + 11'h1e7;
  assign sel_268472 = $signed({1'h0, add_268158, array_index_261210[0]}) < $signed({1'h0, sel_268160}) ? {add_268158, array_index_261210[0]} : sel_268160;
  assign add_268482 = array_index_262439[11:0] + 12'h141;
  assign sel_268484 = $signed({1'h0, add_268170}) < $signed({1'h0, sel_268172}) ? add_268170 : sel_268172;
  assign add_268486 = array_index_262442[11:0] + 12'h141;
  assign sel_268488 = $signed({1'h0, add_268174}) < $signed({1'h0, sel_268176}) ? add_268174 : sel_268176;
  assign add_268490 = array_index_262871[11:1] + 11'h079;
  assign sel_268492 = $signed({1'h0, add_268178, array_index_262439[0]}) < $signed({1'h0, sel_268180}) ? {add_268178, array_index_262439[0]} : sel_268180;
  assign add_268494 = array_index_262874[11:1] + 11'h079;
  assign sel_268496 = $signed({1'h0, add_268182, array_index_262442[0]}) < $signed({1'h0, sel_268184}) ? {add_268182, array_index_262442[0]} : sel_268184;
  assign add_268498 = array_index_263303[11:0] + 12'h59d;
  assign sel_268500 = $signed({1'h0, add_268186}) < $signed({1'h0, sel_268188}) ? add_268186 : sel_268188;
  assign add_268502 = array_index_263306[11:0] + 12'h59d;
  assign sel_268504 = $signed({1'h0, add_268190}) < $signed({1'h0, sel_268192}) ? add_268190 : sel_268192;
  assign add_268506 = array_index_263735[11:0] + 12'ha6f;
  assign sel_268508 = $signed({1'h0, add_268194}) < $signed({1'h0, sel_268196}) ? add_268194 : sel_268196;
  assign add_268510 = array_index_263738[11:0] + 12'ha6f;
  assign sel_268512 = $signed({1'h0, add_268198}) < $signed({1'h0, sel_268200}) ? add_268198 : sel_268200;
  assign add_268514 = array_index_264167[11:1] + 11'h499;
  assign sel_268516 = $signed({1'h0, add_268202, array_index_263735[0]}) < $signed({1'h0, sel_268204}) ? {add_268202, array_index_263735[0]} : sel_268204;
  assign add_268518 = array_index_264170[11:1] + 11'h499;
  assign sel_268520 = $signed({1'h0, add_268206, array_index_263738[0]}) < $signed({1'h0, sel_268208}) ? {add_268206, array_index_263738[0]} : sel_268208;
  assign add_268522 = array_index_264599[11:1] + 11'h345;
  assign sel_268525 = $signed({1'h0, add_268210, array_index_264167[0]}) < $signed({1'h0, sel_268213}) ? {add_268210, array_index_264167[0]} : sel_268213;
  assign add_268527 = array_index_264602[11:1] + 11'h345;
  assign sel_268530 = $signed({1'h0, add_268215, array_index_264170[0]}) < $signed({1'h0, sel_268218}) ? {add_268215, array_index_264170[0]} : sel_268218;
  assign add_268532 = array_index_265031[11:0] + 12'h30f;
  assign sel_268534 = $signed({1'h0, add_268220}) < $signed({1'h0, sel_268222}) ? add_268220 : sel_268222;
  assign add_268536 = array_index_265034[11:0] + 12'h30f;
  assign sel_268538 = $signed({1'h0, add_268224}) < $signed({1'h0, sel_268226}) ? add_268224 : sel_268226;
  assign add_268540 = array_index_265463[11:0] + 12'hb55;
  assign sel_268542 = $signed({1'h0, add_268228}) < $signed({1'h0, sel_268230}) ? add_268228 : sel_268230;
  assign add_268544 = array_index_265466[11:0] + 12'hb55;
  assign sel_268546 = $signed({1'h0, add_268232}) < $signed({1'h0, sel_268234}) ? add_268232 : sel_268234;
  assign concat_268549 = {1'h0, ($signed({1'h0, add_267916}) < $signed({1'h0, sel_267918}) ? add_267916 : sel_267918) == ($signed({1'h0, add_267920}) < $signed({1'h0, sel_267922}) ? add_267920 : sel_267922) ? add_268334 : concat_268245};
  assign add_268556 = array_index_260507[11:2] + 10'h29b;
  assign sel_268558 = $signed({1'h0, add_268252, array_index_260195[1:0]}) < $signed({1'h0, sel_268254}) ? {add_268252, array_index_260195[1:0]} : sel_268254;
  assign add_268560 = array_index_260510[11:2] + 10'h29b;
  assign sel_268562 = $signed({1'h0, add_268256, array_index_260198[1:0]}) < $signed({1'h0, sel_268258}) ? {add_268256, array_index_260198[1:0]} : sel_268258;
  assign add_268572 = array_index_261207[11:0] + 12'h9cf;
  assign sel_268574 = $signed({1'h0, add_268268}) < $signed({1'h0, sel_268270}) ? add_268268 : sel_268270;
  assign add_268576 = array_index_261210[11:0] + 12'h9cf;
  assign sel_268578 = $signed({1'h0, add_268272}) < $signed({1'h0, sel_268274}) ? add_268272 : sel_268274;
  assign add_268588 = array_index_262007[11:0] + 12'h30b;
  assign sel_268590 = $signed({1'h0, add_268284}) < $signed({1'h0, sel_268286}) ? add_268284 : sel_268286;
  assign add_268592 = array_index_262010[11:0] + 12'h30b;
  assign sel_268594 = $signed({1'h0, add_268288}) < $signed({1'h0, sel_268290}) ? add_268288 : sel_268290;
  assign add_268634 = concat_268549 + 8'h01;
  assign add_268644 = array_index_260845[11:0] + 12'hc05;
  assign sel_268646 = $signed({1'h0, add_268344}) < $signed({1'h0, sel_268346}) ? add_268344 : sel_268346;
  assign add_268648 = array_index_260848[11:0] + 12'hc05;
  assign sel_268650 = $signed({1'h0, add_268348}) < $signed({1'h0, sel_268350}) ? add_268348 : sel_268350;
  assign add_268662 = array_index_261595[11:0] + 12'h83f;
  assign sel_268664 = $signed({1'h0, add_268362}) < $signed({1'h0, sel_268364}) ? add_268362 : sel_268364;
  assign add_268666 = array_index_261598[11:0] + 12'h83f;
  assign sel_268668 = $signed({1'h0, add_268366}) < $signed({1'h0, sel_268368}) ? add_268366 : sel_268368;
  assign add_268680 = array_index_262439[11:1] + 11'h7b5;
  assign sel_268682 = $signed({1'h0, add_268380, array_index_262007[0]}) < $signed({1'h0, sel_268382}) ? {add_268380, array_index_262007[0]} : sel_268382;
  assign add_268684 = array_index_262442[11:1] + 11'h7b5;
  assign sel_268686 = $signed({1'h0, add_268384, array_index_262010[0]}) < $signed({1'h0, sel_268386}) ? {add_268384, array_index_262010[0]} : sel_268386;
  assign add_268728 = array_index_260507[11:0] + 12'hdab;
  assign sel_268730 = $signed({1'h0, add_268432}) < $signed({1'h0, sel_268434}) ? add_268432 : sel_268434;
  assign add_268732 = array_index_260510[11:0] + 12'hdab;
  assign sel_268734 = $signed({1'h0, add_268436}) < $signed({1'h0, sel_268438}) ? add_268436 : sel_268438;
  assign add_268746 = array_index_261207[11:2] + 10'h2b3;
  assign sel_268748 = $signed({1'h0, add_268450, array_index_260845[1:0]}) < $signed({1'h0, sel_268452}) ? {add_268450, array_index_260845[1:0]} : sel_268452;
  assign add_268750 = array_index_261210[11:2] + 10'h2b3;
  assign sel_268752 = $signed({1'h0, add_268454, array_index_260848[1:0]}) < $signed({1'h0, sel_268456}) ? {add_268454, array_index_260848[1:0]} : sel_268456;
  assign add_268762 = array_index_262007[11:1] + 11'h1e7;
  assign sel_268764 = $signed({1'h0, add_268466, array_index_261595[0]}) < $signed({1'h0, sel_268468}) ? {add_268466, array_index_261595[0]} : sel_268468;
  assign add_268766 = array_index_262010[11:1] + 11'h1e7;
  assign sel_268768 = $signed({1'h0, add_268470, array_index_261598[0]}) < $signed({1'h0, sel_268472}) ? {add_268470, array_index_261598[0]} : sel_268472;
  assign add_268778 = array_index_262871[11:0] + 12'h141;
  assign sel_268780 = $signed({1'h0, add_268482}) < $signed({1'h0, sel_268484}) ? add_268482 : sel_268484;
  assign add_268782 = array_index_262874[11:0] + 12'h141;
  assign sel_268784 = $signed({1'h0, add_268486}) < $signed({1'h0, sel_268488}) ? add_268486 : sel_268488;
  assign add_268786 = array_index_263303[11:1] + 11'h079;
  assign sel_268788 = $signed({1'h0, add_268490, array_index_262871[0]}) < $signed({1'h0, sel_268492}) ? {add_268490, array_index_262871[0]} : sel_268492;
  assign add_268790 = array_index_263306[11:1] + 11'h079;
  assign sel_268792 = $signed({1'h0, add_268494, array_index_262874[0]}) < $signed({1'h0, sel_268496}) ? {add_268494, array_index_262874[0]} : sel_268496;
  assign add_268794 = array_index_263735[11:0] + 12'h59d;
  assign sel_268796 = $signed({1'h0, add_268498}) < $signed({1'h0, sel_268500}) ? add_268498 : sel_268500;
  assign add_268798 = array_index_263738[11:0] + 12'h59d;
  assign sel_268800 = $signed({1'h0, add_268502}) < $signed({1'h0, sel_268504}) ? add_268502 : sel_268504;
  assign add_268802 = array_index_264167[11:0] + 12'ha6f;
  assign sel_268804 = $signed({1'h0, add_268506}) < $signed({1'h0, sel_268508}) ? add_268506 : sel_268508;
  assign add_268806 = array_index_264170[11:0] + 12'ha6f;
  assign sel_268808 = $signed({1'h0, add_268510}) < $signed({1'h0, sel_268512}) ? add_268510 : sel_268512;
  assign add_268810 = array_index_264599[11:1] + 11'h499;
  assign sel_268812 = $signed({1'h0, add_268514, array_index_264167[0]}) < $signed({1'h0, sel_268516}) ? {add_268514, array_index_264167[0]} : sel_268516;
  assign add_268814 = array_index_264602[11:1] + 11'h499;
  assign sel_268816 = $signed({1'h0, add_268518, array_index_264170[0]}) < $signed({1'h0, sel_268520}) ? {add_268518, array_index_264170[0]} : sel_268520;
  assign add_268818 = array_index_265031[11:1] + 11'h345;
  assign sel_268821 = $signed({1'h0, add_268522, array_index_264599[0]}) < $signed({1'h0, sel_268525}) ? {add_268522, array_index_264599[0]} : sel_268525;
  assign add_268823 = array_index_265034[11:1] + 11'h345;
  assign sel_268826 = $signed({1'h0, add_268527, array_index_264602[0]}) < $signed({1'h0, sel_268530}) ? {add_268527, array_index_264602[0]} : sel_268530;
  assign add_268828 = array_index_265463[11:0] + 12'h30f;
  assign sel_268830 = $signed({1'h0, add_268532}) < $signed({1'h0, sel_268534}) ? add_268532 : sel_268534;
  assign add_268832 = array_index_265466[11:0] + 12'h30f;
  assign sel_268834 = $signed({1'h0, add_268536}) < $signed({1'h0, sel_268538}) ? add_268536 : sel_268538;
  assign concat_268837 = {1'h0, ($signed({1'h0, add_268236}) < $signed({1'h0, sel_268238}) ? add_268236 : sel_268238) == ($signed({1'h0, add_268240}) < $signed({1'h0, sel_268242}) ? add_268240 : sel_268242) ? add_268634 : concat_268549};
  assign add_268844 = array_index_260845[11:2] + 10'h29b;
  assign sel_268846 = $signed({1'h0, add_268556, array_index_260507[1:0]}) < $signed({1'h0, sel_268558}) ? {add_268556, array_index_260507[1:0]} : sel_268558;
  assign add_268848 = array_index_260848[11:2] + 10'h29b;
  assign sel_268850 = $signed({1'h0, add_268560, array_index_260510[1:0]}) < $signed({1'h0, sel_268562}) ? {add_268560, array_index_260510[1:0]} : sel_268562;
  assign add_268860 = array_index_261595[11:0] + 12'h9cf;
  assign sel_268862 = $signed({1'h0, add_268572}) < $signed({1'h0, sel_268574}) ? add_268572 : sel_268574;
  assign add_268864 = array_index_261598[11:0] + 12'h9cf;
  assign sel_268866 = $signed({1'h0, add_268576}) < $signed({1'h0, sel_268578}) ? add_268576 : sel_268578;
  assign add_268876 = array_index_262439[11:0] + 12'h30b;
  assign sel_268878 = $signed({1'h0, add_268588}) < $signed({1'h0, sel_268590}) ? add_268588 : sel_268590;
  assign add_268880 = array_index_262442[11:0] + 12'h30b;
  assign sel_268882 = $signed({1'h0, add_268592}) < $signed({1'h0, sel_268594}) ? add_268592 : sel_268594;
  assign add_268918 = concat_268837 + 9'h001;
  assign add_268928 = array_index_261207[11:0] + 12'hc05;
  assign sel_268930 = $signed({1'h0, add_268644}) < $signed({1'h0, sel_268646}) ? add_268644 : sel_268646;
  assign add_268932 = array_index_261210[11:0] + 12'hc05;
  assign sel_268934 = $signed({1'h0, add_268648}) < $signed({1'h0, sel_268650}) ? add_268648 : sel_268650;
  assign add_268946 = array_index_262007[11:0] + 12'h83f;
  assign sel_268948 = $signed({1'h0, add_268662}) < $signed({1'h0, sel_268664}) ? add_268662 : sel_268664;
  assign add_268950 = array_index_262010[11:0] + 12'h83f;
  assign sel_268952 = $signed({1'h0, add_268666}) < $signed({1'h0, sel_268668}) ? add_268666 : sel_268668;
  assign add_268964 = array_index_262871[11:1] + 11'h7b5;
  assign sel_268966 = $signed({1'h0, add_268680, array_index_262439[0]}) < $signed({1'h0, sel_268682}) ? {add_268680, array_index_262439[0]} : sel_268682;
  assign add_268968 = array_index_262874[11:1] + 11'h7b5;
  assign sel_268970 = $signed({1'h0, add_268684, array_index_262442[0]}) < $signed({1'h0, sel_268686}) ? {add_268684, array_index_262442[0]} : sel_268686;
  assign add_269008 = array_index_260845[11:0] + 12'hdab;
  assign sel_269010 = $signed({1'h0, add_268728}) < $signed({1'h0, sel_268730}) ? add_268728 : sel_268730;
  assign add_269012 = array_index_260848[11:0] + 12'hdab;
  assign sel_269014 = $signed({1'h0, add_268732}) < $signed({1'h0, sel_268734}) ? add_268732 : sel_268734;
  assign add_269026 = array_index_261595[11:2] + 10'h2b3;
  assign sel_269028 = $signed({1'h0, add_268746, array_index_261207[1:0]}) < $signed({1'h0, sel_268748}) ? {add_268746, array_index_261207[1:0]} : sel_268748;
  assign add_269030 = array_index_261598[11:2] + 10'h2b3;
  assign sel_269032 = $signed({1'h0, add_268750, array_index_261210[1:0]}) < $signed({1'h0, sel_268752}) ? {add_268750, array_index_261210[1:0]} : sel_268752;
  assign add_269042 = array_index_262439[11:1] + 11'h1e7;
  assign sel_269044 = $signed({1'h0, add_268762, array_index_262007[0]}) < $signed({1'h0, sel_268764}) ? {add_268762, array_index_262007[0]} : sel_268764;
  assign add_269046 = array_index_262442[11:1] + 11'h1e7;
  assign sel_269048 = $signed({1'h0, add_268766, array_index_262010[0]}) < $signed({1'h0, sel_268768}) ? {add_268766, array_index_262010[0]} : sel_268768;
  assign add_269058 = array_index_263303[11:0] + 12'h141;
  assign sel_269060 = $signed({1'h0, add_268778}) < $signed({1'h0, sel_268780}) ? add_268778 : sel_268780;
  assign add_269062 = array_index_263306[11:0] + 12'h141;
  assign sel_269064 = $signed({1'h0, add_268782}) < $signed({1'h0, sel_268784}) ? add_268782 : sel_268784;
  assign add_269066 = array_index_263735[11:1] + 11'h079;
  assign sel_269068 = $signed({1'h0, add_268786, array_index_263303[0]}) < $signed({1'h0, sel_268788}) ? {add_268786, array_index_263303[0]} : sel_268788;
  assign add_269070 = array_index_263738[11:1] + 11'h079;
  assign sel_269072 = $signed({1'h0, add_268790, array_index_263306[0]}) < $signed({1'h0, sel_268792}) ? {add_268790, array_index_263306[0]} : sel_268792;
  assign add_269074 = array_index_264167[11:0] + 12'h59d;
  assign sel_269076 = $signed({1'h0, add_268794}) < $signed({1'h0, sel_268796}) ? add_268794 : sel_268796;
  assign add_269078 = array_index_264170[11:0] + 12'h59d;
  assign sel_269080 = $signed({1'h0, add_268798}) < $signed({1'h0, sel_268800}) ? add_268798 : sel_268800;
  assign add_269082 = array_index_264599[11:0] + 12'ha6f;
  assign sel_269084 = $signed({1'h0, add_268802}) < $signed({1'h0, sel_268804}) ? add_268802 : sel_268804;
  assign add_269086 = array_index_264602[11:0] + 12'ha6f;
  assign sel_269088 = $signed({1'h0, add_268806}) < $signed({1'h0, sel_268808}) ? add_268806 : sel_268808;
  assign add_269090 = array_index_265031[11:1] + 11'h499;
  assign sel_269092 = $signed({1'h0, add_268810, array_index_264599[0]}) < $signed({1'h0, sel_268812}) ? {add_268810, array_index_264599[0]} : sel_268812;
  assign add_269094 = array_index_265034[11:1] + 11'h499;
  assign sel_269096 = $signed({1'h0, add_268814, array_index_264602[0]}) < $signed({1'h0, sel_268816}) ? {add_268814, array_index_264602[0]} : sel_268816;
  assign add_269098 = array_index_265463[11:1] + 11'h345;
  assign sel_269101 = $signed({1'h0, add_268818, array_index_265031[0]}) < $signed({1'h0, sel_268821}) ? {add_268818, array_index_265031[0]} : sel_268821;
  assign add_269103 = array_index_265466[11:1] + 11'h345;
  assign sel_269106 = $signed({1'h0, add_268823, array_index_265034[0]}) < $signed({1'h0, sel_268826}) ? {add_268823, array_index_265034[0]} : sel_268826;
  assign concat_269109 = {1'h0, ($signed({1'h0, add_268540}) < $signed({1'h0, sel_268542}) ? add_268540 : sel_268542) == ($signed({1'h0, add_268544}) < $signed({1'h0, sel_268546}) ? add_268544 : sel_268546) ? add_268918 : concat_268837};
  assign add_269116 = array_index_261207[11:2] + 10'h29b;
  assign sel_269118 = $signed({1'h0, add_268844, array_index_260845[1:0]}) < $signed({1'h0, sel_268846}) ? {add_268844, array_index_260845[1:0]} : sel_268846;
  assign add_269120 = array_index_261210[11:2] + 10'h29b;
  assign sel_269122 = $signed({1'h0, add_268848, array_index_260848[1:0]}) < $signed({1'h0, sel_268850}) ? {add_268848, array_index_260848[1:0]} : sel_268850;
  assign add_269132 = array_index_262007[11:0] + 12'h9cf;
  assign sel_269134 = $signed({1'h0, add_268860}) < $signed({1'h0, sel_268862}) ? add_268860 : sel_268862;
  assign add_269136 = array_index_262010[11:0] + 12'h9cf;
  assign sel_269138 = $signed({1'h0, add_268864}) < $signed({1'h0, sel_268866}) ? add_268864 : sel_268866;
  assign add_269148 = array_index_262871[11:0] + 12'h30b;
  assign sel_269150 = $signed({1'h0, add_268876}) < $signed({1'h0, sel_268878}) ? add_268876 : sel_268878;
  assign add_269152 = array_index_262874[11:0] + 12'h30b;
  assign sel_269154 = $signed({1'h0, add_268880}) < $signed({1'h0, sel_268882}) ? add_268880 : sel_268882;
  assign add_269186 = concat_269109 + 10'h001;
  assign add_269196 = array_index_261595[11:0] + 12'hc05;
  assign sel_269198 = $signed({1'h0, add_268928}) < $signed({1'h0, sel_268930}) ? add_268928 : sel_268930;
  assign add_269200 = array_index_261598[11:0] + 12'hc05;
  assign sel_269202 = $signed({1'h0, add_268932}) < $signed({1'h0, sel_268934}) ? add_268932 : sel_268934;
  assign add_269214 = array_index_262439[11:0] + 12'h83f;
  assign sel_269216 = $signed({1'h0, add_268946}) < $signed({1'h0, sel_268948}) ? add_268946 : sel_268948;
  assign add_269218 = array_index_262442[11:0] + 12'h83f;
  assign sel_269220 = $signed({1'h0, add_268950}) < $signed({1'h0, sel_268952}) ? add_268950 : sel_268952;
  assign add_269232 = array_index_263303[11:1] + 11'h7b5;
  assign sel_269234 = $signed({1'h0, add_268964, array_index_262871[0]}) < $signed({1'h0, sel_268966}) ? {add_268964, array_index_262871[0]} : sel_268966;
  assign add_269236 = array_index_263306[11:1] + 11'h7b5;
  assign sel_269238 = $signed({1'h0, add_268968, array_index_262874[0]}) < $signed({1'h0, sel_268970}) ? {add_268968, array_index_262874[0]} : sel_268970;
  assign add_269270 = array_index_261207[11:0] + 12'hdab;
  assign sel_269272 = $signed({1'h0, add_269008}) < $signed({1'h0, sel_269010}) ? add_269008 : sel_269010;
  assign add_269274 = array_index_261210[11:0] + 12'hdab;
  assign sel_269276 = $signed({1'h0, add_269012}) < $signed({1'h0, sel_269014}) ? add_269012 : sel_269014;
  assign add_269288 = array_index_262007[11:2] + 10'h2b3;
  assign sel_269290 = $signed({1'h0, add_269026, array_index_261595[1:0]}) < $signed({1'h0, sel_269028}) ? {add_269026, array_index_261595[1:0]} : sel_269028;
  assign add_269292 = array_index_262010[11:2] + 10'h2b3;
  assign sel_269294 = $signed({1'h0, add_269030, array_index_261598[1:0]}) < $signed({1'h0, sel_269032}) ? {add_269030, array_index_261598[1:0]} : sel_269032;
  assign add_269304 = array_index_262871[11:1] + 11'h1e7;
  assign sel_269306 = $signed({1'h0, add_269042, array_index_262439[0]}) < $signed({1'h0, sel_269044}) ? {add_269042, array_index_262439[0]} : sel_269044;
  assign add_269308 = array_index_262874[11:1] + 11'h1e7;
  assign sel_269310 = $signed({1'h0, add_269046, array_index_262442[0]}) < $signed({1'h0, sel_269048}) ? {add_269046, array_index_262442[0]} : sel_269048;
  assign add_269320 = array_index_263735[11:0] + 12'h141;
  assign sel_269322 = $signed({1'h0, add_269058}) < $signed({1'h0, sel_269060}) ? add_269058 : sel_269060;
  assign add_269324 = array_index_263738[11:0] + 12'h141;
  assign sel_269326 = $signed({1'h0, add_269062}) < $signed({1'h0, sel_269064}) ? add_269062 : sel_269064;
  assign add_269328 = array_index_264167[11:1] + 11'h079;
  assign sel_269330 = $signed({1'h0, add_269066, array_index_263735[0]}) < $signed({1'h0, sel_269068}) ? {add_269066, array_index_263735[0]} : sel_269068;
  assign add_269332 = array_index_264170[11:1] + 11'h079;
  assign sel_269334 = $signed({1'h0, add_269070, array_index_263738[0]}) < $signed({1'h0, sel_269072}) ? {add_269070, array_index_263738[0]} : sel_269072;
  assign add_269336 = array_index_264599[11:0] + 12'h59d;
  assign sel_269338 = $signed({1'h0, add_269074}) < $signed({1'h0, sel_269076}) ? add_269074 : sel_269076;
  assign add_269340 = array_index_264602[11:0] + 12'h59d;
  assign sel_269342 = $signed({1'h0, add_269078}) < $signed({1'h0, sel_269080}) ? add_269078 : sel_269080;
  assign add_269344 = array_index_265031[11:0] + 12'ha6f;
  assign sel_269346 = $signed({1'h0, add_269082}) < $signed({1'h0, sel_269084}) ? add_269082 : sel_269084;
  assign add_269348 = array_index_265034[11:0] + 12'ha6f;
  assign sel_269350 = $signed({1'h0, add_269086}) < $signed({1'h0, sel_269088}) ? add_269086 : sel_269088;
  assign add_269352 = array_index_265463[11:1] + 11'h499;
  assign sel_269354 = $signed({1'h0, add_269090, array_index_265031[0]}) < $signed({1'h0, sel_269092}) ? {add_269090, array_index_265031[0]} : sel_269092;
  assign add_269356 = array_index_265466[11:1] + 11'h499;
  assign sel_269358 = $signed({1'h0, add_269094, array_index_265034[0]}) < $signed({1'h0, sel_269096}) ? {add_269094, array_index_265034[0]} : sel_269096;
  assign concat_269361 = {1'h0, ($signed({1'h0, add_268828}) < $signed({1'h0, sel_268830}) ? add_268828 : sel_268830) == ($signed({1'h0, add_268832}) < $signed({1'h0, sel_268834}) ? add_268832 : sel_268834) ? add_269186 : concat_269109};
  assign add_269368 = array_index_261595[11:2] + 10'h29b;
  assign sel_269370 = $signed({1'h0, add_269116, array_index_261207[1:0]}) < $signed({1'h0, sel_269118}) ? {add_269116, array_index_261207[1:0]} : sel_269118;
  assign add_269372 = array_index_261598[11:2] + 10'h29b;
  assign sel_269374 = $signed({1'h0, add_269120, array_index_261210[1:0]}) < $signed({1'h0, sel_269122}) ? {add_269120, array_index_261210[1:0]} : sel_269122;
  assign add_269384 = array_index_262439[11:0] + 12'h9cf;
  assign sel_269386 = $signed({1'h0, add_269132}) < $signed({1'h0, sel_269134}) ? add_269132 : sel_269134;
  assign add_269388 = array_index_262442[11:0] + 12'h9cf;
  assign sel_269390 = $signed({1'h0, add_269136}) < $signed({1'h0, sel_269138}) ? add_269136 : sel_269138;
  assign add_269400 = array_index_263303[11:0] + 12'h30b;
  assign sel_269402 = $signed({1'h0, add_269148}) < $signed({1'h0, sel_269150}) ? add_269148 : sel_269150;
  assign add_269404 = array_index_263306[11:0] + 12'h30b;
  assign sel_269406 = $signed({1'h0, add_269152}) < $signed({1'h0, sel_269154}) ? add_269152 : sel_269154;
  assign add_269434 = concat_269361 + 11'h001;
  assign add_269444 = array_index_262007[11:0] + 12'hc05;
  assign sel_269446 = $signed({1'h0, add_269196}) < $signed({1'h0, sel_269198}) ? add_269196 : sel_269198;
  assign add_269448 = array_index_262010[11:0] + 12'hc05;
  assign sel_269450 = $signed({1'h0, add_269200}) < $signed({1'h0, sel_269202}) ? add_269200 : sel_269202;
  assign add_269462 = array_index_262871[11:0] + 12'h83f;
  assign sel_269464 = $signed({1'h0, add_269214}) < $signed({1'h0, sel_269216}) ? add_269214 : sel_269216;
  assign add_269466 = array_index_262874[11:0] + 12'h83f;
  assign sel_269468 = $signed({1'h0, add_269218}) < $signed({1'h0, sel_269220}) ? add_269218 : sel_269220;
  assign add_269480 = array_index_263735[11:1] + 11'h7b5;
  assign sel_269482 = $signed({1'h0, add_269232, array_index_263303[0]}) < $signed({1'h0, sel_269234}) ? {add_269232, array_index_263303[0]} : sel_269234;
  assign add_269484 = array_index_263738[11:1] + 11'h7b5;
  assign sel_269486 = $signed({1'h0, add_269236, array_index_263306[0]}) < $signed({1'h0, sel_269238}) ? {add_269236, array_index_263306[0]} : sel_269238;
  assign add_269512 = array_index_261595[11:0] + 12'hdab;
  assign sel_269514 = $signed({1'h0, add_269270}) < $signed({1'h0, sel_269272}) ? add_269270 : sel_269272;
  assign add_269516 = array_index_261598[11:0] + 12'hdab;
  assign sel_269518 = $signed({1'h0, add_269274}) < $signed({1'h0, sel_269276}) ? add_269274 : sel_269276;
  assign add_269530 = array_index_262439[11:2] + 10'h2b3;
  assign sel_269532 = $signed({1'h0, add_269288, array_index_262007[1:0]}) < $signed({1'h0, sel_269290}) ? {add_269288, array_index_262007[1:0]} : sel_269290;
  assign add_269534 = array_index_262442[11:2] + 10'h2b3;
  assign sel_269536 = $signed({1'h0, add_269292, array_index_262010[1:0]}) < $signed({1'h0, sel_269294}) ? {add_269292, array_index_262010[1:0]} : sel_269294;
  assign add_269546 = array_index_263303[11:1] + 11'h1e7;
  assign sel_269548 = $signed({1'h0, add_269304, array_index_262871[0]}) < $signed({1'h0, sel_269306}) ? {add_269304, array_index_262871[0]} : sel_269306;
  assign add_269550 = array_index_263306[11:1] + 11'h1e7;
  assign sel_269552 = $signed({1'h0, add_269308, array_index_262874[0]}) < $signed({1'h0, sel_269310}) ? {add_269308, array_index_262874[0]} : sel_269310;
  assign add_269562 = array_index_264167[11:0] + 12'h141;
  assign sel_269564 = $signed({1'h0, add_269320}) < $signed({1'h0, sel_269322}) ? add_269320 : sel_269322;
  assign add_269566 = array_index_264170[11:0] + 12'h141;
  assign sel_269568 = $signed({1'h0, add_269324}) < $signed({1'h0, sel_269326}) ? add_269324 : sel_269326;
  assign add_269570 = array_index_264599[11:1] + 11'h079;
  assign sel_269572 = $signed({1'h0, add_269328, array_index_264167[0]}) < $signed({1'h0, sel_269330}) ? {add_269328, array_index_264167[0]} : sel_269330;
  assign add_269574 = array_index_264602[11:1] + 11'h079;
  assign sel_269576 = $signed({1'h0, add_269332, array_index_264170[0]}) < $signed({1'h0, sel_269334}) ? {add_269332, array_index_264170[0]} : sel_269334;
  assign add_269578 = array_index_265031[11:0] + 12'h59d;
  assign sel_269580 = $signed({1'h0, add_269336}) < $signed({1'h0, sel_269338}) ? add_269336 : sel_269338;
  assign add_269582 = array_index_265034[11:0] + 12'h59d;
  assign sel_269584 = $signed({1'h0, add_269340}) < $signed({1'h0, sel_269342}) ? add_269340 : sel_269342;
  assign add_269586 = array_index_265463[11:0] + 12'ha6f;
  assign sel_269588 = $signed({1'h0, add_269344}) < $signed({1'h0, sel_269346}) ? add_269344 : sel_269346;
  assign add_269590 = array_index_265466[11:0] + 12'ha6f;
  assign sel_269592 = $signed({1'h0, add_269348}) < $signed({1'h0, sel_269350}) ? add_269348 : sel_269350;
  assign concat_269595 = {1'h0, ($signed({1'h0, add_269098, array_index_265463[0]}) < $signed({1'h0, sel_269101}) ? {add_269098, array_index_265463[0]} : sel_269101) == ($signed({1'h0, add_269103, array_index_265466[0]}) < $signed({1'h0, sel_269106}) ? {add_269103, array_index_265466[0]} : sel_269106) ? add_269434 : concat_269361};
  assign add_269602 = array_index_262007[11:2] + 10'h29b;
  assign sel_269604 = $signed({1'h0, add_269368, array_index_261595[1:0]}) < $signed({1'h0, sel_269370}) ? {add_269368, array_index_261595[1:0]} : sel_269370;
  assign add_269606 = array_index_262010[11:2] + 10'h29b;
  assign sel_269608 = $signed({1'h0, add_269372, array_index_261598[1:0]}) < $signed({1'h0, sel_269374}) ? {add_269372, array_index_261598[1:0]} : sel_269374;
  assign add_269618 = array_index_262871[11:0] + 12'h9cf;
  assign sel_269620 = $signed({1'h0, add_269384}) < $signed({1'h0, sel_269386}) ? add_269384 : sel_269386;
  assign add_269622 = array_index_262874[11:0] + 12'h9cf;
  assign sel_269624 = $signed({1'h0, add_269388}) < $signed({1'h0, sel_269390}) ? add_269388 : sel_269390;
  assign add_269634 = array_index_263735[11:0] + 12'h30b;
  assign sel_269636 = $signed({1'h0, add_269400}) < $signed({1'h0, sel_269402}) ? add_269400 : sel_269402;
  assign add_269638 = array_index_263738[11:0] + 12'h30b;
  assign sel_269640 = $signed({1'h0, add_269404}) < $signed({1'h0, sel_269406}) ? add_269404 : sel_269406;
  assign add_269664 = concat_269595 + 12'h001;
  assign add_269674 = array_index_262439[11:0] + 12'hc05;
  assign sel_269676 = $signed({1'h0, add_269444}) < $signed({1'h0, sel_269446}) ? add_269444 : sel_269446;
  assign add_269678 = array_index_262442[11:0] + 12'hc05;
  assign sel_269680 = $signed({1'h0, add_269448}) < $signed({1'h0, sel_269450}) ? add_269448 : sel_269450;
  assign add_269692 = array_index_263303[11:0] + 12'h83f;
  assign sel_269694 = $signed({1'h0, add_269462}) < $signed({1'h0, sel_269464}) ? add_269462 : sel_269464;
  assign add_269696 = array_index_263306[11:0] + 12'h83f;
  assign sel_269698 = $signed({1'h0, add_269466}) < $signed({1'h0, sel_269468}) ? add_269466 : sel_269468;
  assign add_269710 = array_index_264167[11:1] + 11'h7b5;
  assign sel_269712 = $signed({1'h0, add_269480, array_index_263735[0]}) < $signed({1'h0, sel_269482}) ? {add_269480, array_index_263735[0]} : sel_269482;
  assign add_269714 = array_index_264170[11:1] + 11'h7b5;
  assign sel_269716 = $signed({1'h0, add_269484, array_index_263738[0]}) < $signed({1'h0, sel_269486}) ? {add_269484, array_index_263738[0]} : sel_269486;
  assign add_269736 = array_index_262007[11:0] + 12'hdab;
  assign sel_269738 = $signed({1'h0, add_269512}) < $signed({1'h0, sel_269514}) ? add_269512 : sel_269514;
  assign add_269740 = array_index_262010[11:0] + 12'hdab;
  assign sel_269742 = $signed({1'h0, add_269516}) < $signed({1'h0, sel_269518}) ? add_269516 : sel_269518;
  assign add_269754 = array_index_262871[11:2] + 10'h2b3;
  assign sel_269756 = $signed({1'h0, add_269530, array_index_262439[1:0]}) < $signed({1'h0, sel_269532}) ? {add_269530, array_index_262439[1:0]} : sel_269532;
  assign add_269758 = array_index_262874[11:2] + 10'h2b3;
  assign sel_269760 = $signed({1'h0, add_269534, array_index_262442[1:0]}) < $signed({1'h0, sel_269536}) ? {add_269534, array_index_262442[1:0]} : sel_269536;
  assign add_269770 = array_index_263735[11:1] + 11'h1e7;
  assign sel_269772 = $signed({1'h0, add_269546, array_index_263303[0]}) < $signed({1'h0, sel_269548}) ? {add_269546, array_index_263303[0]} : sel_269548;
  assign add_269774 = array_index_263738[11:1] + 11'h1e7;
  assign sel_269776 = $signed({1'h0, add_269550, array_index_263306[0]}) < $signed({1'h0, sel_269552}) ? {add_269550, array_index_263306[0]} : sel_269552;
  assign add_269786 = array_index_264599[11:0] + 12'h141;
  assign sel_269788 = $signed({1'h0, add_269562}) < $signed({1'h0, sel_269564}) ? add_269562 : sel_269564;
  assign add_269790 = array_index_264602[11:0] + 12'h141;
  assign sel_269792 = $signed({1'h0, add_269566}) < $signed({1'h0, sel_269568}) ? add_269566 : sel_269568;
  assign add_269794 = array_index_265031[11:1] + 11'h079;
  assign sel_269796 = $signed({1'h0, add_269570, array_index_264599[0]}) < $signed({1'h0, sel_269572}) ? {add_269570, array_index_264599[0]} : sel_269572;
  assign add_269798 = array_index_265034[11:1] + 11'h079;
  assign sel_269800 = $signed({1'h0, add_269574, array_index_264602[0]}) < $signed({1'h0, sel_269576}) ? {add_269574, array_index_264602[0]} : sel_269576;
  assign add_269802 = array_index_265463[11:0] + 12'h59d;
  assign sel_269804 = $signed({1'h0, add_269578}) < $signed({1'h0, sel_269580}) ? add_269578 : sel_269580;
  assign add_269806 = array_index_265466[11:0] + 12'h59d;
  assign sel_269808 = $signed({1'h0, add_269582}) < $signed({1'h0, sel_269584}) ? add_269582 : sel_269584;
  assign concat_269811 = {1'h0, ($signed({1'h0, add_269352, array_index_265463[0]}) < $signed({1'h0, sel_269354}) ? {add_269352, array_index_265463[0]} : sel_269354) == ($signed({1'h0, add_269356, array_index_265466[0]}) < $signed({1'h0, sel_269358}) ? {add_269356, array_index_265466[0]} : sel_269358) ? add_269664 : concat_269595};
  assign add_269818 = array_index_262439[11:2] + 10'h29b;
  assign sel_269820 = $signed({1'h0, add_269602, array_index_262007[1:0]}) < $signed({1'h0, sel_269604}) ? {add_269602, array_index_262007[1:0]} : sel_269604;
  assign add_269822 = array_index_262442[11:2] + 10'h29b;
  assign sel_269824 = $signed({1'h0, add_269606, array_index_262010[1:0]}) < $signed({1'h0, sel_269608}) ? {add_269606, array_index_262010[1:0]} : sel_269608;
  assign add_269834 = array_index_263303[11:0] + 12'h9cf;
  assign sel_269836 = $signed({1'h0, add_269618}) < $signed({1'h0, sel_269620}) ? add_269618 : sel_269620;
  assign add_269838 = array_index_263306[11:0] + 12'h9cf;
  assign sel_269840 = $signed({1'h0, add_269622}) < $signed({1'h0, sel_269624}) ? add_269622 : sel_269624;
  assign add_269850 = array_index_264167[11:0] + 12'h30b;
  assign sel_269852 = $signed({1'h0, add_269634}) < $signed({1'h0, sel_269636}) ? add_269634 : sel_269636;
  assign add_269854 = array_index_264170[11:0] + 12'h30b;
  assign sel_269856 = $signed({1'h0, add_269638}) < $signed({1'h0, sel_269640}) ? add_269638 : sel_269640;
  assign add_269876 = concat_269811 + 13'h0001;
  assign add_269886 = array_index_262871[11:0] + 12'hc05;
  assign sel_269888 = $signed({1'h0, add_269674}) < $signed({1'h0, sel_269676}) ? add_269674 : sel_269676;
  assign add_269890 = array_index_262874[11:0] + 12'hc05;
  assign sel_269892 = $signed({1'h0, add_269678}) < $signed({1'h0, sel_269680}) ? add_269678 : sel_269680;
  assign add_269904 = array_index_263735[11:0] + 12'h83f;
  assign sel_269906 = $signed({1'h0, add_269692}) < $signed({1'h0, sel_269694}) ? add_269692 : sel_269694;
  assign add_269908 = array_index_263738[11:0] + 12'h83f;
  assign sel_269910 = $signed({1'h0, add_269696}) < $signed({1'h0, sel_269698}) ? add_269696 : sel_269698;
  assign add_269922 = array_index_264599[11:1] + 11'h7b5;
  assign sel_269924 = $signed({1'h0, add_269710, array_index_264167[0]}) < $signed({1'h0, sel_269712}) ? {add_269710, array_index_264167[0]} : sel_269712;
  assign add_269926 = array_index_264602[11:1] + 11'h7b5;
  assign sel_269928 = $signed({1'h0, add_269714, array_index_264170[0]}) < $signed({1'h0, sel_269716}) ? {add_269714, array_index_264170[0]} : sel_269716;
  assign add_269944 = array_index_262439[11:0] + 12'hdab;
  assign sel_269946 = $signed({1'h0, add_269736}) < $signed({1'h0, sel_269738}) ? add_269736 : sel_269738;
  assign add_269948 = array_index_262442[11:0] + 12'hdab;
  assign sel_269950 = $signed({1'h0, add_269740}) < $signed({1'h0, sel_269742}) ? add_269740 : sel_269742;
  assign add_269962 = array_index_263303[11:2] + 10'h2b3;
  assign sel_269964 = $signed({1'h0, add_269754, array_index_262871[1:0]}) < $signed({1'h0, sel_269756}) ? {add_269754, array_index_262871[1:0]} : sel_269756;
  assign add_269966 = array_index_263306[11:2] + 10'h2b3;
  assign sel_269968 = $signed({1'h0, add_269758, array_index_262874[1:0]}) < $signed({1'h0, sel_269760}) ? {add_269758, array_index_262874[1:0]} : sel_269760;
  assign add_269978 = array_index_264167[11:1] + 11'h1e7;
  assign sel_269980 = $signed({1'h0, add_269770, array_index_263735[0]}) < $signed({1'h0, sel_269772}) ? {add_269770, array_index_263735[0]} : sel_269772;
  assign add_269982 = array_index_264170[11:1] + 11'h1e7;
  assign sel_269984 = $signed({1'h0, add_269774, array_index_263738[0]}) < $signed({1'h0, sel_269776}) ? {add_269774, array_index_263738[0]} : sel_269776;
  assign add_269994 = array_index_265031[11:0] + 12'h141;
  assign sel_269996 = $signed({1'h0, add_269786}) < $signed({1'h0, sel_269788}) ? add_269786 : sel_269788;
  assign add_269998 = array_index_265034[11:0] + 12'h141;
  assign sel_270000 = $signed({1'h0, add_269790}) < $signed({1'h0, sel_269792}) ? add_269790 : sel_269792;
  assign add_270002 = array_index_265463[11:1] + 11'h079;
  assign sel_270004 = $signed({1'h0, add_269794, array_index_265031[0]}) < $signed({1'h0, sel_269796}) ? {add_269794, array_index_265031[0]} : sel_269796;
  assign add_270006 = array_index_265466[11:1] + 11'h079;
  assign sel_270008 = $signed({1'h0, add_269798, array_index_265034[0]}) < $signed({1'h0, sel_269800}) ? {add_269798, array_index_265034[0]} : sel_269800;
  assign concat_270011 = {1'h0, ($signed({1'h0, add_269586}) < $signed({1'h0, sel_269588}) ? add_269586 : sel_269588) == ($signed({1'h0, add_269590}) < $signed({1'h0, sel_269592}) ? add_269590 : sel_269592) ? add_269876 : concat_269811};
  assign add_270018 = array_index_262871[11:2] + 10'h29b;
  assign sel_270020 = $signed({1'h0, add_269818, array_index_262439[1:0]}) < $signed({1'h0, sel_269820}) ? {add_269818, array_index_262439[1:0]} : sel_269820;
  assign add_270022 = array_index_262874[11:2] + 10'h29b;
  assign sel_270024 = $signed({1'h0, add_269822, array_index_262442[1:0]}) < $signed({1'h0, sel_269824}) ? {add_269822, array_index_262442[1:0]} : sel_269824;
  assign add_270034 = array_index_263735[11:0] + 12'h9cf;
  assign sel_270036 = $signed({1'h0, add_269834}) < $signed({1'h0, sel_269836}) ? add_269834 : sel_269836;
  assign add_270038 = array_index_263738[11:0] + 12'h9cf;
  assign sel_270040 = $signed({1'h0, add_269838}) < $signed({1'h0, sel_269840}) ? add_269838 : sel_269840;
  assign add_270050 = array_index_264599[11:0] + 12'h30b;
  assign sel_270052 = $signed({1'h0, add_269850}) < $signed({1'h0, sel_269852}) ? add_269850 : sel_269852;
  assign add_270054 = array_index_264602[11:0] + 12'h30b;
  assign sel_270056 = $signed({1'h0, add_269854}) < $signed({1'h0, sel_269856}) ? add_269854 : sel_269856;
  assign add_270072 = concat_270011 + 14'h0001;
  assign add_270082 = array_index_263303[11:0] + 12'hc05;
  assign sel_270084 = $signed({1'h0, add_269886}) < $signed({1'h0, sel_269888}) ? add_269886 : sel_269888;
  assign add_270086 = array_index_263306[11:0] + 12'hc05;
  assign sel_270088 = $signed({1'h0, add_269890}) < $signed({1'h0, sel_269892}) ? add_269890 : sel_269892;
  assign add_270100 = array_index_264167[11:0] + 12'h83f;
  assign sel_270102 = $signed({1'h0, add_269904}) < $signed({1'h0, sel_269906}) ? add_269904 : sel_269906;
  assign add_270104 = array_index_264170[11:0] + 12'h83f;
  assign sel_270106 = $signed({1'h0, add_269908}) < $signed({1'h0, sel_269910}) ? add_269908 : sel_269910;
  assign add_270118 = array_index_265031[11:1] + 11'h7b5;
  assign sel_270120 = $signed({1'h0, add_269922, array_index_264599[0]}) < $signed({1'h0, sel_269924}) ? {add_269922, array_index_264599[0]} : sel_269924;
  assign add_270122 = array_index_265034[11:1] + 11'h7b5;
  assign sel_270124 = $signed({1'h0, add_269926, array_index_264602[0]}) < $signed({1'h0, sel_269928}) ? {add_269926, array_index_264602[0]} : sel_269928;
  assign add_270136 = array_index_262871[11:0] + 12'hdab;
  assign sel_270138 = $signed({1'h0, add_269944}) < $signed({1'h0, sel_269946}) ? add_269944 : sel_269946;
  assign add_270140 = array_index_262874[11:0] + 12'hdab;
  assign sel_270142 = $signed({1'h0, add_269948}) < $signed({1'h0, sel_269950}) ? add_269948 : sel_269950;
  assign add_270154 = array_index_263735[11:2] + 10'h2b3;
  assign sel_270156 = $signed({1'h0, add_269962, array_index_263303[1:0]}) < $signed({1'h0, sel_269964}) ? {add_269962, array_index_263303[1:0]} : sel_269964;
  assign add_270158 = array_index_263738[11:2] + 10'h2b3;
  assign sel_270160 = $signed({1'h0, add_269966, array_index_263306[1:0]}) < $signed({1'h0, sel_269968}) ? {add_269966, array_index_263306[1:0]} : sel_269968;
  assign add_270170 = array_index_264599[11:1] + 11'h1e7;
  assign sel_270172 = $signed({1'h0, add_269978, array_index_264167[0]}) < $signed({1'h0, sel_269980}) ? {add_269978, array_index_264167[0]} : sel_269980;
  assign add_270174 = array_index_264602[11:1] + 11'h1e7;
  assign sel_270176 = $signed({1'h0, add_269982, array_index_264170[0]}) < $signed({1'h0, sel_269984}) ? {add_269982, array_index_264170[0]} : sel_269984;
  assign add_270186 = array_index_265463[11:0] + 12'h141;
  assign sel_270188 = $signed({1'h0, add_269994}) < $signed({1'h0, sel_269996}) ? add_269994 : sel_269996;
  assign add_270190 = array_index_265466[11:0] + 12'h141;
  assign sel_270192 = $signed({1'h0, add_269998}) < $signed({1'h0, sel_270000}) ? add_269998 : sel_270000;
  assign concat_270195 = {1'h0, ($signed({1'h0, add_269802}) < $signed({1'h0, sel_269804}) ? add_269802 : sel_269804) == ($signed({1'h0, add_269806}) < $signed({1'h0, sel_269808}) ? add_269806 : sel_269808) ? add_270072 : concat_270011};
  assign add_270202 = array_index_263303[11:2] + 10'h29b;
  assign sel_270204 = $signed({1'h0, add_270018, array_index_262871[1:0]}) < $signed({1'h0, sel_270020}) ? {add_270018, array_index_262871[1:0]} : sel_270020;
  assign add_270206 = array_index_263306[11:2] + 10'h29b;
  assign sel_270208 = $signed({1'h0, add_270022, array_index_262874[1:0]}) < $signed({1'h0, sel_270024}) ? {add_270022, array_index_262874[1:0]} : sel_270024;
  assign add_270218 = array_index_264167[11:0] + 12'h9cf;
  assign sel_270220 = $signed({1'h0, add_270034}) < $signed({1'h0, sel_270036}) ? add_270034 : sel_270036;
  assign add_270222 = array_index_264170[11:0] + 12'h9cf;
  assign sel_270224 = $signed({1'h0, add_270038}) < $signed({1'h0, sel_270040}) ? add_270038 : sel_270040;
  assign add_270234 = array_index_265031[11:0] + 12'h30b;
  assign sel_270236 = $signed({1'h0, add_270050}) < $signed({1'h0, sel_270052}) ? add_270050 : sel_270052;
  assign add_270238 = array_index_265034[11:0] + 12'h30b;
  assign sel_270240 = $signed({1'h0, add_270054}) < $signed({1'h0, sel_270056}) ? add_270054 : sel_270056;
  assign add_270252 = concat_270195 + 15'h0001;
  assign add_270262 = array_index_263735[11:0] + 12'hc05;
  assign sel_270264 = $signed({1'h0, add_270082}) < $signed({1'h0, sel_270084}) ? add_270082 : sel_270084;
  assign add_270266 = array_index_263738[11:0] + 12'hc05;
  assign sel_270268 = $signed({1'h0, add_270086}) < $signed({1'h0, sel_270088}) ? add_270086 : sel_270088;
  assign add_270280 = array_index_264599[11:0] + 12'h83f;
  assign sel_270282 = $signed({1'h0, add_270100}) < $signed({1'h0, sel_270102}) ? add_270100 : sel_270102;
  assign add_270284 = array_index_264602[11:0] + 12'h83f;
  assign sel_270286 = $signed({1'h0, add_270104}) < $signed({1'h0, sel_270106}) ? add_270104 : sel_270106;
  assign add_270298 = array_index_265463[11:1] + 11'h7b5;
  assign sel_270300 = $signed({1'h0, add_270118, array_index_265031[0]}) < $signed({1'h0, sel_270120}) ? {add_270118, array_index_265031[0]} : sel_270120;
  assign add_270302 = array_index_265466[11:1] + 11'h7b5;
  assign sel_270304 = $signed({1'h0, add_270122, array_index_265034[0]}) < $signed({1'h0, sel_270124}) ? {add_270122, array_index_265034[0]} : sel_270124;
  assign add_270310 = array_index_263303[11:0] + 12'hdab;
  assign sel_270312 = $signed({1'h0, add_270136}) < $signed({1'h0, sel_270138}) ? add_270136 : sel_270138;
  assign add_270314 = array_index_263306[11:0] + 12'hdab;
  assign sel_270316 = $signed({1'h0, add_270140}) < $signed({1'h0, sel_270142}) ? add_270140 : sel_270142;
  assign add_270328 = array_index_264167[11:2] + 10'h2b3;
  assign sel_270330 = $signed({1'h0, add_270154, array_index_263735[1:0]}) < $signed({1'h0, sel_270156}) ? {add_270154, array_index_263735[1:0]} : sel_270156;
  assign add_270332 = array_index_264170[11:2] + 10'h2b3;
  assign sel_270334 = $signed({1'h0, add_270158, array_index_263738[1:0]}) < $signed({1'h0, sel_270160}) ? {add_270158, array_index_263738[1:0]} : sel_270160;
  assign add_270344 = array_index_265031[11:1] + 11'h1e7;
  assign sel_270346 = $signed({1'h0, add_270170, array_index_264599[0]}) < $signed({1'h0, sel_270172}) ? {add_270170, array_index_264599[0]} : sel_270172;
  assign add_270348 = array_index_265034[11:1] + 11'h1e7;
  assign sel_270350 = $signed({1'h0, add_270174, array_index_264602[0]}) < $signed({1'h0, sel_270176}) ? {add_270174, array_index_264602[0]} : sel_270176;
  assign concat_270361 = {1'h0, ($signed({1'h0, add_270002, array_index_265463[0]}) < $signed({1'h0, sel_270004}) ? {add_270002, array_index_265463[0]} : sel_270004) == ($signed({1'h0, add_270006, array_index_265466[0]}) < $signed({1'h0, sel_270008}) ? {add_270006, array_index_265466[0]} : sel_270008) ? add_270252 : concat_270195};
  assign add_270368 = array_index_263735[11:2] + 10'h29b;
  assign sel_270370 = $signed({1'h0, add_270202, array_index_263303[1:0]}) < $signed({1'h0, sel_270204}) ? {add_270202, array_index_263303[1:0]} : sel_270204;
  assign add_270372 = array_index_263738[11:2] + 10'h29b;
  assign sel_270374 = $signed({1'h0, add_270206, array_index_263306[1:0]}) < $signed({1'h0, sel_270208}) ? {add_270206, array_index_263306[1:0]} : sel_270208;
  assign add_270384 = array_index_264599[11:0] + 12'h9cf;
  assign sel_270386 = $signed({1'h0, add_270218}) < $signed({1'h0, sel_270220}) ? add_270218 : sel_270220;
  assign add_270388 = array_index_264602[11:0] + 12'h9cf;
  assign sel_270390 = $signed({1'h0, add_270222}) < $signed({1'h0, sel_270224}) ? add_270222 : sel_270224;
  assign add_270400 = array_index_265463[11:0] + 12'h30b;
  assign sel_270402 = $signed({1'h0, add_270234}) < $signed({1'h0, sel_270236}) ? add_270234 : sel_270236;
  assign add_270404 = array_index_265466[11:0] + 12'h30b;
  assign sel_270406 = $signed({1'h0, add_270238}) < $signed({1'h0, sel_270240}) ? add_270238 : sel_270240;
  assign add_270412 = concat_270361 + 16'h0001;
  assign add_270422 = array_index_264167[11:0] + 12'hc05;
  assign sel_270424 = $signed({1'h0, add_270262}) < $signed({1'h0, sel_270264}) ? add_270262 : sel_270264;
  assign add_270426 = array_index_264170[11:0] + 12'hc05;
  assign sel_270428 = $signed({1'h0, add_270266}) < $signed({1'h0, sel_270268}) ? add_270266 : sel_270268;
  assign add_270440 = array_index_265031[11:0] + 12'h83f;
  assign sel_270442 = $signed({1'h0, add_270280}) < $signed({1'h0, sel_270282}) ? add_270280 : sel_270282;
  assign add_270444 = array_index_265034[11:0] + 12'h83f;
  assign sel_270446 = $signed({1'h0, add_270284}) < $signed({1'h0, sel_270286}) ? add_270284 : sel_270286;
  assign sel_270459 = ($signed({1'h0, add_270186}) < $signed({1'h0, sel_270188}) ? add_270186 : sel_270188) == ($signed({1'h0, add_270190}) < $signed({1'h0, sel_270192}) ? add_270190 : sel_270192) ? add_270412 : concat_270361;
  assign add_270462 = array_index_263735[11:0] + 12'hdab;
  assign sel_270464 = $signed({1'h0, add_270310}) < $signed({1'h0, sel_270312}) ? add_270310 : sel_270312;
  assign add_270466 = array_index_263738[11:0] + 12'hdab;
  assign sel_270468 = $signed({1'h0, add_270314}) < $signed({1'h0, sel_270316}) ? add_270314 : sel_270316;
  assign add_270480 = array_index_264599[11:2] + 10'h2b3;
  assign sel_270482 = $signed({1'h0, add_270328, array_index_264167[1:0]}) < $signed({1'h0, sel_270330}) ? {add_270328, array_index_264167[1:0]} : sel_270330;
  assign add_270484 = array_index_264602[11:2] + 10'h2b3;
  assign sel_270486 = $signed({1'h0, add_270332, array_index_264170[1:0]}) < $signed({1'h0, sel_270334}) ? {add_270332, array_index_264170[1:0]} : sel_270334;
  assign add_270496 = array_index_265463[11:1] + 11'h1e7;
  assign sel_270498 = $signed({1'h0, add_270344, array_index_265031[0]}) < $signed({1'h0, sel_270346}) ? {add_270344, array_index_265031[0]} : sel_270346;
  assign add_270500 = array_index_265466[11:1] + 11'h1e7;
  assign sel_270502 = $signed({1'h0, add_270348, array_index_265034[0]}) < $signed({1'h0, sel_270350}) ? {add_270348, array_index_265034[0]} : sel_270350;
  assign add_270506 = sel_270459 + 16'h0001;
  assign add_270512 = array_index_264167[11:2] + 10'h29b;
  assign sel_270514 = $signed({1'h0, add_270368, array_index_263735[1:0]}) < $signed({1'h0, sel_270370}) ? {add_270368, array_index_263735[1:0]} : sel_270370;
  assign add_270516 = array_index_264170[11:2] + 10'h29b;
  assign sel_270518 = $signed({1'h0, add_270372, array_index_263738[1:0]}) < $signed({1'h0, sel_270374}) ? {add_270372, array_index_263738[1:0]} : sel_270374;
  assign add_270528 = array_index_265031[11:0] + 12'h9cf;
  assign sel_270530 = $signed({1'h0, add_270384}) < $signed({1'h0, sel_270386}) ? add_270384 : sel_270386;
  assign add_270532 = array_index_265034[11:0] + 12'h9cf;
  assign sel_270534 = $signed({1'h0, add_270388}) < $signed({1'h0, sel_270390}) ? add_270388 : sel_270390;
  assign sel_270545 = ($signed({1'h0, add_270298, array_index_265463[0]}) < $signed({1'h0, sel_270300}) ? {add_270298, array_index_265463[0]} : sel_270300) == ($signed({1'h0, add_270302, array_index_265466[0]}) < $signed({1'h0, sel_270304}) ? {add_270302, array_index_265466[0]} : sel_270304) ? add_270506 : sel_270459;
  assign add_270556 = array_index_264599[11:0] + 12'hc05;
  assign sel_270558 = $signed({1'h0, add_270422}) < $signed({1'h0, sel_270424}) ? add_270422 : sel_270424;
  assign add_270560 = array_index_264602[11:0] + 12'hc05;
  assign sel_270562 = $signed({1'h0, add_270426}) < $signed({1'h0, sel_270428}) ? add_270426 : sel_270428;
  assign add_270574 = array_index_265463[11:0] + 12'h83f;
  assign sel_270576 = $signed({1'h0, add_270440}) < $signed({1'h0, sel_270442}) ? add_270440 : sel_270442;
  assign add_270578 = array_index_265466[11:0] + 12'h83f;
  assign sel_270580 = $signed({1'h0, add_270444}) < $signed({1'h0, sel_270446}) ? add_270444 : sel_270446;
  assign add_270586 = sel_270545 + 16'h0001;
  assign add_270588 = array_index_264167[11:0] + 12'hdab;
  assign sel_270590 = $signed({1'h0, add_270462}) < $signed({1'h0, sel_270464}) ? add_270462 : sel_270464;
  assign add_270592 = array_index_264170[11:0] + 12'hdab;
  assign sel_270594 = $signed({1'h0, add_270466}) < $signed({1'h0, sel_270468}) ? add_270466 : sel_270468;
  assign add_270606 = array_index_265031[11:2] + 10'h2b3;
  assign sel_270608 = $signed({1'h0, add_270480, array_index_264599[1:0]}) < $signed({1'h0, sel_270482}) ? {add_270480, array_index_264599[1:0]} : sel_270482;
  assign add_270610 = array_index_265034[11:2] + 10'h2b3;
  assign sel_270612 = $signed({1'h0, add_270484, array_index_264602[1:0]}) < $signed({1'h0, sel_270486}) ? {add_270484, array_index_264602[1:0]} : sel_270486;
  assign sel_270623 = ($signed({1'h0, add_270400}) < $signed({1'h0, sel_270402}) ? add_270400 : sel_270402) == ($signed({1'h0, add_270404}) < $signed({1'h0, sel_270406}) ? add_270404 : sel_270406) ? add_270586 : sel_270545;
  assign add_270630 = array_index_264599[11:2] + 10'h29b;
  assign sel_270632 = $signed({1'h0, add_270512, array_index_264167[1:0]}) < $signed({1'h0, sel_270514}) ? {add_270512, array_index_264167[1:0]} : sel_270514;
  assign add_270634 = array_index_264602[11:2] + 10'h29b;
  assign sel_270636 = $signed({1'h0, add_270516, array_index_264170[1:0]}) < $signed({1'h0, sel_270518}) ? {add_270516, array_index_264170[1:0]} : sel_270518;
  assign add_270646 = array_index_265463[11:0] + 12'h9cf;
  assign sel_270648 = $signed({1'h0, add_270528}) < $signed({1'h0, sel_270530}) ? add_270528 : sel_270530;
  assign add_270650 = array_index_265466[11:0] + 12'h9cf;
  assign sel_270652 = $signed({1'h0, add_270532}) < $signed({1'h0, sel_270534}) ? add_270532 : sel_270534;
  assign add_270656 = sel_270623 + 16'h0001;
  assign add_270666 = array_index_265031[11:0] + 12'hc05;
  assign sel_270668 = $signed({1'h0, add_270556}) < $signed({1'h0, sel_270558}) ? add_270556 : sel_270558;
  assign add_270670 = array_index_265034[11:0] + 12'hc05;
  assign sel_270672 = $signed({1'h0, add_270560}) < $signed({1'h0, sel_270562}) ? add_270560 : sel_270562;
  assign sel_270685 = ($signed({1'h0, add_270496, array_index_265463[0]}) < $signed({1'h0, sel_270498}) ? {add_270496, array_index_265463[0]} : sel_270498) == ($signed({1'h0, add_270500, array_index_265466[0]}) < $signed({1'h0, sel_270502}) ? {add_270500, array_index_265466[0]} : sel_270502) ? add_270656 : sel_270623;
  assign add_270688 = array_index_264599[11:0] + 12'hdab;
  assign sel_270690 = $signed({1'h0, add_270588}) < $signed({1'h0, sel_270590}) ? add_270588 : sel_270590;
  assign add_270692 = array_index_264602[11:0] + 12'hdab;
  assign sel_270694 = $signed({1'h0, add_270592}) < $signed({1'h0, sel_270594}) ? add_270592 : sel_270594;
  assign add_270706 = array_index_265463[11:2] + 10'h2b3;
  assign sel_270708 = $signed({1'h0, add_270606, array_index_265031[1:0]}) < $signed({1'h0, sel_270608}) ? {add_270606, array_index_265031[1:0]} : sel_270608;
  assign add_270710 = array_index_265466[11:2] + 10'h2b3;
  assign sel_270712 = $signed({1'h0, add_270610, array_index_265034[1:0]}) < $signed({1'h0, sel_270612}) ? {add_270610, array_index_265034[1:0]} : sel_270612;
  assign add_270716 = sel_270685 + 16'h0001;
  assign add_270722 = array_index_265031[11:2] + 10'h29b;
  assign sel_270724 = $signed({1'h0, add_270630, array_index_264599[1:0]}) < $signed({1'h0, sel_270632}) ? {add_270630, array_index_264599[1:0]} : sel_270632;
  assign add_270726 = array_index_265034[11:2] + 10'h29b;
  assign sel_270728 = $signed({1'h0, add_270634, array_index_264602[1:0]}) < $signed({1'h0, sel_270636}) ? {add_270634, array_index_264602[1:0]} : sel_270636;
  assign sel_270739 = ($signed({1'h0, add_270574}) < $signed({1'h0, sel_270576}) ? add_270574 : sel_270576) == ($signed({1'h0, add_270578}) < $signed({1'h0, sel_270580}) ? add_270578 : sel_270580) ? add_270716 : sel_270685;
  assign add_270750 = array_index_265463[11:0] + 12'hc05;
  assign sel_270752 = $signed({1'h0, add_270666}) < $signed({1'h0, sel_270668}) ? add_270666 : sel_270668;
  assign add_270754 = array_index_265466[11:0] + 12'hc05;
  assign sel_270756 = $signed({1'h0, add_270670}) < $signed({1'h0, sel_270672}) ? add_270670 : sel_270672;
  assign add_270762 = sel_270739 + 16'h0001;
  assign add_270764 = array_index_265031[11:0] + 12'hdab;
  assign sel_270766 = $signed({1'h0, add_270688}) < $signed({1'h0, sel_270690}) ? add_270688 : sel_270690;
  assign add_270768 = array_index_265034[11:0] + 12'hdab;
  assign sel_270770 = $signed({1'h0, add_270692}) < $signed({1'h0, sel_270694}) ? add_270692 : sel_270694;
  assign sel_270783 = ($signed({1'h0, add_270646}) < $signed({1'h0, sel_270648}) ? add_270646 : sel_270648) == ($signed({1'h0, add_270650}) < $signed({1'h0, sel_270652}) ? add_270650 : sel_270652) ? add_270762 : sel_270739;
  assign add_270790 = array_index_265463[11:2] + 10'h29b;
  assign sel_270792 = $signed({1'h0, add_270722, array_index_265031[1:0]}) < $signed({1'h0, sel_270724}) ? {add_270722, array_index_265031[1:0]} : sel_270724;
  assign add_270794 = array_index_265466[11:2] + 10'h29b;
  assign sel_270796 = $signed({1'h0, add_270726, array_index_265034[1:0]}) < $signed({1'h0, sel_270728}) ? {add_270726, array_index_265034[1:0]} : sel_270728;
  assign add_270800 = sel_270783 + 16'h0001;
  assign sel_270811 = ($signed({1'h0, add_270706, array_index_265463[1:0]}) < $signed({1'h0, sel_270708}) ? {add_270706, array_index_265463[1:0]} : sel_270708) == ($signed({1'h0, add_270710, array_index_265466[1:0]}) < $signed({1'h0, sel_270712}) ? {add_270710, array_index_265466[1:0]} : sel_270712) ? add_270800 : sel_270783;
  assign add_270814 = array_index_265463[11:0] + 12'hdab;
  assign sel_270816 = $signed({1'h0, add_270764}) < $signed({1'h0, sel_270766}) ? add_270764 : sel_270766;
  assign add_270818 = array_index_265466[11:0] + 12'hdab;
  assign sel_270820 = $signed({1'h0, add_270768}) < $signed({1'h0, sel_270770}) ? add_270768 : sel_270770;
  assign add_270826 = sel_270811 + 16'h0001;
  assign sel_270833 = ($signed({1'h0, add_270750}) < $signed({1'h0, sel_270752}) ? add_270750 : sel_270752) == ($signed({1'h0, add_270754}) < $signed({1'h0, sel_270756}) ? add_270754 : sel_270756) ? add_270826 : sel_270811;
  assign add_270838 = sel_270833 + 16'h0001;
  assign sel_270841 = ($signed({1'h0, add_270790, array_index_265463[1:0]}) < $signed({1'h0, sel_270792}) ? {add_270790, array_index_265463[1:0]} : sel_270792) == ($signed({1'h0, add_270794, array_index_265466[1:0]}) < $signed({1'h0, sel_270796}) ? {add_270794, array_index_265466[1:0]} : sel_270796) ? add_270838 : sel_270833;
  assign add_270844 = sel_270841 + 16'h0001;
  assign out = {($signed({1'h0, add_270814}) < $signed({1'h0, sel_270816}) ? add_270814 : sel_270816) == ($signed({1'h0, add_270818}) < $signed({1'h0, sel_270820}) ? add_270818 : sel_270820) ? add_270844 : sel_270841, {set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
