module min_hash(
  input wire [1599:0] set1,
  input wire [1599:0] set2,
  output wire [3215:0] out
);
  wire [15:0] set1_unflattened[100];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  assign set1_unflattened[50] = set1[815:800];
  assign set1_unflattened[51] = set1[831:816];
  assign set1_unflattened[52] = set1[847:832];
  assign set1_unflattened[53] = set1[863:848];
  assign set1_unflattened[54] = set1[879:864];
  assign set1_unflattened[55] = set1[895:880];
  assign set1_unflattened[56] = set1[911:896];
  assign set1_unflattened[57] = set1[927:912];
  assign set1_unflattened[58] = set1[943:928];
  assign set1_unflattened[59] = set1[959:944];
  assign set1_unflattened[60] = set1[975:960];
  assign set1_unflattened[61] = set1[991:976];
  assign set1_unflattened[62] = set1[1007:992];
  assign set1_unflattened[63] = set1[1023:1008];
  assign set1_unflattened[64] = set1[1039:1024];
  assign set1_unflattened[65] = set1[1055:1040];
  assign set1_unflattened[66] = set1[1071:1056];
  assign set1_unflattened[67] = set1[1087:1072];
  assign set1_unflattened[68] = set1[1103:1088];
  assign set1_unflattened[69] = set1[1119:1104];
  assign set1_unflattened[70] = set1[1135:1120];
  assign set1_unflattened[71] = set1[1151:1136];
  assign set1_unflattened[72] = set1[1167:1152];
  assign set1_unflattened[73] = set1[1183:1168];
  assign set1_unflattened[74] = set1[1199:1184];
  assign set1_unflattened[75] = set1[1215:1200];
  assign set1_unflattened[76] = set1[1231:1216];
  assign set1_unflattened[77] = set1[1247:1232];
  assign set1_unflattened[78] = set1[1263:1248];
  assign set1_unflattened[79] = set1[1279:1264];
  assign set1_unflattened[80] = set1[1295:1280];
  assign set1_unflattened[81] = set1[1311:1296];
  assign set1_unflattened[82] = set1[1327:1312];
  assign set1_unflattened[83] = set1[1343:1328];
  assign set1_unflattened[84] = set1[1359:1344];
  assign set1_unflattened[85] = set1[1375:1360];
  assign set1_unflattened[86] = set1[1391:1376];
  assign set1_unflattened[87] = set1[1407:1392];
  assign set1_unflattened[88] = set1[1423:1408];
  assign set1_unflattened[89] = set1[1439:1424];
  assign set1_unflattened[90] = set1[1455:1440];
  assign set1_unflattened[91] = set1[1471:1456];
  assign set1_unflattened[92] = set1[1487:1472];
  assign set1_unflattened[93] = set1[1503:1488];
  assign set1_unflattened[94] = set1[1519:1504];
  assign set1_unflattened[95] = set1[1535:1520];
  assign set1_unflattened[96] = set1[1551:1536];
  assign set1_unflattened[97] = set1[1567:1552];
  assign set1_unflattened[98] = set1[1583:1568];
  assign set1_unflattened[99] = set1[1599:1584];
  wire [15:0] set2_unflattened[100];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  assign set2_unflattened[50] = set2[815:800];
  assign set2_unflattened[51] = set2[831:816];
  assign set2_unflattened[52] = set2[847:832];
  assign set2_unflattened[53] = set2[863:848];
  assign set2_unflattened[54] = set2[879:864];
  assign set2_unflattened[55] = set2[895:880];
  assign set2_unflattened[56] = set2[911:896];
  assign set2_unflattened[57] = set2[927:912];
  assign set2_unflattened[58] = set2[943:928];
  assign set2_unflattened[59] = set2[959:944];
  assign set2_unflattened[60] = set2[975:960];
  assign set2_unflattened[61] = set2[991:976];
  assign set2_unflattened[62] = set2[1007:992];
  assign set2_unflattened[63] = set2[1023:1008];
  assign set2_unflattened[64] = set2[1039:1024];
  assign set2_unflattened[65] = set2[1055:1040];
  assign set2_unflattened[66] = set2[1071:1056];
  assign set2_unflattened[67] = set2[1087:1072];
  assign set2_unflattened[68] = set2[1103:1088];
  assign set2_unflattened[69] = set2[1119:1104];
  assign set2_unflattened[70] = set2[1135:1120];
  assign set2_unflattened[71] = set2[1151:1136];
  assign set2_unflattened[72] = set2[1167:1152];
  assign set2_unflattened[73] = set2[1183:1168];
  assign set2_unflattened[74] = set2[1199:1184];
  assign set2_unflattened[75] = set2[1215:1200];
  assign set2_unflattened[76] = set2[1231:1216];
  assign set2_unflattened[77] = set2[1247:1232];
  assign set2_unflattened[78] = set2[1263:1248];
  assign set2_unflattened[79] = set2[1279:1264];
  assign set2_unflattened[80] = set2[1295:1280];
  assign set2_unflattened[81] = set2[1311:1296];
  assign set2_unflattened[82] = set2[1327:1312];
  assign set2_unflattened[83] = set2[1343:1328];
  assign set2_unflattened[84] = set2[1359:1344];
  assign set2_unflattened[85] = set2[1375:1360];
  assign set2_unflattened[86] = set2[1391:1376];
  assign set2_unflattened[87] = set2[1407:1392];
  assign set2_unflattened[88] = set2[1423:1408];
  assign set2_unflattened[89] = set2[1439:1424];
  assign set2_unflattened[90] = set2[1455:1440];
  assign set2_unflattened[91] = set2[1471:1456];
  assign set2_unflattened[92] = set2[1487:1472];
  assign set2_unflattened[93] = set2[1503:1488];
  assign set2_unflattened[94] = set2[1519:1504];
  assign set2_unflattened[95] = set2[1535:1520];
  assign set2_unflattened[96] = set2[1551:1536];
  assign set2_unflattened[97] = set2[1567:1552];
  assign set2_unflattened[98] = set2[1583:1568];
  assign set2_unflattened[99] = set2[1599:1584];
  wire [15:0] array_index_172855;
  wire [15:0] array_index_172856;
  wire [11:0] add_172863;
  wire [11:0] add_172866;
  wire [15:0] array_index_172871;
  wire [15:0] array_index_172874;
  wire [10:0] add_172878;
  wire [10:0] add_172881;
  wire [11:0] add_172897;
  wire [11:0] sel_172899;
  wire [11:0] add_172902;
  wire [11:0] sel_172904;
  wire [15:0] array_index_172919;
  wire [15:0] array_index_172922;
  wire [8:0] add_172926;
  wire [8:0] add_172929;
  wire [10:0] add_172932;
  wire [11:0] sel_172935;
  wire [10:0] add_172937;
  wire [11:0] sel_172940;
  wire [11:0] add_172957;
  wire [11:0] sel_172959;
  wire [11:0] add_172962;
  wire [11:0] sel_172964;
  wire [15:0] array_index_172985;
  wire [15:0] array_index_172988;
  wire [10:0] add_172992;
  wire [10:0] add_172994;
  wire [8:0] add_172996;
  wire [11:0] sel_172999;
  wire [8:0] add_173001;
  wire [11:0] sel_173004;
  wire [10:0] add_173006;
  wire [11:0] sel_173009;
  wire [10:0] add_173011;
  wire [11:0] sel_173014;
  wire [11:0] add_173035;
  wire [11:0] sel_173037;
  wire [11:0] add_173040;
  wire [11:0] sel_173042;
  wire [15:0] array_index_173069;
  wire [15:0] array_index_173072;
  wire [10:0] add_173076;
  wire [10:0] add_173078;
  wire [10:0] add_173080;
  wire [11:0] sel_173082;
  wire [10:0] add_173084;
  wire [11:0] sel_173086;
  wire [8:0] add_173088;
  wire [11:0] sel_173091;
  wire [8:0] add_173093;
  wire [11:0] sel_173096;
  wire [10:0] add_173098;
  wire [11:0] sel_173101;
  wire [10:0] add_173103;
  wire [11:0] sel_173106;
  wire [11:0] add_173131;
  wire [11:0] sel_173133;
  wire [11:0] add_173136;
  wire [11:0] sel_173138;
  wire [15:0] array_index_173169;
  wire [15:0] array_index_173172;
  wire [10:0] add_173176;
  wire [11:0] sel_173178;
  wire [10:0] add_173180;
  wire [11:0] sel_173182;
  wire [10:0] add_173184;
  wire [11:0] sel_173186;
  wire [10:0] add_173188;
  wire [11:0] sel_173190;
  wire [8:0] add_173192;
  wire [11:0] sel_173195;
  wire [8:0] add_173197;
  wire [11:0] sel_173200;
  wire [10:0] add_173202;
  wire [11:0] sel_173205;
  wire [10:0] add_173207;
  wire [11:0] sel_173210;
  wire [11:0] add_173235;
  wire [11:0] sel_173237;
  wire [11:0] add_173240;
  wire [11:0] sel_173242;
  wire [15:0] array_index_173271;
  wire [15:0] array_index_173274;
  wire [10:0] add_173278;
  wire [11:0] sel_173280;
  wire [10:0] add_173282;
  wire [11:0] sel_173284;
  wire [10:0] add_173286;
  wire [11:0] sel_173288;
  wire [10:0] add_173290;
  wire [11:0] sel_173292;
  wire [8:0] add_173294;
  wire [11:0] sel_173297;
  wire [8:0] add_173299;
  wire [11:0] sel_173302;
  wire [10:0] add_173304;
  wire [11:0] sel_173307;
  wire [10:0] add_173309;
  wire [11:0] sel_173312;
  wire [11:0] add_173337;
  wire [11:0] sel_173339;
  wire [11:0] add_173342;
  wire [11:0] sel_173344;
  wire [15:0] array_index_173373;
  wire [15:0] array_index_173376;
  wire [10:0] add_173380;
  wire [11:0] sel_173382;
  wire [10:0] add_173384;
  wire [11:0] sel_173386;
  wire [10:0] add_173388;
  wire [11:0] sel_173390;
  wire [10:0] add_173392;
  wire [11:0] sel_173394;
  wire [8:0] add_173396;
  wire [11:0] sel_173399;
  wire [8:0] add_173401;
  wire [11:0] sel_173404;
  wire [10:0] add_173406;
  wire [11:0] sel_173409;
  wire [10:0] add_173411;
  wire [11:0] sel_173414;
  wire [11:0] add_173439;
  wire [11:0] sel_173441;
  wire [11:0] add_173444;
  wire [11:0] sel_173446;
  wire [15:0] array_index_173475;
  wire [15:0] array_index_173478;
  wire [10:0] add_173482;
  wire [11:0] sel_173484;
  wire [10:0] add_173486;
  wire [11:0] sel_173488;
  wire [10:0] add_173490;
  wire [11:0] sel_173492;
  wire [10:0] add_173494;
  wire [11:0] sel_173496;
  wire [8:0] add_173498;
  wire [11:0] sel_173501;
  wire [8:0] add_173503;
  wire [11:0] sel_173506;
  wire [10:0] add_173508;
  wire [11:0] sel_173511;
  wire [10:0] add_173513;
  wire [11:0] sel_173516;
  wire [11:0] add_173541;
  wire [11:0] sel_173543;
  wire [11:0] add_173546;
  wire [11:0] sel_173548;
  wire [15:0] array_index_173577;
  wire [15:0] array_index_173580;
  wire [10:0] add_173584;
  wire [11:0] sel_173586;
  wire [10:0] add_173588;
  wire [11:0] sel_173590;
  wire [10:0] add_173592;
  wire [11:0] sel_173594;
  wire [10:0] add_173596;
  wire [11:0] sel_173598;
  wire [8:0] add_173600;
  wire [11:0] sel_173603;
  wire [8:0] add_173605;
  wire [11:0] sel_173608;
  wire [10:0] add_173610;
  wire [11:0] sel_173613;
  wire [10:0] add_173615;
  wire [11:0] sel_173618;
  wire [11:0] add_173643;
  wire [11:0] sel_173645;
  wire [11:0] add_173648;
  wire [11:0] sel_173650;
  wire [15:0] array_index_173679;
  wire [15:0] array_index_173682;
  wire [10:0] add_173686;
  wire [11:0] sel_173688;
  wire [10:0] add_173690;
  wire [11:0] sel_173692;
  wire [10:0] add_173694;
  wire [11:0] sel_173696;
  wire [10:0] add_173698;
  wire [11:0] sel_173700;
  wire [8:0] add_173702;
  wire [11:0] sel_173705;
  wire [8:0] add_173707;
  wire [11:0] sel_173710;
  wire [10:0] add_173712;
  wire [11:0] sel_173715;
  wire [10:0] add_173717;
  wire [11:0] sel_173720;
  wire [11:0] add_173745;
  wire [11:0] sel_173747;
  wire [11:0] add_173750;
  wire [11:0] sel_173752;
  wire [15:0] array_index_173781;
  wire [15:0] array_index_173784;
  wire [10:0] add_173788;
  wire [11:0] sel_173790;
  wire [10:0] add_173792;
  wire [11:0] sel_173794;
  wire [10:0] add_173796;
  wire [11:0] sel_173798;
  wire [10:0] add_173800;
  wire [11:0] sel_173802;
  wire [8:0] add_173804;
  wire [11:0] sel_173807;
  wire [8:0] add_173809;
  wire [11:0] sel_173812;
  wire [10:0] add_173814;
  wire [11:0] sel_173817;
  wire [10:0] add_173819;
  wire [11:0] sel_173822;
  wire [11:0] add_173847;
  wire [11:0] sel_173849;
  wire [11:0] add_173852;
  wire [11:0] sel_173854;
  wire [15:0] array_index_173883;
  wire [15:0] array_index_173886;
  wire [10:0] add_173890;
  wire [11:0] sel_173892;
  wire [10:0] add_173894;
  wire [11:0] sel_173896;
  wire [10:0] add_173898;
  wire [11:0] sel_173900;
  wire [10:0] add_173902;
  wire [11:0] sel_173904;
  wire [8:0] add_173906;
  wire [11:0] sel_173909;
  wire [8:0] add_173911;
  wire [11:0] sel_173914;
  wire [10:0] add_173916;
  wire [11:0] sel_173919;
  wire [10:0] add_173921;
  wire [11:0] sel_173924;
  wire [11:0] add_173949;
  wire [11:0] sel_173951;
  wire [11:0] add_173954;
  wire [11:0] sel_173956;
  wire [15:0] array_index_173985;
  wire [15:0] array_index_173988;
  wire [10:0] add_173992;
  wire [11:0] sel_173994;
  wire [10:0] add_173996;
  wire [11:0] sel_173998;
  wire [10:0] add_174000;
  wire [11:0] sel_174002;
  wire [10:0] add_174004;
  wire [11:0] sel_174006;
  wire [8:0] add_174008;
  wire [11:0] sel_174011;
  wire [8:0] add_174013;
  wire [11:0] sel_174016;
  wire [10:0] add_174018;
  wire [11:0] sel_174021;
  wire [10:0] add_174023;
  wire [11:0] sel_174026;
  wire [11:0] add_174051;
  wire [11:0] sel_174053;
  wire [11:0] add_174056;
  wire [11:0] sel_174058;
  wire [15:0] array_index_174087;
  wire [15:0] array_index_174090;
  wire [10:0] add_174094;
  wire [11:0] sel_174096;
  wire [10:0] add_174098;
  wire [11:0] sel_174100;
  wire [10:0] add_174102;
  wire [11:0] sel_174104;
  wire [10:0] add_174106;
  wire [11:0] sel_174108;
  wire [8:0] add_174110;
  wire [11:0] sel_174113;
  wire [8:0] add_174115;
  wire [11:0] sel_174118;
  wire [10:0] add_174120;
  wire [11:0] sel_174123;
  wire [10:0] add_174125;
  wire [11:0] sel_174128;
  wire [11:0] add_174153;
  wire [11:0] sel_174155;
  wire [11:0] add_174158;
  wire [11:0] sel_174160;
  wire [15:0] array_index_174189;
  wire [15:0] array_index_174192;
  wire [10:0] add_174196;
  wire [11:0] sel_174198;
  wire [10:0] add_174200;
  wire [11:0] sel_174202;
  wire [10:0] add_174204;
  wire [11:0] sel_174206;
  wire [10:0] add_174208;
  wire [11:0] sel_174210;
  wire [8:0] add_174212;
  wire [11:0] sel_174215;
  wire [8:0] add_174217;
  wire [11:0] sel_174220;
  wire [10:0] add_174222;
  wire [11:0] sel_174225;
  wire [10:0] add_174227;
  wire [11:0] sel_174230;
  wire [11:0] add_174255;
  wire [11:0] sel_174257;
  wire [11:0] add_174260;
  wire [11:0] sel_174262;
  wire [15:0] array_index_174291;
  wire [15:0] array_index_174294;
  wire [10:0] add_174298;
  wire [11:0] sel_174300;
  wire [10:0] add_174302;
  wire [11:0] sel_174304;
  wire [10:0] add_174306;
  wire [11:0] sel_174308;
  wire [10:0] add_174310;
  wire [11:0] sel_174312;
  wire [8:0] add_174314;
  wire [11:0] sel_174317;
  wire [8:0] add_174319;
  wire [11:0] sel_174322;
  wire [10:0] add_174324;
  wire [11:0] sel_174327;
  wire [10:0] add_174329;
  wire [11:0] sel_174332;
  wire [11:0] add_174357;
  wire [11:0] sel_174359;
  wire [11:0] add_174362;
  wire [11:0] sel_174364;
  wire [15:0] array_index_174393;
  wire [15:0] array_index_174396;
  wire [10:0] add_174400;
  wire [11:0] sel_174402;
  wire [10:0] add_174404;
  wire [11:0] sel_174406;
  wire [10:0] add_174408;
  wire [11:0] sel_174410;
  wire [10:0] add_174412;
  wire [11:0] sel_174414;
  wire [8:0] add_174416;
  wire [11:0] sel_174419;
  wire [8:0] add_174421;
  wire [11:0] sel_174424;
  wire [10:0] add_174426;
  wire [11:0] sel_174429;
  wire [10:0] add_174431;
  wire [11:0] sel_174434;
  wire [11:0] add_174459;
  wire [11:0] sel_174461;
  wire [11:0] add_174464;
  wire [11:0] sel_174466;
  wire [15:0] array_index_174495;
  wire [15:0] array_index_174498;
  wire [10:0] add_174502;
  wire [11:0] sel_174504;
  wire [10:0] add_174506;
  wire [11:0] sel_174508;
  wire [10:0] add_174510;
  wire [11:0] sel_174512;
  wire [10:0] add_174514;
  wire [11:0] sel_174516;
  wire [8:0] add_174518;
  wire [11:0] sel_174521;
  wire [8:0] add_174523;
  wire [11:0] sel_174526;
  wire [10:0] add_174528;
  wire [11:0] sel_174531;
  wire [10:0] add_174533;
  wire [11:0] sel_174536;
  wire [11:0] add_174561;
  wire [11:0] sel_174563;
  wire [11:0] add_174566;
  wire [11:0] sel_174568;
  wire [15:0] array_index_174597;
  wire [15:0] array_index_174600;
  wire [10:0] add_174604;
  wire [11:0] sel_174606;
  wire [10:0] add_174608;
  wire [11:0] sel_174610;
  wire [10:0] add_174612;
  wire [11:0] sel_174614;
  wire [10:0] add_174616;
  wire [11:0] sel_174618;
  wire [8:0] add_174620;
  wire [11:0] sel_174623;
  wire [8:0] add_174625;
  wire [11:0] sel_174628;
  wire [10:0] add_174630;
  wire [11:0] sel_174633;
  wire [10:0] add_174635;
  wire [11:0] sel_174638;
  wire [11:0] add_174663;
  wire [11:0] sel_174665;
  wire [11:0] add_174668;
  wire [11:0] sel_174670;
  wire [15:0] array_index_174699;
  wire [15:0] array_index_174702;
  wire [10:0] add_174706;
  wire [11:0] sel_174708;
  wire [10:0] add_174710;
  wire [11:0] sel_174712;
  wire [10:0] add_174714;
  wire [11:0] sel_174716;
  wire [10:0] add_174718;
  wire [11:0] sel_174720;
  wire [8:0] add_174722;
  wire [11:0] sel_174725;
  wire [8:0] add_174727;
  wire [11:0] sel_174730;
  wire [10:0] add_174732;
  wire [11:0] sel_174735;
  wire [10:0] add_174737;
  wire [11:0] sel_174740;
  wire [11:0] add_174765;
  wire [11:0] sel_174767;
  wire [11:0] add_174770;
  wire [11:0] sel_174772;
  wire [15:0] array_index_174801;
  wire [15:0] array_index_174804;
  wire [10:0] add_174808;
  wire [11:0] sel_174810;
  wire [10:0] add_174812;
  wire [11:0] sel_174814;
  wire [10:0] add_174816;
  wire [11:0] sel_174818;
  wire [10:0] add_174820;
  wire [11:0] sel_174822;
  wire [8:0] add_174824;
  wire [11:0] sel_174827;
  wire [8:0] add_174829;
  wire [11:0] sel_174832;
  wire [10:0] add_174834;
  wire [11:0] sel_174837;
  wire [10:0] add_174839;
  wire [11:0] sel_174842;
  wire [11:0] add_174867;
  wire [11:0] sel_174869;
  wire [11:0] add_174872;
  wire [11:0] sel_174874;
  wire [15:0] array_index_174903;
  wire [15:0] array_index_174906;
  wire [10:0] add_174910;
  wire [11:0] sel_174912;
  wire [10:0] add_174914;
  wire [11:0] sel_174916;
  wire [10:0] add_174918;
  wire [11:0] sel_174920;
  wire [10:0] add_174922;
  wire [11:0] sel_174924;
  wire [8:0] add_174926;
  wire [11:0] sel_174929;
  wire [8:0] add_174931;
  wire [11:0] sel_174934;
  wire [10:0] add_174936;
  wire [11:0] sel_174939;
  wire [10:0] add_174941;
  wire [11:0] sel_174944;
  wire [11:0] add_174969;
  wire [11:0] sel_174971;
  wire [11:0] add_174974;
  wire [11:0] sel_174976;
  wire [15:0] array_index_175005;
  wire [15:0] array_index_175008;
  wire [10:0] add_175012;
  wire [11:0] sel_175014;
  wire [10:0] add_175016;
  wire [11:0] sel_175018;
  wire [10:0] add_175020;
  wire [11:0] sel_175022;
  wire [10:0] add_175024;
  wire [11:0] sel_175026;
  wire [8:0] add_175028;
  wire [11:0] sel_175031;
  wire [8:0] add_175033;
  wire [11:0] sel_175036;
  wire [10:0] add_175038;
  wire [11:0] sel_175041;
  wire [10:0] add_175043;
  wire [11:0] sel_175046;
  wire [11:0] add_175071;
  wire [11:0] sel_175073;
  wire [11:0] add_175076;
  wire [11:0] sel_175078;
  wire [15:0] array_index_175107;
  wire [15:0] array_index_175110;
  wire [10:0] add_175114;
  wire [11:0] sel_175116;
  wire [10:0] add_175118;
  wire [11:0] sel_175120;
  wire [10:0] add_175122;
  wire [11:0] sel_175124;
  wire [10:0] add_175126;
  wire [11:0] sel_175128;
  wire [8:0] add_175130;
  wire [11:0] sel_175133;
  wire [8:0] add_175135;
  wire [11:0] sel_175138;
  wire [10:0] add_175140;
  wire [11:0] sel_175143;
  wire [10:0] add_175145;
  wire [11:0] sel_175148;
  wire [11:0] add_175173;
  wire [11:0] sel_175175;
  wire [11:0] add_175178;
  wire [11:0] sel_175180;
  wire [15:0] array_index_175209;
  wire [15:0] array_index_175212;
  wire [10:0] add_175216;
  wire [11:0] sel_175218;
  wire [10:0] add_175220;
  wire [11:0] sel_175222;
  wire [10:0] add_175224;
  wire [11:0] sel_175226;
  wire [10:0] add_175228;
  wire [11:0] sel_175230;
  wire [8:0] add_175232;
  wire [11:0] sel_175235;
  wire [8:0] add_175237;
  wire [11:0] sel_175240;
  wire [10:0] add_175242;
  wire [11:0] sel_175245;
  wire [10:0] add_175247;
  wire [11:0] sel_175250;
  wire [11:0] add_175275;
  wire [11:0] sel_175277;
  wire [11:0] add_175280;
  wire [11:0] sel_175282;
  wire [15:0] array_index_175311;
  wire [15:0] array_index_175314;
  wire [10:0] add_175318;
  wire [11:0] sel_175320;
  wire [10:0] add_175322;
  wire [11:0] sel_175324;
  wire [10:0] add_175326;
  wire [11:0] sel_175328;
  wire [10:0] add_175330;
  wire [11:0] sel_175332;
  wire [8:0] add_175334;
  wire [11:0] sel_175337;
  wire [8:0] add_175339;
  wire [11:0] sel_175342;
  wire [10:0] add_175344;
  wire [11:0] sel_175347;
  wire [10:0] add_175349;
  wire [11:0] sel_175352;
  wire [11:0] add_175377;
  wire [11:0] sel_175379;
  wire [11:0] add_175382;
  wire [11:0] sel_175384;
  wire [15:0] array_index_175413;
  wire [15:0] array_index_175416;
  wire [10:0] add_175420;
  wire [11:0] sel_175422;
  wire [10:0] add_175424;
  wire [11:0] sel_175426;
  wire [10:0] add_175428;
  wire [11:0] sel_175430;
  wire [10:0] add_175432;
  wire [11:0] sel_175434;
  wire [8:0] add_175436;
  wire [11:0] sel_175439;
  wire [8:0] add_175441;
  wire [11:0] sel_175444;
  wire [10:0] add_175446;
  wire [11:0] sel_175449;
  wire [10:0] add_175451;
  wire [11:0] sel_175454;
  wire [11:0] add_175479;
  wire [11:0] sel_175481;
  wire [11:0] add_175484;
  wire [11:0] sel_175486;
  wire [15:0] array_index_175515;
  wire [15:0] array_index_175518;
  wire [10:0] add_175522;
  wire [11:0] sel_175524;
  wire [10:0] add_175526;
  wire [11:0] sel_175528;
  wire [10:0] add_175530;
  wire [11:0] sel_175532;
  wire [10:0] add_175534;
  wire [11:0] sel_175536;
  wire [8:0] add_175538;
  wire [11:0] sel_175541;
  wire [8:0] add_175543;
  wire [11:0] sel_175546;
  wire [10:0] add_175548;
  wire [11:0] sel_175551;
  wire [10:0] add_175553;
  wire [11:0] sel_175556;
  wire [11:0] add_175581;
  wire [11:0] sel_175583;
  wire [11:0] add_175586;
  wire [11:0] sel_175588;
  wire [15:0] array_index_175617;
  wire [15:0] array_index_175620;
  wire [10:0] add_175624;
  wire [11:0] sel_175626;
  wire [10:0] add_175628;
  wire [11:0] sel_175630;
  wire [10:0] add_175632;
  wire [11:0] sel_175634;
  wire [10:0] add_175636;
  wire [11:0] sel_175638;
  wire [8:0] add_175640;
  wire [11:0] sel_175643;
  wire [8:0] add_175645;
  wire [11:0] sel_175648;
  wire [10:0] add_175650;
  wire [11:0] sel_175653;
  wire [10:0] add_175655;
  wire [11:0] sel_175658;
  wire [11:0] add_175683;
  wire [11:0] sel_175685;
  wire [11:0] add_175688;
  wire [11:0] sel_175690;
  wire [15:0] array_index_175719;
  wire [15:0] array_index_175722;
  wire [10:0] add_175726;
  wire [11:0] sel_175728;
  wire [10:0] add_175730;
  wire [11:0] sel_175732;
  wire [10:0] add_175734;
  wire [11:0] sel_175736;
  wire [10:0] add_175738;
  wire [11:0] sel_175740;
  wire [8:0] add_175742;
  wire [11:0] sel_175745;
  wire [8:0] add_175747;
  wire [11:0] sel_175750;
  wire [10:0] add_175752;
  wire [11:0] sel_175755;
  wire [10:0] add_175757;
  wire [11:0] sel_175760;
  wire [11:0] add_175785;
  wire [11:0] sel_175787;
  wire [11:0] add_175790;
  wire [11:0] sel_175792;
  wire [15:0] array_index_175821;
  wire [15:0] array_index_175824;
  wire [10:0] add_175828;
  wire [11:0] sel_175830;
  wire [10:0] add_175832;
  wire [11:0] sel_175834;
  wire [10:0] add_175836;
  wire [11:0] sel_175838;
  wire [10:0] add_175840;
  wire [11:0] sel_175842;
  wire [8:0] add_175844;
  wire [11:0] sel_175847;
  wire [8:0] add_175849;
  wire [11:0] sel_175852;
  wire [10:0] add_175854;
  wire [11:0] sel_175857;
  wire [10:0] add_175859;
  wire [11:0] sel_175862;
  wire [11:0] add_175887;
  wire [11:0] sel_175889;
  wire [11:0] add_175892;
  wire [11:0] sel_175894;
  wire [15:0] array_index_175923;
  wire [15:0] array_index_175926;
  wire [10:0] add_175930;
  wire [11:0] sel_175932;
  wire [10:0] add_175934;
  wire [11:0] sel_175936;
  wire [10:0] add_175938;
  wire [11:0] sel_175940;
  wire [10:0] add_175942;
  wire [11:0] sel_175944;
  wire [8:0] add_175946;
  wire [11:0] sel_175949;
  wire [8:0] add_175951;
  wire [11:0] sel_175954;
  wire [10:0] add_175956;
  wire [11:0] sel_175959;
  wire [10:0] add_175961;
  wire [11:0] sel_175964;
  wire [11:0] add_175989;
  wire [11:0] sel_175991;
  wire [11:0] add_175994;
  wire [11:0] sel_175996;
  wire [15:0] array_index_176025;
  wire [15:0] array_index_176028;
  wire [10:0] add_176032;
  wire [11:0] sel_176034;
  wire [10:0] add_176036;
  wire [11:0] sel_176038;
  wire [10:0] add_176040;
  wire [11:0] sel_176042;
  wire [10:0] add_176044;
  wire [11:0] sel_176046;
  wire [8:0] add_176048;
  wire [11:0] sel_176051;
  wire [8:0] add_176053;
  wire [11:0] sel_176056;
  wire [10:0] add_176058;
  wire [11:0] sel_176061;
  wire [10:0] add_176063;
  wire [11:0] sel_176066;
  wire [11:0] add_176091;
  wire [11:0] sel_176093;
  wire [11:0] add_176096;
  wire [11:0] sel_176098;
  wire [15:0] array_index_176127;
  wire [15:0] array_index_176130;
  wire [10:0] add_176134;
  wire [11:0] sel_176136;
  wire [10:0] add_176138;
  wire [11:0] sel_176140;
  wire [10:0] add_176142;
  wire [11:0] sel_176144;
  wire [10:0] add_176146;
  wire [11:0] sel_176148;
  wire [8:0] add_176150;
  wire [11:0] sel_176153;
  wire [8:0] add_176155;
  wire [11:0] sel_176158;
  wire [10:0] add_176160;
  wire [11:0] sel_176163;
  wire [10:0] add_176165;
  wire [11:0] sel_176168;
  wire [11:0] add_176193;
  wire [11:0] sel_176195;
  wire [11:0] add_176198;
  wire [11:0] sel_176200;
  wire [15:0] array_index_176229;
  wire [15:0] array_index_176232;
  wire [10:0] add_176236;
  wire [11:0] sel_176238;
  wire [10:0] add_176240;
  wire [11:0] sel_176242;
  wire [10:0] add_176244;
  wire [11:0] sel_176246;
  wire [10:0] add_176248;
  wire [11:0] sel_176250;
  wire [8:0] add_176252;
  wire [11:0] sel_176255;
  wire [8:0] add_176257;
  wire [11:0] sel_176260;
  wire [10:0] add_176262;
  wire [11:0] sel_176265;
  wire [10:0] add_176267;
  wire [11:0] sel_176270;
  wire [11:0] add_176295;
  wire [11:0] sel_176297;
  wire [11:0] add_176300;
  wire [11:0] sel_176302;
  wire [15:0] array_index_176331;
  wire [15:0] array_index_176334;
  wire [10:0] add_176338;
  wire [11:0] sel_176340;
  wire [10:0] add_176342;
  wire [11:0] sel_176344;
  wire [10:0] add_176346;
  wire [11:0] sel_176348;
  wire [10:0] add_176350;
  wire [11:0] sel_176352;
  wire [8:0] add_176354;
  wire [11:0] sel_176357;
  wire [8:0] add_176359;
  wire [11:0] sel_176362;
  wire [10:0] add_176364;
  wire [11:0] sel_176367;
  wire [10:0] add_176369;
  wire [11:0] sel_176372;
  wire [11:0] add_176397;
  wire [11:0] sel_176399;
  wire [11:0] add_176402;
  wire [11:0] sel_176404;
  wire [15:0] array_index_176433;
  wire [15:0] array_index_176436;
  wire [10:0] add_176440;
  wire [11:0] sel_176442;
  wire [10:0] add_176444;
  wire [11:0] sel_176446;
  wire [10:0] add_176448;
  wire [11:0] sel_176450;
  wire [10:0] add_176452;
  wire [11:0] sel_176454;
  wire [8:0] add_176456;
  wire [11:0] sel_176459;
  wire [8:0] add_176461;
  wire [11:0] sel_176464;
  wire [10:0] add_176466;
  wire [11:0] sel_176469;
  wire [10:0] add_176471;
  wire [11:0] sel_176474;
  wire [11:0] add_176499;
  wire [11:0] sel_176501;
  wire [11:0] add_176504;
  wire [11:0] sel_176506;
  wire [15:0] array_index_176535;
  wire [15:0] array_index_176538;
  wire [10:0] add_176542;
  wire [11:0] sel_176544;
  wire [10:0] add_176546;
  wire [11:0] sel_176548;
  wire [10:0] add_176550;
  wire [11:0] sel_176552;
  wire [10:0] add_176554;
  wire [11:0] sel_176556;
  wire [8:0] add_176558;
  wire [11:0] sel_176561;
  wire [8:0] add_176563;
  wire [11:0] sel_176566;
  wire [10:0] add_176568;
  wire [11:0] sel_176571;
  wire [10:0] add_176573;
  wire [11:0] sel_176576;
  wire [11:0] add_176601;
  wire [11:0] sel_176603;
  wire [11:0] add_176606;
  wire [11:0] sel_176608;
  wire [15:0] array_index_176637;
  wire [15:0] array_index_176640;
  wire [10:0] add_176644;
  wire [11:0] sel_176646;
  wire [10:0] add_176648;
  wire [11:0] sel_176650;
  wire [10:0] add_176652;
  wire [11:0] sel_176654;
  wire [10:0] add_176656;
  wire [11:0] sel_176658;
  wire [8:0] add_176660;
  wire [11:0] sel_176663;
  wire [8:0] add_176665;
  wire [11:0] sel_176668;
  wire [10:0] add_176670;
  wire [11:0] sel_176673;
  wire [10:0] add_176675;
  wire [11:0] sel_176678;
  wire [11:0] add_176703;
  wire [11:0] sel_176705;
  wire [11:0] add_176708;
  wire [11:0] sel_176710;
  wire [15:0] array_index_176739;
  wire [15:0] array_index_176742;
  wire [10:0] add_176746;
  wire [11:0] sel_176748;
  wire [10:0] add_176750;
  wire [11:0] sel_176752;
  wire [10:0] add_176754;
  wire [11:0] sel_176756;
  wire [10:0] add_176758;
  wire [11:0] sel_176760;
  wire [8:0] add_176762;
  wire [11:0] sel_176765;
  wire [8:0] add_176767;
  wire [11:0] sel_176770;
  wire [10:0] add_176772;
  wire [11:0] sel_176775;
  wire [10:0] add_176777;
  wire [11:0] sel_176780;
  wire [11:0] add_176805;
  wire [11:0] sel_176807;
  wire [11:0] add_176810;
  wire [11:0] sel_176812;
  wire [15:0] array_index_176841;
  wire [15:0] array_index_176844;
  wire [10:0] add_176848;
  wire [11:0] sel_176850;
  wire [10:0] add_176852;
  wire [11:0] sel_176854;
  wire [10:0] add_176856;
  wire [11:0] sel_176858;
  wire [10:0] add_176860;
  wire [11:0] sel_176862;
  wire [8:0] add_176864;
  wire [11:0] sel_176867;
  wire [8:0] add_176869;
  wire [11:0] sel_176872;
  wire [10:0] add_176874;
  wire [11:0] sel_176877;
  wire [10:0] add_176879;
  wire [11:0] sel_176882;
  wire [11:0] add_176907;
  wire [11:0] sel_176909;
  wire [11:0] add_176912;
  wire [11:0] sel_176914;
  wire [15:0] array_index_176943;
  wire [15:0] array_index_176946;
  wire [10:0] add_176950;
  wire [11:0] sel_176952;
  wire [10:0] add_176954;
  wire [11:0] sel_176956;
  wire [10:0] add_176958;
  wire [11:0] sel_176960;
  wire [10:0] add_176962;
  wire [11:0] sel_176964;
  wire [8:0] add_176966;
  wire [11:0] sel_176969;
  wire [8:0] add_176971;
  wire [11:0] sel_176974;
  wire [10:0] add_176976;
  wire [11:0] sel_176979;
  wire [10:0] add_176981;
  wire [11:0] sel_176984;
  wire [11:0] add_177009;
  wire [11:0] sel_177011;
  wire [11:0] add_177014;
  wire [11:0] sel_177016;
  wire [15:0] array_index_177045;
  wire [15:0] array_index_177048;
  wire [10:0] add_177052;
  wire [11:0] sel_177054;
  wire [10:0] add_177056;
  wire [11:0] sel_177058;
  wire [10:0] add_177060;
  wire [11:0] sel_177062;
  wire [10:0] add_177064;
  wire [11:0] sel_177066;
  wire [8:0] add_177068;
  wire [11:0] sel_177071;
  wire [8:0] add_177073;
  wire [11:0] sel_177076;
  wire [10:0] add_177078;
  wire [11:0] sel_177081;
  wire [10:0] add_177083;
  wire [11:0] sel_177086;
  wire [11:0] add_177111;
  wire [11:0] sel_177113;
  wire [11:0] add_177116;
  wire [11:0] sel_177118;
  wire [15:0] array_index_177147;
  wire [15:0] array_index_177150;
  wire [10:0] add_177154;
  wire [11:0] sel_177156;
  wire [10:0] add_177158;
  wire [11:0] sel_177160;
  wire [10:0] add_177162;
  wire [11:0] sel_177164;
  wire [10:0] add_177166;
  wire [11:0] sel_177168;
  wire [8:0] add_177170;
  wire [11:0] sel_177173;
  wire [8:0] add_177175;
  wire [11:0] sel_177178;
  wire [10:0] add_177180;
  wire [11:0] sel_177183;
  wire [10:0] add_177185;
  wire [11:0] sel_177188;
  wire [11:0] add_177213;
  wire [11:0] sel_177215;
  wire [11:0] add_177218;
  wire [11:0] sel_177220;
  wire [15:0] array_index_177249;
  wire [15:0] array_index_177252;
  wire [10:0] add_177256;
  wire [11:0] sel_177258;
  wire [10:0] add_177260;
  wire [11:0] sel_177262;
  wire [10:0] add_177264;
  wire [11:0] sel_177266;
  wire [10:0] add_177268;
  wire [11:0] sel_177270;
  wire [8:0] add_177272;
  wire [11:0] sel_177275;
  wire [8:0] add_177277;
  wire [11:0] sel_177280;
  wire [10:0] add_177282;
  wire [11:0] sel_177285;
  wire [10:0] add_177287;
  wire [11:0] sel_177290;
  wire [11:0] add_177315;
  wire [11:0] sel_177317;
  wire [11:0] add_177320;
  wire [11:0] sel_177322;
  wire [15:0] array_index_177351;
  wire [15:0] array_index_177354;
  wire [10:0] add_177358;
  wire [11:0] sel_177360;
  wire [10:0] add_177362;
  wire [11:0] sel_177364;
  wire [10:0] add_177366;
  wire [11:0] sel_177368;
  wire [10:0] add_177370;
  wire [11:0] sel_177372;
  wire [8:0] add_177374;
  wire [11:0] sel_177377;
  wire [8:0] add_177379;
  wire [11:0] sel_177382;
  wire [10:0] add_177384;
  wire [11:0] sel_177387;
  wire [10:0] add_177389;
  wire [11:0] sel_177392;
  wire [11:0] add_177417;
  wire [11:0] sel_177419;
  wire [11:0] add_177422;
  wire [11:0] sel_177424;
  wire [15:0] array_index_177453;
  wire [15:0] array_index_177456;
  wire [10:0] add_177460;
  wire [11:0] sel_177462;
  wire [10:0] add_177464;
  wire [11:0] sel_177466;
  wire [10:0] add_177468;
  wire [11:0] sel_177470;
  wire [10:0] add_177472;
  wire [11:0] sel_177474;
  wire [8:0] add_177476;
  wire [11:0] sel_177479;
  wire [8:0] add_177481;
  wire [11:0] sel_177484;
  wire [10:0] add_177486;
  wire [11:0] sel_177489;
  wire [10:0] add_177491;
  wire [11:0] sel_177494;
  wire [11:0] add_177519;
  wire [11:0] sel_177521;
  wire [11:0] add_177524;
  wire [11:0] sel_177526;
  wire [15:0] array_index_177555;
  wire [15:0] array_index_177558;
  wire [10:0] add_177562;
  wire [11:0] sel_177564;
  wire [10:0] add_177566;
  wire [11:0] sel_177568;
  wire [10:0] add_177570;
  wire [11:0] sel_177572;
  wire [10:0] add_177574;
  wire [11:0] sel_177576;
  wire [8:0] add_177578;
  wire [11:0] sel_177581;
  wire [8:0] add_177583;
  wire [11:0] sel_177586;
  wire [10:0] add_177588;
  wire [11:0] sel_177591;
  wire [10:0] add_177593;
  wire [11:0] sel_177596;
  wire [11:0] add_177621;
  wire [11:0] sel_177623;
  wire [11:0] add_177626;
  wire [11:0] sel_177628;
  wire [15:0] array_index_177657;
  wire [15:0] array_index_177660;
  wire [10:0] add_177664;
  wire [11:0] sel_177666;
  wire [10:0] add_177668;
  wire [11:0] sel_177670;
  wire [10:0] add_177672;
  wire [11:0] sel_177674;
  wire [10:0] add_177676;
  wire [11:0] sel_177678;
  wire [8:0] add_177680;
  wire [11:0] sel_177683;
  wire [8:0] add_177685;
  wire [11:0] sel_177688;
  wire [10:0] add_177690;
  wire [11:0] sel_177693;
  wire [10:0] add_177695;
  wire [11:0] sel_177698;
  wire [11:0] add_177723;
  wire [11:0] sel_177725;
  wire [11:0] add_177728;
  wire [11:0] sel_177730;
  wire [15:0] array_index_177759;
  wire [15:0] array_index_177762;
  wire [10:0] add_177766;
  wire [11:0] sel_177768;
  wire [10:0] add_177770;
  wire [11:0] sel_177772;
  wire [10:0] add_177774;
  wire [11:0] sel_177776;
  wire [10:0] add_177778;
  wire [11:0] sel_177780;
  wire [8:0] add_177782;
  wire [11:0] sel_177785;
  wire [8:0] add_177787;
  wire [11:0] sel_177790;
  wire [10:0] add_177792;
  wire [11:0] sel_177795;
  wire [10:0] add_177797;
  wire [11:0] sel_177800;
  wire [11:0] add_177825;
  wire [11:0] sel_177827;
  wire [11:0] add_177830;
  wire [11:0] sel_177832;
  wire [15:0] array_index_177861;
  wire [15:0] array_index_177864;
  wire [10:0] add_177868;
  wire [11:0] sel_177870;
  wire [10:0] add_177872;
  wire [11:0] sel_177874;
  wire [10:0] add_177876;
  wire [11:0] sel_177878;
  wire [10:0] add_177880;
  wire [11:0] sel_177882;
  wire [8:0] add_177884;
  wire [11:0] sel_177887;
  wire [8:0] add_177889;
  wire [11:0] sel_177892;
  wire [10:0] add_177894;
  wire [11:0] sel_177897;
  wire [10:0] add_177899;
  wire [11:0] sel_177902;
  wire [11:0] add_177927;
  wire [11:0] sel_177929;
  wire [11:0] add_177932;
  wire [11:0] sel_177934;
  wire [15:0] array_index_177963;
  wire [15:0] array_index_177966;
  wire [10:0] add_177970;
  wire [11:0] sel_177972;
  wire [10:0] add_177974;
  wire [11:0] sel_177976;
  wire [10:0] add_177978;
  wire [11:0] sel_177980;
  wire [10:0] add_177982;
  wire [11:0] sel_177984;
  wire [8:0] add_177986;
  wire [11:0] sel_177989;
  wire [8:0] add_177991;
  wire [11:0] sel_177994;
  wire [10:0] add_177996;
  wire [11:0] sel_177999;
  wire [10:0] add_178001;
  wire [11:0] sel_178004;
  wire [11:0] add_178029;
  wire [11:0] sel_178031;
  wire [11:0] add_178034;
  wire [11:0] sel_178036;
  wire [15:0] array_index_178065;
  wire [15:0] array_index_178068;
  wire [10:0] add_178072;
  wire [11:0] sel_178074;
  wire [10:0] add_178076;
  wire [11:0] sel_178078;
  wire [10:0] add_178080;
  wire [11:0] sel_178082;
  wire [10:0] add_178084;
  wire [11:0] sel_178086;
  wire [8:0] add_178088;
  wire [11:0] sel_178091;
  wire [8:0] add_178093;
  wire [11:0] sel_178096;
  wire [10:0] add_178098;
  wire [11:0] sel_178101;
  wire [10:0] add_178103;
  wire [11:0] sel_178106;
  wire [11:0] add_178131;
  wire [11:0] sel_178133;
  wire [11:0] add_178136;
  wire [11:0] sel_178138;
  wire [15:0] array_index_178167;
  wire [15:0] array_index_178170;
  wire [10:0] add_178174;
  wire [11:0] sel_178176;
  wire [10:0] add_178178;
  wire [11:0] sel_178180;
  wire [10:0] add_178182;
  wire [11:0] sel_178184;
  wire [10:0] add_178186;
  wire [11:0] sel_178188;
  wire [8:0] add_178190;
  wire [11:0] sel_178193;
  wire [8:0] add_178195;
  wire [11:0] sel_178198;
  wire [10:0] add_178200;
  wire [11:0] sel_178203;
  wire [10:0] add_178205;
  wire [11:0] sel_178208;
  wire [11:0] add_178233;
  wire [11:0] sel_178235;
  wire [11:0] add_178238;
  wire [11:0] sel_178240;
  wire [15:0] array_index_178269;
  wire [15:0] array_index_178272;
  wire [10:0] add_178276;
  wire [11:0] sel_178278;
  wire [10:0] add_178280;
  wire [11:0] sel_178282;
  wire [10:0] add_178284;
  wire [11:0] sel_178286;
  wire [10:0] add_178288;
  wire [11:0] sel_178290;
  wire [8:0] add_178292;
  wire [11:0] sel_178295;
  wire [8:0] add_178297;
  wire [11:0] sel_178300;
  wire [10:0] add_178302;
  wire [11:0] sel_178305;
  wire [10:0] add_178307;
  wire [11:0] sel_178310;
  wire [11:0] add_178335;
  wire [11:0] sel_178337;
  wire [11:0] add_178340;
  wire [11:0] sel_178342;
  wire [15:0] array_index_178371;
  wire [15:0] array_index_178374;
  wire [10:0] add_178378;
  wire [11:0] sel_178380;
  wire [10:0] add_178382;
  wire [11:0] sel_178384;
  wire [10:0] add_178386;
  wire [11:0] sel_178388;
  wire [10:0] add_178390;
  wire [11:0] sel_178392;
  wire [8:0] add_178394;
  wire [11:0] sel_178397;
  wire [8:0] add_178399;
  wire [11:0] sel_178402;
  wire [10:0] add_178404;
  wire [11:0] sel_178407;
  wire [10:0] add_178409;
  wire [11:0] sel_178412;
  wire [11:0] add_178437;
  wire [11:0] sel_178439;
  wire [11:0] add_178442;
  wire [11:0] sel_178444;
  wire [15:0] array_index_178473;
  wire [15:0] array_index_178476;
  wire [10:0] add_178480;
  wire [11:0] sel_178482;
  wire [10:0] add_178484;
  wire [11:0] sel_178486;
  wire [10:0] add_178488;
  wire [11:0] sel_178490;
  wire [10:0] add_178492;
  wire [11:0] sel_178494;
  wire [8:0] add_178496;
  wire [11:0] sel_178499;
  wire [8:0] add_178501;
  wire [11:0] sel_178504;
  wire [10:0] add_178506;
  wire [11:0] sel_178509;
  wire [10:0] add_178511;
  wire [11:0] sel_178514;
  wire [11:0] add_178539;
  wire [11:0] sel_178541;
  wire [11:0] add_178544;
  wire [11:0] sel_178546;
  wire [15:0] array_index_178575;
  wire [15:0] array_index_178578;
  wire [10:0] add_178582;
  wire [11:0] sel_178584;
  wire [10:0] add_178586;
  wire [11:0] sel_178588;
  wire [10:0] add_178590;
  wire [11:0] sel_178592;
  wire [10:0] add_178594;
  wire [11:0] sel_178596;
  wire [8:0] add_178598;
  wire [11:0] sel_178601;
  wire [8:0] add_178603;
  wire [11:0] sel_178606;
  wire [10:0] add_178608;
  wire [11:0] sel_178611;
  wire [10:0] add_178613;
  wire [11:0] sel_178616;
  wire [11:0] add_178641;
  wire [11:0] sel_178643;
  wire [11:0] add_178646;
  wire [11:0] sel_178648;
  wire [15:0] array_index_178677;
  wire [15:0] array_index_178680;
  wire [10:0] add_178684;
  wire [11:0] sel_178686;
  wire [10:0] add_178688;
  wire [11:0] sel_178690;
  wire [10:0] add_178692;
  wire [11:0] sel_178694;
  wire [10:0] add_178696;
  wire [11:0] sel_178698;
  wire [8:0] add_178700;
  wire [11:0] sel_178703;
  wire [8:0] add_178705;
  wire [11:0] sel_178708;
  wire [10:0] add_178710;
  wire [11:0] sel_178713;
  wire [10:0] add_178715;
  wire [11:0] sel_178718;
  wire [11:0] add_178743;
  wire [11:0] sel_178745;
  wire [11:0] add_178748;
  wire [11:0] sel_178750;
  wire [15:0] array_index_178779;
  wire [15:0] array_index_178782;
  wire [10:0] add_178786;
  wire [11:0] sel_178788;
  wire [10:0] add_178790;
  wire [11:0] sel_178792;
  wire [10:0] add_178794;
  wire [11:0] sel_178796;
  wire [10:0] add_178798;
  wire [11:0] sel_178800;
  wire [8:0] add_178802;
  wire [11:0] sel_178805;
  wire [8:0] add_178807;
  wire [11:0] sel_178810;
  wire [10:0] add_178812;
  wire [11:0] sel_178815;
  wire [10:0] add_178817;
  wire [11:0] sel_178820;
  wire [11:0] add_178845;
  wire [11:0] sel_178847;
  wire [11:0] add_178850;
  wire [11:0] sel_178852;
  wire [15:0] array_index_178881;
  wire [15:0] array_index_178884;
  wire [10:0] add_178888;
  wire [11:0] sel_178890;
  wire [10:0] add_178892;
  wire [11:0] sel_178894;
  wire [10:0] add_178896;
  wire [11:0] sel_178898;
  wire [10:0] add_178900;
  wire [11:0] sel_178902;
  wire [8:0] add_178904;
  wire [11:0] sel_178907;
  wire [8:0] add_178909;
  wire [11:0] sel_178912;
  wire [10:0] add_178914;
  wire [11:0] sel_178917;
  wire [10:0] add_178919;
  wire [11:0] sel_178922;
  wire [11:0] add_178947;
  wire [11:0] sel_178949;
  wire [11:0] add_178952;
  wire [11:0] sel_178954;
  wire [15:0] array_index_178983;
  wire [15:0] array_index_178986;
  wire [10:0] add_178990;
  wire [11:0] sel_178992;
  wire [10:0] add_178994;
  wire [11:0] sel_178996;
  wire [10:0] add_178998;
  wire [11:0] sel_179000;
  wire [10:0] add_179002;
  wire [11:0] sel_179004;
  wire [8:0] add_179006;
  wire [11:0] sel_179009;
  wire [8:0] add_179011;
  wire [11:0] sel_179014;
  wire [10:0] add_179016;
  wire [11:0] sel_179019;
  wire [10:0] add_179021;
  wire [11:0] sel_179024;
  wire [11:0] add_179049;
  wire [11:0] sel_179051;
  wire [11:0] add_179054;
  wire [11:0] sel_179056;
  wire [15:0] array_index_179085;
  wire [15:0] array_index_179088;
  wire [10:0] add_179092;
  wire [11:0] sel_179094;
  wire [10:0] add_179096;
  wire [11:0] sel_179098;
  wire [10:0] add_179100;
  wire [11:0] sel_179102;
  wire [10:0] add_179104;
  wire [11:0] sel_179106;
  wire [8:0] add_179108;
  wire [11:0] sel_179111;
  wire [8:0] add_179113;
  wire [11:0] sel_179116;
  wire [10:0] add_179118;
  wire [11:0] sel_179121;
  wire [10:0] add_179123;
  wire [11:0] sel_179126;
  wire [11:0] add_179151;
  wire [11:0] sel_179153;
  wire [11:0] add_179156;
  wire [11:0] sel_179158;
  wire [15:0] array_index_179187;
  wire [15:0] array_index_179190;
  wire [10:0] add_179194;
  wire [11:0] sel_179196;
  wire [10:0] add_179198;
  wire [11:0] sel_179200;
  wire [10:0] add_179202;
  wire [11:0] sel_179204;
  wire [10:0] add_179206;
  wire [11:0] sel_179208;
  wire [8:0] add_179210;
  wire [11:0] sel_179213;
  wire [8:0] add_179215;
  wire [11:0] sel_179218;
  wire [10:0] add_179220;
  wire [11:0] sel_179223;
  wire [10:0] add_179225;
  wire [11:0] sel_179228;
  wire [11:0] add_179253;
  wire [11:0] sel_179255;
  wire [11:0] add_179258;
  wire [11:0] sel_179260;
  wire [15:0] array_index_179289;
  wire [15:0] array_index_179292;
  wire [10:0] add_179296;
  wire [11:0] sel_179298;
  wire [10:0] add_179300;
  wire [11:0] sel_179302;
  wire [10:0] add_179304;
  wire [11:0] sel_179306;
  wire [10:0] add_179308;
  wire [11:0] sel_179310;
  wire [8:0] add_179312;
  wire [11:0] sel_179315;
  wire [8:0] add_179317;
  wire [11:0] sel_179320;
  wire [10:0] add_179322;
  wire [11:0] sel_179325;
  wire [10:0] add_179327;
  wire [11:0] sel_179330;
  wire [11:0] add_179355;
  wire [11:0] sel_179357;
  wire [11:0] add_179360;
  wire [11:0] sel_179362;
  wire [15:0] array_index_179391;
  wire [15:0] array_index_179394;
  wire [10:0] add_179398;
  wire [11:0] sel_179400;
  wire [10:0] add_179402;
  wire [11:0] sel_179404;
  wire [10:0] add_179406;
  wire [11:0] sel_179408;
  wire [10:0] add_179410;
  wire [11:0] sel_179412;
  wire [8:0] add_179414;
  wire [11:0] sel_179417;
  wire [8:0] add_179419;
  wire [11:0] sel_179422;
  wire [10:0] add_179424;
  wire [11:0] sel_179427;
  wire [10:0] add_179429;
  wire [11:0] sel_179432;
  wire [11:0] add_179457;
  wire [11:0] sel_179459;
  wire [11:0] add_179462;
  wire [11:0] sel_179464;
  wire [15:0] array_index_179493;
  wire [15:0] array_index_179496;
  wire [10:0] add_179500;
  wire [11:0] sel_179502;
  wire [10:0] add_179504;
  wire [11:0] sel_179506;
  wire [10:0] add_179508;
  wire [11:0] sel_179510;
  wire [10:0] add_179512;
  wire [11:0] sel_179514;
  wire [8:0] add_179516;
  wire [11:0] sel_179519;
  wire [8:0] add_179521;
  wire [11:0] sel_179524;
  wire [10:0] add_179526;
  wire [11:0] sel_179529;
  wire [10:0] add_179531;
  wire [11:0] sel_179534;
  wire [11:0] add_179559;
  wire [11:0] sel_179561;
  wire [11:0] add_179564;
  wire [11:0] sel_179566;
  wire [15:0] array_index_179595;
  wire [15:0] array_index_179598;
  wire [10:0] add_179602;
  wire [11:0] sel_179604;
  wire [10:0] add_179606;
  wire [11:0] sel_179608;
  wire [10:0] add_179610;
  wire [11:0] sel_179612;
  wire [10:0] add_179614;
  wire [11:0] sel_179616;
  wire [8:0] add_179618;
  wire [11:0] sel_179621;
  wire [8:0] add_179623;
  wire [11:0] sel_179626;
  wire [10:0] add_179628;
  wire [11:0] sel_179631;
  wire [10:0] add_179633;
  wire [11:0] sel_179636;
  wire [11:0] add_179661;
  wire [11:0] sel_179663;
  wire [11:0] add_179666;
  wire [11:0] sel_179668;
  wire [15:0] array_index_179697;
  wire [15:0] array_index_179700;
  wire [10:0] add_179704;
  wire [11:0] sel_179706;
  wire [10:0] add_179708;
  wire [11:0] sel_179710;
  wire [10:0] add_179712;
  wire [11:0] sel_179714;
  wire [10:0] add_179716;
  wire [11:0] sel_179718;
  wire [8:0] add_179720;
  wire [11:0] sel_179723;
  wire [8:0] add_179725;
  wire [11:0] sel_179728;
  wire [10:0] add_179730;
  wire [11:0] sel_179733;
  wire [10:0] add_179735;
  wire [11:0] sel_179738;
  wire [11:0] add_179763;
  wire [11:0] sel_179765;
  wire [11:0] add_179768;
  wire [11:0] sel_179770;
  wire [15:0] array_index_179799;
  wire [15:0] array_index_179802;
  wire [10:0] add_179806;
  wire [11:0] sel_179808;
  wire [10:0] add_179810;
  wire [11:0] sel_179812;
  wire [10:0] add_179814;
  wire [11:0] sel_179816;
  wire [10:0] add_179818;
  wire [11:0] sel_179820;
  wire [8:0] add_179822;
  wire [11:0] sel_179825;
  wire [8:0] add_179827;
  wire [11:0] sel_179830;
  wire [10:0] add_179832;
  wire [11:0] sel_179835;
  wire [10:0] add_179837;
  wire [11:0] sel_179840;
  wire [11:0] add_179865;
  wire [11:0] sel_179867;
  wire [11:0] add_179870;
  wire [11:0] sel_179872;
  wire [15:0] array_index_179901;
  wire [15:0] array_index_179904;
  wire [10:0] add_179908;
  wire [11:0] sel_179910;
  wire [10:0] add_179912;
  wire [11:0] sel_179914;
  wire [10:0] add_179916;
  wire [11:0] sel_179918;
  wire [10:0] add_179920;
  wire [11:0] sel_179922;
  wire [8:0] add_179924;
  wire [11:0] sel_179927;
  wire [8:0] add_179929;
  wire [11:0] sel_179932;
  wire [10:0] add_179934;
  wire [11:0] sel_179937;
  wire [10:0] add_179939;
  wire [11:0] sel_179942;
  wire [11:0] add_179967;
  wire [11:0] sel_179969;
  wire [11:0] add_179972;
  wire [11:0] sel_179974;
  wire [15:0] array_index_180003;
  wire [15:0] array_index_180006;
  wire [10:0] add_180010;
  wire [11:0] sel_180012;
  wire [10:0] add_180014;
  wire [11:0] sel_180016;
  wire [10:0] add_180018;
  wire [11:0] sel_180020;
  wire [10:0] add_180022;
  wire [11:0] sel_180024;
  wire [8:0] add_180026;
  wire [11:0] sel_180029;
  wire [8:0] add_180031;
  wire [11:0] sel_180034;
  wire [10:0] add_180036;
  wire [11:0] sel_180039;
  wire [10:0] add_180041;
  wire [11:0] sel_180044;
  wire [11:0] add_180069;
  wire [11:0] sel_180071;
  wire [11:0] add_180074;
  wire [11:0] sel_180076;
  wire [15:0] array_index_180105;
  wire [15:0] array_index_180108;
  wire [10:0] add_180112;
  wire [11:0] sel_180114;
  wire [10:0] add_180116;
  wire [11:0] sel_180118;
  wire [10:0] add_180120;
  wire [11:0] sel_180122;
  wire [10:0] add_180124;
  wire [11:0] sel_180126;
  wire [8:0] add_180128;
  wire [11:0] sel_180131;
  wire [8:0] add_180133;
  wire [11:0] sel_180136;
  wire [10:0] add_180138;
  wire [11:0] sel_180141;
  wire [10:0] add_180143;
  wire [11:0] sel_180146;
  wire [11:0] add_180171;
  wire [11:0] sel_180173;
  wire [11:0] add_180176;
  wire [11:0] sel_180178;
  wire [15:0] array_index_180207;
  wire [15:0] array_index_180210;
  wire [10:0] add_180214;
  wire [11:0] sel_180216;
  wire [10:0] add_180218;
  wire [11:0] sel_180220;
  wire [10:0] add_180222;
  wire [11:0] sel_180224;
  wire [10:0] add_180226;
  wire [11:0] sel_180228;
  wire [8:0] add_180230;
  wire [11:0] sel_180233;
  wire [8:0] add_180235;
  wire [11:0] sel_180238;
  wire [10:0] add_180240;
  wire [11:0] sel_180243;
  wire [10:0] add_180245;
  wire [11:0] sel_180248;
  wire [11:0] add_180273;
  wire [11:0] sel_180275;
  wire [11:0] add_180278;
  wire [11:0] sel_180280;
  wire [15:0] array_index_180309;
  wire [15:0] array_index_180312;
  wire [10:0] add_180316;
  wire [11:0] sel_180318;
  wire [10:0] add_180320;
  wire [11:0] sel_180322;
  wire [10:0] add_180324;
  wire [11:0] sel_180326;
  wire [10:0] add_180328;
  wire [11:0] sel_180330;
  wire [8:0] add_180332;
  wire [11:0] sel_180335;
  wire [8:0] add_180337;
  wire [11:0] sel_180340;
  wire [10:0] add_180342;
  wire [11:0] sel_180345;
  wire [10:0] add_180347;
  wire [11:0] sel_180350;
  wire [11:0] add_180375;
  wire [11:0] sel_180377;
  wire [11:0] add_180380;
  wire [11:0] sel_180382;
  wire [15:0] array_index_180411;
  wire [15:0] array_index_180414;
  wire [10:0] add_180418;
  wire [11:0] sel_180420;
  wire [10:0] add_180422;
  wire [11:0] sel_180424;
  wire [10:0] add_180426;
  wire [11:0] sel_180428;
  wire [10:0] add_180430;
  wire [11:0] sel_180432;
  wire [8:0] add_180434;
  wire [11:0] sel_180437;
  wire [8:0] add_180439;
  wire [11:0] sel_180442;
  wire [10:0] add_180444;
  wire [11:0] sel_180447;
  wire [10:0] add_180449;
  wire [11:0] sel_180452;
  wire [11:0] add_180477;
  wire [11:0] sel_180479;
  wire [11:0] add_180482;
  wire [11:0] sel_180484;
  wire [15:0] array_index_180513;
  wire [15:0] array_index_180516;
  wire [10:0] add_180520;
  wire [11:0] sel_180522;
  wire [10:0] add_180524;
  wire [11:0] sel_180526;
  wire [10:0] add_180528;
  wire [11:0] sel_180530;
  wire [10:0] add_180532;
  wire [11:0] sel_180534;
  wire [8:0] add_180536;
  wire [11:0] sel_180539;
  wire [8:0] add_180541;
  wire [11:0] sel_180544;
  wire [10:0] add_180546;
  wire [11:0] sel_180549;
  wire [10:0] add_180551;
  wire [11:0] sel_180554;
  wire [11:0] add_180579;
  wire [11:0] sel_180581;
  wire [11:0] add_180584;
  wire [11:0] sel_180586;
  wire [15:0] array_index_180615;
  wire [15:0] array_index_180618;
  wire [10:0] add_180622;
  wire [11:0] sel_180624;
  wire [10:0] add_180626;
  wire [11:0] sel_180628;
  wire [10:0] add_180630;
  wire [11:0] sel_180632;
  wire [10:0] add_180634;
  wire [11:0] sel_180636;
  wire [8:0] add_180638;
  wire [11:0] sel_180641;
  wire [8:0] add_180643;
  wire [11:0] sel_180646;
  wire [10:0] add_180648;
  wire [11:0] sel_180651;
  wire [10:0] add_180653;
  wire [11:0] sel_180656;
  wire [11:0] add_180681;
  wire [11:0] sel_180683;
  wire [11:0] add_180686;
  wire [11:0] sel_180688;
  wire [15:0] array_index_180717;
  wire [15:0] array_index_180720;
  wire [10:0] add_180724;
  wire [11:0] sel_180726;
  wire [10:0] add_180728;
  wire [11:0] sel_180730;
  wire [10:0] add_180732;
  wire [11:0] sel_180734;
  wire [10:0] add_180736;
  wire [11:0] sel_180738;
  wire [8:0] add_180740;
  wire [11:0] sel_180743;
  wire [8:0] add_180745;
  wire [11:0] sel_180748;
  wire [10:0] add_180750;
  wire [11:0] sel_180753;
  wire [10:0] add_180755;
  wire [11:0] sel_180758;
  wire [11:0] add_180783;
  wire [11:0] sel_180785;
  wire [11:0] add_180788;
  wire [11:0] sel_180790;
  wire [15:0] array_index_180819;
  wire [15:0] array_index_180822;
  wire [10:0] add_180826;
  wire [11:0] sel_180828;
  wire [10:0] add_180830;
  wire [11:0] sel_180832;
  wire [10:0] add_180834;
  wire [11:0] sel_180836;
  wire [10:0] add_180838;
  wire [11:0] sel_180840;
  wire [8:0] add_180842;
  wire [11:0] sel_180845;
  wire [8:0] add_180847;
  wire [11:0] sel_180850;
  wire [10:0] add_180852;
  wire [11:0] sel_180855;
  wire [10:0] add_180857;
  wire [11:0] sel_180860;
  wire [11:0] add_180885;
  wire [11:0] sel_180887;
  wire [11:0] add_180890;
  wire [11:0] sel_180892;
  wire [15:0] array_index_180921;
  wire [15:0] array_index_180924;
  wire [10:0] add_180928;
  wire [11:0] sel_180930;
  wire [10:0] add_180932;
  wire [11:0] sel_180934;
  wire [10:0] add_180936;
  wire [11:0] sel_180938;
  wire [10:0] add_180940;
  wire [11:0] sel_180942;
  wire [8:0] add_180944;
  wire [11:0] sel_180947;
  wire [8:0] add_180949;
  wire [11:0] sel_180952;
  wire [10:0] add_180954;
  wire [11:0] sel_180957;
  wire [10:0] add_180959;
  wire [11:0] sel_180962;
  wire [11:0] add_180987;
  wire [11:0] sel_180989;
  wire [11:0] add_180992;
  wire [11:0] sel_180994;
  wire [15:0] array_index_181023;
  wire [15:0] array_index_181026;
  wire [10:0] add_181030;
  wire [11:0] sel_181032;
  wire [10:0] add_181034;
  wire [11:0] sel_181036;
  wire [10:0] add_181038;
  wire [11:0] sel_181040;
  wire [10:0] add_181042;
  wire [11:0] sel_181044;
  wire [8:0] add_181046;
  wire [11:0] sel_181049;
  wire [8:0] add_181051;
  wire [11:0] sel_181054;
  wire [10:0] add_181056;
  wire [11:0] sel_181059;
  wire [10:0] add_181061;
  wire [11:0] sel_181064;
  wire [11:0] add_181089;
  wire [11:0] sel_181091;
  wire [11:0] add_181094;
  wire [11:0] sel_181096;
  wire [15:0] array_index_181125;
  wire [15:0] array_index_181128;
  wire [10:0] add_181132;
  wire [11:0] sel_181134;
  wire [10:0] add_181136;
  wire [11:0] sel_181138;
  wire [10:0] add_181140;
  wire [11:0] sel_181142;
  wire [10:0] add_181144;
  wire [11:0] sel_181146;
  wire [8:0] add_181148;
  wire [11:0] sel_181151;
  wire [8:0] add_181153;
  wire [11:0] sel_181156;
  wire [10:0] add_181158;
  wire [11:0] sel_181161;
  wire [10:0] add_181163;
  wire [11:0] sel_181166;
  wire [11:0] add_181191;
  wire [11:0] sel_181193;
  wire [11:0] add_181196;
  wire [11:0] sel_181198;
  wire [15:0] array_index_181227;
  wire [15:0] array_index_181230;
  wire [10:0] add_181234;
  wire [11:0] sel_181236;
  wire [10:0] add_181238;
  wire [11:0] sel_181240;
  wire [10:0] add_181242;
  wire [11:0] sel_181244;
  wire [10:0] add_181246;
  wire [11:0] sel_181248;
  wire [8:0] add_181250;
  wire [11:0] sel_181253;
  wire [8:0] add_181255;
  wire [11:0] sel_181258;
  wire [10:0] add_181260;
  wire [11:0] sel_181263;
  wire [10:0] add_181265;
  wire [11:0] sel_181268;
  wire [11:0] add_181293;
  wire [11:0] sel_181295;
  wire [11:0] add_181298;
  wire [11:0] sel_181300;
  wire [15:0] array_index_181329;
  wire [15:0] array_index_181332;
  wire [10:0] add_181336;
  wire [11:0] sel_181338;
  wire [10:0] add_181340;
  wire [11:0] sel_181342;
  wire [10:0] add_181344;
  wire [11:0] sel_181346;
  wire [10:0] add_181348;
  wire [11:0] sel_181350;
  wire [8:0] add_181352;
  wire [11:0] sel_181355;
  wire [8:0] add_181357;
  wire [11:0] sel_181360;
  wire [10:0] add_181362;
  wire [11:0] sel_181365;
  wire [10:0] add_181367;
  wire [11:0] sel_181370;
  wire [11:0] add_181395;
  wire [11:0] sel_181397;
  wire [11:0] add_181400;
  wire [11:0] sel_181402;
  wire [15:0] array_index_181431;
  wire [15:0] array_index_181434;
  wire [10:0] add_181438;
  wire [11:0] sel_181440;
  wire [10:0] add_181442;
  wire [11:0] sel_181444;
  wire [10:0] add_181446;
  wire [11:0] sel_181448;
  wire [10:0] add_181450;
  wire [11:0] sel_181452;
  wire [8:0] add_181454;
  wire [11:0] sel_181457;
  wire [8:0] add_181459;
  wire [11:0] sel_181462;
  wire [10:0] add_181464;
  wire [11:0] sel_181467;
  wire [10:0] add_181469;
  wire [11:0] sel_181472;
  wire [11:0] add_181497;
  wire [11:0] sel_181499;
  wire [11:0] add_181502;
  wire [11:0] sel_181504;
  wire [15:0] array_index_181533;
  wire [15:0] array_index_181536;
  wire [10:0] add_181540;
  wire [11:0] sel_181542;
  wire [10:0] add_181544;
  wire [11:0] sel_181546;
  wire [10:0] add_181548;
  wire [11:0] sel_181550;
  wire [10:0] add_181552;
  wire [11:0] sel_181554;
  wire [8:0] add_181556;
  wire [11:0] sel_181559;
  wire [8:0] add_181561;
  wire [11:0] sel_181564;
  wire [10:0] add_181566;
  wire [11:0] sel_181569;
  wire [10:0] add_181571;
  wire [11:0] sel_181574;
  wire [11:0] add_181599;
  wire [11:0] sel_181601;
  wire [11:0] add_181604;
  wire [11:0] sel_181606;
  wire [15:0] array_index_181635;
  wire [15:0] array_index_181638;
  wire [10:0] add_181642;
  wire [11:0] sel_181644;
  wire [10:0] add_181646;
  wire [11:0] sel_181648;
  wire [10:0] add_181650;
  wire [11:0] sel_181652;
  wire [10:0] add_181654;
  wire [11:0] sel_181656;
  wire [8:0] add_181658;
  wire [11:0] sel_181661;
  wire [8:0] add_181663;
  wire [11:0] sel_181666;
  wire [10:0] add_181668;
  wire [11:0] sel_181671;
  wire [10:0] add_181673;
  wire [11:0] sel_181676;
  wire [11:0] add_181701;
  wire [11:0] sel_181703;
  wire [11:0] add_181706;
  wire [11:0] sel_181708;
  wire [15:0] array_index_181737;
  wire [15:0] array_index_181740;
  wire [10:0] add_181744;
  wire [11:0] sel_181746;
  wire [10:0] add_181748;
  wire [11:0] sel_181750;
  wire [10:0] add_181752;
  wire [11:0] sel_181754;
  wire [10:0] add_181756;
  wire [11:0] sel_181758;
  wire [8:0] add_181760;
  wire [11:0] sel_181763;
  wire [8:0] add_181765;
  wire [11:0] sel_181768;
  wire [10:0] add_181770;
  wire [11:0] sel_181773;
  wire [10:0] add_181775;
  wire [11:0] sel_181778;
  wire [11:0] add_181803;
  wire [11:0] sel_181805;
  wire [11:0] add_181808;
  wire [11:0] sel_181810;
  wire [15:0] array_index_181839;
  wire [15:0] array_index_181842;
  wire [10:0] add_181846;
  wire [11:0] sel_181848;
  wire [10:0] add_181850;
  wire [11:0] sel_181852;
  wire [10:0] add_181854;
  wire [11:0] sel_181856;
  wire [10:0] add_181858;
  wire [11:0] sel_181860;
  wire [8:0] add_181862;
  wire [11:0] sel_181865;
  wire [8:0] add_181867;
  wire [11:0] sel_181870;
  wire [10:0] add_181872;
  wire [11:0] sel_181875;
  wire [10:0] add_181877;
  wire [11:0] sel_181880;
  wire [11:0] add_181905;
  wire [11:0] sel_181907;
  wire [11:0] add_181910;
  wire [11:0] sel_181912;
  wire [15:0] array_index_181941;
  wire [15:0] array_index_181944;
  wire [10:0] add_181948;
  wire [11:0] sel_181950;
  wire [10:0] add_181952;
  wire [11:0] sel_181954;
  wire [10:0] add_181956;
  wire [11:0] sel_181958;
  wire [10:0] add_181960;
  wire [11:0] sel_181962;
  wire [8:0] add_181964;
  wire [11:0] sel_181967;
  wire [8:0] add_181969;
  wire [11:0] sel_181972;
  wire [10:0] add_181974;
  wire [11:0] sel_181977;
  wire [10:0] add_181979;
  wire [11:0] sel_181982;
  wire [11:0] add_182007;
  wire [11:0] sel_182009;
  wire [11:0] add_182012;
  wire [11:0] sel_182014;
  wire [15:0] array_index_182043;
  wire [15:0] array_index_182046;
  wire [10:0] add_182050;
  wire [11:0] sel_182052;
  wire [10:0] add_182054;
  wire [11:0] sel_182056;
  wire [10:0] add_182058;
  wire [11:0] sel_182060;
  wire [10:0] add_182062;
  wire [11:0] sel_182064;
  wire [8:0] add_182066;
  wire [11:0] sel_182069;
  wire [8:0] add_182071;
  wire [11:0] sel_182074;
  wire [10:0] add_182076;
  wire [11:0] sel_182079;
  wire [10:0] add_182081;
  wire [11:0] sel_182084;
  wire [11:0] add_182109;
  wire [11:0] sel_182111;
  wire [11:0] add_182114;
  wire [11:0] sel_182116;
  wire [15:0] array_index_182145;
  wire [15:0] array_index_182148;
  wire [10:0] add_182152;
  wire [11:0] sel_182154;
  wire [10:0] add_182156;
  wire [11:0] sel_182158;
  wire [10:0] add_182160;
  wire [11:0] sel_182162;
  wire [10:0] add_182164;
  wire [11:0] sel_182166;
  wire [8:0] add_182168;
  wire [11:0] sel_182171;
  wire [8:0] add_182173;
  wire [11:0] sel_182176;
  wire [10:0] add_182178;
  wire [11:0] sel_182181;
  wire [10:0] add_182183;
  wire [11:0] sel_182186;
  wire [11:0] add_182211;
  wire [11:0] sel_182213;
  wire [11:0] add_182216;
  wire [11:0] sel_182218;
  wire [15:0] array_index_182247;
  wire [15:0] array_index_182250;
  wire [10:0] add_182254;
  wire [11:0] sel_182256;
  wire [10:0] add_182258;
  wire [11:0] sel_182260;
  wire [10:0] add_182262;
  wire [11:0] sel_182264;
  wire [10:0] add_182266;
  wire [11:0] sel_182268;
  wire [8:0] add_182270;
  wire [11:0] sel_182273;
  wire [8:0] add_182275;
  wire [11:0] sel_182278;
  wire [10:0] add_182280;
  wire [11:0] sel_182283;
  wire [10:0] add_182285;
  wire [11:0] sel_182288;
  wire [11:0] add_182313;
  wire [11:0] sel_182315;
  wire [11:0] add_182318;
  wire [11:0] sel_182320;
  wire [15:0] array_index_182349;
  wire [15:0] array_index_182352;
  wire [10:0] add_182356;
  wire [11:0] sel_182358;
  wire [10:0] add_182360;
  wire [11:0] sel_182362;
  wire [10:0] add_182364;
  wire [11:0] sel_182366;
  wire [10:0] add_182368;
  wire [11:0] sel_182370;
  wire [8:0] add_182372;
  wire [11:0] sel_182375;
  wire [8:0] add_182377;
  wire [11:0] sel_182380;
  wire [10:0] add_182382;
  wire [11:0] sel_182385;
  wire [10:0] add_182387;
  wire [11:0] sel_182390;
  wire [11:0] add_182415;
  wire [11:0] sel_182417;
  wire [11:0] add_182420;
  wire [11:0] sel_182422;
  wire [15:0] array_index_182451;
  wire [15:0] array_index_182454;
  wire [10:0] add_182458;
  wire [11:0] sel_182460;
  wire [10:0] add_182462;
  wire [11:0] sel_182464;
  wire [10:0] add_182466;
  wire [11:0] sel_182468;
  wire [10:0] add_182470;
  wire [11:0] sel_182472;
  wire [8:0] add_182474;
  wire [11:0] sel_182477;
  wire [8:0] add_182479;
  wire [11:0] sel_182482;
  wire [10:0] add_182484;
  wire [11:0] sel_182487;
  wire [10:0] add_182489;
  wire [11:0] sel_182492;
  wire [11:0] add_182517;
  wire [11:0] sel_182519;
  wire [11:0] add_182522;
  wire [11:0] sel_182524;
  wire [15:0] array_index_182553;
  wire [15:0] array_index_182556;
  wire [10:0] add_182560;
  wire [11:0] sel_182562;
  wire [10:0] add_182564;
  wire [11:0] sel_182566;
  wire [10:0] add_182568;
  wire [11:0] sel_182570;
  wire [10:0] add_182572;
  wire [11:0] sel_182574;
  wire [8:0] add_182576;
  wire [11:0] sel_182579;
  wire [8:0] add_182581;
  wire [11:0] sel_182584;
  wire [10:0] add_182586;
  wire [11:0] sel_182589;
  wire [10:0] add_182591;
  wire [11:0] sel_182594;
  wire [11:0] add_182619;
  wire [11:0] sel_182621;
  wire [11:0] add_182624;
  wire [11:0] sel_182626;
  wire [15:0] array_index_182655;
  wire [15:0] array_index_182658;
  wire [10:0] add_182662;
  wire [11:0] sel_182664;
  wire [10:0] add_182666;
  wire [11:0] sel_182668;
  wire [10:0] add_182670;
  wire [11:0] sel_182672;
  wire [10:0] add_182674;
  wire [11:0] sel_182676;
  wire [8:0] add_182678;
  wire [11:0] sel_182681;
  wire [8:0] add_182683;
  wire [11:0] sel_182686;
  wire [10:0] add_182688;
  wire [11:0] sel_182691;
  wire [10:0] add_182693;
  wire [11:0] sel_182696;
  wire [11:0] add_182721;
  wire [11:0] sel_182723;
  wire [11:0] add_182726;
  wire [11:0] sel_182728;
  wire [15:0] array_index_182757;
  wire [15:0] array_index_182760;
  wire [10:0] add_182764;
  wire [11:0] sel_182766;
  wire [10:0] add_182768;
  wire [11:0] sel_182770;
  wire [10:0] add_182772;
  wire [11:0] sel_182774;
  wire [10:0] add_182776;
  wire [11:0] sel_182778;
  wire [8:0] add_182780;
  wire [11:0] sel_182783;
  wire [8:0] add_182785;
  wire [11:0] sel_182788;
  wire [10:0] add_182790;
  wire [11:0] sel_182793;
  wire [10:0] add_182795;
  wire [11:0] sel_182798;
  wire [11:0] add_182822;
  wire [11:0] sel_182824;
  wire [11:0] add_182826;
  wire [11:0] sel_182828;
  wire [10:0] add_182862;
  wire [11:0] sel_182864;
  wire [10:0] add_182866;
  wire [11:0] sel_182868;
  wire [10:0] add_182870;
  wire [11:0] sel_182872;
  wire [10:0] add_182874;
  wire [11:0] sel_182876;
  wire [8:0] add_182878;
  wire [11:0] sel_182881;
  wire [8:0] add_182883;
  wire [11:0] sel_182886;
  wire [10:0] add_182888;
  wire [11:0] sel_182891;
  wire [10:0] add_182893;
  wire [11:0] sel_182896;
  wire [10:0] add_182944;
  wire [11:0] sel_182946;
  wire [10:0] add_182948;
  wire [11:0] sel_182950;
  wire [10:0] add_182952;
  wire [11:0] sel_182954;
  wire [10:0] add_182956;
  wire [11:0] sel_182958;
  wire [8:0] add_182960;
  wire [11:0] sel_182963;
  wire [8:0] add_182965;
  wire [11:0] sel_182968;
  wire [1:0] concat_182971;
  wire [1:0] add_182986;
  wire [10:0] add_183006;
  wire [11:0] sel_183008;
  wire [10:0] add_183010;
  wire [11:0] sel_183012;
  wire [10:0] add_183014;
  wire [11:0] sel_183016;
  wire [10:0] add_183018;
  wire [11:0] sel_183020;
  wire [2:0] concat_183023;
  wire [2:0] add_183034;
  wire [10:0] add_183048;
  wire [11:0] sel_183050;
  wire [10:0] add_183052;
  wire [11:0] sel_183054;
  wire [3:0] concat_183057;
  wire [3:0] add_183064;
  wire [4:0] concat_183073;
  wire [4:0] add_183076;
  assign array_index_172855 = set1_unflattened[7'h00];
  assign array_index_172856 = set2_unflattened[7'h00];
  assign add_172863 = array_index_172855[11:0] + 12'h247;
  assign add_172866 = array_index_172856[11:0] + 12'h247;
  assign array_index_172871 = set1_unflattened[7'h01];
  assign array_index_172874 = set2_unflattened[7'h01];
  assign add_172878 = array_index_172855[11:1] + 11'h247;
  assign add_172881 = array_index_172856[11:1] + 11'h247;
  assign add_172897 = array_index_172871[11:0] + 12'h247;
  assign sel_172899 = $signed({1'h0, add_172863}) < $signed(13'h0fff) ? add_172863 : 12'hfff;
  assign add_172902 = array_index_172874[11:0] + 12'h247;
  assign sel_172904 = $signed({1'h0, add_172866}) < $signed(13'h0fff) ? add_172866 : 12'hfff;
  assign array_index_172919 = set1_unflattened[7'h02];
  assign array_index_172922 = set2_unflattened[7'h02];
  assign add_172926 = array_index_172855[11:3] + 9'h0bd;
  assign add_172929 = array_index_172856[11:3] + 9'h0bd;
  assign add_172932 = array_index_172871[11:1] + 11'h247;
  assign sel_172935 = $signed({1'h0, add_172878, array_index_172855[0]}) < $signed(13'h0fff) ? {add_172878, array_index_172855[0]} : 12'hfff;
  assign add_172937 = array_index_172874[11:1] + 11'h247;
  assign sel_172940 = $signed({1'h0, add_172881, array_index_172856[0]}) < $signed(13'h0fff) ? {add_172881, array_index_172856[0]} : 12'hfff;
  assign add_172957 = array_index_172919[11:0] + 12'h247;
  assign sel_172959 = $signed({1'h0, add_172897}) < $signed({1'h0, sel_172899}) ? add_172897 : sel_172899;
  assign add_172962 = array_index_172922[11:0] + 12'h247;
  assign sel_172964 = $signed({1'h0, add_172902}) < $signed({1'h0, sel_172904}) ? add_172902 : sel_172904;
  assign array_index_172985 = set1_unflattened[7'h03];
  assign array_index_172988 = set2_unflattened[7'h03];
  assign add_172992 = array_index_172855[11:1] + 11'h347;
  assign add_172994 = array_index_172856[11:1] + 11'h347;
  assign add_172996 = array_index_172871[11:3] + 9'h0bd;
  assign sel_172999 = $signed({1'h0, add_172926, array_index_172855[2:0]}) < $signed(13'h0fff) ? {add_172926, array_index_172855[2:0]} : 12'hfff;
  assign add_173001 = array_index_172874[11:3] + 9'h0bd;
  assign sel_173004 = $signed({1'h0, add_172929, array_index_172856[2:0]}) < $signed(13'h0fff) ? {add_172929, array_index_172856[2:0]} : 12'hfff;
  assign add_173006 = array_index_172919[11:1] + 11'h247;
  assign sel_173009 = $signed({1'h0, add_172932, array_index_172871[0]}) < $signed({1'h0, sel_172935}) ? {add_172932, array_index_172871[0]} : sel_172935;
  assign add_173011 = array_index_172922[11:1] + 11'h247;
  assign sel_173014 = $signed({1'h0, add_172937, array_index_172874[0]}) < $signed({1'h0, sel_172940}) ? {add_172937, array_index_172874[0]} : sel_172940;
  assign add_173035 = array_index_172985[11:0] + 12'h247;
  assign sel_173037 = $signed({1'h0, add_172957}) < $signed({1'h0, sel_172959}) ? add_172957 : sel_172959;
  assign add_173040 = array_index_172988[11:0] + 12'h247;
  assign sel_173042 = $signed({1'h0, add_172962}) < $signed({1'h0, sel_172964}) ? add_172962 : sel_172964;
  assign array_index_173069 = set1_unflattened[7'h04];
  assign array_index_173072 = set2_unflattened[7'h04];
  assign add_173076 = array_index_172855[11:1] + 11'h79d;
  assign add_173078 = array_index_172856[11:1] + 11'h79d;
  assign add_173080 = array_index_172871[11:1] + 11'h347;
  assign sel_173082 = $signed({1'h0, add_172992, array_index_172855[0]}) < $signed(13'h0fff) ? {add_172992, array_index_172855[0]} : 12'hfff;
  assign add_173084 = array_index_172874[11:1] + 11'h347;
  assign sel_173086 = $signed({1'h0, add_172994, array_index_172856[0]}) < $signed(13'h0fff) ? {add_172994, array_index_172856[0]} : 12'hfff;
  assign add_173088 = array_index_172919[11:3] + 9'h0bd;
  assign sel_173091 = $signed({1'h0, add_172996, array_index_172871[2:0]}) < $signed({1'h0, sel_172999}) ? {add_172996, array_index_172871[2:0]} : sel_172999;
  assign add_173093 = array_index_172922[11:3] + 9'h0bd;
  assign sel_173096 = $signed({1'h0, add_173001, array_index_172874[2:0]}) < $signed({1'h0, sel_173004}) ? {add_173001, array_index_172874[2:0]} : sel_173004;
  assign add_173098 = array_index_172985[11:1] + 11'h247;
  assign sel_173101 = $signed({1'h0, add_173006, array_index_172919[0]}) < $signed({1'h0, sel_173009}) ? {add_173006, array_index_172919[0]} : sel_173009;
  assign add_173103 = array_index_172988[11:1] + 11'h247;
  assign sel_173106 = $signed({1'h0, add_173011, array_index_172922[0]}) < $signed({1'h0, sel_173014}) ? {add_173011, array_index_172922[0]} : sel_173014;
  assign add_173131 = array_index_173069[11:0] + 12'h247;
  assign sel_173133 = $signed({1'h0, add_173035}) < $signed({1'h0, sel_173037}) ? add_173035 : sel_173037;
  assign add_173136 = array_index_173072[11:0] + 12'h247;
  assign sel_173138 = $signed({1'h0, add_173040}) < $signed({1'h0, sel_173042}) ? add_173040 : sel_173042;
  assign array_index_173169 = set1_unflattened[7'h05];
  assign array_index_173172 = set2_unflattened[7'h05];
  assign add_173176 = array_index_172871[11:1] + 11'h79d;
  assign sel_173178 = $signed({1'h0, add_173076, array_index_172855[0]}) < $signed(13'h0fff) ? {add_173076, array_index_172855[0]} : 12'hfff;
  assign add_173180 = array_index_172874[11:1] + 11'h79d;
  assign sel_173182 = $signed({1'h0, add_173078, array_index_172856[0]}) < $signed(13'h0fff) ? {add_173078, array_index_172856[0]} : 12'hfff;
  assign add_173184 = array_index_172919[11:1] + 11'h347;
  assign sel_173186 = $signed({1'h0, add_173080, array_index_172871[0]}) < $signed({1'h0, sel_173082}) ? {add_173080, array_index_172871[0]} : sel_173082;
  assign add_173188 = array_index_172922[11:1] + 11'h347;
  assign sel_173190 = $signed({1'h0, add_173084, array_index_172874[0]}) < $signed({1'h0, sel_173086}) ? {add_173084, array_index_172874[0]} : sel_173086;
  assign add_173192 = array_index_172985[11:3] + 9'h0bd;
  assign sel_173195 = $signed({1'h0, add_173088, array_index_172919[2:0]}) < $signed({1'h0, sel_173091}) ? {add_173088, array_index_172919[2:0]} : sel_173091;
  assign add_173197 = array_index_172988[11:3] + 9'h0bd;
  assign sel_173200 = $signed({1'h0, add_173093, array_index_172922[2:0]}) < $signed({1'h0, sel_173096}) ? {add_173093, array_index_172922[2:0]} : sel_173096;
  assign add_173202 = array_index_173069[11:1] + 11'h247;
  assign sel_173205 = $signed({1'h0, add_173098, array_index_172985[0]}) < $signed({1'h0, sel_173101}) ? {add_173098, array_index_172985[0]} : sel_173101;
  assign add_173207 = array_index_173072[11:1] + 11'h247;
  assign sel_173210 = $signed({1'h0, add_173103, array_index_172988[0]}) < $signed({1'h0, sel_173106}) ? {add_173103, array_index_172988[0]} : sel_173106;
  assign add_173235 = array_index_173169[11:0] + 12'h247;
  assign sel_173237 = $signed({1'h0, add_173131}) < $signed({1'h0, sel_173133}) ? add_173131 : sel_173133;
  assign add_173240 = array_index_173172[11:0] + 12'h247;
  assign sel_173242 = $signed({1'h0, add_173136}) < $signed({1'h0, sel_173138}) ? add_173136 : sel_173138;
  assign array_index_173271 = set1_unflattened[7'h06];
  assign array_index_173274 = set2_unflattened[7'h06];
  assign add_173278 = array_index_172919[11:1] + 11'h79d;
  assign sel_173280 = $signed({1'h0, add_173176, array_index_172871[0]}) < $signed({1'h0, sel_173178}) ? {add_173176, array_index_172871[0]} : sel_173178;
  assign add_173282 = array_index_172922[11:1] + 11'h79d;
  assign sel_173284 = $signed({1'h0, add_173180, array_index_172874[0]}) < $signed({1'h0, sel_173182}) ? {add_173180, array_index_172874[0]} : sel_173182;
  assign add_173286 = array_index_172985[11:1] + 11'h347;
  assign sel_173288 = $signed({1'h0, add_173184, array_index_172919[0]}) < $signed({1'h0, sel_173186}) ? {add_173184, array_index_172919[0]} : sel_173186;
  assign add_173290 = array_index_172988[11:1] + 11'h347;
  assign sel_173292 = $signed({1'h0, add_173188, array_index_172922[0]}) < $signed({1'h0, sel_173190}) ? {add_173188, array_index_172922[0]} : sel_173190;
  assign add_173294 = array_index_173069[11:3] + 9'h0bd;
  assign sel_173297 = $signed({1'h0, add_173192, array_index_172985[2:0]}) < $signed({1'h0, sel_173195}) ? {add_173192, array_index_172985[2:0]} : sel_173195;
  assign add_173299 = array_index_173072[11:3] + 9'h0bd;
  assign sel_173302 = $signed({1'h0, add_173197, array_index_172988[2:0]}) < $signed({1'h0, sel_173200}) ? {add_173197, array_index_172988[2:0]} : sel_173200;
  assign add_173304 = array_index_173169[11:1] + 11'h247;
  assign sel_173307 = $signed({1'h0, add_173202, array_index_173069[0]}) < $signed({1'h0, sel_173205}) ? {add_173202, array_index_173069[0]} : sel_173205;
  assign add_173309 = array_index_173172[11:1] + 11'h247;
  assign sel_173312 = $signed({1'h0, add_173207, array_index_173072[0]}) < $signed({1'h0, sel_173210}) ? {add_173207, array_index_173072[0]} : sel_173210;
  assign add_173337 = array_index_173271[11:0] + 12'h247;
  assign sel_173339 = $signed({1'h0, add_173235}) < $signed({1'h0, sel_173237}) ? add_173235 : sel_173237;
  assign add_173342 = array_index_173274[11:0] + 12'h247;
  assign sel_173344 = $signed({1'h0, add_173240}) < $signed({1'h0, sel_173242}) ? add_173240 : sel_173242;
  assign array_index_173373 = set1_unflattened[7'h07];
  assign array_index_173376 = set2_unflattened[7'h07];
  assign add_173380 = array_index_172985[11:1] + 11'h79d;
  assign sel_173382 = $signed({1'h0, add_173278, array_index_172919[0]}) < $signed({1'h0, sel_173280}) ? {add_173278, array_index_172919[0]} : sel_173280;
  assign add_173384 = array_index_172988[11:1] + 11'h79d;
  assign sel_173386 = $signed({1'h0, add_173282, array_index_172922[0]}) < $signed({1'h0, sel_173284}) ? {add_173282, array_index_172922[0]} : sel_173284;
  assign add_173388 = array_index_173069[11:1] + 11'h347;
  assign sel_173390 = $signed({1'h0, add_173286, array_index_172985[0]}) < $signed({1'h0, sel_173288}) ? {add_173286, array_index_172985[0]} : sel_173288;
  assign add_173392 = array_index_173072[11:1] + 11'h347;
  assign sel_173394 = $signed({1'h0, add_173290, array_index_172988[0]}) < $signed({1'h0, sel_173292}) ? {add_173290, array_index_172988[0]} : sel_173292;
  assign add_173396 = array_index_173169[11:3] + 9'h0bd;
  assign sel_173399 = $signed({1'h0, add_173294, array_index_173069[2:0]}) < $signed({1'h0, sel_173297}) ? {add_173294, array_index_173069[2:0]} : sel_173297;
  assign add_173401 = array_index_173172[11:3] + 9'h0bd;
  assign sel_173404 = $signed({1'h0, add_173299, array_index_173072[2:0]}) < $signed({1'h0, sel_173302}) ? {add_173299, array_index_173072[2:0]} : sel_173302;
  assign add_173406 = array_index_173271[11:1] + 11'h247;
  assign sel_173409 = $signed({1'h0, add_173304, array_index_173169[0]}) < $signed({1'h0, sel_173307}) ? {add_173304, array_index_173169[0]} : sel_173307;
  assign add_173411 = array_index_173274[11:1] + 11'h247;
  assign sel_173414 = $signed({1'h0, add_173309, array_index_173172[0]}) < $signed({1'h0, sel_173312}) ? {add_173309, array_index_173172[0]} : sel_173312;
  assign add_173439 = array_index_173373[11:0] + 12'h247;
  assign sel_173441 = $signed({1'h0, add_173337}) < $signed({1'h0, sel_173339}) ? add_173337 : sel_173339;
  assign add_173444 = array_index_173376[11:0] + 12'h247;
  assign sel_173446 = $signed({1'h0, add_173342}) < $signed({1'h0, sel_173344}) ? add_173342 : sel_173344;
  assign array_index_173475 = set1_unflattened[7'h08];
  assign array_index_173478 = set2_unflattened[7'h08];
  assign add_173482 = array_index_173069[11:1] + 11'h79d;
  assign sel_173484 = $signed({1'h0, add_173380, array_index_172985[0]}) < $signed({1'h0, sel_173382}) ? {add_173380, array_index_172985[0]} : sel_173382;
  assign add_173486 = array_index_173072[11:1] + 11'h79d;
  assign sel_173488 = $signed({1'h0, add_173384, array_index_172988[0]}) < $signed({1'h0, sel_173386}) ? {add_173384, array_index_172988[0]} : sel_173386;
  assign add_173490 = array_index_173169[11:1] + 11'h347;
  assign sel_173492 = $signed({1'h0, add_173388, array_index_173069[0]}) < $signed({1'h0, sel_173390}) ? {add_173388, array_index_173069[0]} : sel_173390;
  assign add_173494 = array_index_173172[11:1] + 11'h347;
  assign sel_173496 = $signed({1'h0, add_173392, array_index_173072[0]}) < $signed({1'h0, sel_173394}) ? {add_173392, array_index_173072[0]} : sel_173394;
  assign add_173498 = array_index_173271[11:3] + 9'h0bd;
  assign sel_173501 = $signed({1'h0, add_173396, array_index_173169[2:0]}) < $signed({1'h0, sel_173399}) ? {add_173396, array_index_173169[2:0]} : sel_173399;
  assign add_173503 = array_index_173274[11:3] + 9'h0bd;
  assign sel_173506 = $signed({1'h0, add_173401, array_index_173172[2:0]}) < $signed({1'h0, sel_173404}) ? {add_173401, array_index_173172[2:0]} : sel_173404;
  assign add_173508 = array_index_173373[11:1] + 11'h247;
  assign sel_173511 = $signed({1'h0, add_173406, array_index_173271[0]}) < $signed({1'h0, sel_173409}) ? {add_173406, array_index_173271[0]} : sel_173409;
  assign add_173513 = array_index_173376[11:1] + 11'h247;
  assign sel_173516 = $signed({1'h0, add_173411, array_index_173274[0]}) < $signed({1'h0, sel_173414}) ? {add_173411, array_index_173274[0]} : sel_173414;
  assign add_173541 = array_index_173475[11:0] + 12'h247;
  assign sel_173543 = $signed({1'h0, add_173439}) < $signed({1'h0, sel_173441}) ? add_173439 : sel_173441;
  assign add_173546 = array_index_173478[11:0] + 12'h247;
  assign sel_173548 = $signed({1'h0, add_173444}) < $signed({1'h0, sel_173446}) ? add_173444 : sel_173446;
  assign array_index_173577 = set1_unflattened[7'h09];
  assign array_index_173580 = set2_unflattened[7'h09];
  assign add_173584 = array_index_173169[11:1] + 11'h79d;
  assign sel_173586 = $signed({1'h0, add_173482, array_index_173069[0]}) < $signed({1'h0, sel_173484}) ? {add_173482, array_index_173069[0]} : sel_173484;
  assign add_173588 = array_index_173172[11:1] + 11'h79d;
  assign sel_173590 = $signed({1'h0, add_173486, array_index_173072[0]}) < $signed({1'h0, sel_173488}) ? {add_173486, array_index_173072[0]} : sel_173488;
  assign add_173592 = array_index_173271[11:1] + 11'h347;
  assign sel_173594 = $signed({1'h0, add_173490, array_index_173169[0]}) < $signed({1'h0, sel_173492}) ? {add_173490, array_index_173169[0]} : sel_173492;
  assign add_173596 = array_index_173274[11:1] + 11'h347;
  assign sel_173598 = $signed({1'h0, add_173494, array_index_173172[0]}) < $signed({1'h0, sel_173496}) ? {add_173494, array_index_173172[0]} : sel_173496;
  assign add_173600 = array_index_173373[11:3] + 9'h0bd;
  assign sel_173603 = $signed({1'h0, add_173498, array_index_173271[2:0]}) < $signed({1'h0, sel_173501}) ? {add_173498, array_index_173271[2:0]} : sel_173501;
  assign add_173605 = array_index_173376[11:3] + 9'h0bd;
  assign sel_173608 = $signed({1'h0, add_173503, array_index_173274[2:0]}) < $signed({1'h0, sel_173506}) ? {add_173503, array_index_173274[2:0]} : sel_173506;
  assign add_173610 = array_index_173475[11:1] + 11'h247;
  assign sel_173613 = $signed({1'h0, add_173508, array_index_173373[0]}) < $signed({1'h0, sel_173511}) ? {add_173508, array_index_173373[0]} : sel_173511;
  assign add_173615 = array_index_173478[11:1] + 11'h247;
  assign sel_173618 = $signed({1'h0, add_173513, array_index_173376[0]}) < $signed({1'h0, sel_173516}) ? {add_173513, array_index_173376[0]} : sel_173516;
  assign add_173643 = array_index_173577[11:0] + 12'h247;
  assign sel_173645 = $signed({1'h0, add_173541}) < $signed({1'h0, sel_173543}) ? add_173541 : sel_173543;
  assign add_173648 = array_index_173580[11:0] + 12'h247;
  assign sel_173650 = $signed({1'h0, add_173546}) < $signed({1'h0, sel_173548}) ? add_173546 : sel_173548;
  assign array_index_173679 = set1_unflattened[7'h0a];
  assign array_index_173682 = set2_unflattened[7'h0a];
  assign add_173686 = array_index_173271[11:1] + 11'h79d;
  assign sel_173688 = $signed({1'h0, add_173584, array_index_173169[0]}) < $signed({1'h0, sel_173586}) ? {add_173584, array_index_173169[0]} : sel_173586;
  assign add_173690 = array_index_173274[11:1] + 11'h79d;
  assign sel_173692 = $signed({1'h0, add_173588, array_index_173172[0]}) < $signed({1'h0, sel_173590}) ? {add_173588, array_index_173172[0]} : sel_173590;
  assign add_173694 = array_index_173373[11:1] + 11'h347;
  assign sel_173696 = $signed({1'h0, add_173592, array_index_173271[0]}) < $signed({1'h0, sel_173594}) ? {add_173592, array_index_173271[0]} : sel_173594;
  assign add_173698 = array_index_173376[11:1] + 11'h347;
  assign sel_173700 = $signed({1'h0, add_173596, array_index_173274[0]}) < $signed({1'h0, sel_173598}) ? {add_173596, array_index_173274[0]} : sel_173598;
  assign add_173702 = array_index_173475[11:3] + 9'h0bd;
  assign sel_173705 = $signed({1'h0, add_173600, array_index_173373[2:0]}) < $signed({1'h0, sel_173603}) ? {add_173600, array_index_173373[2:0]} : sel_173603;
  assign add_173707 = array_index_173478[11:3] + 9'h0bd;
  assign sel_173710 = $signed({1'h0, add_173605, array_index_173376[2:0]}) < $signed({1'h0, sel_173608}) ? {add_173605, array_index_173376[2:0]} : sel_173608;
  assign add_173712 = array_index_173577[11:1] + 11'h247;
  assign sel_173715 = $signed({1'h0, add_173610, array_index_173475[0]}) < $signed({1'h0, sel_173613}) ? {add_173610, array_index_173475[0]} : sel_173613;
  assign add_173717 = array_index_173580[11:1] + 11'h247;
  assign sel_173720 = $signed({1'h0, add_173615, array_index_173478[0]}) < $signed({1'h0, sel_173618}) ? {add_173615, array_index_173478[0]} : sel_173618;
  assign add_173745 = array_index_173679[11:0] + 12'h247;
  assign sel_173747 = $signed({1'h0, add_173643}) < $signed({1'h0, sel_173645}) ? add_173643 : sel_173645;
  assign add_173750 = array_index_173682[11:0] + 12'h247;
  assign sel_173752 = $signed({1'h0, add_173648}) < $signed({1'h0, sel_173650}) ? add_173648 : sel_173650;
  assign array_index_173781 = set1_unflattened[7'h0b];
  assign array_index_173784 = set2_unflattened[7'h0b];
  assign add_173788 = array_index_173373[11:1] + 11'h79d;
  assign sel_173790 = $signed({1'h0, add_173686, array_index_173271[0]}) < $signed({1'h0, sel_173688}) ? {add_173686, array_index_173271[0]} : sel_173688;
  assign add_173792 = array_index_173376[11:1] + 11'h79d;
  assign sel_173794 = $signed({1'h0, add_173690, array_index_173274[0]}) < $signed({1'h0, sel_173692}) ? {add_173690, array_index_173274[0]} : sel_173692;
  assign add_173796 = array_index_173475[11:1] + 11'h347;
  assign sel_173798 = $signed({1'h0, add_173694, array_index_173373[0]}) < $signed({1'h0, sel_173696}) ? {add_173694, array_index_173373[0]} : sel_173696;
  assign add_173800 = array_index_173478[11:1] + 11'h347;
  assign sel_173802 = $signed({1'h0, add_173698, array_index_173376[0]}) < $signed({1'h0, sel_173700}) ? {add_173698, array_index_173376[0]} : sel_173700;
  assign add_173804 = array_index_173577[11:3] + 9'h0bd;
  assign sel_173807 = $signed({1'h0, add_173702, array_index_173475[2:0]}) < $signed({1'h0, sel_173705}) ? {add_173702, array_index_173475[2:0]} : sel_173705;
  assign add_173809 = array_index_173580[11:3] + 9'h0bd;
  assign sel_173812 = $signed({1'h0, add_173707, array_index_173478[2:0]}) < $signed({1'h0, sel_173710}) ? {add_173707, array_index_173478[2:0]} : sel_173710;
  assign add_173814 = array_index_173679[11:1] + 11'h247;
  assign sel_173817 = $signed({1'h0, add_173712, array_index_173577[0]}) < $signed({1'h0, sel_173715}) ? {add_173712, array_index_173577[0]} : sel_173715;
  assign add_173819 = array_index_173682[11:1] + 11'h247;
  assign sel_173822 = $signed({1'h0, add_173717, array_index_173580[0]}) < $signed({1'h0, sel_173720}) ? {add_173717, array_index_173580[0]} : sel_173720;
  assign add_173847 = array_index_173781[11:0] + 12'h247;
  assign sel_173849 = $signed({1'h0, add_173745}) < $signed({1'h0, sel_173747}) ? add_173745 : sel_173747;
  assign add_173852 = array_index_173784[11:0] + 12'h247;
  assign sel_173854 = $signed({1'h0, add_173750}) < $signed({1'h0, sel_173752}) ? add_173750 : sel_173752;
  assign array_index_173883 = set1_unflattened[7'h0c];
  assign array_index_173886 = set2_unflattened[7'h0c];
  assign add_173890 = array_index_173475[11:1] + 11'h79d;
  assign sel_173892 = $signed({1'h0, add_173788, array_index_173373[0]}) < $signed({1'h0, sel_173790}) ? {add_173788, array_index_173373[0]} : sel_173790;
  assign add_173894 = array_index_173478[11:1] + 11'h79d;
  assign sel_173896 = $signed({1'h0, add_173792, array_index_173376[0]}) < $signed({1'h0, sel_173794}) ? {add_173792, array_index_173376[0]} : sel_173794;
  assign add_173898 = array_index_173577[11:1] + 11'h347;
  assign sel_173900 = $signed({1'h0, add_173796, array_index_173475[0]}) < $signed({1'h0, sel_173798}) ? {add_173796, array_index_173475[0]} : sel_173798;
  assign add_173902 = array_index_173580[11:1] + 11'h347;
  assign sel_173904 = $signed({1'h0, add_173800, array_index_173478[0]}) < $signed({1'h0, sel_173802}) ? {add_173800, array_index_173478[0]} : sel_173802;
  assign add_173906 = array_index_173679[11:3] + 9'h0bd;
  assign sel_173909 = $signed({1'h0, add_173804, array_index_173577[2:0]}) < $signed({1'h0, sel_173807}) ? {add_173804, array_index_173577[2:0]} : sel_173807;
  assign add_173911 = array_index_173682[11:3] + 9'h0bd;
  assign sel_173914 = $signed({1'h0, add_173809, array_index_173580[2:0]}) < $signed({1'h0, sel_173812}) ? {add_173809, array_index_173580[2:0]} : sel_173812;
  assign add_173916 = array_index_173781[11:1] + 11'h247;
  assign sel_173919 = $signed({1'h0, add_173814, array_index_173679[0]}) < $signed({1'h0, sel_173817}) ? {add_173814, array_index_173679[0]} : sel_173817;
  assign add_173921 = array_index_173784[11:1] + 11'h247;
  assign sel_173924 = $signed({1'h0, add_173819, array_index_173682[0]}) < $signed({1'h0, sel_173822}) ? {add_173819, array_index_173682[0]} : sel_173822;
  assign add_173949 = array_index_173883[11:0] + 12'h247;
  assign sel_173951 = $signed({1'h0, add_173847}) < $signed({1'h0, sel_173849}) ? add_173847 : sel_173849;
  assign add_173954 = array_index_173886[11:0] + 12'h247;
  assign sel_173956 = $signed({1'h0, add_173852}) < $signed({1'h0, sel_173854}) ? add_173852 : sel_173854;
  assign array_index_173985 = set1_unflattened[7'h0d];
  assign array_index_173988 = set2_unflattened[7'h0d];
  assign add_173992 = array_index_173577[11:1] + 11'h79d;
  assign sel_173994 = $signed({1'h0, add_173890, array_index_173475[0]}) < $signed({1'h0, sel_173892}) ? {add_173890, array_index_173475[0]} : sel_173892;
  assign add_173996 = array_index_173580[11:1] + 11'h79d;
  assign sel_173998 = $signed({1'h0, add_173894, array_index_173478[0]}) < $signed({1'h0, sel_173896}) ? {add_173894, array_index_173478[0]} : sel_173896;
  assign add_174000 = array_index_173679[11:1] + 11'h347;
  assign sel_174002 = $signed({1'h0, add_173898, array_index_173577[0]}) < $signed({1'h0, sel_173900}) ? {add_173898, array_index_173577[0]} : sel_173900;
  assign add_174004 = array_index_173682[11:1] + 11'h347;
  assign sel_174006 = $signed({1'h0, add_173902, array_index_173580[0]}) < $signed({1'h0, sel_173904}) ? {add_173902, array_index_173580[0]} : sel_173904;
  assign add_174008 = array_index_173781[11:3] + 9'h0bd;
  assign sel_174011 = $signed({1'h0, add_173906, array_index_173679[2:0]}) < $signed({1'h0, sel_173909}) ? {add_173906, array_index_173679[2:0]} : sel_173909;
  assign add_174013 = array_index_173784[11:3] + 9'h0bd;
  assign sel_174016 = $signed({1'h0, add_173911, array_index_173682[2:0]}) < $signed({1'h0, sel_173914}) ? {add_173911, array_index_173682[2:0]} : sel_173914;
  assign add_174018 = array_index_173883[11:1] + 11'h247;
  assign sel_174021 = $signed({1'h0, add_173916, array_index_173781[0]}) < $signed({1'h0, sel_173919}) ? {add_173916, array_index_173781[0]} : sel_173919;
  assign add_174023 = array_index_173886[11:1] + 11'h247;
  assign sel_174026 = $signed({1'h0, add_173921, array_index_173784[0]}) < $signed({1'h0, sel_173924}) ? {add_173921, array_index_173784[0]} : sel_173924;
  assign add_174051 = array_index_173985[11:0] + 12'h247;
  assign sel_174053 = $signed({1'h0, add_173949}) < $signed({1'h0, sel_173951}) ? add_173949 : sel_173951;
  assign add_174056 = array_index_173988[11:0] + 12'h247;
  assign sel_174058 = $signed({1'h0, add_173954}) < $signed({1'h0, sel_173956}) ? add_173954 : sel_173956;
  assign array_index_174087 = set1_unflattened[7'h0e];
  assign array_index_174090 = set2_unflattened[7'h0e];
  assign add_174094 = array_index_173679[11:1] + 11'h79d;
  assign sel_174096 = $signed({1'h0, add_173992, array_index_173577[0]}) < $signed({1'h0, sel_173994}) ? {add_173992, array_index_173577[0]} : sel_173994;
  assign add_174098 = array_index_173682[11:1] + 11'h79d;
  assign sel_174100 = $signed({1'h0, add_173996, array_index_173580[0]}) < $signed({1'h0, sel_173998}) ? {add_173996, array_index_173580[0]} : sel_173998;
  assign add_174102 = array_index_173781[11:1] + 11'h347;
  assign sel_174104 = $signed({1'h0, add_174000, array_index_173679[0]}) < $signed({1'h0, sel_174002}) ? {add_174000, array_index_173679[0]} : sel_174002;
  assign add_174106 = array_index_173784[11:1] + 11'h347;
  assign sel_174108 = $signed({1'h0, add_174004, array_index_173682[0]}) < $signed({1'h0, sel_174006}) ? {add_174004, array_index_173682[0]} : sel_174006;
  assign add_174110 = array_index_173883[11:3] + 9'h0bd;
  assign sel_174113 = $signed({1'h0, add_174008, array_index_173781[2:0]}) < $signed({1'h0, sel_174011}) ? {add_174008, array_index_173781[2:0]} : sel_174011;
  assign add_174115 = array_index_173886[11:3] + 9'h0bd;
  assign sel_174118 = $signed({1'h0, add_174013, array_index_173784[2:0]}) < $signed({1'h0, sel_174016}) ? {add_174013, array_index_173784[2:0]} : sel_174016;
  assign add_174120 = array_index_173985[11:1] + 11'h247;
  assign sel_174123 = $signed({1'h0, add_174018, array_index_173883[0]}) < $signed({1'h0, sel_174021}) ? {add_174018, array_index_173883[0]} : sel_174021;
  assign add_174125 = array_index_173988[11:1] + 11'h247;
  assign sel_174128 = $signed({1'h0, add_174023, array_index_173886[0]}) < $signed({1'h0, sel_174026}) ? {add_174023, array_index_173886[0]} : sel_174026;
  assign add_174153 = array_index_174087[11:0] + 12'h247;
  assign sel_174155 = $signed({1'h0, add_174051}) < $signed({1'h0, sel_174053}) ? add_174051 : sel_174053;
  assign add_174158 = array_index_174090[11:0] + 12'h247;
  assign sel_174160 = $signed({1'h0, add_174056}) < $signed({1'h0, sel_174058}) ? add_174056 : sel_174058;
  assign array_index_174189 = set1_unflattened[7'h0f];
  assign array_index_174192 = set2_unflattened[7'h0f];
  assign add_174196 = array_index_173781[11:1] + 11'h79d;
  assign sel_174198 = $signed({1'h0, add_174094, array_index_173679[0]}) < $signed({1'h0, sel_174096}) ? {add_174094, array_index_173679[0]} : sel_174096;
  assign add_174200 = array_index_173784[11:1] + 11'h79d;
  assign sel_174202 = $signed({1'h0, add_174098, array_index_173682[0]}) < $signed({1'h0, sel_174100}) ? {add_174098, array_index_173682[0]} : sel_174100;
  assign add_174204 = array_index_173883[11:1] + 11'h347;
  assign sel_174206 = $signed({1'h0, add_174102, array_index_173781[0]}) < $signed({1'h0, sel_174104}) ? {add_174102, array_index_173781[0]} : sel_174104;
  assign add_174208 = array_index_173886[11:1] + 11'h347;
  assign sel_174210 = $signed({1'h0, add_174106, array_index_173784[0]}) < $signed({1'h0, sel_174108}) ? {add_174106, array_index_173784[0]} : sel_174108;
  assign add_174212 = array_index_173985[11:3] + 9'h0bd;
  assign sel_174215 = $signed({1'h0, add_174110, array_index_173883[2:0]}) < $signed({1'h0, sel_174113}) ? {add_174110, array_index_173883[2:0]} : sel_174113;
  assign add_174217 = array_index_173988[11:3] + 9'h0bd;
  assign sel_174220 = $signed({1'h0, add_174115, array_index_173886[2:0]}) < $signed({1'h0, sel_174118}) ? {add_174115, array_index_173886[2:0]} : sel_174118;
  assign add_174222 = array_index_174087[11:1] + 11'h247;
  assign sel_174225 = $signed({1'h0, add_174120, array_index_173985[0]}) < $signed({1'h0, sel_174123}) ? {add_174120, array_index_173985[0]} : sel_174123;
  assign add_174227 = array_index_174090[11:1] + 11'h247;
  assign sel_174230 = $signed({1'h0, add_174125, array_index_173988[0]}) < $signed({1'h0, sel_174128}) ? {add_174125, array_index_173988[0]} : sel_174128;
  assign add_174255 = array_index_174189[11:0] + 12'h247;
  assign sel_174257 = $signed({1'h0, add_174153}) < $signed({1'h0, sel_174155}) ? add_174153 : sel_174155;
  assign add_174260 = array_index_174192[11:0] + 12'h247;
  assign sel_174262 = $signed({1'h0, add_174158}) < $signed({1'h0, sel_174160}) ? add_174158 : sel_174160;
  assign array_index_174291 = set1_unflattened[7'h10];
  assign array_index_174294 = set2_unflattened[7'h10];
  assign add_174298 = array_index_173883[11:1] + 11'h79d;
  assign sel_174300 = $signed({1'h0, add_174196, array_index_173781[0]}) < $signed({1'h0, sel_174198}) ? {add_174196, array_index_173781[0]} : sel_174198;
  assign add_174302 = array_index_173886[11:1] + 11'h79d;
  assign sel_174304 = $signed({1'h0, add_174200, array_index_173784[0]}) < $signed({1'h0, sel_174202}) ? {add_174200, array_index_173784[0]} : sel_174202;
  assign add_174306 = array_index_173985[11:1] + 11'h347;
  assign sel_174308 = $signed({1'h0, add_174204, array_index_173883[0]}) < $signed({1'h0, sel_174206}) ? {add_174204, array_index_173883[0]} : sel_174206;
  assign add_174310 = array_index_173988[11:1] + 11'h347;
  assign sel_174312 = $signed({1'h0, add_174208, array_index_173886[0]}) < $signed({1'h0, sel_174210}) ? {add_174208, array_index_173886[0]} : sel_174210;
  assign add_174314 = array_index_174087[11:3] + 9'h0bd;
  assign sel_174317 = $signed({1'h0, add_174212, array_index_173985[2:0]}) < $signed({1'h0, sel_174215}) ? {add_174212, array_index_173985[2:0]} : sel_174215;
  assign add_174319 = array_index_174090[11:3] + 9'h0bd;
  assign sel_174322 = $signed({1'h0, add_174217, array_index_173988[2:0]}) < $signed({1'h0, sel_174220}) ? {add_174217, array_index_173988[2:0]} : sel_174220;
  assign add_174324 = array_index_174189[11:1] + 11'h247;
  assign sel_174327 = $signed({1'h0, add_174222, array_index_174087[0]}) < $signed({1'h0, sel_174225}) ? {add_174222, array_index_174087[0]} : sel_174225;
  assign add_174329 = array_index_174192[11:1] + 11'h247;
  assign sel_174332 = $signed({1'h0, add_174227, array_index_174090[0]}) < $signed({1'h0, sel_174230}) ? {add_174227, array_index_174090[0]} : sel_174230;
  assign add_174357 = array_index_174291[11:0] + 12'h247;
  assign sel_174359 = $signed({1'h0, add_174255}) < $signed({1'h0, sel_174257}) ? add_174255 : sel_174257;
  assign add_174362 = array_index_174294[11:0] + 12'h247;
  assign sel_174364 = $signed({1'h0, add_174260}) < $signed({1'h0, sel_174262}) ? add_174260 : sel_174262;
  assign array_index_174393 = set1_unflattened[7'h11];
  assign array_index_174396 = set2_unflattened[7'h11];
  assign add_174400 = array_index_173985[11:1] + 11'h79d;
  assign sel_174402 = $signed({1'h0, add_174298, array_index_173883[0]}) < $signed({1'h0, sel_174300}) ? {add_174298, array_index_173883[0]} : sel_174300;
  assign add_174404 = array_index_173988[11:1] + 11'h79d;
  assign sel_174406 = $signed({1'h0, add_174302, array_index_173886[0]}) < $signed({1'h0, sel_174304}) ? {add_174302, array_index_173886[0]} : sel_174304;
  assign add_174408 = array_index_174087[11:1] + 11'h347;
  assign sel_174410 = $signed({1'h0, add_174306, array_index_173985[0]}) < $signed({1'h0, sel_174308}) ? {add_174306, array_index_173985[0]} : sel_174308;
  assign add_174412 = array_index_174090[11:1] + 11'h347;
  assign sel_174414 = $signed({1'h0, add_174310, array_index_173988[0]}) < $signed({1'h0, sel_174312}) ? {add_174310, array_index_173988[0]} : sel_174312;
  assign add_174416 = array_index_174189[11:3] + 9'h0bd;
  assign sel_174419 = $signed({1'h0, add_174314, array_index_174087[2:0]}) < $signed({1'h0, sel_174317}) ? {add_174314, array_index_174087[2:0]} : sel_174317;
  assign add_174421 = array_index_174192[11:3] + 9'h0bd;
  assign sel_174424 = $signed({1'h0, add_174319, array_index_174090[2:0]}) < $signed({1'h0, sel_174322}) ? {add_174319, array_index_174090[2:0]} : sel_174322;
  assign add_174426 = array_index_174291[11:1] + 11'h247;
  assign sel_174429 = $signed({1'h0, add_174324, array_index_174189[0]}) < $signed({1'h0, sel_174327}) ? {add_174324, array_index_174189[0]} : sel_174327;
  assign add_174431 = array_index_174294[11:1] + 11'h247;
  assign sel_174434 = $signed({1'h0, add_174329, array_index_174192[0]}) < $signed({1'h0, sel_174332}) ? {add_174329, array_index_174192[0]} : sel_174332;
  assign add_174459 = array_index_174393[11:0] + 12'h247;
  assign sel_174461 = $signed({1'h0, add_174357}) < $signed({1'h0, sel_174359}) ? add_174357 : sel_174359;
  assign add_174464 = array_index_174396[11:0] + 12'h247;
  assign sel_174466 = $signed({1'h0, add_174362}) < $signed({1'h0, sel_174364}) ? add_174362 : sel_174364;
  assign array_index_174495 = set1_unflattened[7'h12];
  assign array_index_174498 = set2_unflattened[7'h12];
  assign add_174502 = array_index_174087[11:1] + 11'h79d;
  assign sel_174504 = $signed({1'h0, add_174400, array_index_173985[0]}) < $signed({1'h0, sel_174402}) ? {add_174400, array_index_173985[0]} : sel_174402;
  assign add_174506 = array_index_174090[11:1] + 11'h79d;
  assign sel_174508 = $signed({1'h0, add_174404, array_index_173988[0]}) < $signed({1'h0, sel_174406}) ? {add_174404, array_index_173988[0]} : sel_174406;
  assign add_174510 = array_index_174189[11:1] + 11'h347;
  assign sel_174512 = $signed({1'h0, add_174408, array_index_174087[0]}) < $signed({1'h0, sel_174410}) ? {add_174408, array_index_174087[0]} : sel_174410;
  assign add_174514 = array_index_174192[11:1] + 11'h347;
  assign sel_174516 = $signed({1'h0, add_174412, array_index_174090[0]}) < $signed({1'h0, sel_174414}) ? {add_174412, array_index_174090[0]} : sel_174414;
  assign add_174518 = array_index_174291[11:3] + 9'h0bd;
  assign sel_174521 = $signed({1'h0, add_174416, array_index_174189[2:0]}) < $signed({1'h0, sel_174419}) ? {add_174416, array_index_174189[2:0]} : sel_174419;
  assign add_174523 = array_index_174294[11:3] + 9'h0bd;
  assign sel_174526 = $signed({1'h0, add_174421, array_index_174192[2:0]}) < $signed({1'h0, sel_174424}) ? {add_174421, array_index_174192[2:0]} : sel_174424;
  assign add_174528 = array_index_174393[11:1] + 11'h247;
  assign sel_174531 = $signed({1'h0, add_174426, array_index_174291[0]}) < $signed({1'h0, sel_174429}) ? {add_174426, array_index_174291[0]} : sel_174429;
  assign add_174533 = array_index_174396[11:1] + 11'h247;
  assign sel_174536 = $signed({1'h0, add_174431, array_index_174294[0]}) < $signed({1'h0, sel_174434}) ? {add_174431, array_index_174294[0]} : sel_174434;
  assign add_174561 = array_index_174495[11:0] + 12'h247;
  assign sel_174563 = $signed({1'h0, add_174459}) < $signed({1'h0, sel_174461}) ? add_174459 : sel_174461;
  assign add_174566 = array_index_174498[11:0] + 12'h247;
  assign sel_174568 = $signed({1'h0, add_174464}) < $signed({1'h0, sel_174466}) ? add_174464 : sel_174466;
  assign array_index_174597 = set1_unflattened[7'h13];
  assign array_index_174600 = set2_unflattened[7'h13];
  assign add_174604 = array_index_174189[11:1] + 11'h79d;
  assign sel_174606 = $signed({1'h0, add_174502, array_index_174087[0]}) < $signed({1'h0, sel_174504}) ? {add_174502, array_index_174087[0]} : sel_174504;
  assign add_174608 = array_index_174192[11:1] + 11'h79d;
  assign sel_174610 = $signed({1'h0, add_174506, array_index_174090[0]}) < $signed({1'h0, sel_174508}) ? {add_174506, array_index_174090[0]} : sel_174508;
  assign add_174612 = array_index_174291[11:1] + 11'h347;
  assign sel_174614 = $signed({1'h0, add_174510, array_index_174189[0]}) < $signed({1'h0, sel_174512}) ? {add_174510, array_index_174189[0]} : sel_174512;
  assign add_174616 = array_index_174294[11:1] + 11'h347;
  assign sel_174618 = $signed({1'h0, add_174514, array_index_174192[0]}) < $signed({1'h0, sel_174516}) ? {add_174514, array_index_174192[0]} : sel_174516;
  assign add_174620 = array_index_174393[11:3] + 9'h0bd;
  assign sel_174623 = $signed({1'h0, add_174518, array_index_174291[2:0]}) < $signed({1'h0, sel_174521}) ? {add_174518, array_index_174291[2:0]} : sel_174521;
  assign add_174625 = array_index_174396[11:3] + 9'h0bd;
  assign sel_174628 = $signed({1'h0, add_174523, array_index_174294[2:0]}) < $signed({1'h0, sel_174526}) ? {add_174523, array_index_174294[2:0]} : sel_174526;
  assign add_174630 = array_index_174495[11:1] + 11'h247;
  assign sel_174633 = $signed({1'h0, add_174528, array_index_174393[0]}) < $signed({1'h0, sel_174531}) ? {add_174528, array_index_174393[0]} : sel_174531;
  assign add_174635 = array_index_174498[11:1] + 11'h247;
  assign sel_174638 = $signed({1'h0, add_174533, array_index_174396[0]}) < $signed({1'h0, sel_174536}) ? {add_174533, array_index_174396[0]} : sel_174536;
  assign add_174663 = array_index_174597[11:0] + 12'h247;
  assign sel_174665 = $signed({1'h0, add_174561}) < $signed({1'h0, sel_174563}) ? add_174561 : sel_174563;
  assign add_174668 = array_index_174600[11:0] + 12'h247;
  assign sel_174670 = $signed({1'h0, add_174566}) < $signed({1'h0, sel_174568}) ? add_174566 : sel_174568;
  assign array_index_174699 = set1_unflattened[7'h14];
  assign array_index_174702 = set2_unflattened[7'h14];
  assign add_174706 = array_index_174291[11:1] + 11'h79d;
  assign sel_174708 = $signed({1'h0, add_174604, array_index_174189[0]}) < $signed({1'h0, sel_174606}) ? {add_174604, array_index_174189[0]} : sel_174606;
  assign add_174710 = array_index_174294[11:1] + 11'h79d;
  assign sel_174712 = $signed({1'h0, add_174608, array_index_174192[0]}) < $signed({1'h0, sel_174610}) ? {add_174608, array_index_174192[0]} : sel_174610;
  assign add_174714 = array_index_174393[11:1] + 11'h347;
  assign sel_174716 = $signed({1'h0, add_174612, array_index_174291[0]}) < $signed({1'h0, sel_174614}) ? {add_174612, array_index_174291[0]} : sel_174614;
  assign add_174718 = array_index_174396[11:1] + 11'h347;
  assign sel_174720 = $signed({1'h0, add_174616, array_index_174294[0]}) < $signed({1'h0, sel_174618}) ? {add_174616, array_index_174294[0]} : sel_174618;
  assign add_174722 = array_index_174495[11:3] + 9'h0bd;
  assign sel_174725 = $signed({1'h0, add_174620, array_index_174393[2:0]}) < $signed({1'h0, sel_174623}) ? {add_174620, array_index_174393[2:0]} : sel_174623;
  assign add_174727 = array_index_174498[11:3] + 9'h0bd;
  assign sel_174730 = $signed({1'h0, add_174625, array_index_174396[2:0]}) < $signed({1'h0, sel_174628}) ? {add_174625, array_index_174396[2:0]} : sel_174628;
  assign add_174732 = array_index_174597[11:1] + 11'h247;
  assign sel_174735 = $signed({1'h0, add_174630, array_index_174495[0]}) < $signed({1'h0, sel_174633}) ? {add_174630, array_index_174495[0]} : sel_174633;
  assign add_174737 = array_index_174600[11:1] + 11'h247;
  assign sel_174740 = $signed({1'h0, add_174635, array_index_174498[0]}) < $signed({1'h0, sel_174638}) ? {add_174635, array_index_174498[0]} : sel_174638;
  assign add_174765 = array_index_174699[11:0] + 12'h247;
  assign sel_174767 = $signed({1'h0, add_174663}) < $signed({1'h0, sel_174665}) ? add_174663 : sel_174665;
  assign add_174770 = array_index_174702[11:0] + 12'h247;
  assign sel_174772 = $signed({1'h0, add_174668}) < $signed({1'h0, sel_174670}) ? add_174668 : sel_174670;
  assign array_index_174801 = set1_unflattened[7'h15];
  assign array_index_174804 = set2_unflattened[7'h15];
  assign add_174808 = array_index_174393[11:1] + 11'h79d;
  assign sel_174810 = $signed({1'h0, add_174706, array_index_174291[0]}) < $signed({1'h0, sel_174708}) ? {add_174706, array_index_174291[0]} : sel_174708;
  assign add_174812 = array_index_174396[11:1] + 11'h79d;
  assign sel_174814 = $signed({1'h0, add_174710, array_index_174294[0]}) < $signed({1'h0, sel_174712}) ? {add_174710, array_index_174294[0]} : sel_174712;
  assign add_174816 = array_index_174495[11:1] + 11'h347;
  assign sel_174818 = $signed({1'h0, add_174714, array_index_174393[0]}) < $signed({1'h0, sel_174716}) ? {add_174714, array_index_174393[0]} : sel_174716;
  assign add_174820 = array_index_174498[11:1] + 11'h347;
  assign sel_174822 = $signed({1'h0, add_174718, array_index_174396[0]}) < $signed({1'h0, sel_174720}) ? {add_174718, array_index_174396[0]} : sel_174720;
  assign add_174824 = array_index_174597[11:3] + 9'h0bd;
  assign sel_174827 = $signed({1'h0, add_174722, array_index_174495[2:0]}) < $signed({1'h0, sel_174725}) ? {add_174722, array_index_174495[2:0]} : sel_174725;
  assign add_174829 = array_index_174600[11:3] + 9'h0bd;
  assign sel_174832 = $signed({1'h0, add_174727, array_index_174498[2:0]}) < $signed({1'h0, sel_174730}) ? {add_174727, array_index_174498[2:0]} : sel_174730;
  assign add_174834 = array_index_174699[11:1] + 11'h247;
  assign sel_174837 = $signed({1'h0, add_174732, array_index_174597[0]}) < $signed({1'h0, sel_174735}) ? {add_174732, array_index_174597[0]} : sel_174735;
  assign add_174839 = array_index_174702[11:1] + 11'h247;
  assign sel_174842 = $signed({1'h0, add_174737, array_index_174600[0]}) < $signed({1'h0, sel_174740}) ? {add_174737, array_index_174600[0]} : sel_174740;
  assign add_174867 = array_index_174801[11:0] + 12'h247;
  assign sel_174869 = $signed({1'h0, add_174765}) < $signed({1'h0, sel_174767}) ? add_174765 : sel_174767;
  assign add_174872 = array_index_174804[11:0] + 12'h247;
  assign sel_174874 = $signed({1'h0, add_174770}) < $signed({1'h0, sel_174772}) ? add_174770 : sel_174772;
  assign array_index_174903 = set1_unflattened[7'h16];
  assign array_index_174906 = set2_unflattened[7'h16];
  assign add_174910 = array_index_174495[11:1] + 11'h79d;
  assign sel_174912 = $signed({1'h0, add_174808, array_index_174393[0]}) < $signed({1'h0, sel_174810}) ? {add_174808, array_index_174393[0]} : sel_174810;
  assign add_174914 = array_index_174498[11:1] + 11'h79d;
  assign sel_174916 = $signed({1'h0, add_174812, array_index_174396[0]}) < $signed({1'h0, sel_174814}) ? {add_174812, array_index_174396[0]} : sel_174814;
  assign add_174918 = array_index_174597[11:1] + 11'h347;
  assign sel_174920 = $signed({1'h0, add_174816, array_index_174495[0]}) < $signed({1'h0, sel_174818}) ? {add_174816, array_index_174495[0]} : sel_174818;
  assign add_174922 = array_index_174600[11:1] + 11'h347;
  assign sel_174924 = $signed({1'h0, add_174820, array_index_174498[0]}) < $signed({1'h0, sel_174822}) ? {add_174820, array_index_174498[0]} : sel_174822;
  assign add_174926 = array_index_174699[11:3] + 9'h0bd;
  assign sel_174929 = $signed({1'h0, add_174824, array_index_174597[2:0]}) < $signed({1'h0, sel_174827}) ? {add_174824, array_index_174597[2:0]} : sel_174827;
  assign add_174931 = array_index_174702[11:3] + 9'h0bd;
  assign sel_174934 = $signed({1'h0, add_174829, array_index_174600[2:0]}) < $signed({1'h0, sel_174832}) ? {add_174829, array_index_174600[2:0]} : sel_174832;
  assign add_174936 = array_index_174801[11:1] + 11'h247;
  assign sel_174939 = $signed({1'h0, add_174834, array_index_174699[0]}) < $signed({1'h0, sel_174837}) ? {add_174834, array_index_174699[0]} : sel_174837;
  assign add_174941 = array_index_174804[11:1] + 11'h247;
  assign sel_174944 = $signed({1'h0, add_174839, array_index_174702[0]}) < $signed({1'h0, sel_174842}) ? {add_174839, array_index_174702[0]} : sel_174842;
  assign add_174969 = array_index_174903[11:0] + 12'h247;
  assign sel_174971 = $signed({1'h0, add_174867}) < $signed({1'h0, sel_174869}) ? add_174867 : sel_174869;
  assign add_174974 = array_index_174906[11:0] + 12'h247;
  assign sel_174976 = $signed({1'h0, add_174872}) < $signed({1'h0, sel_174874}) ? add_174872 : sel_174874;
  assign array_index_175005 = set1_unflattened[7'h17];
  assign array_index_175008 = set2_unflattened[7'h17];
  assign add_175012 = array_index_174597[11:1] + 11'h79d;
  assign sel_175014 = $signed({1'h0, add_174910, array_index_174495[0]}) < $signed({1'h0, sel_174912}) ? {add_174910, array_index_174495[0]} : sel_174912;
  assign add_175016 = array_index_174600[11:1] + 11'h79d;
  assign sel_175018 = $signed({1'h0, add_174914, array_index_174498[0]}) < $signed({1'h0, sel_174916}) ? {add_174914, array_index_174498[0]} : sel_174916;
  assign add_175020 = array_index_174699[11:1] + 11'h347;
  assign sel_175022 = $signed({1'h0, add_174918, array_index_174597[0]}) < $signed({1'h0, sel_174920}) ? {add_174918, array_index_174597[0]} : sel_174920;
  assign add_175024 = array_index_174702[11:1] + 11'h347;
  assign sel_175026 = $signed({1'h0, add_174922, array_index_174600[0]}) < $signed({1'h0, sel_174924}) ? {add_174922, array_index_174600[0]} : sel_174924;
  assign add_175028 = array_index_174801[11:3] + 9'h0bd;
  assign sel_175031 = $signed({1'h0, add_174926, array_index_174699[2:0]}) < $signed({1'h0, sel_174929}) ? {add_174926, array_index_174699[2:0]} : sel_174929;
  assign add_175033 = array_index_174804[11:3] + 9'h0bd;
  assign sel_175036 = $signed({1'h0, add_174931, array_index_174702[2:0]}) < $signed({1'h0, sel_174934}) ? {add_174931, array_index_174702[2:0]} : sel_174934;
  assign add_175038 = array_index_174903[11:1] + 11'h247;
  assign sel_175041 = $signed({1'h0, add_174936, array_index_174801[0]}) < $signed({1'h0, sel_174939}) ? {add_174936, array_index_174801[0]} : sel_174939;
  assign add_175043 = array_index_174906[11:1] + 11'h247;
  assign sel_175046 = $signed({1'h0, add_174941, array_index_174804[0]}) < $signed({1'h0, sel_174944}) ? {add_174941, array_index_174804[0]} : sel_174944;
  assign add_175071 = array_index_175005[11:0] + 12'h247;
  assign sel_175073 = $signed({1'h0, add_174969}) < $signed({1'h0, sel_174971}) ? add_174969 : sel_174971;
  assign add_175076 = array_index_175008[11:0] + 12'h247;
  assign sel_175078 = $signed({1'h0, add_174974}) < $signed({1'h0, sel_174976}) ? add_174974 : sel_174976;
  assign array_index_175107 = set1_unflattened[7'h18];
  assign array_index_175110 = set2_unflattened[7'h18];
  assign add_175114 = array_index_174699[11:1] + 11'h79d;
  assign sel_175116 = $signed({1'h0, add_175012, array_index_174597[0]}) < $signed({1'h0, sel_175014}) ? {add_175012, array_index_174597[0]} : sel_175014;
  assign add_175118 = array_index_174702[11:1] + 11'h79d;
  assign sel_175120 = $signed({1'h0, add_175016, array_index_174600[0]}) < $signed({1'h0, sel_175018}) ? {add_175016, array_index_174600[0]} : sel_175018;
  assign add_175122 = array_index_174801[11:1] + 11'h347;
  assign sel_175124 = $signed({1'h0, add_175020, array_index_174699[0]}) < $signed({1'h0, sel_175022}) ? {add_175020, array_index_174699[0]} : sel_175022;
  assign add_175126 = array_index_174804[11:1] + 11'h347;
  assign sel_175128 = $signed({1'h0, add_175024, array_index_174702[0]}) < $signed({1'h0, sel_175026}) ? {add_175024, array_index_174702[0]} : sel_175026;
  assign add_175130 = array_index_174903[11:3] + 9'h0bd;
  assign sel_175133 = $signed({1'h0, add_175028, array_index_174801[2:0]}) < $signed({1'h0, sel_175031}) ? {add_175028, array_index_174801[2:0]} : sel_175031;
  assign add_175135 = array_index_174906[11:3] + 9'h0bd;
  assign sel_175138 = $signed({1'h0, add_175033, array_index_174804[2:0]}) < $signed({1'h0, sel_175036}) ? {add_175033, array_index_174804[2:0]} : sel_175036;
  assign add_175140 = array_index_175005[11:1] + 11'h247;
  assign sel_175143 = $signed({1'h0, add_175038, array_index_174903[0]}) < $signed({1'h0, sel_175041}) ? {add_175038, array_index_174903[0]} : sel_175041;
  assign add_175145 = array_index_175008[11:1] + 11'h247;
  assign sel_175148 = $signed({1'h0, add_175043, array_index_174906[0]}) < $signed({1'h0, sel_175046}) ? {add_175043, array_index_174906[0]} : sel_175046;
  assign add_175173 = array_index_175107[11:0] + 12'h247;
  assign sel_175175 = $signed({1'h0, add_175071}) < $signed({1'h0, sel_175073}) ? add_175071 : sel_175073;
  assign add_175178 = array_index_175110[11:0] + 12'h247;
  assign sel_175180 = $signed({1'h0, add_175076}) < $signed({1'h0, sel_175078}) ? add_175076 : sel_175078;
  assign array_index_175209 = set1_unflattened[7'h19];
  assign array_index_175212 = set2_unflattened[7'h19];
  assign add_175216 = array_index_174801[11:1] + 11'h79d;
  assign sel_175218 = $signed({1'h0, add_175114, array_index_174699[0]}) < $signed({1'h0, sel_175116}) ? {add_175114, array_index_174699[0]} : sel_175116;
  assign add_175220 = array_index_174804[11:1] + 11'h79d;
  assign sel_175222 = $signed({1'h0, add_175118, array_index_174702[0]}) < $signed({1'h0, sel_175120}) ? {add_175118, array_index_174702[0]} : sel_175120;
  assign add_175224 = array_index_174903[11:1] + 11'h347;
  assign sel_175226 = $signed({1'h0, add_175122, array_index_174801[0]}) < $signed({1'h0, sel_175124}) ? {add_175122, array_index_174801[0]} : sel_175124;
  assign add_175228 = array_index_174906[11:1] + 11'h347;
  assign sel_175230 = $signed({1'h0, add_175126, array_index_174804[0]}) < $signed({1'h0, sel_175128}) ? {add_175126, array_index_174804[0]} : sel_175128;
  assign add_175232 = array_index_175005[11:3] + 9'h0bd;
  assign sel_175235 = $signed({1'h0, add_175130, array_index_174903[2:0]}) < $signed({1'h0, sel_175133}) ? {add_175130, array_index_174903[2:0]} : sel_175133;
  assign add_175237 = array_index_175008[11:3] + 9'h0bd;
  assign sel_175240 = $signed({1'h0, add_175135, array_index_174906[2:0]}) < $signed({1'h0, sel_175138}) ? {add_175135, array_index_174906[2:0]} : sel_175138;
  assign add_175242 = array_index_175107[11:1] + 11'h247;
  assign sel_175245 = $signed({1'h0, add_175140, array_index_175005[0]}) < $signed({1'h0, sel_175143}) ? {add_175140, array_index_175005[0]} : sel_175143;
  assign add_175247 = array_index_175110[11:1] + 11'h247;
  assign sel_175250 = $signed({1'h0, add_175145, array_index_175008[0]}) < $signed({1'h0, sel_175148}) ? {add_175145, array_index_175008[0]} : sel_175148;
  assign add_175275 = array_index_175209[11:0] + 12'h247;
  assign sel_175277 = $signed({1'h0, add_175173}) < $signed({1'h0, sel_175175}) ? add_175173 : sel_175175;
  assign add_175280 = array_index_175212[11:0] + 12'h247;
  assign sel_175282 = $signed({1'h0, add_175178}) < $signed({1'h0, sel_175180}) ? add_175178 : sel_175180;
  assign array_index_175311 = set1_unflattened[7'h1a];
  assign array_index_175314 = set2_unflattened[7'h1a];
  assign add_175318 = array_index_174903[11:1] + 11'h79d;
  assign sel_175320 = $signed({1'h0, add_175216, array_index_174801[0]}) < $signed({1'h0, sel_175218}) ? {add_175216, array_index_174801[0]} : sel_175218;
  assign add_175322 = array_index_174906[11:1] + 11'h79d;
  assign sel_175324 = $signed({1'h0, add_175220, array_index_174804[0]}) < $signed({1'h0, sel_175222}) ? {add_175220, array_index_174804[0]} : sel_175222;
  assign add_175326 = array_index_175005[11:1] + 11'h347;
  assign sel_175328 = $signed({1'h0, add_175224, array_index_174903[0]}) < $signed({1'h0, sel_175226}) ? {add_175224, array_index_174903[0]} : sel_175226;
  assign add_175330 = array_index_175008[11:1] + 11'h347;
  assign sel_175332 = $signed({1'h0, add_175228, array_index_174906[0]}) < $signed({1'h0, sel_175230}) ? {add_175228, array_index_174906[0]} : sel_175230;
  assign add_175334 = array_index_175107[11:3] + 9'h0bd;
  assign sel_175337 = $signed({1'h0, add_175232, array_index_175005[2:0]}) < $signed({1'h0, sel_175235}) ? {add_175232, array_index_175005[2:0]} : sel_175235;
  assign add_175339 = array_index_175110[11:3] + 9'h0bd;
  assign sel_175342 = $signed({1'h0, add_175237, array_index_175008[2:0]}) < $signed({1'h0, sel_175240}) ? {add_175237, array_index_175008[2:0]} : sel_175240;
  assign add_175344 = array_index_175209[11:1] + 11'h247;
  assign sel_175347 = $signed({1'h0, add_175242, array_index_175107[0]}) < $signed({1'h0, sel_175245}) ? {add_175242, array_index_175107[0]} : sel_175245;
  assign add_175349 = array_index_175212[11:1] + 11'h247;
  assign sel_175352 = $signed({1'h0, add_175247, array_index_175110[0]}) < $signed({1'h0, sel_175250}) ? {add_175247, array_index_175110[0]} : sel_175250;
  assign add_175377 = array_index_175311[11:0] + 12'h247;
  assign sel_175379 = $signed({1'h0, add_175275}) < $signed({1'h0, sel_175277}) ? add_175275 : sel_175277;
  assign add_175382 = array_index_175314[11:0] + 12'h247;
  assign sel_175384 = $signed({1'h0, add_175280}) < $signed({1'h0, sel_175282}) ? add_175280 : sel_175282;
  assign array_index_175413 = set1_unflattened[7'h1b];
  assign array_index_175416 = set2_unflattened[7'h1b];
  assign add_175420 = array_index_175005[11:1] + 11'h79d;
  assign sel_175422 = $signed({1'h0, add_175318, array_index_174903[0]}) < $signed({1'h0, sel_175320}) ? {add_175318, array_index_174903[0]} : sel_175320;
  assign add_175424 = array_index_175008[11:1] + 11'h79d;
  assign sel_175426 = $signed({1'h0, add_175322, array_index_174906[0]}) < $signed({1'h0, sel_175324}) ? {add_175322, array_index_174906[0]} : sel_175324;
  assign add_175428 = array_index_175107[11:1] + 11'h347;
  assign sel_175430 = $signed({1'h0, add_175326, array_index_175005[0]}) < $signed({1'h0, sel_175328}) ? {add_175326, array_index_175005[0]} : sel_175328;
  assign add_175432 = array_index_175110[11:1] + 11'h347;
  assign sel_175434 = $signed({1'h0, add_175330, array_index_175008[0]}) < $signed({1'h0, sel_175332}) ? {add_175330, array_index_175008[0]} : sel_175332;
  assign add_175436 = array_index_175209[11:3] + 9'h0bd;
  assign sel_175439 = $signed({1'h0, add_175334, array_index_175107[2:0]}) < $signed({1'h0, sel_175337}) ? {add_175334, array_index_175107[2:0]} : sel_175337;
  assign add_175441 = array_index_175212[11:3] + 9'h0bd;
  assign sel_175444 = $signed({1'h0, add_175339, array_index_175110[2:0]}) < $signed({1'h0, sel_175342}) ? {add_175339, array_index_175110[2:0]} : sel_175342;
  assign add_175446 = array_index_175311[11:1] + 11'h247;
  assign sel_175449 = $signed({1'h0, add_175344, array_index_175209[0]}) < $signed({1'h0, sel_175347}) ? {add_175344, array_index_175209[0]} : sel_175347;
  assign add_175451 = array_index_175314[11:1] + 11'h247;
  assign sel_175454 = $signed({1'h0, add_175349, array_index_175212[0]}) < $signed({1'h0, sel_175352}) ? {add_175349, array_index_175212[0]} : sel_175352;
  assign add_175479 = array_index_175413[11:0] + 12'h247;
  assign sel_175481 = $signed({1'h0, add_175377}) < $signed({1'h0, sel_175379}) ? add_175377 : sel_175379;
  assign add_175484 = array_index_175416[11:0] + 12'h247;
  assign sel_175486 = $signed({1'h0, add_175382}) < $signed({1'h0, sel_175384}) ? add_175382 : sel_175384;
  assign array_index_175515 = set1_unflattened[7'h1c];
  assign array_index_175518 = set2_unflattened[7'h1c];
  assign add_175522 = array_index_175107[11:1] + 11'h79d;
  assign sel_175524 = $signed({1'h0, add_175420, array_index_175005[0]}) < $signed({1'h0, sel_175422}) ? {add_175420, array_index_175005[0]} : sel_175422;
  assign add_175526 = array_index_175110[11:1] + 11'h79d;
  assign sel_175528 = $signed({1'h0, add_175424, array_index_175008[0]}) < $signed({1'h0, sel_175426}) ? {add_175424, array_index_175008[0]} : sel_175426;
  assign add_175530 = array_index_175209[11:1] + 11'h347;
  assign sel_175532 = $signed({1'h0, add_175428, array_index_175107[0]}) < $signed({1'h0, sel_175430}) ? {add_175428, array_index_175107[0]} : sel_175430;
  assign add_175534 = array_index_175212[11:1] + 11'h347;
  assign sel_175536 = $signed({1'h0, add_175432, array_index_175110[0]}) < $signed({1'h0, sel_175434}) ? {add_175432, array_index_175110[0]} : sel_175434;
  assign add_175538 = array_index_175311[11:3] + 9'h0bd;
  assign sel_175541 = $signed({1'h0, add_175436, array_index_175209[2:0]}) < $signed({1'h0, sel_175439}) ? {add_175436, array_index_175209[2:0]} : sel_175439;
  assign add_175543 = array_index_175314[11:3] + 9'h0bd;
  assign sel_175546 = $signed({1'h0, add_175441, array_index_175212[2:0]}) < $signed({1'h0, sel_175444}) ? {add_175441, array_index_175212[2:0]} : sel_175444;
  assign add_175548 = array_index_175413[11:1] + 11'h247;
  assign sel_175551 = $signed({1'h0, add_175446, array_index_175311[0]}) < $signed({1'h0, sel_175449}) ? {add_175446, array_index_175311[0]} : sel_175449;
  assign add_175553 = array_index_175416[11:1] + 11'h247;
  assign sel_175556 = $signed({1'h0, add_175451, array_index_175314[0]}) < $signed({1'h0, sel_175454}) ? {add_175451, array_index_175314[0]} : sel_175454;
  assign add_175581 = array_index_175515[11:0] + 12'h247;
  assign sel_175583 = $signed({1'h0, add_175479}) < $signed({1'h0, sel_175481}) ? add_175479 : sel_175481;
  assign add_175586 = array_index_175518[11:0] + 12'h247;
  assign sel_175588 = $signed({1'h0, add_175484}) < $signed({1'h0, sel_175486}) ? add_175484 : sel_175486;
  assign array_index_175617 = set1_unflattened[7'h1d];
  assign array_index_175620 = set2_unflattened[7'h1d];
  assign add_175624 = array_index_175209[11:1] + 11'h79d;
  assign sel_175626 = $signed({1'h0, add_175522, array_index_175107[0]}) < $signed({1'h0, sel_175524}) ? {add_175522, array_index_175107[0]} : sel_175524;
  assign add_175628 = array_index_175212[11:1] + 11'h79d;
  assign sel_175630 = $signed({1'h0, add_175526, array_index_175110[0]}) < $signed({1'h0, sel_175528}) ? {add_175526, array_index_175110[0]} : sel_175528;
  assign add_175632 = array_index_175311[11:1] + 11'h347;
  assign sel_175634 = $signed({1'h0, add_175530, array_index_175209[0]}) < $signed({1'h0, sel_175532}) ? {add_175530, array_index_175209[0]} : sel_175532;
  assign add_175636 = array_index_175314[11:1] + 11'h347;
  assign sel_175638 = $signed({1'h0, add_175534, array_index_175212[0]}) < $signed({1'h0, sel_175536}) ? {add_175534, array_index_175212[0]} : sel_175536;
  assign add_175640 = array_index_175413[11:3] + 9'h0bd;
  assign sel_175643 = $signed({1'h0, add_175538, array_index_175311[2:0]}) < $signed({1'h0, sel_175541}) ? {add_175538, array_index_175311[2:0]} : sel_175541;
  assign add_175645 = array_index_175416[11:3] + 9'h0bd;
  assign sel_175648 = $signed({1'h0, add_175543, array_index_175314[2:0]}) < $signed({1'h0, sel_175546}) ? {add_175543, array_index_175314[2:0]} : sel_175546;
  assign add_175650 = array_index_175515[11:1] + 11'h247;
  assign sel_175653 = $signed({1'h0, add_175548, array_index_175413[0]}) < $signed({1'h0, sel_175551}) ? {add_175548, array_index_175413[0]} : sel_175551;
  assign add_175655 = array_index_175518[11:1] + 11'h247;
  assign sel_175658 = $signed({1'h0, add_175553, array_index_175416[0]}) < $signed({1'h0, sel_175556}) ? {add_175553, array_index_175416[0]} : sel_175556;
  assign add_175683 = array_index_175617[11:0] + 12'h247;
  assign sel_175685 = $signed({1'h0, add_175581}) < $signed({1'h0, sel_175583}) ? add_175581 : sel_175583;
  assign add_175688 = array_index_175620[11:0] + 12'h247;
  assign sel_175690 = $signed({1'h0, add_175586}) < $signed({1'h0, sel_175588}) ? add_175586 : sel_175588;
  assign array_index_175719 = set1_unflattened[7'h1e];
  assign array_index_175722 = set2_unflattened[7'h1e];
  assign add_175726 = array_index_175311[11:1] + 11'h79d;
  assign sel_175728 = $signed({1'h0, add_175624, array_index_175209[0]}) < $signed({1'h0, sel_175626}) ? {add_175624, array_index_175209[0]} : sel_175626;
  assign add_175730 = array_index_175314[11:1] + 11'h79d;
  assign sel_175732 = $signed({1'h0, add_175628, array_index_175212[0]}) < $signed({1'h0, sel_175630}) ? {add_175628, array_index_175212[0]} : sel_175630;
  assign add_175734 = array_index_175413[11:1] + 11'h347;
  assign sel_175736 = $signed({1'h0, add_175632, array_index_175311[0]}) < $signed({1'h0, sel_175634}) ? {add_175632, array_index_175311[0]} : sel_175634;
  assign add_175738 = array_index_175416[11:1] + 11'h347;
  assign sel_175740 = $signed({1'h0, add_175636, array_index_175314[0]}) < $signed({1'h0, sel_175638}) ? {add_175636, array_index_175314[0]} : sel_175638;
  assign add_175742 = array_index_175515[11:3] + 9'h0bd;
  assign sel_175745 = $signed({1'h0, add_175640, array_index_175413[2:0]}) < $signed({1'h0, sel_175643}) ? {add_175640, array_index_175413[2:0]} : sel_175643;
  assign add_175747 = array_index_175518[11:3] + 9'h0bd;
  assign sel_175750 = $signed({1'h0, add_175645, array_index_175416[2:0]}) < $signed({1'h0, sel_175648}) ? {add_175645, array_index_175416[2:0]} : sel_175648;
  assign add_175752 = array_index_175617[11:1] + 11'h247;
  assign sel_175755 = $signed({1'h0, add_175650, array_index_175515[0]}) < $signed({1'h0, sel_175653}) ? {add_175650, array_index_175515[0]} : sel_175653;
  assign add_175757 = array_index_175620[11:1] + 11'h247;
  assign sel_175760 = $signed({1'h0, add_175655, array_index_175518[0]}) < $signed({1'h0, sel_175658}) ? {add_175655, array_index_175518[0]} : sel_175658;
  assign add_175785 = array_index_175719[11:0] + 12'h247;
  assign sel_175787 = $signed({1'h0, add_175683}) < $signed({1'h0, sel_175685}) ? add_175683 : sel_175685;
  assign add_175790 = array_index_175722[11:0] + 12'h247;
  assign sel_175792 = $signed({1'h0, add_175688}) < $signed({1'h0, sel_175690}) ? add_175688 : sel_175690;
  assign array_index_175821 = set1_unflattened[7'h1f];
  assign array_index_175824 = set2_unflattened[7'h1f];
  assign add_175828 = array_index_175413[11:1] + 11'h79d;
  assign sel_175830 = $signed({1'h0, add_175726, array_index_175311[0]}) < $signed({1'h0, sel_175728}) ? {add_175726, array_index_175311[0]} : sel_175728;
  assign add_175832 = array_index_175416[11:1] + 11'h79d;
  assign sel_175834 = $signed({1'h0, add_175730, array_index_175314[0]}) < $signed({1'h0, sel_175732}) ? {add_175730, array_index_175314[0]} : sel_175732;
  assign add_175836 = array_index_175515[11:1] + 11'h347;
  assign sel_175838 = $signed({1'h0, add_175734, array_index_175413[0]}) < $signed({1'h0, sel_175736}) ? {add_175734, array_index_175413[0]} : sel_175736;
  assign add_175840 = array_index_175518[11:1] + 11'h347;
  assign sel_175842 = $signed({1'h0, add_175738, array_index_175416[0]}) < $signed({1'h0, sel_175740}) ? {add_175738, array_index_175416[0]} : sel_175740;
  assign add_175844 = array_index_175617[11:3] + 9'h0bd;
  assign sel_175847 = $signed({1'h0, add_175742, array_index_175515[2:0]}) < $signed({1'h0, sel_175745}) ? {add_175742, array_index_175515[2:0]} : sel_175745;
  assign add_175849 = array_index_175620[11:3] + 9'h0bd;
  assign sel_175852 = $signed({1'h0, add_175747, array_index_175518[2:0]}) < $signed({1'h0, sel_175750}) ? {add_175747, array_index_175518[2:0]} : sel_175750;
  assign add_175854 = array_index_175719[11:1] + 11'h247;
  assign sel_175857 = $signed({1'h0, add_175752, array_index_175617[0]}) < $signed({1'h0, sel_175755}) ? {add_175752, array_index_175617[0]} : sel_175755;
  assign add_175859 = array_index_175722[11:1] + 11'h247;
  assign sel_175862 = $signed({1'h0, add_175757, array_index_175620[0]}) < $signed({1'h0, sel_175760}) ? {add_175757, array_index_175620[0]} : sel_175760;
  assign add_175887 = array_index_175821[11:0] + 12'h247;
  assign sel_175889 = $signed({1'h0, add_175785}) < $signed({1'h0, sel_175787}) ? add_175785 : sel_175787;
  assign add_175892 = array_index_175824[11:0] + 12'h247;
  assign sel_175894 = $signed({1'h0, add_175790}) < $signed({1'h0, sel_175792}) ? add_175790 : sel_175792;
  assign array_index_175923 = set1_unflattened[7'h20];
  assign array_index_175926 = set2_unflattened[7'h20];
  assign add_175930 = array_index_175515[11:1] + 11'h79d;
  assign sel_175932 = $signed({1'h0, add_175828, array_index_175413[0]}) < $signed({1'h0, sel_175830}) ? {add_175828, array_index_175413[0]} : sel_175830;
  assign add_175934 = array_index_175518[11:1] + 11'h79d;
  assign sel_175936 = $signed({1'h0, add_175832, array_index_175416[0]}) < $signed({1'h0, sel_175834}) ? {add_175832, array_index_175416[0]} : sel_175834;
  assign add_175938 = array_index_175617[11:1] + 11'h347;
  assign sel_175940 = $signed({1'h0, add_175836, array_index_175515[0]}) < $signed({1'h0, sel_175838}) ? {add_175836, array_index_175515[0]} : sel_175838;
  assign add_175942 = array_index_175620[11:1] + 11'h347;
  assign sel_175944 = $signed({1'h0, add_175840, array_index_175518[0]}) < $signed({1'h0, sel_175842}) ? {add_175840, array_index_175518[0]} : sel_175842;
  assign add_175946 = array_index_175719[11:3] + 9'h0bd;
  assign sel_175949 = $signed({1'h0, add_175844, array_index_175617[2:0]}) < $signed({1'h0, sel_175847}) ? {add_175844, array_index_175617[2:0]} : sel_175847;
  assign add_175951 = array_index_175722[11:3] + 9'h0bd;
  assign sel_175954 = $signed({1'h0, add_175849, array_index_175620[2:0]}) < $signed({1'h0, sel_175852}) ? {add_175849, array_index_175620[2:0]} : sel_175852;
  assign add_175956 = array_index_175821[11:1] + 11'h247;
  assign sel_175959 = $signed({1'h0, add_175854, array_index_175719[0]}) < $signed({1'h0, sel_175857}) ? {add_175854, array_index_175719[0]} : sel_175857;
  assign add_175961 = array_index_175824[11:1] + 11'h247;
  assign sel_175964 = $signed({1'h0, add_175859, array_index_175722[0]}) < $signed({1'h0, sel_175862}) ? {add_175859, array_index_175722[0]} : sel_175862;
  assign add_175989 = array_index_175923[11:0] + 12'h247;
  assign sel_175991 = $signed({1'h0, add_175887}) < $signed({1'h0, sel_175889}) ? add_175887 : sel_175889;
  assign add_175994 = array_index_175926[11:0] + 12'h247;
  assign sel_175996 = $signed({1'h0, add_175892}) < $signed({1'h0, sel_175894}) ? add_175892 : sel_175894;
  assign array_index_176025 = set1_unflattened[7'h21];
  assign array_index_176028 = set2_unflattened[7'h21];
  assign add_176032 = array_index_175617[11:1] + 11'h79d;
  assign sel_176034 = $signed({1'h0, add_175930, array_index_175515[0]}) < $signed({1'h0, sel_175932}) ? {add_175930, array_index_175515[0]} : sel_175932;
  assign add_176036 = array_index_175620[11:1] + 11'h79d;
  assign sel_176038 = $signed({1'h0, add_175934, array_index_175518[0]}) < $signed({1'h0, sel_175936}) ? {add_175934, array_index_175518[0]} : sel_175936;
  assign add_176040 = array_index_175719[11:1] + 11'h347;
  assign sel_176042 = $signed({1'h0, add_175938, array_index_175617[0]}) < $signed({1'h0, sel_175940}) ? {add_175938, array_index_175617[0]} : sel_175940;
  assign add_176044 = array_index_175722[11:1] + 11'h347;
  assign sel_176046 = $signed({1'h0, add_175942, array_index_175620[0]}) < $signed({1'h0, sel_175944}) ? {add_175942, array_index_175620[0]} : sel_175944;
  assign add_176048 = array_index_175821[11:3] + 9'h0bd;
  assign sel_176051 = $signed({1'h0, add_175946, array_index_175719[2:0]}) < $signed({1'h0, sel_175949}) ? {add_175946, array_index_175719[2:0]} : sel_175949;
  assign add_176053 = array_index_175824[11:3] + 9'h0bd;
  assign sel_176056 = $signed({1'h0, add_175951, array_index_175722[2:0]}) < $signed({1'h0, sel_175954}) ? {add_175951, array_index_175722[2:0]} : sel_175954;
  assign add_176058 = array_index_175923[11:1] + 11'h247;
  assign sel_176061 = $signed({1'h0, add_175956, array_index_175821[0]}) < $signed({1'h0, sel_175959}) ? {add_175956, array_index_175821[0]} : sel_175959;
  assign add_176063 = array_index_175926[11:1] + 11'h247;
  assign sel_176066 = $signed({1'h0, add_175961, array_index_175824[0]}) < $signed({1'h0, sel_175964}) ? {add_175961, array_index_175824[0]} : sel_175964;
  assign add_176091 = array_index_176025[11:0] + 12'h247;
  assign sel_176093 = $signed({1'h0, add_175989}) < $signed({1'h0, sel_175991}) ? add_175989 : sel_175991;
  assign add_176096 = array_index_176028[11:0] + 12'h247;
  assign sel_176098 = $signed({1'h0, add_175994}) < $signed({1'h0, sel_175996}) ? add_175994 : sel_175996;
  assign array_index_176127 = set1_unflattened[7'h22];
  assign array_index_176130 = set2_unflattened[7'h22];
  assign add_176134 = array_index_175719[11:1] + 11'h79d;
  assign sel_176136 = $signed({1'h0, add_176032, array_index_175617[0]}) < $signed({1'h0, sel_176034}) ? {add_176032, array_index_175617[0]} : sel_176034;
  assign add_176138 = array_index_175722[11:1] + 11'h79d;
  assign sel_176140 = $signed({1'h0, add_176036, array_index_175620[0]}) < $signed({1'h0, sel_176038}) ? {add_176036, array_index_175620[0]} : sel_176038;
  assign add_176142 = array_index_175821[11:1] + 11'h347;
  assign sel_176144 = $signed({1'h0, add_176040, array_index_175719[0]}) < $signed({1'h0, sel_176042}) ? {add_176040, array_index_175719[0]} : sel_176042;
  assign add_176146 = array_index_175824[11:1] + 11'h347;
  assign sel_176148 = $signed({1'h0, add_176044, array_index_175722[0]}) < $signed({1'h0, sel_176046}) ? {add_176044, array_index_175722[0]} : sel_176046;
  assign add_176150 = array_index_175923[11:3] + 9'h0bd;
  assign sel_176153 = $signed({1'h0, add_176048, array_index_175821[2:0]}) < $signed({1'h0, sel_176051}) ? {add_176048, array_index_175821[2:0]} : sel_176051;
  assign add_176155 = array_index_175926[11:3] + 9'h0bd;
  assign sel_176158 = $signed({1'h0, add_176053, array_index_175824[2:0]}) < $signed({1'h0, sel_176056}) ? {add_176053, array_index_175824[2:0]} : sel_176056;
  assign add_176160 = array_index_176025[11:1] + 11'h247;
  assign sel_176163 = $signed({1'h0, add_176058, array_index_175923[0]}) < $signed({1'h0, sel_176061}) ? {add_176058, array_index_175923[0]} : sel_176061;
  assign add_176165 = array_index_176028[11:1] + 11'h247;
  assign sel_176168 = $signed({1'h0, add_176063, array_index_175926[0]}) < $signed({1'h0, sel_176066}) ? {add_176063, array_index_175926[0]} : sel_176066;
  assign add_176193 = array_index_176127[11:0] + 12'h247;
  assign sel_176195 = $signed({1'h0, add_176091}) < $signed({1'h0, sel_176093}) ? add_176091 : sel_176093;
  assign add_176198 = array_index_176130[11:0] + 12'h247;
  assign sel_176200 = $signed({1'h0, add_176096}) < $signed({1'h0, sel_176098}) ? add_176096 : sel_176098;
  assign array_index_176229 = set1_unflattened[7'h23];
  assign array_index_176232 = set2_unflattened[7'h23];
  assign add_176236 = array_index_175821[11:1] + 11'h79d;
  assign sel_176238 = $signed({1'h0, add_176134, array_index_175719[0]}) < $signed({1'h0, sel_176136}) ? {add_176134, array_index_175719[0]} : sel_176136;
  assign add_176240 = array_index_175824[11:1] + 11'h79d;
  assign sel_176242 = $signed({1'h0, add_176138, array_index_175722[0]}) < $signed({1'h0, sel_176140}) ? {add_176138, array_index_175722[0]} : sel_176140;
  assign add_176244 = array_index_175923[11:1] + 11'h347;
  assign sel_176246 = $signed({1'h0, add_176142, array_index_175821[0]}) < $signed({1'h0, sel_176144}) ? {add_176142, array_index_175821[0]} : sel_176144;
  assign add_176248 = array_index_175926[11:1] + 11'h347;
  assign sel_176250 = $signed({1'h0, add_176146, array_index_175824[0]}) < $signed({1'h0, sel_176148}) ? {add_176146, array_index_175824[0]} : sel_176148;
  assign add_176252 = array_index_176025[11:3] + 9'h0bd;
  assign sel_176255 = $signed({1'h0, add_176150, array_index_175923[2:0]}) < $signed({1'h0, sel_176153}) ? {add_176150, array_index_175923[2:0]} : sel_176153;
  assign add_176257 = array_index_176028[11:3] + 9'h0bd;
  assign sel_176260 = $signed({1'h0, add_176155, array_index_175926[2:0]}) < $signed({1'h0, sel_176158}) ? {add_176155, array_index_175926[2:0]} : sel_176158;
  assign add_176262 = array_index_176127[11:1] + 11'h247;
  assign sel_176265 = $signed({1'h0, add_176160, array_index_176025[0]}) < $signed({1'h0, sel_176163}) ? {add_176160, array_index_176025[0]} : sel_176163;
  assign add_176267 = array_index_176130[11:1] + 11'h247;
  assign sel_176270 = $signed({1'h0, add_176165, array_index_176028[0]}) < $signed({1'h0, sel_176168}) ? {add_176165, array_index_176028[0]} : sel_176168;
  assign add_176295 = array_index_176229[11:0] + 12'h247;
  assign sel_176297 = $signed({1'h0, add_176193}) < $signed({1'h0, sel_176195}) ? add_176193 : sel_176195;
  assign add_176300 = array_index_176232[11:0] + 12'h247;
  assign sel_176302 = $signed({1'h0, add_176198}) < $signed({1'h0, sel_176200}) ? add_176198 : sel_176200;
  assign array_index_176331 = set1_unflattened[7'h24];
  assign array_index_176334 = set2_unflattened[7'h24];
  assign add_176338 = array_index_175923[11:1] + 11'h79d;
  assign sel_176340 = $signed({1'h0, add_176236, array_index_175821[0]}) < $signed({1'h0, sel_176238}) ? {add_176236, array_index_175821[0]} : sel_176238;
  assign add_176342 = array_index_175926[11:1] + 11'h79d;
  assign sel_176344 = $signed({1'h0, add_176240, array_index_175824[0]}) < $signed({1'h0, sel_176242}) ? {add_176240, array_index_175824[0]} : sel_176242;
  assign add_176346 = array_index_176025[11:1] + 11'h347;
  assign sel_176348 = $signed({1'h0, add_176244, array_index_175923[0]}) < $signed({1'h0, sel_176246}) ? {add_176244, array_index_175923[0]} : sel_176246;
  assign add_176350 = array_index_176028[11:1] + 11'h347;
  assign sel_176352 = $signed({1'h0, add_176248, array_index_175926[0]}) < $signed({1'h0, sel_176250}) ? {add_176248, array_index_175926[0]} : sel_176250;
  assign add_176354 = array_index_176127[11:3] + 9'h0bd;
  assign sel_176357 = $signed({1'h0, add_176252, array_index_176025[2:0]}) < $signed({1'h0, sel_176255}) ? {add_176252, array_index_176025[2:0]} : sel_176255;
  assign add_176359 = array_index_176130[11:3] + 9'h0bd;
  assign sel_176362 = $signed({1'h0, add_176257, array_index_176028[2:0]}) < $signed({1'h0, sel_176260}) ? {add_176257, array_index_176028[2:0]} : sel_176260;
  assign add_176364 = array_index_176229[11:1] + 11'h247;
  assign sel_176367 = $signed({1'h0, add_176262, array_index_176127[0]}) < $signed({1'h0, sel_176265}) ? {add_176262, array_index_176127[0]} : sel_176265;
  assign add_176369 = array_index_176232[11:1] + 11'h247;
  assign sel_176372 = $signed({1'h0, add_176267, array_index_176130[0]}) < $signed({1'h0, sel_176270}) ? {add_176267, array_index_176130[0]} : sel_176270;
  assign add_176397 = array_index_176331[11:0] + 12'h247;
  assign sel_176399 = $signed({1'h0, add_176295}) < $signed({1'h0, sel_176297}) ? add_176295 : sel_176297;
  assign add_176402 = array_index_176334[11:0] + 12'h247;
  assign sel_176404 = $signed({1'h0, add_176300}) < $signed({1'h0, sel_176302}) ? add_176300 : sel_176302;
  assign array_index_176433 = set1_unflattened[7'h25];
  assign array_index_176436 = set2_unflattened[7'h25];
  assign add_176440 = array_index_176025[11:1] + 11'h79d;
  assign sel_176442 = $signed({1'h0, add_176338, array_index_175923[0]}) < $signed({1'h0, sel_176340}) ? {add_176338, array_index_175923[0]} : sel_176340;
  assign add_176444 = array_index_176028[11:1] + 11'h79d;
  assign sel_176446 = $signed({1'h0, add_176342, array_index_175926[0]}) < $signed({1'h0, sel_176344}) ? {add_176342, array_index_175926[0]} : sel_176344;
  assign add_176448 = array_index_176127[11:1] + 11'h347;
  assign sel_176450 = $signed({1'h0, add_176346, array_index_176025[0]}) < $signed({1'h0, sel_176348}) ? {add_176346, array_index_176025[0]} : sel_176348;
  assign add_176452 = array_index_176130[11:1] + 11'h347;
  assign sel_176454 = $signed({1'h0, add_176350, array_index_176028[0]}) < $signed({1'h0, sel_176352}) ? {add_176350, array_index_176028[0]} : sel_176352;
  assign add_176456 = array_index_176229[11:3] + 9'h0bd;
  assign sel_176459 = $signed({1'h0, add_176354, array_index_176127[2:0]}) < $signed({1'h0, sel_176357}) ? {add_176354, array_index_176127[2:0]} : sel_176357;
  assign add_176461 = array_index_176232[11:3] + 9'h0bd;
  assign sel_176464 = $signed({1'h0, add_176359, array_index_176130[2:0]}) < $signed({1'h0, sel_176362}) ? {add_176359, array_index_176130[2:0]} : sel_176362;
  assign add_176466 = array_index_176331[11:1] + 11'h247;
  assign sel_176469 = $signed({1'h0, add_176364, array_index_176229[0]}) < $signed({1'h0, sel_176367}) ? {add_176364, array_index_176229[0]} : sel_176367;
  assign add_176471 = array_index_176334[11:1] + 11'h247;
  assign sel_176474 = $signed({1'h0, add_176369, array_index_176232[0]}) < $signed({1'h0, sel_176372}) ? {add_176369, array_index_176232[0]} : sel_176372;
  assign add_176499 = array_index_176433[11:0] + 12'h247;
  assign sel_176501 = $signed({1'h0, add_176397}) < $signed({1'h0, sel_176399}) ? add_176397 : sel_176399;
  assign add_176504 = array_index_176436[11:0] + 12'h247;
  assign sel_176506 = $signed({1'h0, add_176402}) < $signed({1'h0, sel_176404}) ? add_176402 : sel_176404;
  assign array_index_176535 = set1_unflattened[7'h26];
  assign array_index_176538 = set2_unflattened[7'h26];
  assign add_176542 = array_index_176127[11:1] + 11'h79d;
  assign sel_176544 = $signed({1'h0, add_176440, array_index_176025[0]}) < $signed({1'h0, sel_176442}) ? {add_176440, array_index_176025[0]} : sel_176442;
  assign add_176546 = array_index_176130[11:1] + 11'h79d;
  assign sel_176548 = $signed({1'h0, add_176444, array_index_176028[0]}) < $signed({1'h0, sel_176446}) ? {add_176444, array_index_176028[0]} : sel_176446;
  assign add_176550 = array_index_176229[11:1] + 11'h347;
  assign sel_176552 = $signed({1'h0, add_176448, array_index_176127[0]}) < $signed({1'h0, sel_176450}) ? {add_176448, array_index_176127[0]} : sel_176450;
  assign add_176554 = array_index_176232[11:1] + 11'h347;
  assign sel_176556 = $signed({1'h0, add_176452, array_index_176130[0]}) < $signed({1'h0, sel_176454}) ? {add_176452, array_index_176130[0]} : sel_176454;
  assign add_176558 = array_index_176331[11:3] + 9'h0bd;
  assign sel_176561 = $signed({1'h0, add_176456, array_index_176229[2:0]}) < $signed({1'h0, sel_176459}) ? {add_176456, array_index_176229[2:0]} : sel_176459;
  assign add_176563 = array_index_176334[11:3] + 9'h0bd;
  assign sel_176566 = $signed({1'h0, add_176461, array_index_176232[2:0]}) < $signed({1'h0, sel_176464}) ? {add_176461, array_index_176232[2:0]} : sel_176464;
  assign add_176568 = array_index_176433[11:1] + 11'h247;
  assign sel_176571 = $signed({1'h0, add_176466, array_index_176331[0]}) < $signed({1'h0, sel_176469}) ? {add_176466, array_index_176331[0]} : sel_176469;
  assign add_176573 = array_index_176436[11:1] + 11'h247;
  assign sel_176576 = $signed({1'h0, add_176471, array_index_176334[0]}) < $signed({1'h0, sel_176474}) ? {add_176471, array_index_176334[0]} : sel_176474;
  assign add_176601 = array_index_176535[11:0] + 12'h247;
  assign sel_176603 = $signed({1'h0, add_176499}) < $signed({1'h0, sel_176501}) ? add_176499 : sel_176501;
  assign add_176606 = array_index_176538[11:0] + 12'h247;
  assign sel_176608 = $signed({1'h0, add_176504}) < $signed({1'h0, sel_176506}) ? add_176504 : sel_176506;
  assign array_index_176637 = set1_unflattened[7'h27];
  assign array_index_176640 = set2_unflattened[7'h27];
  assign add_176644 = array_index_176229[11:1] + 11'h79d;
  assign sel_176646 = $signed({1'h0, add_176542, array_index_176127[0]}) < $signed({1'h0, sel_176544}) ? {add_176542, array_index_176127[0]} : sel_176544;
  assign add_176648 = array_index_176232[11:1] + 11'h79d;
  assign sel_176650 = $signed({1'h0, add_176546, array_index_176130[0]}) < $signed({1'h0, sel_176548}) ? {add_176546, array_index_176130[0]} : sel_176548;
  assign add_176652 = array_index_176331[11:1] + 11'h347;
  assign sel_176654 = $signed({1'h0, add_176550, array_index_176229[0]}) < $signed({1'h0, sel_176552}) ? {add_176550, array_index_176229[0]} : sel_176552;
  assign add_176656 = array_index_176334[11:1] + 11'h347;
  assign sel_176658 = $signed({1'h0, add_176554, array_index_176232[0]}) < $signed({1'h0, sel_176556}) ? {add_176554, array_index_176232[0]} : sel_176556;
  assign add_176660 = array_index_176433[11:3] + 9'h0bd;
  assign sel_176663 = $signed({1'h0, add_176558, array_index_176331[2:0]}) < $signed({1'h0, sel_176561}) ? {add_176558, array_index_176331[2:0]} : sel_176561;
  assign add_176665 = array_index_176436[11:3] + 9'h0bd;
  assign sel_176668 = $signed({1'h0, add_176563, array_index_176334[2:0]}) < $signed({1'h0, sel_176566}) ? {add_176563, array_index_176334[2:0]} : sel_176566;
  assign add_176670 = array_index_176535[11:1] + 11'h247;
  assign sel_176673 = $signed({1'h0, add_176568, array_index_176433[0]}) < $signed({1'h0, sel_176571}) ? {add_176568, array_index_176433[0]} : sel_176571;
  assign add_176675 = array_index_176538[11:1] + 11'h247;
  assign sel_176678 = $signed({1'h0, add_176573, array_index_176436[0]}) < $signed({1'h0, sel_176576}) ? {add_176573, array_index_176436[0]} : sel_176576;
  assign add_176703 = array_index_176637[11:0] + 12'h247;
  assign sel_176705 = $signed({1'h0, add_176601}) < $signed({1'h0, sel_176603}) ? add_176601 : sel_176603;
  assign add_176708 = array_index_176640[11:0] + 12'h247;
  assign sel_176710 = $signed({1'h0, add_176606}) < $signed({1'h0, sel_176608}) ? add_176606 : sel_176608;
  assign array_index_176739 = set1_unflattened[7'h28];
  assign array_index_176742 = set2_unflattened[7'h28];
  assign add_176746 = array_index_176331[11:1] + 11'h79d;
  assign sel_176748 = $signed({1'h0, add_176644, array_index_176229[0]}) < $signed({1'h0, sel_176646}) ? {add_176644, array_index_176229[0]} : sel_176646;
  assign add_176750 = array_index_176334[11:1] + 11'h79d;
  assign sel_176752 = $signed({1'h0, add_176648, array_index_176232[0]}) < $signed({1'h0, sel_176650}) ? {add_176648, array_index_176232[0]} : sel_176650;
  assign add_176754 = array_index_176433[11:1] + 11'h347;
  assign sel_176756 = $signed({1'h0, add_176652, array_index_176331[0]}) < $signed({1'h0, sel_176654}) ? {add_176652, array_index_176331[0]} : sel_176654;
  assign add_176758 = array_index_176436[11:1] + 11'h347;
  assign sel_176760 = $signed({1'h0, add_176656, array_index_176334[0]}) < $signed({1'h0, sel_176658}) ? {add_176656, array_index_176334[0]} : sel_176658;
  assign add_176762 = array_index_176535[11:3] + 9'h0bd;
  assign sel_176765 = $signed({1'h0, add_176660, array_index_176433[2:0]}) < $signed({1'h0, sel_176663}) ? {add_176660, array_index_176433[2:0]} : sel_176663;
  assign add_176767 = array_index_176538[11:3] + 9'h0bd;
  assign sel_176770 = $signed({1'h0, add_176665, array_index_176436[2:0]}) < $signed({1'h0, sel_176668}) ? {add_176665, array_index_176436[2:0]} : sel_176668;
  assign add_176772 = array_index_176637[11:1] + 11'h247;
  assign sel_176775 = $signed({1'h0, add_176670, array_index_176535[0]}) < $signed({1'h0, sel_176673}) ? {add_176670, array_index_176535[0]} : sel_176673;
  assign add_176777 = array_index_176640[11:1] + 11'h247;
  assign sel_176780 = $signed({1'h0, add_176675, array_index_176538[0]}) < $signed({1'h0, sel_176678}) ? {add_176675, array_index_176538[0]} : sel_176678;
  assign add_176805 = array_index_176739[11:0] + 12'h247;
  assign sel_176807 = $signed({1'h0, add_176703}) < $signed({1'h0, sel_176705}) ? add_176703 : sel_176705;
  assign add_176810 = array_index_176742[11:0] + 12'h247;
  assign sel_176812 = $signed({1'h0, add_176708}) < $signed({1'h0, sel_176710}) ? add_176708 : sel_176710;
  assign array_index_176841 = set1_unflattened[7'h29];
  assign array_index_176844 = set2_unflattened[7'h29];
  assign add_176848 = array_index_176433[11:1] + 11'h79d;
  assign sel_176850 = $signed({1'h0, add_176746, array_index_176331[0]}) < $signed({1'h0, sel_176748}) ? {add_176746, array_index_176331[0]} : sel_176748;
  assign add_176852 = array_index_176436[11:1] + 11'h79d;
  assign sel_176854 = $signed({1'h0, add_176750, array_index_176334[0]}) < $signed({1'h0, sel_176752}) ? {add_176750, array_index_176334[0]} : sel_176752;
  assign add_176856 = array_index_176535[11:1] + 11'h347;
  assign sel_176858 = $signed({1'h0, add_176754, array_index_176433[0]}) < $signed({1'h0, sel_176756}) ? {add_176754, array_index_176433[0]} : sel_176756;
  assign add_176860 = array_index_176538[11:1] + 11'h347;
  assign sel_176862 = $signed({1'h0, add_176758, array_index_176436[0]}) < $signed({1'h0, sel_176760}) ? {add_176758, array_index_176436[0]} : sel_176760;
  assign add_176864 = array_index_176637[11:3] + 9'h0bd;
  assign sel_176867 = $signed({1'h0, add_176762, array_index_176535[2:0]}) < $signed({1'h0, sel_176765}) ? {add_176762, array_index_176535[2:0]} : sel_176765;
  assign add_176869 = array_index_176640[11:3] + 9'h0bd;
  assign sel_176872 = $signed({1'h0, add_176767, array_index_176538[2:0]}) < $signed({1'h0, sel_176770}) ? {add_176767, array_index_176538[2:0]} : sel_176770;
  assign add_176874 = array_index_176739[11:1] + 11'h247;
  assign sel_176877 = $signed({1'h0, add_176772, array_index_176637[0]}) < $signed({1'h0, sel_176775}) ? {add_176772, array_index_176637[0]} : sel_176775;
  assign add_176879 = array_index_176742[11:1] + 11'h247;
  assign sel_176882 = $signed({1'h0, add_176777, array_index_176640[0]}) < $signed({1'h0, sel_176780}) ? {add_176777, array_index_176640[0]} : sel_176780;
  assign add_176907 = array_index_176841[11:0] + 12'h247;
  assign sel_176909 = $signed({1'h0, add_176805}) < $signed({1'h0, sel_176807}) ? add_176805 : sel_176807;
  assign add_176912 = array_index_176844[11:0] + 12'h247;
  assign sel_176914 = $signed({1'h0, add_176810}) < $signed({1'h0, sel_176812}) ? add_176810 : sel_176812;
  assign array_index_176943 = set1_unflattened[7'h2a];
  assign array_index_176946 = set2_unflattened[7'h2a];
  assign add_176950 = array_index_176535[11:1] + 11'h79d;
  assign sel_176952 = $signed({1'h0, add_176848, array_index_176433[0]}) < $signed({1'h0, sel_176850}) ? {add_176848, array_index_176433[0]} : sel_176850;
  assign add_176954 = array_index_176538[11:1] + 11'h79d;
  assign sel_176956 = $signed({1'h0, add_176852, array_index_176436[0]}) < $signed({1'h0, sel_176854}) ? {add_176852, array_index_176436[0]} : sel_176854;
  assign add_176958 = array_index_176637[11:1] + 11'h347;
  assign sel_176960 = $signed({1'h0, add_176856, array_index_176535[0]}) < $signed({1'h0, sel_176858}) ? {add_176856, array_index_176535[0]} : sel_176858;
  assign add_176962 = array_index_176640[11:1] + 11'h347;
  assign sel_176964 = $signed({1'h0, add_176860, array_index_176538[0]}) < $signed({1'h0, sel_176862}) ? {add_176860, array_index_176538[0]} : sel_176862;
  assign add_176966 = array_index_176739[11:3] + 9'h0bd;
  assign sel_176969 = $signed({1'h0, add_176864, array_index_176637[2:0]}) < $signed({1'h0, sel_176867}) ? {add_176864, array_index_176637[2:0]} : sel_176867;
  assign add_176971 = array_index_176742[11:3] + 9'h0bd;
  assign sel_176974 = $signed({1'h0, add_176869, array_index_176640[2:0]}) < $signed({1'h0, sel_176872}) ? {add_176869, array_index_176640[2:0]} : sel_176872;
  assign add_176976 = array_index_176841[11:1] + 11'h247;
  assign sel_176979 = $signed({1'h0, add_176874, array_index_176739[0]}) < $signed({1'h0, sel_176877}) ? {add_176874, array_index_176739[0]} : sel_176877;
  assign add_176981 = array_index_176844[11:1] + 11'h247;
  assign sel_176984 = $signed({1'h0, add_176879, array_index_176742[0]}) < $signed({1'h0, sel_176882}) ? {add_176879, array_index_176742[0]} : sel_176882;
  assign add_177009 = array_index_176943[11:0] + 12'h247;
  assign sel_177011 = $signed({1'h0, add_176907}) < $signed({1'h0, sel_176909}) ? add_176907 : sel_176909;
  assign add_177014 = array_index_176946[11:0] + 12'h247;
  assign sel_177016 = $signed({1'h0, add_176912}) < $signed({1'h0, sel_176914}) ? add_176912 : sel_176914;
  assign array_index_177045 = set1_unflattened[7'h2b];
  assign array_index_177048 = set2_unflattened[7'h2b];
  assign add_177052 = array_index_176637[11:1] + 11'h79d;
  assign sel_177054 = $signed({1'h0, add_176950, array_index_176535[0]}) < $signed({1'h0, sel_176952}) ? {add_176950, array_index_176535[0]} : sel_176952;
  assign add_177056 = array_index_176640[11:1] + 11'h79d;
  assign sel_177058 = $signed({1'h0, add_176954, array_index_176538[0]}) < $signed({1'h0, sel_176956}) ? {add_176954, array_index_176538[0]} : sel_176956;
  assign add_177060 = array_index_176739[11:1] + 11'h347;
  assign sel_177062 = $signed({1'h0, add_176958, array_index_176637[0]}) < $signed({1'h0, sel_176960}) ? {add_176958, array_index_176637[0]} : sel_176960;
  assign add_177064 = array_index_176742[11:1] + 11'h347;
  assign sel_177066 = $signed({1'h0, add_176962, array_index_176640[0]}) < $signed({1'h0, sel_176964}) ? {add_176962, array_index_176640[0]} : sel_176964;
  assign add_177068 = array_index_176841[11:3] + 9'h0bd;
  assign sel_177071 = $signed({1'h0, add_176966, array_index_176739[2:0]}) < $signed({1'h0, sel_176969}) ? {add_176966, array_index_176739[2:0]} : sel_176969;
  assign add_177073 = array_index_176844[11:3] + 9'h0bd;
  assign sel_177076 = $signed({1'h0, add_176971, array_index_176742[2:0]}) < $signed({1'h0, sel_176974}) ? {add_176971, array_index_176742[2:0]} : sel_176974;
  assign add_177078 = array_index_176943[11:1] + 11'h247;
  assign sel_177081 = $signed({1'h0, add_176976, array_index_176841[0]}) < $signed({1'h0, sel_176979}) ? {add_176976, array_index_176841[0]} : sel_176979;
  assign add_177083 = array_index_176946[11:1] + 11'h247;
  assign sel_177086 = $signed({1'h0, add_176981, array_index_176844[0]}) < $signed({1'h0, sel_176984}) ? {add_176981, array_index_176844[0]} : sel_176984;
  assign add_177111 = array_index_177045[11:0] + 12'h247;
  assign sel_177113 = $signed({1'h0, add_177009}) < $signed({1'h0, sel_177011}) ? add_177009 : sel_177011;
  assign add_177116 = array_index_177048[11:0] + 12'h247;
  assign sel_177118 = $signed({1'h0, add_177014}) < $signed({1'h0, sel_177016}) ? add_177014 : sel_177016;
  assign array_index_177147 = set1_unflattened[7'h2c];
  assign array_index_177150 = set2_unflattened[7'h2c];
  assign add_177154 = array_index_176739[11:1] + 11'h79d;
  assign sel_177156 = $signed({1'h0, add_177052, array_index_176637[0]}) < $signed({1'h0, sel_177054}) ? {add_177052, array_index_176637[0]} : sel_177054;
  assign add_177158 = array_index_176742[11:1] + 11'h79d;
  assign sel_177160 = $signed({1'h0, add_177056, array_index_176640[0]}) < $signed({1'h0, sel_177058}) ? {add_177056, array_index_176640[0]} : sel_177058;
  assign add_177162 = array_index_176841[11:1] + 11'h347;
  assign sel_177164 = $signed({1'h0, add_177060, array_index_176739[0]}) < $signed({1'h0, sel_177062}) ? {add_177060, array_index_176739[0]} : sel_177062;
  assign add_177166 = array_index_176844[11:1] + 11'h347;
  assign sel_177168 = $signed({1'h0, add_177064, array_index_176742[0]}) < $signed({1'h0, sel_177066}) ? {add_177064, array_index_176742[0]} : sel_177066;
  assign add_177170 = array_index_176943[11:3] + 9'h0bd;
  assign sel_177173 = $signed({1'h0, add_177068, array_index_176841[2:0]}) < $signed({1'h0, sel_177071}) ? {add_177068, array_index_176841[2:0]} : sel_177071;
  assign add_177175 = array_index_176946[11:3] + 9'h0bd;
  assign sel_177178 = $signed({1'h0, add_177073, array_index_176844[2:0]}) < $signed({1'h0, sel_177076}) ? {add_177073, array_index_176844[2:0]} : sel_177076;
  assign add_177180 = array_index_177045[11:1] + 11'h247;
  assign sel_177183 = $signed({1'h0, add_177078, array_index_176943[0]}) < $signed({1'h0, sel_177081}) ? {add_177078, array_index_176943[0]} : sel_177081;
  assign add_177185 = array_index_177048[11:1] + 11'h247;
  assign sel_177188 = $signed({1'h0, add_177083, array_index_176946[0]}) < $signed({1'h0, sel_177086}) ? {add_177083, array_index_176946[0]} : sel_177086;
  assign add_177213 = array_index_177147[11:0] + 12'h247;
  assign sel_177215 = $signed({1'h0, add_177111}) < $signed({1'h0, sel_177113}) ? add_177111 : sel_177113;
  assign add_177218 = array_index_177150[11:0] + 12'h247;
  assign sel_177220 = $signed({1'h0, add_177116}) < $signed({1'h0, sel_177118}) ? add_177116 : sel_177118;
  assign array_index_177249 = set1_unflattened[7'h2d];
  assign array_index_177252 = set2_unflattened[7'h2d];
  assign add_177256 = array_index_176841[11:1] + 11'h79d;
  assign sel_177258 = $signed({1'h0, add_177154, array_index_176739[0]}) < $signed({1'h0, sel_177156}) ? {add_177154, array_index_176739[0]} : sel_177156;
  assign add_177260 = array_index_176844[11:1] + 11'h79d;
  assign sel_177262 = $signed({1'h0, add_177158, array_index_176742[0]}) < $signed({1'h0, sel_177160}) ? {add_177158, array_index_176742[0]} : sel_177160;
  assign add_177264 = array_index_176943[11:1] + 11'h347;
  assign sel_177266 = $signed({1'h0, add_177162, array_index_176841[0]}) < $signed({1'h0, sel_177164}) ? {add_177162, array_index_176841[0]} : sel_177164;
  assign add_177268 = array_index_176946[11:1] + 11'h347;
  assign sel_177270 = $signed({1'h0, add_177166, array_index_176844[0]}) < $signed({1'h0, sel_177168}) ? {add_177166, array_index_176844[0]} : sel_177168;
  assign add_177272 = array_index_177045[11:3] + 9'h0bd;
  assign sel_177275 = $signed({1'h0, add_177170, array_index_176943[2:0]}) < $signed({1'h0, sel_177173}) ? {add_177170, array_index_176943[2:0]} : sel_177173;
  assign add_177277 = array_index_177048[11:3] + 9'h0bd;
  assign sel_177280 = $signed({1'h0, add_177175, array_index_176946[2:0]}) < $signed({1'h0, sel_177178}) ? {add_177175, array_index_176946[2:0]} : sel_177178;
  assign add_177282 = array_index_177147[11:1] + 11'h247;
  assign sel_177285 = $signed({1'h0, add_177180, array_index_177045[0]}) < $signed({1'h0, sel_177183}) ? {add_177180, array_index_177045[0]} : sel_177183;
  assign add_177287 = array_index_177150[11:1] + 11'h247;
  assign sel_177290 = $signed({1'h0, add_177185, array_index_177048[0]}) < $signed({1'h0, sel_177188}) ? {add_177185, array_index_177048[0]} : sel_177188;
  assign add_177315 = array_index_177249[11:0] + 12'h247;
  assign sel_177317 = $signed({1'h0, add_177213}) < $signed({1'h0, sel_177215}) ? add_177213 : sel_177215;
  assign add_177320 = array_index_177252[11:0] + 12'h247;
  assign sel_177322 = $signed({1'h0, add_177218}) < $signed({1'h0, sel_177220}) ? add_177218 : sel_177220;
  assign array_index_177351 = set1_unflattened[7'h2e];
  assign array_index_177354 = set2_unflattened[7'h2e];
  assign add_177358 = array_index_176943[11:1] + 11'h79d;
  assign sel_177360 = $signed({1'h0, add_177256, array_index_176841[0]}) < $signed({1'h0, sel_177258}) ? {add_177256, array_index_176841[0]} : sel_177258;
  assign add_177362 = array_index_176946[11:1] + 11'h79d;
  assign sel_177364 = $signed({1'h0, add_177260, array_index_176844[0]}) < $signed({1'h0, sel_177262}) ? {add_177260, array_index_176844[0]} : sel_177262;
  assign add_177366 = array_index_177045[11:1] + 11'h347;
  assign sel_177368 = $signed({1'h0, add_177264, array_index_176943[0]}) < $signed({1'h0, sel_177266}) ? {add_177264, array_index_176943[0]} : sel_177266;
  assign add_177370 = array_index_177048[11:1] + 11'h347;
  assign sel_177372 = $signed({1'h0, add_177268, array_index_176946[0]}) < $signed({1'h0, sel_177270}) ? {add_177268, array_index_176946[0]} : sel_177270;
  assign add_177374 = array_index_177147[11:3] + 9'h0bd;
  assign sel_177377 = $signed({1'h0, add_177272, array_index_177045[2:0]}) < $signed({1'h0, sel_177275}) ? {add_177272, array_index_177045[2:0]} : sel_177275;
  assign add_177379 = array_index_177150[11:3] + 9'h0bd;
  assign sel_177382 = $signed({1'h0, add_177277, array_index_177048[2:0]}) < $signed({1'h0, sel_177280}) ? {add_177277, array_index_177048[2:0]} : sel_177280;
  assign add_177384 = array_index_177249[11:1] + 11'h247;
  assign sel_177387 = $signed({1'h0, add_177282, array_index_177147[0]}) < $signed({1'h0, sel_177285}) ? {add_177282, array_index_177147[0]} : sel_177285;
  assign add_177389 = array_index_177252[11:1] + 11'h247;
  assign sel_177392 = $signed({1'h0, add_177287, array_index_177150[0]}) < $signed({1'h0, sel_177290}) ? {add_177287, array_index_177150[0]} : sel_177290;
  assign add_177417 = array_index_177351[11:0] + 12'h247;
  assign sel_177419 = $signed({1'h0, add_177315}) < $signed({1'h0, sel_177317}) ? add_177315 : sel_177317;
  assign add_177422 = array_index_177354[11:0] + 12'h247;
  assign sel_177424 = $signed({1'h0, add_177320}) < $signed({1'h0, sel_177322}) ? add_177320 : sel_177322;
  assign array_index_177453 = set1_unflattened[7'h2f];
  assign array_index_177456 = set2_unflattened[7'h2f];
  assign add_177460 = array_index_177045[11:1] + 11'h79d;
  assign sel_177462 = $signed({1'h0, add_177358, array_index_176943[0]}) < $signed({1'h0, sel_177360}) ? {add_177358, array_index_176943[0]} : sel_177360;
  assign add_177464 = array_index_177048[11:1] + 11'h79d;
  assign sel_177466 = $signed({1'h0, add_177362, array_index_176946[0]}) < $signed({1'h0, sel_177364}) ? {add_177362, array_index_176946[0]} : sel_177364;
  assign add_177468 = array_index_177147[11:1] + 11'h347;
  assign sel_177470 = $signed({1'h0, add_177366, array_index_177045[0]}) < $signed({1'h0, sel_177368}) ? {add_177366, array_index_177045[0]} : sel_177368;
  assign add_177472 = array_index_177150[11:1] + 11'h347;
  assign sel_177474 = $signed({1'h0, add_177370, array_index_177048[0]}) < $signed({1'h0, sel_177372}) ? {add_177370, array_index_177048[0]} : sel_177372;
  assign add_177476 = array_index_177249[11:3] + 9'h0bd;
  assign sel_177479 = $signed({1'h0, add_177374, array_index_177147[2:0]}) < $signed({1'h0, sel_177377}) ? {add_177374, array_index_177147[2:0]} : sel_177377;
  assign add_177481 = array_index_177252[11:3] + 9'h0bd;
  assign sel_177484 = $signed({1'h0, add_177379, array_index_177150[2:0]}) < $signed({1'h0, sel_177382}) ? {add_177379, array_index_177150[2:0]} : sel_177382;
  assign add_177486 = array_index_177351[11:1] + 11'h247;
  assign sel_177489 = $signed({1'h0, add_177384, array_index_177249[0]}) < $signed({1'h0, sel_177387}) ? {add_177384, array_index_177249[0]} : sel_177387;
  assign add_177491 = array_index_177354[11:1] + 11'h247;
  assign sel_177494 = $signed({1'h0, add_177389, array_index_177252[0]}) < $signed({1'h0, sel_177392}) ? {add_177389, array_index_177252[0]} : sel_177392;
  assign add_177519 = array_index_177453[11:0] + 12'h247;
  assign sel_177521 = $signed({1'h0, add_177417}) < $signed({1'h0, sel_177419}) ? add_177417 : sel_177419;
  assign add_177524 = array_index_177456[11:0] + 12'h247;
  assign sel_177526 = $signed({1'h0, add_177422}) < $signed({1'h0, sel_177424}) ? add_177422 : sel_177424;
  assign array_index_177555 = set1_unflattened[7'h30];
  assign array_index_177558 = set2_unflattened[7'h30];
  assign add_177562 = array_index_177147[11:1] + 11'h79d;
  assign sel_177564 = $signed({1'h0, add_177460, array_index_177045[0]}) < $signed({1'h0, sel_177462}) ? {add_177460, array_index_177045[0]} : sel_177462;
  assign add_177566 = array_index_177150[11:1] + 11'h79d;
  assign sel_177568 = $signed({1'h0, add_177464, array_index_177048[0]}) < $signed({1'h0, sel_177466}) ? {add_177464, array_index_177048[0]} : sel_177466;
  assign add_177570 = array_index_177249[11:1] + 11'h347;
  assign sel_177572 = $signed({1'h0, add_177468, array_index_177147[0]}) < $signed({1'h0, sel_177470}) ? {add_177468, array_index_177147[0]} : sel_177470;
  assign add_177574 = array_index_177252[11:1] + 11'h347;
  assign sel_177576 = $signed({1'h0, add_177472, array_index_177150[0]}) < $signed({1'h0, sel_177474}) ? {add_177472, array_index_177150[0]} : sel_177474;
  assign add_177578 = array_index_177351[11:3] + 9'h0bd;
  assign sel_177581 = $signed({1'h0, add_177476, array_index_177249[2:0]}) < $signed({1'h0, sel_177479}) ? {add_177476, array_index_177249[2:0]} : sel_177479;
  assign add_177583 = array_index_177354[11:3] + 9'h0bd;
  assign sel_177586 = $signed({1'h0, add_177481, array_index_177252[2:0]}) < $signed({1'h0, sel_177484}) ? {add_177481, array_index_177252[2:0]} : sel_177484;
  assign add_177588 = array_index_177453[11:1] + 11'h247;
  assign sel_177591 = $signed({1'h0, add_177486, array_index_177351[0]}) < $signed({1'h0, sel_177489}) ? {add_177486, array_index_177351[0]} : sel_177489;
  assign add_177593 = array_index_177456[11:1] + 11'h247;
  assign sel_177596 = $signed({1'h0, add_177491, array_index_177354[0]}) < $signed({1'h0, sel_177494}) ? {add_177491, array_index_177354[0]} : sel_177494;
  assign add_177621 = array_index_177555[11:0] + 12'h247;
  assign sel_177623 = $signed({1'h0, add_177519}) < $signed({1'h0, sel_177521}) ? add_177519 : sel_177521;
  assign add_177626 = array_index_177558[11:0] + 12'h247;
  assign sel_177628 = $signed({1'h0, add_177524}) < $signed({1'h0, sel_177526}) ? add_177524 : sel_177526;
  assign array_index_177657 = set1_unflattened[7'h31];
  assign array_index_177660 = set2_unflattened[7'h31];
  assign add_177664 = array_index_177249[11:1] + 11'h79d;
  assign sel_177666 = $signed({1'h0, add_177562, array_index_177147[0]}) < $signed({1'h0, sel_177564}) ? {add_177562, array_index_177147[0]} : sel_177564;
  assign add_177668 = array_index_177252[11:1] + 11'h79d;
  assign sel_177670 = $signed({1'h0, add_177566, array_index_177150[0]}) < $signed({1'h0, sel_177568}) ? {add_177566, array_index_177150[0]} : sel_177568;
  assign add_177672 = array_index_177351[11:1] + 11'h347;
  assign sel_177674 = $signed({1'h0, add_177570, array_index_177249[0]}) < $signed({1'h0, sel_177572}) ? {add_177570, array_index_177249[0]} : sel_177572;
  assign add_177676 = array_index_177354[11:1] + 11'h347;
  assign sel_177678 = $signed({1'h0, add_177574, array_index_177252[0]}) < $signed({1'h0, sel_177576}) ? {add_177574, array_index_177252[0]} : sel_177576;
  assign add_177680 = array_index_177453[11:3] + 9'h0bd;
  assign sel_177683 = $signed({1'h0, add_177578, array_index_177351[2:0]}) < $signed({1'h0, sel_177581}) ? {add_177578, array_index_177351[2:0]} : sel_177581;
  assign add_177685 = array_index_177456[11:3] + 9'h0bd;
  assign sel_177688 = $signed({1'h0, add_177583, array_index_177354[2:0]}) < $signed({1'h0, sel_177586}) ? {add_177583, array_index_177354[2:0]} : sel_177586;
  assign add_177690 = array_index_177555[11:1] + 11'h247;
  assign sel_177693 = $signed({1'h0, add_177588, array_index_177453[0]}) < $signed({1'h0, sel_177591}) ? {add_177588, array_index_177453[0]} : sel_177591;
  assign add_177695 = array_index_177558[11:1] + 11'h247;
  assign sel_177698 = $signed({1'h0, add_177593, array_index_177456[0]}) < $signed({1'h0, sel_177596}) ? {add_177593, array_index_177456[0]} : sel_177596;
  assign add_177723 = array_index_177657[11:0] + 12'h247;
  assign sel_177725 = $signed({1'h0, add_177621}) < $signed({1'h0, sel_177623}) ? add_177621 : sel_177623;
  assign add_177728 = array_index_177660[11:0] + 12'h247;
  assign sel_177730 = $signed({1'h0, add_177626}) < $signed({1'h0, sel_177628}) ? add_177626 : sel_177628;
  assign array_index_177759 = set1_unflattened[7'h32];
  assign array_index_177762 = set2_unflattened[7'h32];
  assign add_177766 = array_index_177351[11:1] + 11'h79d;
  assign sel_177768 = $signed({1'h0, add_177664, array_index_177249[0]}) < $signed({1'h0, sel_177666}) ? {add_177664, array_index_177249[0]} : sel_177666;
  assign add_177770 = array_index_177354[11:1] + 11'h79d;
  assign sel_177772 = $signed({1'h0, add_177668, array_index_177252[0]}) < $signed({1'h0, sel_177670}) ? {add_177668, array_index_177252[0]} : sel_177670;
  assign add_177774 = array_index_177453[11:1] + 11'h347;
  assign sel_177776 = $signed({1'h0, add_177672, array_index_177351[0]}) < $signed({1'h0, sel_177674}) ? {add_177672, array_index_177351[0]} : sel_177674;
  assign add_177778 = array_index_177456[11:1] + 11'h347;
  assign sel_177780 = $signed({1'h0, add_177676, array_index_177354[0]}) < $signed({1'h0, sel_177678}) ? {add_177676, array_index_177354[0]} : sel_177678;
  assign add_177782 = array_index_177555[11:3] + 9'h0bd;
  assign sel_177785 = $signed({1'h0, add_177680, array_index_177453[2:0]}) < $signed({1'h0, sel_177683}) ? {add_177680, array_index_177453[2:0]} : sel_177683;
  assign add_177787 = array_index_177558[11:3] + 9'h0bd;
  assign sel_177790 = $signed({1'h0, add_177685, array_index_177456[2:0]}) < $signed({1'h0, sel_177688}) ? {add_177685, array_index_177456[2:0]} : sel_177688;
  assign add_177792 = array_index_177657[11:1] + 11'h247;
  assign sel_177795 = $signed({1'h0, add_177690, array_index_177555[0]}) < $signed({1'h0, sel_177693}) ? {add_177690, array_index_177555[0]} : sel_177693;
  assign add_177797 = array_index_177660[11:1] + 11'h247;
  assign sel_177800 = $signed({1'h0, add_177695, array_index_177558[0]}) < $signed({1'h0, sel_177698}) ? {add_177695, array_index_177558[0]} : sel_177698;
  assign add_177825 = array_index_177759[11:0] + 12'h247;
  assign sel_177827 = $signed({1'h0, add_177723}) < $signed({1'h0, sel_177725}) ? add_177723 : sel_177725;
  assign add_177830 = array_index_177762[11:0] + 12'h247;
  assign sel_177832 = $signed({1'h0, add_177728}) < $signed({1'h0, sel_177730}) ? add_177728 : sel_177730;
  assign array_index_177861 = set1_unflattened[7'h33];
  assign array_index_177864 = set2_unflattened[7'h33];
  assign add_177868 = array_index_177453[11:1] + 11'h79d;
  assign sel_177870 = $signed({1'h0, add_177766, array_index_177351[0]}) < $signed({1'h0, sel_177768}) ? {add_177766, array_index_177351[0]} : sel_177768;
  assign add_177872 = array_index_177456[11:1] + 11'h79d;
  assign sel_177874 = $signed({1'h0, add_177770, array_index_177354[0]}) < $signed({1'h0, sel_177772}) ? {add_177770, array_index_177354[0]} : sel_177772;
  assign add_177876 = array_index_177555[11:1] + 11'h347;
  assign sel_177878 = $signed({1'h0, add_177774, array_index_177453[0]}) < $signed({1'h0, sel_177776}) ? {add_177774, array_index_177453[0]} : sel_177776;
  assign add_177880 = array_index_177558[11:1] + 11'h347;
  assign sel_177882 = $signed({1'h0, add_177778, array_index_177456[0]}) < $signed({1'h0, sel_177780}) ? {add_177778, array_index_177456[0]} : sel_177780;
  assign add_177884 = array_index_177657[11:3] + 9'h0bd;
  assign sel_177887 = $signed({1'h0, add_177782, array_index_177555[2:0]}) < $signed({1'h0, sel_177785}) ? {add_177782, array_index_177555[2:0]} : sel_177785;
  assign add_177889 = array_index_177660[11:3] + 9'h0bd;
  assign sel_177892 = $signed({1'h0, add_177787, array_index_177558[2:0]}) < $signed({1'h0, sel_177790}) ? {add_177787, array_index_177558[2:0]} : sel_177790;
  assign add_177894 = array_index_177759[11:1] + 11'h247;
  assign sel_177897 = $signed({1'h0, add_177792, array_index_177657[0]}) < $signed({1'h0, sel_177795}) ? {add_177792, array_index_177657[0]} : sel_177795;
  assign add_177899 = array_index_177762[11:1] + 11'h247;
  assign sel_177902 = $signed({1'h0, add_177797, array_index_177660[0]}) < $signed({1'h0, sel_177800}) ? {add_177797, array_index_177660[0]} : sel_177800;
  assign add_177927 = array_index_177861[11:0] + 12'h247;
  assign sel_177929 = $signed({1'h0, add_177825}) < $signed({1'h0, sel_177827}) ? add_177825 : sel_177827;
  assign add_177932 = array_index_177864[11:0] + 12'h247;
  assign sel_177934 = $signed({1'h0, add_177830}) < $signed({1'h0, sel_177832}) ? add_177830 : sel_177832;
  assign array_index_177963 = set1_unflattened[7'h34];
  assign array_index_177966 = set2_unflattened[7'h34];
  assign add_177970 = array_index_177555[11:1] + 11'h79d;
  assign sel_177972 = $signed({1'h0, add_177868, array_index_177453[0]}) < $signed({1'h0, sel_177870}) ? {add_177868, array_index_177453[0]} : sel_177870;
  assign add_177974 = array_index_177558[11:1] + 11'h79d;
  assign sel_177976 = $signed({1'h0, add_177872, array_index_177456[0]}) < $signed({1'h0, sel_177874}) ? {add_177872, array_index_177456[0]} : sel_177874;
  assign add_177978 = array_index_177657[11:1] + 11'h347;
  assign sel_177980 = $signed({1'h0, add_177876, array_index_177555[0]}) < $signed({1'h0, sel_177878}) ? {add_177876, array_index_177555[0]} : sel_177878;
  assign add_177982 = array_index_177660[11:1] + 11'h347;
  assign sel_177984 = $signed({1'h0, add_177880, array_index_177558[0]}) < $signed({1'h0, sel_177882}) ? {add_177880, array_index_177558[0]} : sel_177882;
  assign add_177986 = array_index_177759[11:3] + 9'h0bd;
  assign sel_177989 = $signed({1'h0, add_177884, array_index_177657[2:0]}) < $signed({1'h0, sel_177887}) ? {add_177884, array_index_177657[2:0]} : sel_177887;
  assign add_177991 = array_index_177762[11:3] + 9'h0bd;
  assign sel_177994 = $signed({1'h0, add_177889, array_index_177660[2:0]}) < $signed({1'h0, sel_177892}) ? {add_177889, array_index_177660[2:0]} : sel_177892;
  assign add_177996 = array_index_177861[11:1] + 11'h247;
  assign sel_177999 = $signed({1'h0, add_177894, array_index_177759[0]}) < $signed({1'h0, sel_177897}) ? {add_177894, array_index_177759[0]} : sel_177897;
  assign add_178001 = array_index_177864[11:1] + 11'h247;
  assign sel_178004 = $signed({1'h0, add_177899, array_index_177762[0]}) < $signed({1'h0, sel_177902}) ? {add_177899, array_index_177762[0]} : sel_177902;
  assign add_178029 = array_index_177963[11:0] + 12'h247;
  assign sel_178031 = $signed({1'h0, add_177927}) < $signed({1'h0, sel_177929}) ? add_177927 : sel_177929;
  assign add_178034 = array_index_177966[11:0] + 12'h247;
  assign sel_178036 = $signed({1'h0, add_177932}) < $signed({1'h0, sel_177934}) ? add_177932 : sel_177934;
  assign array_index_178065 = set1_unflattened[7'h35];
  assign array_index_178068 = set2_unflattened[7'h35];
  assign add_178072 = array_index_177657[11:1] + 11'h79d;
  assign sel_178074 = $signed({1'h0, add_177970, array_index_177555[0]}) < $signed({1'h0, sel_177972}) ? {add_177970, array_index_177555[0]} : sel_177972;
  assign add_178076 = array_index_177660[11:1] + 11'h79d;
  assign sel_178078 = $signed({1'h0, add_177974, array_index_177558[0]}) < $signed({1'h0, sel_177976}) ? {add_177974, array_index_177558[0]} : sel_177976;
  assign add_178080 = array_index_177759[11:1] + 11'h347;
  assign sel_178082 = $signed({1'h0, add_177978, array_index_177657[0]}) < $signed({1'h0, sel_177980}) ? {add_177978, array_index_177657[0]} : sel_177980;
  assign add_178084 = array_index_177762[11:1] + 11'h347;
  assign sel_178086 = $signed({1'h0, add_177982, array_index_177660[0]}) < $signed({1'h0, sel_177984}) ? {add_177982, array_index_177660[0]} : sel_177984;
  assign add_178088 = array_index_177861[11:3] + 9'h0bd;
  assign sel_178091 = $signed({1'h0, add_177986, array_index_177759[2:0]}) < $signed({1'h0, sel_177989}) ? {add_177986, array_index_177759[2:0]} : sel_177989;
  assign add_178093 = array_index_177864[11:3] + 9'h0bd;
  assign sel_178096 = $signed({1'h0, add_177991, array_index_177762[2:0]}) < $signed({1'h0, sel_177994}) ? {add_177991, array_index_177762[2:0]} : sel_177994;
  assign add_178098 = array_index_177963[11:1] + 11'h247;
  assign sel_178101 = $signed({1'h0, add_177996, array_index_177861[0]}) < $signed({1'h0, sel_177999}) ? {add_177996, array_index_177861[0]} : sel_177999;
  assign add_178103 = array_index_177966[11:1] + 11'h247;
  assign sel_178106 = $signed({1'h0, add_178001, array_index_177864[0]}) < $signed({1'h0, sel_178004}) ? {add_178001, array_index_177864[0]} : sel_178004;
  assign add_178131 = array_index_178065[11:0] + 12'h247;
  assign sel_178133 = $signed({1'h0, add_178029}) < $signed({1'h0, sel_178031}) ? add_178029 : sel_178031;
  assign add_178136 = array_index_178068[11:0] + 12'h247;
  assign sel_178138 = $signed({1'h0, add_178034}) < $signed({1'h0, sel_178036}) ? add_178034 : sel_178036;
  assign array_index_178167 = set1_unflattened[7'h36];
  assign array_index_178170 = set2_unflattened[7'h36];
  assign add_178174 = array_index_177759[11:1] + 11'h79d;
  assign sel_178176 = $signed({1'h0, add_178072, array_index_177657[0]}) < $signed({1'h0, sel_178074}) ? {add_178072, array_index_177657[0]} : sel_178074;
  assign add_178178 = array_index_177762[11:1] + 11'h79d;
  assign sel_178180 = $signed({1'h0, add_178076, array_index_177660[0]}) < $signed({1'h0, sel_178078}) ? {add_178076, array_index_177660[0]} : sel_178078;
  assign add_178182 = array_index_177861[11:1] + 11'h347;
  assign sel_178184 = $signed({1'h0, add_178080, array_index_177759[0]}) < $signed({1'h0, sel_178082}) ? {add_178080, array_index_177759[0]} : sel_178082;
  assign add_178186 = array_index_177864[11:1] + 11'h347;
  assign sel_178188 = $signed({1'h0, add_178084, array_index_177762[0]}) < $signed({1'h0, sel_178086}) ? {add_178084, array_index_177762[0]} : sel_178086;
  assign add_178190 = array_index_177963[11:3] + 9'h0bd;
  assign sel_178193 = $signed({1'h0, add_178088, array_index_177861[2:0]}) < $signed({1'h0, sel_178091}) ? {add_178088, array_index_177861[2:0]} : sel_178091;
  assign add_178195 = array_index_177966[11:3] + 9'h0bd;
  assign sel_178198 = $signed({1'h0, add_178093, array_index_177864[2:0]}) < $signed({1'h0, sel_178096}) ? {add_178093, array_index_177864[2:0]} : sel_178096;
  assign add_178200 = array_index_178065[11:1] + 11'h247;
  assign sel_178203 = $signed({1'h0, add_178098, array_index_177963[0]}) < $signed({1'h0, sel_178101}) ? {add_178098, array_index_177963[0]} : sel_178101;
  assign add_178205 = array_index_178068[11:1] + 11'h247;
  assign sel_178208 = $signed({1'h0, add_178103, array_index_177966[0]}) < $signed({1'h0, sel_178106}) ? {add_178103, array_index_177966[0]} : sel_178106;
  assign add_178233 = array_index_178167[11:0] + 12'h247;
  assign sel_178235 = $signed({1'h0, add_178131}) < $signed({1'h0, sel_178133}) ? add_178131 : sel_178133;
  assign add_178238 = array_index_178170[11:0] + 12'h247;
  assign sel_178240 = $signed({1'h0, add_178136}) < $signed({1'h0, sel_178138}) ? add_178136 : sel_178138;
  assign array_index_178269 = set1_unflattened[7'h37];
  assign array_index_178272 = set2_unflattened[7'h37];
  assign add_178276 = array_index_177861[11:1] + 11'h79d;
  assign sel_178278 = $signed({1'h0, add_178174, array_index_177759[0]}) < $signed({1'h0, sel_178176}) ? {add_178174, array_index_177759[0]} : sel_178176;
  assign add_178280 = array_index_177864[11:1] + 11'h79d;
  assign sel_178282 = $signed({1'h0, add_178178, array_index_177762[0]}) < $signed({1'h0, sel_178180}) ? {add_178178, array_index_177762[0]} : sel_178180;
  assign add_178284 = array_index_177963[11:1] + 11'h347;
  assign sel_178286 = $signed({1'h0, add_178182, array_index_177861[0]}) < $signed({1'h0, sel_178184}) ? {add_178182, array_index_177861[0]} : sel_178184;
  assign add_178288 = array_index_177966[11:1] + 11'h347;
  assign sel_178290 = $signed({1'h0, add_178186, array_index_177864[0]}) < $signed({1'h0, sel_178188}) ? {add_178186, array_index_177864[0]} : sel_178188;
  assign add_178292 = array_index_178065[11:3] + 9'h0bd;
  assign sel_178295 = $signed({1'h0, add_178190, array_index_177963[2:0]}) < $signed({1'h0, sel_178193}) ? {add_178190, array_index_177963[2:0]} : sel_178193;
  assign add_178297 = array_index_178068[11:3] + 9'h0bd;
  assign sel_178300 = $signed({1'h0, add_178195, array_index_177966[2:0]}) < $signed({1'h0, sel_178198}) ? {add_178195, array_index_177966[2:0]} : sel_178198;
  assign add_178302 = array_index_178167[11:1] + 11'h247;
  assign sel_178305 = $signed({1'h0, add_178200, array_index_178065[0]}) < $signed({1'h0, sel_178203}) ? {add_178200, array_index_178065[0]} : sel_178203;
  assign add_178307 = array_index_178170[11:1] + 11'h247;
  assign sel_178310 = $signed({1'h0, add_178205, array_index_178068[0]}) < $signed({1'h0, sel_178208}) ? {add_178205, array_index_178068[0]} : sel_178208;
  assign add_178335 = array_index_178269[11:0] + 12'h247;
  assign sel_178337 = $signed({1'h0, add_178233}) < $signed({1'h0, sel_178235}) ? add_178233 : sel_178235;
  assign add_178340 = array_index_178272[11:0] + 12'h247;
  assign sel_178342 = $signed({1'h0, add_178238}) < $signed({1'h0, sel_178240}) ? add_178238 : sel_178240;
  assign array_index_178371 = set1_unflattened[7'h38];
  assign array_index_178374 = set2_unflattened[7'h38];
  assign add_178378 = array_index_177963[11:1] + 11'h79d;
  assign sel_178380 = $signed({1'h0, add_178276, array_index_177861[0]}) < $signed({1'h0, sel_178278}) ? {add_178276, array_index_177861[0]} : sel_178278;
  assign add_178382 = array_index_177966[11:1] + 11'h79d;
  assign sel_178384 = $signed({1'h0, add_178280, array_index_177864[0]}) < $signed({1'h0, sel_178282}) ? {add_178280, array_index_177864[0]} : sel_178282;
  assign add_178386 = array_index_178065[11:1] + 11'h347;
  assign sel_178388 = $signed({1'h0, add_178284, array_index_177963[0]}) < $signed({1'h0, sel_178286}) ? {add_178284, array_index_177963[0]} : sel_178286;
  assign add_178390 = array_index_178068[11:1] + 11'h347;
  assign sel_178392 = $signed({1'h0, add_178288, array_index_177966[0]}) < $signed({1'h0, sel_178290}) ? {add_178288, array_index_177966[0]} : sel_178290;
  assign add_178394 = array_index_178167[11:3] + 9'h0bd;
  assign sel_178397 = $signed({1'h0, add_178292, array_index_178065[2:0]}) < $signed({1'h0, sel_178295}) ? {add_178292, array_index_178065[2:0]} : sel_178295;
  assign add_178399 = array_index_178170[11:3] + 9'h0bd;
  assign sel_178402 = $signed({1'h0, add_178297, array_index_178068[2:0]}) < $signed({1'h0, sel_178300}) ? {add_178297, array_index_178068[2:0]} : sel_178300;
  assign add_178404 = array_index_178269[11:1] + 11'h247;
  assign sel_178407 = $signed({1'h0, add_178302, array_index_178167[0]}) < $signed({1'h0, sel_178305}) ? {add_178302, array_index_178167[0]} : sel_178305;
  assign add_178409 = array_index_178272[11:1] + 11'h247;
  assign sel_178412 = $signed({1'h0, add_178307, array_index_178170[0]}) < $signed({1'h0, sel_178310}) ? {add_178307, array_index_178170[0]} : sel_178310;
  assign add_178437 = array_index_178371[11:0] + 12'h247;
  assign sel_178439 = $signed({1'h0, add_178335}) < $signed({1'h0, sel_178337}) ? add_178335 : sel_178337;
  assign add_178442 = array_index_178374[11:0] + 12'h247;
  assign sel_178444 = $signed({1'h0, add_178340}) < $signed({1'h0, sel_178342}) ? add_178340 : sel_178342;
  assign array_index_178473 = set1_unflattened[7'h39];
  assign array_index_178476 = set2_unflattened[7'h39];
  assign add_178480 = array_index_178065[11:1] + 11'h79d;
  assign sel_178482 = $signed({1'h0, add_178378, array_index_177963[0]}) < $signed({1'h0, sel_178380}) ? {add_178378, array_index_177963[0]} : sel_178380;
  assign add_178484 = array_index_178068[11:1] + 11'h79d;
  assign sel_178486 = $signed({1'h0, add_178382, array_index_177966[0]}) < $signed({1'h0, sel_178384}) ? {add_178382, array_index_177966[0]} : sel_178384;
  assign add_178488 = array_index_178167[11:1] + 11'h347;
  assign sel_178490 = $signed({1'h0, add_178386, array_index_178065[0]}) < $signed({1'h0, sel_178388}) ? {add_178386, array_index_178065[0]} : sel_178388;
  assign add_178492 = array_index_178170[11:1] + 11'h347;
  assign sel_178494 = $signed({1'h0, add_178390, array_index_178068[0]}) < $signed({1'h0, sel_178392}) ? {add_178390, array_index_178068[0]} : sel_178392;
  assign add_178496 = array_index_178269[11:3] + 9'h0bd;
  assign sel_178499 = $signed({1'h0, add_178394, array_index_178167[2:0]}) < $signed({1'h0, sel_178397}) ? {add_178394, array_index_178167[2:0]} : sel_178397;
  assign add_178501 = array_index_178272[11:3] + 9'h0bd;
  assign sel_178504 = $signed({1'h0, add_178399, array_index_178170[2:0]}) < $signed({1'h0, sel_178402}) ? {add_178399, array_index_178170[2:0]} : sel_178402;
  assign add_178506 = array_index_178371[11:1] + 11'h247;
  assign sel_178509 = $signed({1'h0, add_178404, array_index_178269[0]}) < $signed({1'h0, sel_178407}) ? {add_178404, array_index_178269[0]} : sel_178407;
  assign add_178511 = array_index_178374[11:1] + 11'h247;
  assign sel_178514 = $signed({1'h0, add_178409, array_index_178272[0]}) < $signed({1'h0, sel_178412}) ? {add_178409, array_index_178272[0]} : sel_178412;
  assign add_178539 = array_index_178473[11:0] + 12'h247;
  assign sel_178541 = $signed({1'h0, add_178437}) < $signed({1'h0, sel_178439}) ? add_178437 : sel_178439;
  assign add_178544 = array_index_178476[11:0] + 12'h247;
  assign sel_178546 = $signed({1'h0, add_178442}) < $signed({1'h0, sel_178444}) ? add_178442 : sel_178444;
  assign array_index_178575 = set1_unflattened[7'h3a];
  assign array_index_178578 = set2_unflattened[7'h3a];
  assign add_178582 = array_index_178167[11:1] + 11'h79d;
  assign sel_178584 = $signed({1'h0, add_178480, array_index_178065[0]}) < $signed({1'h0, sel_178482}) ? {add_178480, array_index_178065[0]} : sel_178482;
  assign add_178586 = array_index_178170[11:1] + 11'h79d;
  assign sel_178588 = $signed({1'h0, add_178484, array_index_178068[0]}) < $signed({1'h0, sel_178486}) ? {add_178484, array_index_178068[0]} : sel_178486;
  assign add_178590 = array_index_178269[11:1] + 11'h347;
  assign sel_178592 = $signed({1'h0, add_178488, array_index_178167[0]}) < $signed({1'h0, sel_178490}) ? {add_178488, array_index_178167[0]} : sel_178490;
  assign add_178594 = array_index_178272[11:1] + 11'h347;
  assign sel_178596 = $signed({1'h0, add_178492, array_index_178170[0]}) < $signed({1'h0, sel_178494}) ? {add_178492, array_index_178170[0]} : sel_178494;
  assign add_178598 = array_index_178371[11:3] + 9'h0bd;
  assign sel_178601 = $signed({1'h0, add_178496, array_index_178269[2:0]}) < $signed({1'h0, sel_178499}) ? {add_178496, array_index_178269[2:0]} : sel_178499;
  assign add_178603 = array_index_178374[11:3] + 9'h0bd;
  assign sel_178606 = $signed({1'h0, add_178501, array_index_178272[2:0]}) < $signed({1'h0, sel_178504}) ? {add_178501, array_index_178272[2:0]} : sel_178504;
  assign add_178608 = array_index_178473[11:1] + 11'h247;
  assign sel_178611 = $signed({1'h0, add_178506, array_index_178371[0]}) < $signed({1'h0, sel_178509}) ? {add_178506, array_index_178371[0]} : sel_178509;
  assign add_178613 = array_index_178476[11:1] + 11'h247;
  assign sel_178616 = $signed({1'h0, add_178511, array_index_178374[0]}) < $signed({1'h0, sel_178514}) ? {add_178511, array_index_178374[0]} : sel_178514;
  assign add_178641 = array_index_178575[11:0] + 12'h247;
  assign sel_178643 = $signed({1'h0, add_178539}) < $signed({1'h0, sel_178541}) ? add_178539 : sel_178541;
  assign add_178646 = array_index_178578[11:0] + 12'h247;
  assign sel_178648 = $signed({1'h0, add_178544}) < $signed({1'h0, sel_178546}) ? add_178544 : sel_178546;
  assign array_index_178677 = set1_unflattened[7'h3b];
  assign array_index_178680 = set2_unflattened[7'h3b];
  assign add_178684 = array_index_178269[11:1] + 11'h79d;
  assign sel_178686 = $signed({1'h0, add_178582, array_index_178167[0]}) < $signed({1'h0, sel_178584}) ? {add_178582, array_index_178167[0]} : sel_178584;
  assign add_178688 = array_index_178272[11:1] + 11'h79d;
  assign sel_178690 = $signed({1'h0, add_178586, array_index_178170[0]}) < $signed({1'h0, sel_178588}) ? {add_178586, array_index_178170[0]} : sel_178588;
  assign add_178692 = array_index_178371[11:1] + 11'h347;
  assign sel_178694 = $signed({1'h0, add_178590, array_index_178269[0]}) < $signed({1'h0, sel_178592}) ? {add_178590, array_index_178269[0]} : sel_178592;
  assign add_178696 = array_index_178374[11:1] + 11'h347;
  assign sel_178698 = $signed({1'h0, add_178594, array_index_178272[0]}) < $signed({1'h0, sel_178596}) ? {add_178594, array_index_178272[0]} : sel_178596;
  assign add_178700 = array_index_178473[11:3] + 9'h0bd;
  assign sel_178703 = $signed({1'h0, add_178598, array_index_178371[2:0]}) < $signed({1'h0, sel_178601}) ? {add_178598, array_index_178371[2:0]} : sel_178601;
  assign add_178705 = array_index_178476[11:3] + 9'h0bd;
  assign sel_178708 = $signed({1'h0, add_178603, array_index_178374[2:0]}) < $signed({1'h0, sel_178606}) ? {add_178603, array_index_178374[2:0]} : sel_178606;
  assign add_178710 = array_index_178575[11:1] + 11'h247;
  assign sel_178713 = $signed({1'h0, add_178608, array_index_178473[0]}) < $signed({1'h0, sel_178611}) ? {add_178608, array_index_178473[0]} : sel_178611;
  assign add_178715 = array_index_178578[11:1] + 11'h247;
  assign sel_178718 = $signed({1'h0, add_178613, array_index_178476[0]}) < $signed({1'h0, sel_178616}) ? {add_178613, array_index_178476[0]} : sel_178616;
  assign add_178743 = array_index_178677[11:0] + 12'h247;
  assign sel_178745 = $signed({1'h0, add_178641}) < $signed({1'h0, sel_178643}) ? add_178641 : sel_178643;
  assign add_178748 = array_index_178680[11:0] + 12'h247;
  assign sel_178750 = $signed({1'h0, add_178646}) < $signed({1'h0, sel_178648}) ? add_178646 : sel_178648;
  assign array_index_178779 = set1_unflattened[7'h3c];
  assign array_index_178782 = set2_unflattened[7'h3c];
  assign add_178786 = array_index_178371[11:1] + 11'h79d;
  assign sel_178788 = $signed({1'h0, add_178684, array_index_178269[0]}) < $signed({1'h0, sel_178686}) ? {add_178684, array_index_178269[0]} : sel_178686;
  assign add_178790 = array_index_178374[11:1] + 11'h79d;
  assign sel_178792 = $signed({1'h0, add_178688, array_index_178272[0]}) < $signed({1'h0, sel_178690}) ? {add_178688, array_index_178272[0]} : sel_178690;
  assign add_178794 = array_index_178473[11:1] + 11'h347;
  assign sel_178796 = $signed({1'h0, add_178692, array_index_178371[0]}) < $signed({1'h0, sel_178694}) ? {add_178692, array_index_178371[0]} : sel_178694;
  assign add_178798 = array_index_178476[11:1] + 11'h347;
  assign sel_178800 = $signed({1'h0, add_178696, array_index_178374[0]}) < $signed({1'h0, sel_178698}) ? {add_178696, array_index_178374[0]} : sel_178698;
  assign add_178802 = array_index_178575[11:3] + 9'h0bd;
  assign sel_178805 = $signed({1'h0, add_178700, array_index_178473[2:0]}) < $signed({1'h0, sel_178703}) ? {add_178700, array_index_178473[2:0]} : sel_178703;
  assign add_178807 = array_index_178578[11:3] + 9'h0bd;
  assign sel_178810 = $signed({1'h0, add_178705, array_index_178476[2:0]}) < $signed({1'h0, sel_178708}) ? {add_178705, array_index_178476[2:0]} : sel_178708;
  assign add_178812 = array_index_178677[11:1] + 11'h247;
  assign sel_178815 = $signed({1'h0, add_178710, array_index_178575[0]}) < $signed({1'h0, sel_178713}) ? {add_178710, array_index_178575[0]} : sel_178713;
  assign add_178817 = array_index_178680[11:1] + 11'h247;
  assign sel_178820 = $signed({1'h0, add_178715, array_index_178578[0]}) < $signed({1'h0, sel_178718}) ? {add_178715, array_index_178578[0]} : sel_178718;
  assign add_178845 = array_index_178779[11:0] + 12'h247;
  assign sel_178847 = $signed({1'h0, add_178743}) < $signed({1'h0, sel_178745}) ? add_178743 : sel_178745;
  assign add_178850 = array_index_178782[11:0] + 12'h247;
  assign sel_178852 = $signed({1'h0, add_178748}) < $signed({1'h0, sel_178750}) ? add_178748 : sel_178750;
  assign array_index_178881 = set1_unflattened[7'h3d];
  assign array_index_178884 = set2_unflattened[7'h3d];
  assign add_178888 = array_index_178473[11:1] + 11'h79d;
  assign sel_178890 = $signed({1'h0, add_178786, array_index_178371[0]}) < $signed({1'h0, sel_178788}) ? {add_178786, array_index_178371[0]} : sel_178788;
  assign add_178892 = array_index_178476[11:1] + 11'h79d;
  assign sel_178894 = $signed({1'h0, add_178790, array_index_178374[0]}) < $signed({1'h0, sel_178792}) ? {add_178790, array_index_178374[0]} : sel_178792;
  assign add_178896 = array_index_178575[11:1] + 11'h347;
  assign sel_178898 = $signed({1'h0, add_178794, array_index_178473[0]}) < $signed({1'h0, sel_178796}) ? {add_178794, array_index_178473[0]} : sel_178796;
  assign add_178900 = array_index_178578[11:1] + 11'h347;
  assign sel_178902 = $signed({1'h0, add_178798, array_index_178476[0]}) < $signed({1'h0, sel_178800}) ? {add_178798, array_index_178476[0]} : sel_178800;
  assign add_178904 = array_index_178677[11:3] + 9'h0bd;
  assign sel_178907 = $signed({1'h0, add_178802, array_index_178575[2:0]}) < $signed({1'h0, sel_178805}) ? {add_178802, array_index_178575[2:0]} : sel_178805;
  assign add_178909 = array_index_178680[11:3] + 9'h0bd;
  assign sel_178912 = $signed({1'h0, add_178807, array_index_178578[2:0]}) < $signed({1'h0, sel_178810}) ? {add_178807, array_index_178578[2:0]} : sel_178810;
  assign add_178914 = array_index_178779[11:1] + 11'h247;
  assign sel_178917 = $signed({1'h0, add_178812, array_index_178677[0]}) < $signed({1'h0, sel_178815}) ? {add_178812, array_index_178677[0]} : sel_178815;
  assign add_178919 = array_index_178782[11:1] + 11'h247;
  assign sel_178922 = $signed({1'h0, add_178817, array_index_178680[0]}) < $signed({1'h0, sel_178820}) ? {add_178817, array_index_178680[0]} : sel_178820;
  assign add_178947 = array_index_178881[11:0] + 12'h247;
  assign sel_178949 = $signed({1'h0, add_178845}) < $signed({1'h0, sel_178847}) ? add_178845 : sel_178847;
  assign add_178952 = array_index_178884[11:0] + 12'h247;
  assign sel_178954 = $signed({1'h0, add_178850}) < $signed({1'h0, sel_178852}) ? add_178850 : sel_178852;
  assign array_index_178983 = set1_unflattened[7'h3e];
  assign array_index_178986 = set2_unflattened[7'h3e];
  assign add_178990 = array_index_178575[11:1] + 11'h79d;
  assign sel_178992 = $signed({1'h0, add_178888, array_index_178473[0]}) < $signed({1'h0, sel_178890}) ? {add_178888, array_index_178473[0]} : sel_178890;
  assign add_178994 = array_index_178578[11:1] + 11'h79d;
  assign sel_178996 = $signed({1'h0, add_178892, array_index_178476[0]}) < $signed({1'h0, sel_178894}) ? {add_178892, array_index_178476[0]} : sel_178894;
  assign add_178998 = array_index_178677[11:1] + 11'h347;
  assign sel_179000 = $signed({1'h0, add_178896, array_index_178575[0]}) < $signed({1'h0, sel_178898}) ? {add_178896, array_index_178575[0]} : sel_178898;
  assign add_179002 = array_index_178680[11:1] + 11'h347;
  assign sel_179004 = $signed({1'h0, add_178900, array_index_178578[0]}) < $signed({1'h0, sel_178902}) ? {add_178900, array_index_178578[0]} : sel_178902;
  assign add_179006 = array_index_178779[11:3] + 9'h0bd;
  assign sel_179009 = $signed({1'h0, add_178904, array_index_178677[2:0]}) < $signed({1'h0, sel_178907}) ? {add_178904, array_index_178677[2:0]} : sel_178907;
  assign add_179011 = array_index_178782[11:3] + 9'h0bd;
  assign sel_179014 = $signed({1'h0, add_178909, array_index_178680[2:0]}) < $signed({1'h0, sel_178912}) ? {add_178909, array_index_178680[2:0]} : sel_178912;
  assign add_179016 = array_index_178881[11:1] + 11'h247;
  assign sel_179019 = $signed({1'h0, add_178914, array_index_178779[0]}) < $signed({1'h0, sel_178917}) ? {add_178914, array_index_178779[0]} : sel_178917;
  assign add_179021 = array_index_178884[11:1] + 11'h247;
  assign sel_179024 = $signed({1'h0, add_178919, array_index_178782[0]}) < $signed({1'h0, sel_178922}) ? {add_178919, array_index_178782[0]} : sel_178922;
  assign add_179049 = array_index_178983[11:0] + 12'h247;
  assign sel_179051 = $signed({1'h0, add_178947}) < $signed({1'h0, sel_178949}) ? add_178947 : sel_178949;
  assign add_179054 = array_index_178986[11:0] + 12'h247;
  assign sel_179056 = $signed({1'h0, add_178952}) < $signed({1'h0, sel_178954}) ? add_178952 : sel_178954;
  assign array_index_179085 = set1_unflattened[7'h3f];
  assign array_index_179088 = set2_unflattened[7'h3f];
  assign add_179092 = array_index_178677[11:1] + 11'h79d;
  assign sel_179094 = $signed({1'h0, add_178990, array_index_178575[0]}) < $signed({1'h0, sel_178992}) ? {add_178990, array_index_178575[0]} : sel_178992;
  assign add_179096 = array_index_178680[11:1] + 11'h79d;
  assign sel_179098 = $signed({1'h0, add_178994, array_index_178578[0]}) < $signed({1'h0, sel_178996}) ? {add_178994, array_index_178578[0]} : sel_178996;
  assign add_179100 = array_index_178779[11:1] + 11'h347;
  assign sel_179102 = $signed({1'h0, add_178998, array_index_178677[0]}) < $signed({1'h0, sel_179000}) ? {add_178998, array_index_178677[0]} : sel_179000;
  assign add_179104 = array_index_178782[11:1] + 11'h347;
  assign sel_179106 = $signed({1'h0, add_179002, array_index_178680[0]}) < $signed({1'h0, sel_179004}) ? {add_179002, array_index_178680[0]} : sel_179004;
  assign add_179108 = array_index_178881[11:3] + 9'h0bd;
  assign sel_179111 = $signed({1'h0, add_179006, array_index_178779[2:0]}) < $signed({1'h0, sel_179009}) ? {add_179006, array_index_178779[2:0]} : sel_179009;
  assign add_179113 = array_index_178884[11:3] + 9'h0bd;
  assign sel_179116 = $signed({1'h0, add_179011, array_index_178782[2:0]}) < $signed({1'h0, sel_179014}) ? {add_179011, array_index_178782[2:0]} : sel_179014;
  assign add_179118 = array_index_178983[11:1] + 11'h247;
  assign sel_179121 = $signed({1'h0, add_179016, array_index_178881[0]}) < $signed({1'h0, sel_179019}) ? {add_179016, array_index_178881[0]} : sel_179019;
  assign add_179123 = array_index_178986[11:1] + 11'h247;
  assign sel_179126 = $signed({1'h0, add_179021, array_index_178884[0]}) < $signed({1'h0, sel_179024}) ? {add_179021, array_index_178884[0]} : sel_179024;
  assign add_179151 = array_index_179085[11:0] + 12'h247;
  assign sel_179153 = $signed({1'h0, add_179049}) < $signed({1'h0, sel_179051}) ? add_179049 : sel_179051;
  assign add_179156 = array_index_179088[11:0] + 12'h247;
  assign sel_179158 = $signed({1'h0, add_179054}) < $signed({1'h0, sel_179056}) ? add_179054 : sel_179056;
  assign array_index_179187 = set1_unflattened[7'h40];
  assign array_index_179190 = set2_unflattened[7'h40];
  assign add_179194 = array_index_178779[11:1] + 11'h79d;
  assign sel_179196 = $signed({1'h0, add_179092, array_index_178677[0]}) < $signed({1'h0, sel_179094}) ? {add_179092, array_index_178677[0]} : sel_179094;
  assign add_179198 = array_index_178782[11:1] + 11'h79d;
  assign sel_179200 = $signed({1'h0, add_179096, array_index_178680[0]}) < $signed({1'h0, sel_179098}) ? {add_179096, array_index_178680[0]} : sel_179098;
  assign add_179202 = array_index_178881[11:1] + 11'h347;
  assign sel_179204 = $signed({1'h0, add_179100, array_index_178779[0]}) < $signed({1'h0, sel_179102}) ? {add_179100, array_index_178779[0]} : sel_179102;
  assign add_179206 = array_index_178884[11:1] + 11'h347;
  assign sel_179208 = $signed({1'h0, add_179104, array_index_178782[0]}) < $signed({1'h0, sel_179106}) ? {add_179104, array_index_178782[0]} : sel_179106;
  assign add_179210 = array_index_178983[11:3] + 9'h0bd;
  assign sel_179213 = $signed({1'h0, add_179108, array_index_178881[2:0]}) < $signed({1'h0, sel_179111}) ? {add_179108, array_index_178881[2:0]} : sel_179111;
  assign add_179215 = array_index_178986[11:3] + 9'h0bd;
  assign sel_179218 = $signed({1'h0, add_179113, array_index_178884[2:0]}) < $signed({1'h0, sel_179116}) ? {add_179113, array_index_178884[2:0]} : sel_179116;
  assign add_179220 = array_index_179085[11:1] + 11'h247;
  assign sel_179223 = $signed({1'h0, add_179118, array_index_178983[0]}) < $signed({1'h0, sel_179121}) ? {add_179118, array_index_178983[0]} : sel_179121;
  assign add_179225 = array_index_179088[11:1] + 11'h247;
  assign sel_179228 = $signed({1'h0, add_179123, array_index_178986[0]}) < $signed({1'h0, sel_179126}) ? {add_179123, array_index_178986[0]} : sel_179126;
  assign add_179253 = array_index_179187[11:0] + 12'h247;
  assign sel_179255 = $signed({1'h0, add_179151}) < $signed({1'h0, sel_179153}) ? add_179151 : sel_179153;
  assign add_179258 = array_index_179190[11:0] + 12'h247;
  assign sel_179260 = $signed({1'h0, add_179156}) < $signed({1'h0, sel_179158}) ? add_179156 : sel_179158;
  assign array_index_179289 = set1_unflattened[7'h41];
  assign array_index_179292 = set2_unflattened[7'h41];
  assign add_179296 = array_index_178881[11:1] + 11'h79d;
  assign sel_179298 = $signed({1'h0, add_179194, array_index_178779[0]}) < $signed({1'h0, sel_179196}) ? {add_179194, array_index_178779[0]} : sel_179196;
  assign add_179300 = array_index_178884[11:1] + 11'h79d;
  assign sel_179302 = $signed({1'h0, add_179198, array_index_178782[0]}) < $signed({1'h0, sel_179200}) ? {add_179198, array_index_178782[0]} : sel_179200;
  assign add_179304 = array_index_178983[11:1] + 11'h347;
  assign sel_179306 = $signed({1'h0, add_179202, array_index_178881[0]}) < $signed({1'h0, sel_179204}) ? {add_179202, array_index_178881[0]} : sel_179204;
  assign add_179308 = array_index_178986[11:1] + 11'h347;
  assign sel_179310 = $signed({1'h0, add_179206, array_index_178884[0]}) < $signed({1'h0, sel_179208}) ? {add_179206, array_index_178884[0]} : sel_179208;
  assign add_179312 = array_index_179085[11:3] + 9'h0bd;
  assign sel_179315 = $signed({1'h0, add_179210, array_index_178983[2:0]}) < $signed({1'h0, sel_179213}) ? {add_179210, array_index_178983[2:0]} : sel_179213;
  assign add_179317 = array_index_179088[11:3] + 9'h0bd;
  assign sel_179320 = $signed({1'h0, add_179215, array_index_178986[2:0]}) < $signed({1'h0, sel_179218}) ? {add_179215, array_index_178986[2:0]} : sel_179218;
  assign add_179322 = array_index_179187[11:1] + 11'h247;
  assign sel_179325 = $signed({1'h0, add_179220, array_index_179085[0]}) < $signed({1'h0, sel_179223}) ? {add_179220, array_index_179085[0]} : sel_179223;
  assign add_179327 = array_index_179190[11:1] + 11'h247;
  assign sel_179330 = $signed({1'h0, add_179225, array_index_179088[0]}) < $signed({1'h0, sel_179228}) ? {add_179225, array_index_179088[0]} : sel_179228;
  assign add_179355 = array_index_179289[11:0] + 12'h247;
  assign sel_179357 = $signed({1'h0, add_179253}) < $signed({1'h0, sel_179255}) ? add_179253 : sel_179255;
  assign add_179360 = array_index_179292[11:0] + 12'h247;
  assign sel_179362 = $signed({1'h0, add_179258}) < $signed({1'h0, sel_179260}) ? add_179258 : sel_179260;
  assign array_index_179391 = set1_unflattened[7'h42];
  assign array_index_179394 = set2_unflattened[7'h42];
  assign add_179398 = array_index_178983[11:1] + 11'h79d;
  assign sel_179400 = $signed({1'h0, add_179296, array_index_178881[0]}) < $signed({1'h0, sel_179298}) ? {add_179296, array_index_178881[0]} : sel_179298;
  assign add_179402 = array_index_178986[11:1] + 11'h79d;
  assign sel_179404 = $signed({1'h0, add_179300, array_index_178884[0]}) < $signed({1'h0, sel_179302}) ? {add_179300, array_index_178884[0]} : sel_179302;
  assign add_179406 = array_index_179085[11:1] + 11'h347;
  assign sel_179408 = $signed({1'h0, add_179304, array_index_178983[0]}) < $signed({1'h0, sel_179306}) ? {add_179304, array_index_178983[0]} : sel_179306;
  assign add_179410 = array_index_179088[11:1] + 11'h347;
  assign sel_179412 = $signed({1'h0, add_179308, array_index_178986[0]}) < $signed({1'h0, sel_179310}) ? {add_179308, array_index_178986[0]} : sel_179310;
  assign add_179414 = array_index_179187[11:3] + 9'h0bd;
  assign sel_179417 = $signed({1'h0, add_179312, array_index_179085[2:0]}) < $signed({1'h0, sel_179315}) ? {add_179312, array_index_179085[2:0]} : sel_179315;
  assign add_179419 = array_index_179190[11:3] + 9'h0bd;
  assign sel_179422 = $signed({1'h0, add_179317, array_index_179088[2:0]}) < $signed({1'h0, sel_179320}) ? {add_179317, array_index_179088[2:0]} : sel_179320;
  assign add_179424 = array_index_179289[11:1] + 11'h247;
  assign sel_179427 = $signed({1'h0, add_179322, array_index_179187[0]}) < $signed({1'h0, sel_179325}) ? {add_179322, array_index_179187[0]} : sel_179325;
  assign add_179429 = array_index_179292[11:1] + 11'h247;
  assign sel_179432 = $signed({1'h0, add_179327, array_index_179190[0]}) < $signed({1'h0, sel_179330}) ? {add_179327, array_index_179190[0]} : sel_179330;
  assign add_179457 = array_index_179391[11:0] + 12'h247;
  assign sel_179459 = $signed({1'h0, add_179355}) < $signed({1'h0, sel_179357}) ? add_179355 : sel_179357;
  assign add_179462 = array_index_179394[11:0] + 12'h247;
  assign sel_179464 = $signed({1'h0, add_179360}) < $signed({1'h0, sel_179362}) ? add_179360 : sel_179362;
  assign array_index_179493 = set1_unflattened[7'h43];
  assign array_index_179496 = set2_unflattened[7'h43];
  assign add_179500 = array_index_179085[11:1] + 11'h79d;
  assign sel_179502 = $signed({1'h0, add_179398, array_index_178983[0]}) < $signed({1'h0, sel_179400}) ? {add_179398, array_index_178983[0]} : sel_179400;
  assign add_179504 = array_index_179088[11:1] + 11'h79d;
  assign sel_179506 = $signed({1'h0, add_179402, array_index_178986[0]}) < $signed({1'h0, sel_179404}) ? {add_179402, array_index_178986[0]} : sel_179404;
  assign add_179508 = array_index_179187[11:1] + 11'h347;
  assign sel_179510 = $signed({1'h0, add_179406, array_index_179085[0]}) < $signed({1'h0, sel_179408}) ? {add_179406, array_index_179085[0]} : sel_179408;
  assign add_179512 = array_index_179190[11:1] + 11'h347;
  assign sel_179514 = $signed({1'h0, add_179410, array_index_179088[0]}) < $signed({1'h0, sel_179412}) ? {add_179410, array_index_179088[0]} : sel_179412;
  assign add_179516 = array_index_179289[11:3] + 9'h0bd;
  assign sel_179519 = $signed({1'h0, add_179414, array_index_179187[2:0]}) < $signed({1'h0, sel_179417}) ? {add_179414, array_index_179187[2:0]} : sel_179417;
  assign add_179521 = array_index_179292[11:3] + 9'h0bd;
  assign sel_179524 = $signed({1'h0, add_179419, array_index_179190[2:0]}) < $signed({1'h0, sel_179422}) ? {add_179419, array_index_179190[2:0]} : sel_179422;
  assign add_179526 = array_index_179391[11:1] + 11'h247;
  assign sel_179529 = $signed({1'h0, add_179424, array_index_179289[0]}) < $signed({1'h0, sel_179427}) ? {add_179424, array_index_179289[0]} : sel_179427;
  assign add_179531 = array_index_179394[11:1] + 11'h247;
  assign sel_179534 = $signed({1'h0, add_179429, array_index_179292[0]}) < $signed({1'h0, sel_179432}) ? {add_179429, array_index_179292[0]} : sel_179432;
  assign add_179559 = array_index_179493[11:0] + 12'h247;
  assign sel_179561 = $signed({1'h0, add_179457}) < $signed({1'h0, sel_179459}) ? add_179457 : sel_179459;
  assign add_179564 = array_index_179496[11:0] + 12'h247;
  assign sel_179566 = $signed({1'h0, add_179462}) < $signed({1'h0, sel_179464}) ? add_179462 : sel_179464;
  assign array_index_179595 = set1_unflattened[7'h44];
  assign array_index_179598 = set2_unflattened[7'h44];
  assign add_179602 = array_index_179187[11:1] + 11'h79d;
  assign sel_179604 = $signed({1'h0, add_179500, array_index_179085[0]}) < $signed({1'h0, sel_179502}) ? {add_179500, array_index_179085[0]} : sel_179502;
  assign add_179606 = array_index_179190[11:1] + 11'h79d;
  assign sel_179608 = $signed({1'h0, add_179504, array_index_179088[0]}) < $signed({1'h0, sel_179506}) ? {add_179504, array_index_179088[0]} : sel_179506;
  assign add_179610 = array_index_179289[11:1] + 11'h347;
  assign sel_179612 = $signed({1'h0, add_179508, array_index_179187[0]}) < $signed({1'h0, sel_179510}) ? {add_179508, array_index_179187[0]} : sel_179510;
  assign add_179614 = array_index_179292[11:1] + 11'h347;
  assign sel_179616 = $signed({1'h0, add_179512, array_index_179190[0]}) < $signed({1'h0, sel_179514}) ? {add_179512, array_index_179190[0]} : sel_179514;
  assign add_179618 = array_index_179391[11:3] + 9'h0bd;
  assign sel_179621 = $signed({1'h0, add_179516, array_index_179289[2:0]}) < $signed({1'h0, sel_179519}) ? {add_179516, array_index_179289[2:0]} : sel_179519;
  assign add_179623 = array_index_179394[11:3] + 9'h0bd;
  assign sel_179626 = $signed({1'h0, add_179521, array_index_179292[2:0]}) < $signed({1'h0, sel_179524}) ? {add_179521, array_index_179292[2:0]} : sel_179524;
  assign add_179628 = array_index_179493[11:1] + 11'h247;
  assign sel_179631 = $signed({1'h0, add_179526, array_index_179391[0]}) < $signed({1'h0, sel_179529}) ? {add_179526, array_index_179391[0]} : sel_179529;
  assign add_179633 = array_index_179496[11:1] + 11'h247;
  assign sel_179636 = $signed({1'h0, add_179531, array_index_179394[0]}) < $signed({1'h0, sel_179534}) ? {add_179531, array_index_179394[0]} : sel_179534;
  assign add_179661 = array_index_179595[11:0] + 12'h247;
  assign sel_179663 = $signed({1'h0, add_179559}) < $signed({1'h0, sel_179561}) ? add_179559 : sel_179561;
  assign add_179666 = array_index_179598[11:0] + 12'h247;
  assign sel_179668 = $signed({1'h0, add_179564}) < $signed({1'h0, sel_179566}) ? add_179564 : sel_179566;
  assign array_index_179697 = set1_unflattened[7'h45];
  assign array_index_179700 = set2_unflattened[7'h45];
  assign add_179704 = array_index_179289[11:1] + 11'h79d;
  assign sel_179706 = $signed({1'h0, add_179602, array_index_179187[0]}) < $signed({1'h0, sel_179604}) ? {add_179602, array_index_179187[0]} : sel_179604;
  assign add_179708 = array_index_179292[11:1] + 11'h79d;
  assign sel_179710 = $signed({1'h0, add_179606, array_index_179190[0]}) < $signed({1'h0, sel_179608}) ? {add_179606, array_index_179190[0]} : sel_179608;
  assign add_179712 = array_index_179391[11:1] + 11'h347;
  assign sel_179714 = $signed({1'h0, add_179610, array_index_179289[0]}) < $signed({1'h0, sel_179612}) ? {add_179610, array_index_179289[0]} : sel_179612;
  assign add_179716 = array_index_179394[11:1] + 11'h347;
  assign sel_179718 = $signed({1'h0, add_179614, array_index_179292[0]}) < $signed({1'h0, sel_179616}) ? {add_179614, array_index_179292[0]} : sel_179616;
  assign add_179720 = array_index_179493[11:3] + 9'h0bd;
  assign sel_179723 = $signed({1'h0, add_179618, array_index_179391[2:0]}) < $signed({1'h0, sel_179621}) ? {add_179618, array_index_179391[2:0]} : sel_179621;
  assign add_179725 = array_index_179496[11:3] + 9'h0bd;
  assign sel_179728 = $signed({1'h0, add_179623, array_index_179394[2:0]}) < $signed({1'h0, sel_179626}) ? {add_179623, array_index_179394[2:0]} : sel_179626;
  assign add_179730 = array_index_179595[11:1] + 11'h247;
  assign sel_179733 = $signed({1'h0, add_179628, array_index_179493[0]}) < $signed({1'h0, sel_179631}) ? {add_179628, array_index_179493[0]} : sel_179631;
  assign add_179735 = array_index_179598[11:1] + 11'h247;
  assign sel_179738 = $signed({1'h0, add_179633, array_index_179496[0]}) < $signed({1'h0, sel_179636}) ? {add_179633, array_index_179496[0]} : sel_179636;
  assign add_179763 = array_index_179697[11:0] + 12'h247;
  assign sel_179765 = $signed({1'h0, add_179661}) < $signed({1'h0, sel_179663}) ? add_179661 : sel_179663;
  assign add_179768 = array_index_179700[11:0] + 12'h247;
  assign sel_179770 = $signed({1'h0, add_179666}) < $signed({1'h0, sel_179668}) ? add_179666 : sel_179668;
  assign array_index_179799 = set1_unflattened[7'h46];
  assign array_index_179802 = set2_unflattened[7'h46];
  assign add_179806 = array_index_179391[11:1] + 11'h79d;
  assign sel_179808 = $signed({1'h0, add_179704, array_index_179289[0]}) < $signed({1'h0, sel_179706}) ? {add_179704, array_index_179289[0]} : sel_179706;
  assign add_179810 = array_index_179394[11:1] + 11'h79d;
  assign sel_179812 = $signed({1'h0, add_179708, array_index_179292[0]}) < $signed({1'h0, sel_179710}) ? {add_179708, array_index_179292[0]} : sel_179710;
  assign add_179814 = array_index_179493[11:1] + 11'h347;
  assign sel_179816 = $signed({1'h0, add_179712, array_index_179391[0]}) < $signed({1'h0, sel_179714}) ? {add_179712, array_index_179391[0]} : sel_179714;
  assign add_179818 = array_index_179496[11:1] + 11'h347;
  assign sel_179820 = $signed({1'h0, add_179716, array_index_179394[0]}) < $signed({1'h0, sel_179718}) ? {add_179716, array_index_179394[0]} : sel_179718;
  assign add_179822 = array_index_179595[11:3] + 9'h0bd;
  assign sel_179825 = $signed({1'h0, add_179720, array_index_179493[2:0]}) < $signed({1'h0, sel_179723}) ? {add_179720, array_index_179493[2:0]} : sel_179723;
  assign add_179827 = array_index_179598[11:3] + 9'h0bd;
  assign sel_179830 = $signed({1'h0, add_179725, array_index_179496[2:0]}) < $signed({1'h0, sel_179728}) ? {add_179725, array_index_179496[2:0]} : sel_179728;
  assign add_179832 = array_index_179697[11:1] + 11'h247;
  assign sel_179835 = $signed({1'h0, add_179730, array_index_179595[0]}) < $signed({1'h0, sel_179733}) ? {add_179730, array_index_179595[0]} : sel_179733;
  assign add_179837 = array_index_179700[11:1] + 11'h247;
  assign sel_179840 = $signed({1'h0, add_179735, array_index_179598[0]}) < $signed({1'h0, sel_179738}) ? {add_179735, array_index_179598[0]} : sel_179738;
  assign add_179865 = array_index_179799[11:0] + 12'h247;
  assign sel_179867 = $signed({1'h0, add_179763}) < $signed({1'h0, sel_179765}) ? add_179763 : sel_179765;
  assign add_179870 = array_index_179802[11:0] + 12'h247;
  assign sel_179872 = $signed({1'h0, add_179768}) < $signed({1'h0, sel_179770}) ? add_179768 : sel_179770;
  assign array_index_179901 = set1_unflattened[7'h47];
  assign array_index_179904 = set2_unflattened[7'h47];
  assign add_179908 = array_index_179493[11:1] + 11'h79d;
  assign sel_179910 = $signed({1'h0, add_179806, array_index_179391[0]}) < $signed({1'h0, sel_179808}) ? {add_179806, array_index_179391[0]} : sel_179808;
  assign add_179912 = array_index_179496[11:1] + 11'h79d;
  assign sel_179914 = $signed({1'h0, add_179810, array_index_179394[0]}) < $signed({1'h0, sel_179812}) ? {add_179810, array_index_179394[0]} : sel_179812;
  assign add_179916 = array_index_179595[11:1] + 11'h347;
  assign sel_179918 = $signed({1'h0, add_179814, array_index_179493[0]}) < $signed({1'h0, sel_179816}) ? {add_179814, array_index_179493[0]} : sel_179816;
  assign add_179920 = array_index_179598[11:1] + 11'h347;
  assign sel_179922 = $signed({1'h0, add_179818, array_index_179496[0]}) < $signed({1'h0, sel_179820}) ? {add_179818, array_index_179496[0]} : sel_179820;
  assign add_179924 = array_index_179697[11:3] + 9'h0bd;
  assign sel_179927 = $signed({1'h0, add_179822, array_index_179595[2:0]}) < $signed({1'h0, sel_179825}) ? {add_179822, array_index_179595[2:0]} : sel_179825;
  assign add_179929 = array_index_179700[11:3] + 9'h0bd;
  assign sel_179932 = $signed({1'h0, add_179827, array_index_179598[2:0]}) < $signed({1'h0, sel_179830}) ? {add_179827, array_index_179598[2:0]} : sel_179830;
  assign add_179934 = array_index_179799[11:1] + 11'h247;
  assign sel_179937 = $signed({1'h0, add_179832, array_index_179697[0]}) < $signed({1'h0, sel_179835}) ? {add_179832, array_index_179697[0]} : sel_179835;
  assign add_179939 = array_index_179802[11:1] + 11'h247;
  assign sel_179942 = $signed({1'h0, add_179837, array_index_179700[0]}) < $signed({1'h0, sel_179840}) ? {add_179837, array_index_179700[0]} : sel_179840;
  assign add_179967 = array_index_179901[11:0] + 12'h247;
  assign sel_179969 = $signed({1'h0, add_179865}) < $signed({1'h0, sel_179867}) ? add_179865 : sel_179867;
  assign add_179972 = array_index_179904[11:0] + 12'h247;
  assign sel_179974 = $signed({1'h0, add_179870}) < $signed({1'h0, sel_179872}) ? add_179870 : sel_179872;
  assign array_index_180003 = set1_unflattened[7'h48];
  assign array_index_180006 = set2_unflattened[7'h48];
  assign add_180010 = array_index_179595[11:1] + 11'h79d;
  assign sel_180012 = $signed({1'h0, add_179908, array_index_179493[0]}) < $signed({1'h0, sel_179910}) ? {add_179908, array_index_179493[0]} : sel_179910;
  assign add_180014 = array_index_179598[11:1] + 11'h79d;
  assign sel_180016 = $signed({1'h0, add_179912, array_index_179496[0]}) < $signed({1'h0, sel_179914}) ? {add_179912, array_index_179496[0]} : sel_179914;
  assign add_180018 = array_index_179697[11:1] + 11'h347;
  assign sel_180020 = $signed({1'h0, add_179916, array_index_179595[0]}) < $signed({1'h0, sel_179918}) ? {add_179916, array_index_179595[0]} : sel_179918;
  assign add_180022 = array_index_179700[11:1] + 11'h347;
  assign sel_180024 = $signed({1'h0, add_179920, array_index_179598[0]}) < $signed({1'h0, sel_179922}) ? {add_179920, array_index_179598[0]} : sel_179922;
  assign add_180026 = array_index_179799[11:3] + 9'h0bd;
  assign sel_180029 = $signed({1'h0, add_179924, array_index_179697[2:0]}) < $signed({1'h0, sel_179927}) ? {add_179924, array_index_179697[2:0]} : sel_179927;
  assign add_180031 = array_index_179802[11:3] + 9'h0bd;
  assign sel_180034 = $signed({1'h0, add_179929, array_index_179700[2:0]}) < $signed({1'h0, sel_179932}) ? {add_179929, array_index_179700[2:0]} : sel_179932;
  assign add_180036 = array_index_179901[11:1] + 11'h247;
  assign sel_180039 = $signed({1'h0, add_179934, array_index_179799[0]}) < $signed({1'h0, sel_179937}) ? {add_179934, array_index_179799[0]} : sel_179937;
  assign add_180041 = array_index_179904[11:1] + 11'h247;
  assign sel_180044 = $signed({1'h0, add_179939, array_index_179802[0]}) < $signed({1'h0, sel_179942}) ? {add_179939, array_index_179802[0]} : sel_179942;
  assign add_180069 = array_index_180003[11:0] + 12'h247;
  assign sel_180071 = $signed({1'h0, add_179967}) < $signed({1'h0, sel_179969}) ? add_179967 : sel_179969;
  assign add_180074 = array_index_180006[11:0] + 12'h247;
  assign sel_180076 = $signed({1'h0, add_179972}) < $signed({1'h0, sel_179974}) ? add_179972 : sel_179974;
  assign array_index_180105 = set1_unflattened[7'h49];
  assign array_index_180108 = set2_unflattened[7'h49];
  assign add_180112 = array_index_179697[11:1] + 11'h79d;
  assign sel_180114 = $signed({1'h0, add_180010, array_index_179595[0]}) < $signed({1'h0, sel_180012}) ? {add_180010, array_index_179595[0]} : sel_180012;
  assign add_180116 = array_index_179700[11:1] + 11'h79d;
  assign sel_180118 = $signed({1'h0, add_180014, array_index_179598[0]}) < $signed({1'h0, sel_180016}) ? {add_180014, array_index_179598[0]} : sel_180016;
  assign add_180120 = array_index_179799[11:1] + 11'h347;
  assign sel_180122 = $signed({1'h0, add_180018, array_index_179697[0]}) < $signed({1'h0, sel_180020}) ? {add_180018, array_index_179697[0]} : sel_180020;
  assign add_180124 = array_index_179802[11:1] + 11'h347;
  assign sel_180126 = $signed({1'h0, add_180022, array_index_179700[0]}) < $signed({1'h0, sel_180024}) ? {add_180022, array_index_179700[0]} : sel_180024;
  assign add_180128 = array_index_179901[11:3] + 9'h0bd;
  assign sel_180131 = $signed({1'h0, add_180026, array_index_179799[2:0]}) < $signed({1'h0, sel_180029}) ? {add_180026, array_index_179799[2:0]} : sel_180029;
  assign add_180133 = array_index_179904[11:3] + 9'h0bd;
  assign sel_180136 = $signed({1'h0, add_180031, array_index_179802[2:0]}) < $signed({1'h0, sel_180034}) ? {add_180031, array_index_179802[2:0]} : sel_180034;
  assign add_180138 = array_index_180003[11:1] + 11'h247;
  assign sel_180141 = $signed({1'h0, add_180036, array_index_179901[0]}) < $signed({1'h0, sel_180039}) ? {add_180036, array_index_179901[0]} : sel_180039;
  assign add_180143 = array_index_180006[11:1] + 11'h247;
  assign sel_180146 = $signed({1'h0, add_180041, array_index_179904[0]}) < $signed({1'h0, sel_180044}) ? {add_180041, array_index_179904[0]} : sel_180044;
  assign add_180171 = array_index_180105[11:0] + 12'h247;
  assign sel_180173 = $signed({1'h0, add_180069}) < $signed({1'h0, sel_180071}) ? add_180069 : sel_180071;
  assign add_180176 = array_index_180108[11:0] + 12'h247;
  assign sel_180178 = $signed({1'h0, add_180074}) < $signed({1'h0, sel_180076}) ? add_180074 : sel_180076;
  assign array_index_180207 = set1_unflattened[7'h4a];
  assign array_index_180210 = set2_unflattened[7'h4a];
  assign add_180214 = array_index_179799[11:1] + 11'h79d;
  assign sel_180216 = $signed({1'h0, add_180112, array_index_179697[0]}) < $signed({1'h0, sel_180114}) ? {add_180112, array_index_179697[0]} : sel_180114;
  assign add_180218 = array_index_179802[11:1] + 11'h79d;
  assign sel_180220 = $signed({1'h0, add_180116, array_index_179700[0]}) < $signed({1'h0, sel_180118}) ? {add_180116, array_index_179700[0]} : sel_180118;
  assign add_180222 = array_index_179901[11:1] + 11'h347;
  assign sel_180224 = $signed({1'h0, add_180120, array_index_179799[0]}) < $signed({1'h0, sel_180122}) ? {add_180120, array_index_179799[0]} : sel_180122;
  assign add_180226 = array_index_179904[11:1] + 11'h347;
  assign sel_180228 = $signed({1'h0, add_180124, array_index_179802[0]}) < $signed({1'h0, sel_180126}) ? {add_180124, array_index_179802[0]} : sel_180126;
  assign add_180230 = array_index_180003[11:3] + 9'h0bd;
  assign sel_180233 = $signed({1'h0, add_180128, array_index_179901[2:0]}) < $signed({1'h0, sel_180131}) ? {add_180128, array_index_179901[2:0]} : sel_180131;
  assign add_180235 = array_index_180006[11:3] + 9'h0bd;
  assign sel_180238 = $signed({1'h0, add_180133, array_index_179904[2:0]}) < $signed({1'h0, sel_180136}) ? {add_180133, array_index_179904[2:0]} : sel_180136;
  assign add_180240 = array_index_180105[11:1] + 11'h247;
  assign sel_180243 = $signed({1'h0, add_180138, array_index_180003[0]}) < $signed({1'h0, sel_180141}) ? {add_180138, array_index_180003[0]} : sel_180141;
  assign add_180245 = array_index_180108[11:1] + 11'h247;
  assign sel_180248 = $signed({1'h0, add_180143, array_index_180006[0]}) < $signed({1'h0, sel_180146}) ? {add_180143, array_index_180006[0]} : sel_180146;
  assign add_180273 = array_index_180207[11:0] + 12'h247;
  assign sel_180275 = $signed({1'h0, add_180171}) < $signed({1'h0, sel_180173}) ? add_180171 : sel_180173;
  assign add_180278 = array_index_180210[11:0] + 12'h247;
  assign sel_180280 = $signed({1'h0, add_180176}) < $signed({1'h0, sel_180178}) ? add_180176 : sel_180178;
  assign array_index_180309 = set1_unflattened[7'h4b];
  assign array_index_180312 = set2_unflattened[7'h4b];
  assign add_180316 = array_index_179901[11:1] + 11'h79d;
  assign sel_180318 = $signed({1'h0, add_180214, array_index_179799[0]}) < $signed({1'h0, sel_180216}) ? {add_180214, array_index_179799[0]} : sel_180216;
  assign add_180320 = array_index_179904[11:1] + 11'h79d;
  assign sel_180322 = $signed({1'h0, add_180218, array_index_179802[0]}) < $signed({1'h0, sel_180220}) ? {add_180218, array_index_179802[0]} : sel_180220;
  assign add_180324 = array_index_180003[11:1] + 11'h347;
  assign sel_180326 = $signed({1'h0, add_180222, array_index_179901[0]}) < $signed({1'h0, sel_180224}) ? {add_180222, array_index_179901[0]} : sel_180224;
  assign add_180328 = array_index_180006[11:1] + 11'h347;
  assign sel_180330 = $signed({1'h0, add_180226, array_index_179904[0]}) < $signed({1'h0, sel_180228}) ? {add_180226, array_index_179904[0]} : sel_180228;
  assign add_180332 = array_index_180105[11:3] + 9'h0bd;
  assign sel_180335 = $signed({1'h0, add_180230, array_index_180003[2:0]}) < $signed({1'h0, sel_180233}) ? {add_180230, array_index_180003[2:0]} : sel_180233;
  assign add_180337 = array_index_180108[11:3] + 9'h0bd;
  assign sel_180340 = $signed({1'h0, add_180235, array_index_180006[2:0]}) < $signed({1'h0, sel_180238}) ? {add_180235, array_index_180006[2:0]} : sel_180238;
  assign add_180342 = array_index_180207[11:1] + 11'h247;
  assign sel_180345 = $signed({1'h0, add_180240, array_index_180105[0]}) < $signed({1'h0, sel_180243}) ? {add_180240, array_index_180105[0]} : sel_180243;
  assign add_180347 = array_index_180210[11:1] + 11'h247;
  assign sel_180350 = $signed({1'h0, add_180245, array_index_180108[0]}) < $signed({1'h0, sel_180248}) ? {add_180245, array_index_180108[0]} : sel_180248;
  assign add_180375 = array_index_180309[11:0] + 12'h247;
  assign sel_180377 = $signed({1'h0, add_180273}) < $signed({1'h0, sel_180275}) ? add_180273 : sel_180275;
  assign add_180380 = array_index_180312[11:0] + 12'h247;
  assign sel_180382 = $signed({1'h0, add_180278}) < $signed({1'h0, sel_180280}) ? add_180278 : sel_180280;
  assign array_index_180411 = set1_unflattened[7'h4c];
  assign array_index_180414 = set2_unflattened[7'h4c];
  assign add_180418 = array_index_180003[11:1] + 11'h79d;
  assign sel_180420 = $signed({1'h0, add_180316, array_index_179901[0]}) < $signed({1'h0, sel_180318}) ? {add_180316, array_index_179901[0]} : sel_180318;
  assign add_180422 = array_index_180006[11:1] + 11'h79d;
  assign sel_180424 = $signed({1'h0, add_180320, array_index_179904[0]}) < $signed({1'h0, sel_180322}) ? {add_180320, array_index_179904[0]} : sel_180322;
  assign add_180426 = array_index_180105[11:1] + 11'h347;
  assign sel_180428 = $signed({1'h0, add_180324, array_index_180003[0]}) < $signed({1'h0, sel_180326}) ? {add_180324, array_index_180003[0]} : sel_180326;
  assign add_180430 = array_index_180108[11:1] + 11'h347;
  assign sel_180432 = $signed({1'h0, add_180328, array_index_180006[0]}) < $signed({1'h0, sel_180330}) ? {add_180328, array_index_180006[0]} : sel_180330;
  assign add_180434 = array_index_180207[11:3] + 9'h0bd;
  assign sel_180437 = $signed({1'h0, add_180332, array_index_180105[2:0]}) < $signed({1'h0, sel_180335}) ? {add_180332, array_index_180105[2:0]} : sel_180335;
  assign add_180439 = array_index_180210[11:3] + 9'h0bd;
  assign sel_180442 = $signed({1'h0, add_180337, array_index_180108[2:0]}) < $signed({1'h0, sel_180340}) ? {add_180337, array_index_180108[2:0]} : sel_180340;
  assign add_180444 = array_index_180309[11:1] + 11'h247;
  assign sel_180447 = $signed({1'h0, add_180342, array_index_180207[0]}) < $signed({1'h0, sel_180345}) ? {add_180342, array_index_180207[0]} : sel_180345;
  assign add_180449 = array_index_180312[11:1] + 11'h247;
  assign sel_180452 = $signed({1'h0, add_180347, array_index_180210[0]}) < $signed({1'h0, sel_180350}) ? {add_180347, array_index_180210[0]} : sel_180350;
  assign add_180477 = array_index_180411[11:0] + 12'h247;
  assign sel_180479 = $signed({1'h0, add_180375}) < $signed({1'h0, sel_180377}) ? add_180375 : sel_180377;
  assign add_180482 = array_index_180414[11:0] + 12'h247;
  assign sel_180484 = $signed({1'h0, add_180380}) < $signed({1'h0, sel_180382}) ? add_180380 : sel_180382;
  assign array_index_180513 = set1_unflattened[7'h4d];
  assign array_index_180516 = set2_unflattened[7'h4d];
  assign add_180520 = array_index_180105[11:1] + 11'h79d;
  assign sel_180522 = $signed({1'h0, add_180418, array_index_180003[0]}) < $signed({1'h0, sel_180420}) ? {add_180418, array_index_180003[0]} : sel_180420;
  assign add_180524 = array_index_180108[11:1] + 11'h79d;
  assign sel_180526 = $signed({1'h0, add_180422, array_index_180006[0]}) < $signed({1'h0, sel_180424}) ? {add_180422, array_index_180006[0]} : sel_180424;
  assign add_180528 = array_index_180207[11:1] + 11'h347;
  assign sel_180530 = $signed({1'h0, add_180426, array_index_180105[0]}) < $signed({1'h0, sel_180428}) ? {add_180426, array_index_180105[0]} : sel_180428;
  assign add_180532 = array_index_180210[11:1] + 11'h347;
  assign sel_180534 = $signed({1'h0, add_180430, array_index_180108[0]}) < $signed({1'h0, sel_180432}) ? {add_180430, array_index_180108[0]} : sel_180432;
  assign add_180536 = array_index_180309[11:3] + 9'h0bd;
  assign sel_180539 = $signed({1'h0, add_180434, array_index_180207[2:0]}) < $signed({1'h0, sel_180437}) ? {add_180434, array_index_180207[2:0]} : sel_180437;
  assign add_180541 = array_index_180312[11:3] + 9'h0bd;
  assign sel_180544 = $signed({1'h0, add_180439, array_index_180210[2:0]}) < $signed({1'h0, sel_180442}) ? {add_180439, array_index_180210[2:0]} : sel_180442;
  assign add_180546 = array_index_180411[11:1] + 11'h247;
  assign sel_180549 = $signed({1'h0, add_180444, array_index_180309[0]}) < $signed({1'h0, sel_180447}) ? {add_180444, array_index_180309[0]} : sel_180447;
  assign add_180551 = array_index_180414[11:1] + 11'h247;
  assign sel_180554 = $signed({1'h0, add_180449, array_index_180312[0]}) < $signed({1'h0, sel_180452}) ? {add_180449, array_index_180312[0]} : sel_180452;
  assign add_180579 = array_index_180513[11:0] + 12'h247;
  assign sel_180581 = $signed({1'h0, add_180477}) < $signed({1'h0, sel_180479}) ? add_180477 : sel_180479;
  assign add_180584 = array_index_180516[11:0] + 12'h247;
  assign sel_180586 = $signed({1'h0, add_180482}) < $signed({1'h0, sel_180484}) ? add_180482 : sel_180484;
  assign array_index_180615 = set1_unflattened[7'h4e];
  assign array_index_180618 = set2_unflattened[7'h4e];
  assign add_180622 = array_index_180207[11:1] + 11'h79d;
  assign sel_180624 = $signed({1'h0, add_180520, array_index_180105[0]}) < $signed({1'h0, sel_180522}) ? {add_180520, array_index_180105[0]} : sel_180522;
  assign add_180626 = array_index_180210[11:1] + 11'h79d;
  assign sel_180628 = $signed({1'h0, add_180524, array_index_180108[0]}) < $signed({1'h0, sel_180526}) ? {add_180524, array_index_180108[0]} : sel_180526;
  assign add_180630 = array_index_180309[11:1] + 11'h347;
  assign sel_180632 = $signed({1'h0, add_180528, array_index_180207[0]}) < $signed({1'h0, sel_180530}) ? {add_180528, array_index_180207[0]} : sel_180530;
  assign add_180634 = array_index_180312[11:1] + 11'h347;
  assign sel_180636 = $signed({1'h0, add_180532, array_index_180210[0]}) < $signed({1'h0, sel_180534}) ? {add_180532, array_index_180210[0]} : sel_180534;
  assign add_180638 = array_index_180411[11:3] + 9'h0bd;
  assign sel_180641 = $signed({1'h0, add_180536, array_index_180309[2:0]}) < $signed({1'h0, sel_180539}) ? {add_180536, array_index_180309[2:0]} : sel_180539;
  assign add_180643 = array_index_180414[11:3] + 9'h0bd;
  assign sel_180646 = $signed({1'h0, add_180541, array_index_180312[2:0]}) < $signed({1'h0, sel_180544}) ? {add_180541, array_index_180312[2:0]} : sel_180544;
  assign add_180648 = array_index_180513[11:1] + 11'h247;
  assign sel_180651 = $signed({1'h0, add_180546, array_index_180411[0]}) < $signed({1'h0, sel_180549}) ? {add_180546, array_index_180411[0]} : sel_180549;
  assign add_180653 = array_index_180516[11:1] + 11'h247;
  assign sel_180656 = $signed({1'h0, add_180551, array_index_180414[0]}) < $signed({1'h0, sel_180554}) ? {add_180551, array_index_180414[0]} : sel_180554;
  assign add_180681 = array_index_180615[11:0] + 12'h247;
  assign sel_180683 = $signed({1'h0, add_180579}) < $signed({1'h0, sel_180581}) ? add_180579 : sel_180581;
  assign add_180686 = array_index_180618[11:0] + 12'h247;
  assign sel_180688 = $signed({1'h0, add_180584}) < $signed({1'h0, sel_180586}) ? add_180584 : sel_180586;
  assign array_index_180717 = set1_unflattened[7'h4f];
  assign array_index_180720 = set2_unflattened[7'h4f];
  assign add_180724 = array_index_180309[11:1] + 11'h79d;
  assign sel_180726 = $signed({1'h0, add_180622, array_index_180207[0]}) < $signed({1'h0, sel_180624}) ? {add_180622, array_index_180207[0]} : sel_180624;
  assign add_180728 = array_index_180312[11:1] + 11'h79d;
  assign sel_180730 = $signed({1'h0, add_180626, array_index_180210[0]}) < $signed({1'h0, sel_180628}) ? {add_180626, array_index_180210[0]} : sel_180628;
  assign add_180732 = array_index_180411[11:1] + 11'h347;
  assign sel_180734 = $signed({1'h0, add_180630, array_index_180309[0]}) < $signed({1'h0, sel_180632}) ? {add_180630, array_index_180309[0]} : sel_180632;
  assign add_180736 = array_index_180414[11:1] + 11'h347;
  assign sel_180738 = $signed({1'h0, add_180634, array_index_180312[0]}) < $signed({1'h0, sel_180636}) ? {add_180634, array_index_180312[0]} : sel_180636;
  assign add_180740 = array_index_180513[11:3] + 9'h0bd;
  assign sel_180743 = $signed({1'h0, add_180638, array_index_180411[2:0]}) < $signed({1'h0, sel_180641}) ? {add_180638, array_index_180411[2:0]} : sel_180641;
  assign add_180745 = array_index_180516[11:3] + 9'h0bd;
  assign sel_180748 = $signed({1'h0, add_180643, array_index_180414[2:0]}) < $signed({1'h0, sel_180646}) ? {add_180643, array_index_180414[2:0]} : sel_180646;
  assign add_180750 = array_index_180615[11:1] + 11'h247;
  assign sel_180753 = $signed({1'h0, add_180648, array_index_180513[0]}) < $signed({1'h0, sel_180651}) ? {add_180648, array_index_180513[0]} : sel_180651;
  assign add_180755 = array_index_180618[11:1] + 11'h247;
  assign sel_180758 = $signed({1'h0, add_180653, array_index_180516[0]}) < $signed({1'h0, sel_180656}) ? {add_180653, array_index_180516[0]} : sel_180656;
  assign add_180783 = array_index_180717[11:0] + 12'h247;
  assign sel_180785 = $signed({1'h0, add_180681}) < $signed({1'h0, sel_180683}) ? add_180681 : sel_180683;
  assign add_180788 = array_index_180720[11:0] + 12'h247;
  assign sel_180790 = $signed({1'h0, add_180686}) < $signed({1'h0, sel_180688}) ? add_180686 : sel_180688;
  assign array_index_180819 = set1_unflattened[7'h50];
  assign array_index_180822 = set2_unflattened[7'h50];
  assign add_180826 = array_index_180411[11:1] + 11'h79d;
  assign sel_180828 = $signed({1'h0, add_180724, array_index_180309[0]}) < $signed({1'h0, sel_180726}) ? {add_180724, array_index_180309[0]} : sel_180726;
  assign add_180830 = array_index_180414[11:1] + 11'h79d;
  assign sel_180832 = $signed({1'h0, add_180728, array_index_180312[0]}) < $signed({1'h0, sel_180730}) ? {add_180728, array_index_180312[0]} : sel_180730;
  assign add_180834 = array_index_180513[11:1] + 11'h347;
  assign sel_180836 = $signed({1'h0, add_180732, array_index_180411[0]}) < $signed({1'h0, sel_180734}) ? {add_180732, array_index_180411[0]} : sel_180734;
  assign add_180838 = array_index_180516[11:1] + 11'h347;
  assign sel_180840 = $signed({1'h0, add_180736, array_index_180414[0]}) < $signed({1'h0, sel_180738}) ? {add_180736, array_index_180414[0]} : sel_180738;
  assign add_180842 = array_index_180615[11:3] + 9'h0bd;
  assign sel_180845 = $signed({1'h0, add_180740, array_index_180513[2:0]}) < $signed({1'h0, sel_180743}) ? {add_180740, array_index_180513[2:0]} : sel_180743;
  assign add_180847 = array_index_180618[11:3] + 9'h0bd;
  assign sel_180850 = $signed({1'h0, add_180745, array_index_180516[2:0]}) < $signed({1'h0, sel_180748}) ? {add_180745, array_index_180516[2:0]} : sel_180748;
  assign add_180852 = array_index_180717[11:1] + 11'h247;
  assign sel_180855 = $signed({1'h0, add_180750, array_index_180615[0]}) < $signed({1'h0, sel_180753}) ? {add_180750, array_index_180615[0]} : sel_180753;
  assign add_180857 = array_index_180720[11:1] + 11'h247;
  assign sel_180860 = $signed({1'h0, add_180755, array_index_180618[0]}) < $signed({1'h0, sel_180758}) ? {add_180755, array_index_180618[0]} : sel_180758;
  assign add_180885 = array_index_180819[11:0] + 12'h247;
  assign sel_180887 = $signed({1'h0, add_180783}) < $signed({1'h0, sel_180785}) ? add_180783 : sel_180785;
  assign add_180890 = array_index_180822[11:0] + 12'h247;
  assign sel_180892 = $signed({1'h0, add_180788}) < $signed({1'h0, sel_180790}) ? add_180788 : sel_180790;
  assign array_index_180921 = set1_unflattened[7'h51];
  assign array_index_180924 = set2_unflattened[7'h51];
  assign add_180928 = array_index_180513[11:1] + 11'h79d;
  assign sel_180930 = $signed({1'h0, add_180826, array_index_180411[0]}) < $signed({1'h0, sel_180828}) ? {add_180826, array_index_180411[0]} : sel_180828;
  assign add_180932 = array_index_180516[11:1] + 11'h79d;
  assign sel_180934 = $signed({1'h0, add_180830, array_index_180414[0]}) < $signed({1'h0, sel_180832}) ? {add_180830, array_index_180414[0]} : sel_180832;
  assign add_180936 = array_index_180615[11:1] + 11'h347;
  assign sel_180938 = $signed({1'h0, add_180834, array_index_180513[0]}) < $signed({1'h0, sel_180836}) ? {add_180834, array_index_180513[0]} : sel_180836;
  assign add_180940 = array_index_180618[11:1] + 11'h347;
  assign sel_180942 = $signed({1'h0, add_180838, array_index_180516[0]}) < $signed({1'h0, sel_180840}) ? {add_180838, array_index_180516[0]} : sel_180840;
  assign add_180944 = array_index_180717[11:3] + 9'h0bd;
  assign sel_180947 = $signed({1'h0, add_180842, array_index_180615[2:0]}) < $signed({1'h0, sel_180845}) ? {add_180842, array_index_180615[2:0]} : sel_180845;
  assign add_180949 = array_index_180720[11:3] + 9'h0bd;
  assign sel_180952 = $signed({1'h0, add_180847, array_index_180618[2:0]}) < $signed({1'h0, sel_180850}) ? {add_180847, array_index_180618[2:0]} : sel_180850;
  assign add_180954 = array_index_180819[11:1] + 11'h247;
  assign sel_180957 = $signed({1'h0, add_180852, array_index_180717[0]}) < $signed({1'h0, sel_180855}) ? {add_180852, array_index_180717[0]} : sel_180855;
  assign add_180959 = array_index_180822[11:1] + 11'h247;
  assign sel_180962 = $signed({1'h0, add_180857, array_index_180720[0]}) < $signed({1'h0, sel_180860}) ? {add_180857, array_index_180720[0]} : sel_180860;
  assign add_180987 = array_index_180921[11:0] + 12'h247;
  assign sel_180989 = $signed({1'h0, add_180885}) < $signed({1'h0, sel_180887}) ? add_180885 : sel_180887;
  assign add_180992 = array_index_180924[11:0] + 12'h247;
  assign sel_180994 = $signed({1'h0, add_180890}) < $signed({1'h0, sel_180892}) ? add_180890 : sel_180892;
  assign array_index_181023 = set1_unflattened[7'h52];
  assign array_index_181026 = set2_unflattened[7'h52];
  assign add_181030 = array_index_180615[11:1] + 11'h79d;
  assign sel_181032 = $signed({1'h0, add_180928, array_index_180513[0]}) < $signed({1'h0, sel_180930}) ? {add_180928, array_index_180513[0]} : sel_180930;
  assign add_181034 = array_index_180618[11:1] + 11'h79d;
  assign sel_181036 = $signed({1'h0, add_180932, array_index_180516[0]}) < $signed({1'h0, sel_180934}) ? {add_180932, array_index_180516[0]} : sel_180934;
  assign add_181038 = array_index_180717[11:1] + 11'h347;
  assign sel_181040 = $signed({1'h0, add_180936, array_index_180615[0]}) < $signed({1'h0, sel_180938}) ? {add_180936, array_index_180615[0]} : sel_180938;
  assign add_181042 = array_index_180720[11:1] + 11'h347;
  assign sel_181044 = $signed({1'h0, add_180940, array_index_180618[0]}) < $signed({1'h0, sel_180942}) ? {add_180940, array_index_180618[0]} : sel_180942;
  assign add_181046 = array_index_180819[11:3] + 9'h0bd;
  assign sel_181049 = $signed({1'h0, add_180944, array_index_180717[2:0]}) < $signed({1'h0, sel_180947}) ? {add_180944, array_index_180717[2:0]} : sel_180947;
  assign add_181051 = array_index_180822[11:3] + 9'h0bd;
  assign sel_181054 = $signed({1'h0, add_180949, array_index_180720[2:0]}) < $signed({1'h0, sel_180952}) ? {add_180949, array_index_180720[2:0]} : sel_180952;
  assign add_181056 = array_index_180921[11:1] + 11'h247;
  assign sel_181059 = $signed({1'h0, add_180954, array_index_180819[0]}) < $signed({1'h0, sel_180957}) ? {add_180954, array_index_180819[0]} : sel_180957;
  assign add_181061 = array_index_180924[11:1] + 11'h247;
  assign sel_181064 = $signed({1'h0, add_180959, array_index_180822[0]}) < $signed({1'h0, sel_180962}) ? {add_180959, array_index_180822[0]} : sel_180962;
  assign add_181089 = array_index_181023[11:0] + 12'h247;
  assign sel_181091 = $signed({1'h0, add_180987}) < $signed({1'h0, sel_180989}) ? add_180987 : sel_180989;
  assign add_181094 = array_index_181026[11:0] + 12'h247;
  assign sel_181096 = $signed({1'h0, add_180992}) < $signed({1'h0, sel_180994}) ? add_180992 : sel_180994;
  assign array_index_181125 = set1_unflattened[7'h53];
  assign array_index_181128 = set2_unflattened[7'h53];
  assign add_181132 = array_index_180717[11:1] + 11'h79d;
  assign sel_181134 = $signed({1'h0, add_181030, array_index_180615[0]}) < $signed({1'h0, sel_181032}) ? {add_181030, array_index_180615[0]} : sel_181032;
  assign add_181136 = array_index_180720[11:1] + 11'h79d;
  assign sel_181138 = $signed({1'h0, add_181034, array_index_180618[0]}) < $signed({1'h0, sel_181036}) ? {add_181034, array_index_180618[0]} : sel_181036;
  assign add_181140 = array_index_180819[11:1] + 11'h347;
  assign sel_181142 = $signed({1'h0, add_181038, array_index_180717[0]}) < $signed({1'h0, sel_181040}) ? {add_181038, array_index_180717[0]} : sel_181040;
  assign add_181144 = array_index_180822[11:1] + 11'h347;
  assign sel_181146 = $signed({1'h0, add_181042, array_index_180720[0]}) < $signed({1'h0, sel_181044}) ? {add_181042, array_index_180720[0]} : sel_181044;
  assign add_181148 = array_index_180921[11:3] + 9'h0bd;
  assign sel_181151 = $signed({1'h0, add_181046, array_index_180819[2:0]}) < $signed({1'h0, sel_181049}) ? {add_181046, array_index_180819[2:0]} : sel_181049;
  assign add_181153 = array_index_180924[11:3] + 9'h0bd;
  assign sel_181156 = $signed({1'h0, add_181051, array_index_180822[2:0]}) < $signed({1'h0, sel_181054}) ? {add_181051, array_index_180822[2:0]} : sel_181054;
  assign add_181158 = array_index_181023[11:1] + 11'h247;
  assign sel_181161 = $signed({1'h0, add_181056, array_index_180921[0]}) < $signed({1'h0, sel_181059}) ? {add_181056, array_index_180921[0]} : sel_181059;
  assign add_181163 = array_index_181026[11:1] + 11'h247;
  assign sel_181166 = $signed({1'h0, add_181061, array_index_180924[0]}) < $signed({1'h0, sel_181064}) ? {add_181061, array_index_180924[0]} : sel_181064;
  assign add_181191 = array_index_181125[11:0] + 12'h247;
  assign sel_181193 = $signed({1'h0, add_181089}) < $signed({1'h0, sel_181091}) ? add_181089 : sel_181091;
  assign add_181196 = array_index_181128[11:0] + 12'h247;
  assign sel_181198 = $signed({1'h0, add_181094}) < $signed({1'h0, sel_181096}) ? add_181094 : sel_181096;
  assign array_index_181227 = set1_unflattened[7'h54];
  assign array_index_181230 = set2_unflattened[7'h54];
  assign add_181234 = array_index_180819[11:1] + 11'h79d;
  assign sel_181236 = $signed({1'h0, add_181132, array_index_180717[0]}) < $signed({1'h0, sel_181134}) ? {add_181132, array_index_180717[0]} : sel_181134;
  assign add_181238 = array_index_180822[11:1] + 11'h79d;
  assign sel_181240 = $signed({1'h0, add_181136, array_index_180720[0]}) < $signed({1'h0, sel_181138}) ? {add_181136, array_index_180720[0]} : sel_181138;
  assign add_181242 = array_index_180921[11:1] + 11'h347;
  assign sel_181244 = $signed({1'h0, add_181140, array_index_180819[0]}) < $signed({1'h0, sel_181142}) ? {add_181140, array_index_180819[0]} : sel_181142;
  assign add_181246 = array_index_180924[11:1] + 11'h347;
  assign sel_181248 = $signed({1'h0, add_181144, array_index_180822[0]}) < $signed({1'h0, sel_181146}) ? {add_181144, array_index_180822[0]} : sel_181146;
  assign add_181250 = array_index_181023[11:3] + 9'h0bd;
  assign sel_181253 = $signed({1'h0, add_181148, array_index_180921[2:0]}) < $signed({1'h0, sel_181151}) ? {add_181148, array_index_180921[2:0]} : sel_181151;
  assign add_181255 = array_index_181026[11:3] + 9'h0bd;
  assign sel_181258 = $signed({1'h0, add_181153, array_index_180924[2:0]}) < $signed({1'h0, sel_181156}) ? {add_181153, array_index_180924[2:0]} : sel_181156;
  assign add_181260 = array_index_181125[11:1] + 11'h247;
  assign sel_181263 = $signed({1'h0, add_181158, array_index_181023[0]}) < $signed({1'h0, sel_181161}) ? {add_181158, array_index_181023[0]} : sel_181161;
  assign add_181265 = array_index_181128[11:1] + 11'h247;
  assign sel_181268 = $signed({1'h0, add_181163, array_index_181026[0]}) < $signed({1'h0, sel_181166}) ? {add_181163, array_index_181026[0]} : sel_181166;
  assign add_181293 = array_index_181227[11:0] + 12'h247;
  assign sel_181295 = $signed({1'h0, add_181191}) < $signed({1'h0, sel_181193}) ? add_181191 : sel_181193;
  assign add_181298 = array_index_181230[11:0] + 12'h247;
  assign sel_181300 = $signed({1'h0, add_181196}) < $signed({1'h0, sel_181198}) ? add_181196 : sel_181198;
  assign array_index_181329 = set1_unflattened[7'h55];
  assign array_index_181332 = set2_unflattened[7'h55];
  assign add_181336 = array_index_180921[11:1] + 11'h79d;
  assign sel_181338 = $signed({1'h0, add_181234, array_index_180819[0]}) < $signed({1'h0, sel_181236}) ? {add_181234, array_index_180819[0]} : sel_181236;
  assign add_181340 = array_index_180924[11:1] + 11'h79d;
  assign sel_181342 = $signed({1'h0, add_181238, array_index_180822[0]}) < $signed({1'h0, sel_181240}) ? {add_181238, array_index_180822[0]} : sel_181240;
  assign add_181344 = array_index_181023[11:1] + 11'h347;
  assign sel_181346 = $signed({1'h0, add_181242, array_index_180921[0]}) < $signed({1'h0, sel_181244}) ? {add_181242, array_index_180921[0]} : sel_181244;
  assign add_181348 = array_index_181026[11:1] + 11'h347;
  assign sel_181350 = $signed({1'h0, add_181246, array_index_180924[0]}) < $signed({1'h0, sel_181248}) ? {add_181246, array_index_180924[0]} : sel_181248;
  assign add_181352 = array_index_181125[11:3] + 9'h0bd;
  assign sel_181355 = $signed({1'h0, add_181250, array_index_181023[2:0]}) < $signed({1'h0, sel_181253}) ? {add_181250, array_index_181023[2:0]} : sel_181253;
  assign add_181357 = array_index_181128[11:3] + 9'h0bd;
  assign sel_181360 = $signed({1'h0, add_181255, array_index_181026[2:0]}) < $signed({1'h0, sel_181258}) ? {add_181255, array_index_181026[2:0]} : sel_181258;
  assign add_181362 = array_index_181227[11:1] + 11'h247;
  assign sel_181365 = $signed({1'h0, add_181260, array_index_181125[0]}) < $signed({1'h0, sel_181263}) ? {add_181260, array_index_181125[0]} : sel_181263;
  assign add_181367 = array_index_181230[11:1] + 11'h247;
  assign sel_181370 = $signed({1'h0, add_181265, array_index_181128[0]}) < $signed({1'h0, sel_181268}) ? {add_181265, array_index_181128[0]} : sel_181268;
  assign add_181395 = array_index_181329[11:0] + 12'h247;
  assign sel_181397 = $signed({1'h0, add_181293}) < $signed({1'h0, sel_181295}) ? add_181293 : sel_181295;
  assign add_181400 = array_index_181332[11:0] + 12'h247;
  assign sel_181402 = $signed({1'h0, add_181298}) < $signed({1'h0, sel_181300}) ? add_181298 : sel_181300;
  assign array_index_181431 = set1_unflattened[7'h56];
  assign array_index_181434 = set2_unflattened[7'h56];
  assign add_181438 = array_index_181023[11:1] + 11'h79d;
  assign sel_181440 = $signed({1'h0, add_181336, array_index_180921[0]}) < $signed({1'h0, sel_181338}) ? {add_181336, array_index_180921[0]} : sel_181338;
  assign add_181442 = array_index_181026[11:1] + 11'h79d;
  assign sel_181444 = $signed({1'h0, add_181340, array_index_180924[0]}) < $signed({1'h0, sel_181342}) ? {add_181340, array_index_180924[0]} : sel_181342;
  assign add_181446 = array_index_181125[11:1] + 11'h347;
  assign sel_181448 = $signed({1'h0, add_181344, array_index_181023[0]}) < $signed({1'h0, sel_181346}) ? {add_181344, array_index_181023[0]} : sel_181346;
  assign add_181450 = array_index_181128[11:1] + 11'h347;
  assign sel_181452 = $signed({1'h0, add_181348, array_index_181026[0]}) < $signed({1'h0, sel_181350}) ? {add_181348, array_index_181026[0]} : sel_181350;
  assign add_181454 = array_index_181227[11:3] + 9'h0bd;
  assign sel_181457 = $signed({1'h0, add_181352, array_index_181125[2:0]}) < $signed({1'h0, sel_181355}) ? {add_181352, array_index_181125[2:0]} : sel_181355;
  assign add_181459 = array_index_181230[11:3] + 9'h0bd;
  assign sel_181462 = $signed({1'h0, add_181357, array_index_181128[2:0]}) < $signed({1'h0, sel_181360}) ? {add_181357, array_index_181128[2:0]} : sel_181360;
  assign add_181464 = array_index_181329[11:1] + 11'h247;
  assign sel_181467 = $signed({1'h0, add_181362, array_index_181227[0]}) < $signed({1'h0, sel_181365}) ? {add_181362, array_index_181227[0]} : sel_181365;
  assign add_181469 = array_index_181332[11:1] + 11'h247;
  assign sel_181472 = $signed({1'h0, add_181367, array_index_181230[0]}) < $signed({1'h0, sel_181370}) ? {add_181367, array_index_181230[0]} : sel_181370;
  assign add_181497 = array_index_181431[11:0] + 12'h247;
  assign sel_181499 = $signed({1'h0, add_181395}) < $signed({1'h0, sel_181397}) ? add_181395 : sel_181397;
  assign add_181502 = array_index_181434[11:0] + 12'h247;
  assign sel_181504 = $signed({1'h0, add_181400}) < $signed({1'h0, sel_181402}) ? add_181400 : sel_181402;
  assign array_index_181533 = set1_unflattened[7'h57];
  assign array_index_181536 = set2_unflattened[7'h57];
  assign add_181540 = array_index_181125[11:1] + 11'h79d;
  assign sel_181542 = $signed({1'h0, add_181438, array_index_181023[0]}) < $signed({1'h0, sel_181440}) ? {add_181438, array_index_181023[0]} : sel_181440;
  assign add_181544 = array_index_181128[11:1] + 11'h79d;
  assign sel_181546 = $signed({1'h0, add_181442, array_index_181026[0]}) < $signed({1'h0, sel_181444}) ? {add_181442, array_index_181026[0]} : sel_181444;
  assign add_181548 = array_index_181227[11:1] + 11'h347;
  assign sel_181550 = $signed({1'h0, add_181446, array_index_181125[0]}) < $signed({1'h0, sel_181448}) ? {add_181446, array_index_181125[0]} : sel_181448;
  assign add_181552 = array_index_181230[11:1] + 11'h347;
  assign sel_181554 = $signed({1'h0, add_181450, array_index_181128[0]}) < $signed({1'h0, sel_181452}) ? {add_181450, array_index_181128[0]} : sel_181452;
  assign add_181556 = array_index_181329[11:3] + 9'h0bd;
  assign sel_181559 = $signed({1'h0, add_181454, array_index_181227[2:0]}) < $signed({1'h0, sel_181457}) ? {add_181454, array_index_181227[2:0]} : sel_181457;
  assign add_181561 = array_index_181332[11:3] + 9'h0bd;
  assign sel_181564 = $signed({1'h0, add_181459, array_index_181230[2:0]}) < $signed({1'h0, sel_181462}) ? {add_181459, array_index_181230[2:0]} : sel_181462;
  assign add_181566 = array_index_181431[11:1] + 11'h247;
  assign sel_181569 = $signed({1'h0, add_181464, array_index_181329[0]}) < $signed({1'h0, sel_181467}) ? {add_181464, array_index_181329[0]} : sel_181467;
  assign add_181571 = array_index_181434[11:1] + 11'h247;
  assign sel_181574 = $signed({1'h0, add_181469, array_index_181332[0]}) < $signed({1'h0, sel_181472}) ? {add_181469, array_index_181332[0]} : sel_181472;
  assign add_181599 = array_index_181533[11:0] + 12'h247;
  assign sel_181601 = $signed({1'h0, add_181497}) < $signed({1'h0, sel_181499}) ? add_181497 : sel_181499;
  assign add_181604 = array_index_181536[11:0] + 12'h247;
  assign sel_181606 = $signed({1'h0, add_181502}) < $signed({1'h0, sel_181504}) ? add_181502 : sel_181504;
  assign array_index_181635 = set1_unflattened[7'h58];
  assign array_index_181638 = set2_unflattened[7'h58];
  assign add_181642 = array_index_181227[11:1] + 11'h79d;
  assign sel_181644 = $signed({1'h0, add_181540, array_index_181125[0]}) < $signed({1'h0, sel_181542}) ? {add_181540, array_index_181125[0]} : sel_181542;
  assign add_181646 = array_index_181230[11:1] + 11'h79d;
  assign sel_181648 = $signed({1'h0, add_181544, array_index_181128[0]}) < $signed({1'h0, sel_181546}) ? {add_181544, array_index_181128[0]} : sel_181546;
  assign add_181650 = array_index_181329[11:1] + 11'h347;
  assign sel_181652 = $signed({1'h0, add_181548, array_index_181227[0]}) < $signed({1'h0, sel_181550}) ? {add_181548, array_index_181227[0]} : sel_181550;
  assign add_181654 = array_index_181332[11:1] + 11'h347;
  assign sel_181656 = $signed({1'h0, add_181552, array_index_181230[0]}) < $signed({1'h0, sel_181554}) ? {add_181552, array_index_181230[0]} : sel_181554;
  assign add_181658 = array_index_181431[11:3] + 9'h0bd;
  assign sel_181661 = $signed({1'h0, add_181556, array_index_181329[2:0]}) < $signed({1'h0, sel_181559}) ? {add_181556, array_index_181329[2:0]} : sel_181559;
  assign add_181663 = array_index_181434[11:3] + 9'h0bd;
  assign sel_181666 = $signed({1'h0, add_181561, array_index_181332[2:0]}) < $signed({1'h0, sel_181564}) ? {add_181561, array_index_181332[2:0]} : sel_181564;
  assign add_181668 = array_index_181533[11:1] + 11'h247;
  assign sel_181671 = $signed({1'h0, add_181566, array_index_181431[0]}) < $signed({1'h0, sel_181569}) ? {add_181566, array_index_181431[0]} : sel_181569;
  assign add_181673 = array_index_181536[11:1] + 11'h247;
  assign sel_181676 = $signed({1'h0, add_181571, array_index_181434[0]}) < $signed({1'h0, sel_181574}) ? {add_181571, array_index_181434[0]} : sel_181574;
  assign add_181701 = array_index_181635[11:0] + 12'h247;
  assign sel_181703 = $signed({1'h0, add_181599}) < $signed({1'h0, sel_181601}) ? add_181599 : sel_181601;
  assign add_181706 = array_index_181638[11:0] + 12'h247;
  assign sel_181708 = $signed({1'h0, add_181604}) < $signed({1'h0, sel_181606}) ? add_181604 : sel_181606;
  assign array_index_181737 = set1_unflattened[7'h59];
  assign array_index_181740 = set2_unflattened[7'h59];
  assign add_181744 = array_index_181329[11:1] + 11'h79d;
  assign sel_181746 = $signed({1'h0, add_181642, array_index_181227[0]}) < $signed({1'h0, sel_181644}) ? {add_181642, array_index_181227[0]} : sel_181644;
  assign add_181748 = array_index_181332[11:1] + 11'h79d;
  assign sel_181750 = $signed({1'h0, add_181646, array_index_181230[0]}) < $signed({1'h0, sel_181648}) ? {add_181646, array_index_181230[0]} : sel_181648;
  assign add_181752 = array_index_181431[11:1] + 11'h347;
  assign sel_181754 = $signed({1'h0, add_181650, array_index_181329[0]}) < $signed({1'h0, sel_181652}) ? {add_181650, array_index_181329[0]} : sel_181652;
  assign add_181756 = array_index_181434[11:1] + 11'h347;
  assign sel_181758 = $signed({1'h0, add_181654, array_index_181332[0]}) < $signed({1'h0, sel_181656}) ? {add_181654, array_index_181332[0]} : sel_181656;
  assign add_181760 = array_index_181533[11:3] + 9'h0bd;
  assign sel_181763 = $signed({1'h0, add_181658, array_index_181431[2:0]}) < $signed({1'h0, sel_181661}) ? {add_181658, array_index_181431[2:0]} : sel_181661;
  assign add_181765 = array_index_181536[11:3] + 9'h0bd;
  assign sel_181768 = $signed({1'h0, add_181663, array_index_181434[2:0]}) < $signed({1'h0, sel_181666}) ? {add_181663, array_index_181434[2:0]} : sel_181666;
  assign add_181770 = array_index_181635[11:1] + 11'h247;
  assign sel_181773 = $signed({1'h0, add_181668, array_index_181533[0]}) < $signed({1'h0, sel_181671}) ? {add_181668, array_index_181533[0]} : sel_181671;
  assign add_181775 = array_index_181638[11:1] + 11'h247;
  assign sel_181778 = $signed({1'h0, add_181673, array_index_181536[0]}) < $signed({1'h0, sel_181676}) ? {add_181673, array_index_181536[0]} : sel_181676;
  assign add_181803 = array_index_181737[11:0] + 12'h247;
  assign sel_181805 = $signed({1'h0, add_181701}) < $signed({1'h0, sel_181703}) ? add_181701 : sel_181703;
  assign add_181808 = array_index_181740[11:0] + 12'h247;
  assign sel_181810 = $signed({1'h0, add_181706}) < $signed({1'h0, sel_181708}) ? add_181706 : sel_181708;
  assign array_index_181839 = set1_unflattened[7'h5a];
  assign array_index_181842 = set2_unflattened[7'h5a];
  assign add_181846 = array_index_181431[11:1] + 11'h79d;
  assign sel_181848 = $signed({1'h0, add_181744, array_index_181329[0]}) < $signed({1'h0, sel_181746}) ? {add_181744, array_index_181329[0]} : sel_181746;
  assign add_181850 = array_index_181434[11:1] + 11'h79d;
  assign sel_181852 = $signed({1'h0, add_181748, array_index_181332[0]}) < $signed({1'h0, sel_181750}) ? {add_181748, array_index_181332[0]} : sel_181750;
  assign add_181854 = array_index_181533[11:1] + 11'h347;
  assign sel_181856 = $signed({1'h0, add_181752, array_index_181431[0]}) < $signed({1'h0, sel_181754}) ? {add_181752, array_index_181431[0]} : sel_181754;
  assign add_181858 = array_index_181536[11:1] + 11'h347;
  assign sel_181860 = $signed({1'h0, add_181756, array_index_181434[0]}) < $signed({1'h0, sel_181758}) ? {add_181756, array_index_181434[0]} : sel_181758;
  assign add_181862 = array_index_181635[11:3] + 9'h0bd;
  assign sel_181865 = $signed({1'h0, add_181760, array_index_181533[2:0]}) < $signed({1'h0, sel_181763}) ? {add_181760, array_index_181533[2:0]} : sel_181763;
  assign add_181867 = array_index_181638[11:3] + 9'h0bd;
  assign sel_181870 = $signed({1'h0, add_181765, array_index_181536[2:0]}) < $signed({1'h0, sel_181768}) ? {add_181765, array_index_181536[2:0]} : sel_181768;
  assign add_181872 = array_index_181737[11:1] + 11'h247;
  assign sel_181875 = $signed({1'h0, add_181770, array_index_181635[0]}) < $signed({1'h0, sel_181773}) ? {add_181770, array_index_181635[0]} : sel_181773;
  assign add_181877 = array_index_181740[11:1] + 11'h247;
  assign sel_181880 = $signed({1'h0, add_181775, array_index_181638[0]}) < $signed({1'h0, sel_181778}) ? {add_181775, array_index_181638[0]} : sel_181778;
  assign add_181905 = array_index_181839[11:0] + 12'h247;
  assign sel_181907 = $signed({1'h0, add_181803}) < $signed({1'h0, sel_181805}) ? add_181803 : sel_181805;
  assign add_181910 = array_index_181842[11:0] + 12'h247;
  assign sel_181912 = $signed({1'h0, add_181808}) < $signed({1'h0, sel_181810}) ? add_181808 : sel_181810;
  assign array_index_181941 = set1_unflattened[7'h5b];
  assign array_index_181944 = set2_unflattened[7'h5b];
  assign add_181948 = array_index_181533[11:1] + 11'h79d;
  assign sel_181950 = $signed({1'h0, add_181846, array_index_181431[0]}) < $signed({1'h0, sel_181848}) ? {add_181846, array_index_181431[0]} : sel_181848;
  assign add_181952 = array_index_181536[11:1] + 11'h79d;
  assign sel_181954 = $signed({1'h0, add_181850, array_index_181434[0]}) < $signed({1'h0, sel_181852}) ? {add_181850, array_index_181434[0]} : sel_181852;
  assign add_181956 = array_index_181635[11:1] + 11'h347;
  assign sel_181958 = $signed({1'h0, add_181854, array_index_181533[0]}) < $signed({1'h0, sel_181856}) ? {add_181854, array_index_181533[0]} : sel_181856;
  assign add_181960 = array_index_181638[11:1] + 11'h347;
  assign sel_181962 = $signed({1'h0, add_181858, array_index_181536[0]}) < $signed({1'h0, sel_181860}) ? {add_181858, array_index_181536[0]} : sel_181860;
  assign add_181964 = array_index_181737[11:3] + 9'h0bd;
  assign sel_181967 = $signed({1'h0, add_181862, array_index_181635[2:0]}) < $signed({1'h0, sel_181865}) ? {add_181862, array_index_181635[2:0]} : sel_181865;
  assign add_181969 = array_index_181740[11:3] + 9'h0bd;
  assign sel_181972 = $signed({1'h0, add_181867, array_index_181638[2:0]}) < $signed({1'h0, sel_181870}) ? {add_181867, array_index_181638[2:0]} : sel_181870;
  assign add_181974 = array_index_181839[11:1] + 11'h247;
  assign sel_181977 = $signed({1'h0, add_181872, array_index_181737[0]}) < $signed({1'h0, sel_181875}) ? {add_181872, array_index_181737[0]} : sel_181875;
  assign add_181979 = array_index_181842[11:1] + 11'h247;
  assign sel_181982 = $signed({1'h0, add_181877, array_index_181740[0]}) < $signed({1'h0, sel_181880}) ? {add_181877, array_index_181740[0]} : sel_181880;
  assign add_182007 = array_index_181941[11:0] + 12'h247;
  assign sel_182009 = $signed({1'h0, add_181905}) < $signed({1'h0, sel_181907}) ? add_181905 : sel_181907;
  assign add_182012 = array_index_181944[11:0] + 12'h247;
  assign sel_182014 = $signed({1'h0, add_181910}) < $signed({1'h0, sel_181912}) ? add_181910 : sel_181912;
  assign array_index_182043 = set1_unflattened[7'h5c];
  assign array_index_182046 = set2_unflattened[7'h5c];
  assign add_182050 = array_index_181635[11:1] + 11'h79d;
  assign sel_182052 = $signed({1'h0, add_181948, array_index_181533[0]}) < $signed({1'h0, sel_181950}) ? {add_181948, array_index_181533[0]} : sel_181950;
  assign add_182054 = array_index_181638[11:1] + 11'h79d;
  assign sel_182056 = $signed({1'h0, add_181952, array_index_181536[0]}) < $signed({1'h0, sel_181954}) ? {add_181952, array_index_181536[0]} : sel_181954;
  assign add_182058 = array_index_181737[11:1] + 11'h347;
  assign sel_182060 = $signed({1'h0, add_181956, array_index_181635[0]}) < $signed({1'h0, sel_181958}) ? {add_181956, array_index_181635[0]} : sel_181958;
  assign add_182062 = array_index_181740[11:1] + 11'h347;
  assign sel_182064 = $signed({1'h0, add_181960, array_index_181638[0]}) < $signed({1'h0, sel_181962}) ? {add_181960, array_index_181638[0]} : sel_181962;
  assign add_182066 = array_index_181839[11:3] + 9'h0bd;
  assign sel_182069 = $signed({1'h0, add_181964, array_index_181737[2:0]}) < $signed({1'h0, sel_181967}) ? {add_181964, array_index_181737[2:0]} : sel_181967;
  assign add_182071 = array_index_181842[11:3] + 9'h0bd;
  assign sel_182074 = $signed({1'h0, add_181969, array_index_181740[2:0]}) < $signed({1'h0, sel_181972}) ? {add_181969, array_index_181740[2:0]} : sel_181972;
  assign add_182076 = array_index_181941[11:1] + 11'h247;
  assign sel_182079 = $signed({1'h0, add_181974, array_index_181839[0]}) < $signed({1'h0, sel_181977}) ? {add_181974, array_index_181839[0]} : sel_181977;
  assign add_182081 = array_index_181944[11:1] + 11'h247;
  assign sel_182084 = $signed({1'h0, add_181979, array_index_181842[0]}) < $signed({1'h0, sel_181982}) ? {add_181979, array_index_181842[0]} : sel_181982;
  assign add_182109 = array_index_182043[11:0] + 12'h247;
  assign sel_182111 = $signed({1'h0, add_182007}) < $signed({1'h0, sel_182009}) ? add_182007 : sel_182009;
  assign add_182114 = array_index_182046[11:0] + 12'h247;
  assign sel_182116 = $signed({1'h0, add_182012}) < $signed({1'h0, sel_182014}) ? add_182012 : sel_182014;
  assign array_index_182145 = set1_unflattened[7'h5d];
  assign array_index_182148 = set2_unflattened[7'h5d];
  assign add_182152 = array_index_181737[11:1] + 11'h79d;
  assign sel_182154 = $signed({1'h0, add_182050, array_index_181635[0]}) < $signed({1'h0, sel_182052}) ? {add_182050, array_index_181635[0]} : sel_182052;
  assign add_182156 = array_index_181740[11:1] + 11'h79d;
  assign sel_182158 = $signed({1'h0, add_182054, array_index_181638[0]}) < $signed({1'h0, sel_182056}) ? {add_182054, array_index_181638[0]} : sel_182056;
  assign add_182160 = array_index_181839[11:1] + 11'h347;
  assign sel_182162 = $signed({1'h0, add_182058, array_index_181737[0]}) < $signed({1'h0, sel_182060}) ? {add_182058, array_index_181737[0]} : sel_182060;
  assign add_182164 = array_index_181842[11:1] + 11'h347;
  assign sel_182166 = $signed({1'h0, add_182062, array_index_181740[0]}) < $signed({1'h0, sel_182064}) ? {add_182062, array_index_181740[0]} : sel_182064;
  assign add_182168 = array_index_181941[11:3] + 9'h0bd;
  assign sel_182171 = $signed({1'h0, add_182066, array_index_181839[2:0]}) < $signed({1'h0, sel_182069}) ? {add_182066, array_index_181839[2:0]} : sel_182069;
  assign add_182173 = array_index_181944[11:3] + 9'h0bd;
  assign sel_182176 = $signed({1'h0, add_182071, array_index_181842[2:0]}) < $signed({1'h0, sel_182074}) ? {add_182071, array_index_181842[2:0]} : sel_182074;
  assign add_182178 = array_index_182043[11:1] + 11'h247;
  assign sel_182181 = $signed({1'h0, add_182076, array_index_181941[0]}) < $signed({1'h0, sel_182079}) ? {add_182076, array_index_181941[0]} : sel_182079;
  assign add_182183 = array_index_182046[11:1] + 11'h247;
  assign sel_182186 = $signed({1'h0, add_182081, array_index_181944[0]}) < $signed({1'h0, sel_182084}) ? {add_182081, array_index_181944[0]} : sel_182084;
  assign add_182211 = array_index_182145[11:0] + 12'h247;
  assign sel_182213 = $signed({1'h0, add_182109}) < $signed({1'h0, sel_182111}) ? add_182109 : sel_182111;
  assign add_182216 = array_index_182148[11:0] + 12'h247;
  assign sel_182218 = $signed({1'h0, add_182114}) < $signed({1'h0, sel_182116}) ? add_182114 : sel_182116;
  assign array_index_182247 = set1_unflattened[7'h5e];
  assign array_index_182250 = set2_unflattened[7'h5e];
  assign add_182254 = array_index_181839[11:1] + 11'h79d;
  assign sel_182256 = $signed({1'h0, add_182152, array_index_181737[0]}) < $signed({1'h0, sel_182154}) ? {add_182152, array_index_181737[0]} : sel_182154;
  assign add_182258 = array_index_181842[11:1] + 11'h79d;
  assign sel_182260 = $signed({1'h0, add_182156, array_index_181740[0]}) < $signed({1'h0, sel_182158}) ? {add_182156, array_index_181740[0]} : sel_182158;
  assign add_182262 = array_index_181941[11:1] + 11'h347;
  assign sel_182264 = $signed({1'h0, add_182160, array_index_181839[0]}) < $signed({1'h0, sel_182162}) ? {add_182160, array_index_181839[0]} : sel_182162;
  assign add_182266 = array_index_181944[11:1] + 11'h347;
  assign sel_182268 = $signed({1'h0, add_182164, array_index_181842[0]}) < $signed({1'h0, sel_182166}) ? {add_182164, array_index_181842[0]} : sel_182166;
  assign add_182270 = array_index_182043[11:3] + 9'h0bd;
  assign sel_182273 = $signed({1'h0, add_182168, array_index_181941[2:0]}) < $signed({1'h0, sel_182171}) ? {add_182168, array_index_181941[2:0]} : sel_182171;
  assign add_182275 = array_index_182046[11:3] + 9'h0bd;
  assign sel_182278 = $signed({1'h0, add_182173, array_index_181944[2:0]}) < $signed({1'h0, sel_182176}) ? {add_182173, array_index_181944[2:0]} : sel_182176;
  assign add_182280 = array_index_182145[11:1] + 11'h247;
  assign sel_182283 = $signed({1'h0, add_182178, array_index_182043[0]}) < $signed({1'h0, sel_182181}) ? {add_182178, array_index_182043[0]} : sel_182181;
  assign add_182285 = array_index_182148[11:1] + 11'h247;
  assign sel_182288 = $signed({1'h0, add_182183, array_index_182046[0]}) < $signed({1'h0, sel_182186}) ? {add_182183, array_index_182046[0]} : sel_182186;
  assign add_182313 = array_index_182247[11:0] + 12'h247;
  assign sel_182315 = $signed({1'h0, add_182211}) < $signed({1'h0, sel_182213}) ? add_182211 : sel_182213;
  assign add_182318 = array_index_182250[11:0] + 12'h247;
  assign sel_182320 = $signed({1'h0, add_182216}) < $signed({1'h0, sel_182218}) ? add_182216 : sel_182218;
  assign array_index_182349 = set1_unflattened[7'h5f];
  assign array_index_182352 = set2_unflattened[7'h5f];
  assign add_182356 = array_index_181941[11:1] + 11'h79d;
  assign sel_182358 = $signed({1'h0, add_182254, array_index_181839[0]}) < $signed({1'h0, sel_182256}) ? {add_182254, array_index_181839[0]} : sel_182256;
  assign add_182360 = array_index_181944[11:1] + 11'h79d;
  assign sel_182362 = $signed({1'h0, add_182258, array_index_181842[0]}) < $signed({1'h0, sel_182260}) ? {add_182258, array_index_181842[0]} : sel_182260;
  assign add_182364 = array_index_182043[11:1] + 11'h347;
  assign sel_182366 = $signed({1'h0, add_182262, array_index_181941[0]}) < $signed({1'h0, sel_182264}) ? {add_182262, array_index_181941[0]} : sel_182264;
  assign add_182368 = array_index_182046[11:1] + 11'h347;
  assign sel_182370 = $signed({1'h0, add_182266, array_index_181944[0]}) < $signed({1'h0, sel_182268}) ? {add_182266, array_index_181944[0]} : sel_182268;
  assign add_182372 = array_index_182145[11:3] + 9'h0bd;
  assign sel_182375 = $signed({1'h0, add_182270, array_index_182043[2:0]}) < $signed({1'h0, sel_182273}) ? {add_182270, array_index_182043[2:0]} : sel_182273;
  assign add_182377 = array_index_182148[11:3] + 9'h0bd;
  assign sel_182380 = $signed({1'h0, add_182275, array_index_182046[2:0]}) < $signed({1'h0, sel_182278}) ? {add_182275, array_index_182046[2:0]} : sel_182278;
  assign add_182382 = array_index_182247[11:1] + 11'h247;
  assign sel_182385 = $signed({1'h0, add_182280, array_index_182145[0]}) < $signed({1'h0, sel_182283}) ? {add_182280, array_index_182145[0]} : sel_182283;
  assign add_182387 = array_index_182250[11:1] + 11'h247;
  assign sel_182390 = $signed({1'h0, add_182285, array_index_182148[0]}) < $signed({1'h0, sel_182288}) ? {add_182285, array_index_182148[0]} : sel_182288;
  assign add_182415 = array_index_182349[11:0] + 12'h247;
  assign sel_182417 = $signed({1'h0, add_182313}) < $signed({1'h0, sel_182315}) ? add_182313 : sel_182315;
  assign add_182420 = array_index_182352[11:0] + 12'h247;
  assign sel_182422 = $signed({1'h0, add_182318}) < $signed({1'h0, sel_182320}) ? add_182318 : sel_182320;
  assign array_index_182451 = set1_unflattened[7'h60];
  assign array_index_182454 = set2_unflattened[7'h60];
  assign add_182458 = array_index_182043[11:1] + 11'h79d;
  assign sel_182460 = $signed({1'h0, add_182356, array_index_181941[0]}) < $signed({1'h0, sel_182358}) ? {add_182356, array_index_181941[0]} : sel_182358;
  assign add_182462 = array_index_182046[11:1] + 11'h79d;
  assign sel_182464 = $signed({1'h0, add_182360, array_index_181944[0]}) < $signed({1'h0, sel_182362}) ? {add_182360, array_index_181944[0]} : sel_182362;
  assign add_182466 = array_index_182145[11:1] + 11'h347;
  assign sel_182468 = $signed({1'h0, add_182364, array_index_182043[0]}) < $signed({1'h0, sel_182366}) ? {add_182364, array_index_182043[0]} : sel_182366;
  assign add_182470 = array_index_182148[11:1] + 11'h347;
  assign sel_182472 = $signed({1'h0, add_182368, array_index_182046[0]}) < $signed({1'h0, sel_182370}) ? {add_182368, array_index_182046[0]} : sel_182370;
  assign add_182474 = array_index_182247[11:3] + 9'h0bd;
  assign sel_182477 = $signed({1'h0, add_182372, array_index_182145[2:0]}) < $signed({1'h0, sel_182375}) ? {add_182372, array_index_182145[2:0]} : sel_182375;
  assign add_182479 = array_index_182250[11:3] + 9'h0bd;
  assign sel_182482 = $signed({1'h0, add_182377, array_index_182148[2:0]}) < $signed({1'h0, sel_182380}) ? {add_182377, array_index_182148[2:0]} : sel_182380;
  assign add_182484 = array_index_182349[11:1] + 11'h247;
  assign sel_182487 = $signed({1'h0, add_182382, array_index_182247[0]}) < $signed({1'h0, sel_182385}) ? {add_182382, array_index_182247[0]} : sel_182385;
  assign add_182489 = array_index_182352[11:1] + 11'h247;
  assign sel_182492 = $signed({1'h0, add_182387, array_index_182250[0]}) < $signed({1'h0, sel_182390}) ? {add_182387, array_index_182250[0]} : sel_182390;
  assign add_182517 = array_index_182451[11:0] + 12'h247;
  assign sel_182519 = $signed({1'h0, add_182415}) < $signed({1'h0, sel_182417}) ? add_182415 : sel_182417;
  assign add_182522 = array_index_182454[11:0] + 12'h247;
  assign sel_182524 = $signed({1'h0, add_182420}) < $signed({1'h0, sel_182422}) ? add_182420 : sel_182422;
  assign array_index_182553 = set1_unflattened[7'h61];
  assign array_index_182556 = set2_unflattened[7'h61];
  assign add_182560 = array_index_182145[11:1] + 11'h79d;
  assign sel_182562 = $signed({1'h0, add_182458, array_index_182043[0]}) < $signed({1'h0, sel_182460}) ? {add_182458, array_index_182043[0]} : sel_182460;
  assign add_182564 = array_index_182148[11:1] + 11'h79d;
  assign sel_182566 = $signed({1'h0, add_182462, array_index_182046[0]}) < $signed({1'h0, sel_182464}) ? {add_182462, array_index_182046[0]} : sel_182464;
  assign add_182568 = array_index_182247[11:1] + 11'h347;
  assign sel_182570 = $signed({1'h0, add_182466, array_index_182145[0]}) < $signed({1'h0, sel_182468}) ? {add_182466, array_index_182145[0]} : sel_182468;
  assign add_182572 = array_index_182250[11:1] + 11'h347;
  assign sel_182574 = $signed({1'h0, add_182470, array_index_182148[0]}) < $signed({1'h0, sel_182472}) ? {add_182470, array_index_182148[0]} : sel_182472;
  assign add_182576 = array_index_182349[11:3] + 9'h0bd;
  assign sel_182579 = $signed({1'h0, add_182474, array_index_182247[2:0]}) < $signed({1'h0, sel_182477}) ? {add_182474, array_index_182247[2:0]} : sel_182477;
  assign add_182581 = array_index_182352[11:3] + 9'h0bd;
  assign sel_182584 = $signed({1'h0, add_182479, array_index_182250[2:0]}) < $signed({1'h0, sel_182482}) ? {add_182479, array_index_182250[2:0]} : sel_182482;
  assign add_182586 = array_index_182451[11:1] + 11'h247;
  assign sel_182589 = $signed({1'h0, add_182484, array_index_182349[0]}) < $signed({1'h0, sel_182487}) ? {add_182484, array_index_182349[0]} : sel_182487;
  assign add_182591 = array_index_182454[11:1] + 11'h247;
  assign sel_182594 = $signed({1'h0, add_182489, array_index_182352[0]}) < $signed({1'h0, sel_182492}) ? {add_182489, array_index_182352[0]} : sel_182492;
  assign add_182619 = array_index_182553[11:0] + 12'h247;
  assign sel_182621 = $signed({1'h0, add_182517}) < $signed({1'h0, sel_182519}) ? add_182517 : sel_182519;
  assign add_182624 = array_index_182556[11:0] + 12'h247;
  assign sel_182626 = $signed({1'h0, add_182522}) < $signed({1'h0, sel_182524}) ? add_182522 : sel_182524;
  assign array_index_182655 = set1_unflattened[7'h62];
  assign array_index_182658 = set2_unflattened[7'h62];
  assign add_182662 = array_index_182247[11:1] + 11'h79d;
  assign sel_182664 = $signed({1'h0, add_182560, array_index_182145[0]}) < $signed({1'h0, sel_182562}) ? {add_182560, array_index_182145[0]} : sel_182562;
  assign add_182666 = array_index_182250[11:1] + 11'h79d;
  assign sel_182668 = $signed({1'h0, add_182564, array_index_182148[0]}) < $signed({1'h0, sel_182566}) ? {add_182564, array_index_182148[0]} : sel_182566;
  assign add_182670 = array_index_182349[11:1] + 11'h347;
  assign sel_182672 = $signed({1'h0, add_182568, array_index_182247[0]}) < $signed({1'h0, sel_182570}) ? {add_182568, array_index_182247[0]} : sel_182570;
  assign add_182674 = array_index_182352[11:1] + 11'h347;
  assign sel_182676 = $signed({1'h0, add_182572, array_index_182250[0]}) < $signed({1'h0, sel_182574}) ? {add_182572, array_index_182250[0]} : sel_182574;
  assign add_182678 = array_index_182451[11:3] + 9'h0bd;
  assign sel_182681 = $signed({1'h0, add_182576, array_index_182349[2:0]}) < $signed({1'h0, sel_182579}) ? {add_182576, array_index_182349[2:0]} : sel_182579;
  assign add_182683 = array_index_182454[11:3] + 9'h0bd;
  assign sel_182686 = $signed({1'h0, add_182581, array_index_182352[2:0]}) < $signed({1'h0, sel_182584}) ? {add_182581, array_index_182352[2:0]} : sel_182584;
  assign add_182688 = array_index_182553[11:1] + 11'h247;
  assign sel_182691 = $signed({1'h0, add_182586, array_index_182451[0]}) < $signed({1'h0, sel_182589}) ? {add_182586, array_index_182451[0]} : sel_182589;
  assign add_182693 = array_index_182556[11:1] + 11'h247;
  assign sel_182696 = $signed({1'h0, add_182591, array_index_182454[0]}) < $signed({1'h0, sel_182594}) ? {add_182591, array_index_182454[0]} : sel_182594;
  assign add_182721 = array_index_182655[11:0] + 12'h247;
  assign sel_182723 = $signed({1'h0, add_182619}) < $signed({1'h0, sel_182621}) ? add_182619 : sel_182621;
  assign add_182726 = array_index_182658[11:0] + 12'h247;
  assign sel_182728 = $signed({1'h0, add_182624}) < $signed({1'h0, sel_182626}) ? add_182624 : sel_182626;
  assign array_index_182757 = set1_unflattened[7'h63];
  assign array_index_182760 = set2_unflattened[7'h63];
  assign add_182764 = array_index_182349[11:1] + 11'h79d;
  assign sel_182766 = $signed({1'h0, add_182662, array_index_182247[0]}) < $signed({1'h0, sel_182664}) ? {add_182662, array_index_182247[0]} : sel_182664;
  assign add_182768 = array_index_182352[11:1] + 11'h79d;
  assign sel_182770 = $signed({1'h0, add_182666, array_index_182250[0]}) < $signed({1'h0, sel_182668}) ? {add_182666, array_index_182250[0]} : sel_182668;
  assign add_182772 = array_index_182451[11:1] + 11'h347;
  assign sel_182774 = $signed({1'h0, add_182670, array_index_182349[0]}) < $signed({1'h0, sel_182672}) ? {add_182670, array_index_182349[0]} : sel_182672;
  assign add_182776 = array_index_182454[11:1] + 11'h347;
  assign sel_182778 = $signed({1'h0, add_182674, array_index_182352[0]}) < $signed({1'h0, sel_182676}) ? {add_182674, array_index_182352[0]} : sel_182676;
  assign add_182780 = array_index_182553[11:3] + 9'h0bd;
  assign sel_182783 = $signed({1'h0, add_182678, array_index_182451[2:0]}) < $signed({1'h0, sel_182681}) ? {add_182678, array_index_182451[2:0]} : sel_182681;
  assign add_182785 = array_index_182556[11:3] + 9'h0bd;
  assign sel_182788 = $signed({1'h0, add_182683, array_index_182454[2:0]}) < $signed({1'h0, sel_182686}) ? {add_182683, array_index_182454[2:0]} : sel_182686;
  assign add_182790 = array_index_182655[11:1] + 11'h247;
  assign sel_182793 = $signed({1'h0, add_182688, array_index_182553[0]}) < $signed({1'h0, sel_182691}) ? {add_182688, array_index_182553[0]} : sel_182691;
  assign add_182795 = array_index_182658[11:1] + 11'h247;
  assign sel_182798 = $signed({1'h0, add_182693, array_index_182556[0]}) < $signed({1'h0, sel_182696}) ? {add_182693, array_index_182556[0]} : sel_182696;
  assign add_182822 = array_index_182757[11:0] + 12'h247;
  assign sel_182824 = $signed({1'h0, add_182721}) < $signed({1'h0, sel_182723}) ? add_182721 : sel_182723;
  assign add_182826 = array_index_182760[11:0] + 12'h247;
  assign sel_182828 = $signed({1'h0, add_182726}) < $signed({1'h0, sel_182728}) ? add_182726 : sel_182728;
  assign add_182862 = array_index_182451[11:1] + 11'h79d;
  assign sel_182864 = $signed({1'h0, add_182764, array_index_182349[0]}) < $signed({1'h0, sel_182766}) ? {add_182764, array_index_182349[0]} : sel_182766;
  assign add_182866 = array_index_182454[11:1] + 11'h79d;
  assign sel_182868 = $signed({1'h0, add_182768, array_index_182352[0]}) < $signed({1'h0, sel_182770}) ? {add_182768, array_index_182352[0]} : sel_182770;
  assign add_182870 = array_index_182553[11:1] + 11'h347;
  assign sel_182872 = $signed({1'h0, add_182772, array_index_182451[0]}) < $signed({1'h0, sel_182774}) ? {add_182772, array_index_182451[0]} : sel_182774;
  assign add_182874 = array_index_182556[11:1] + 11'h347;
  assign sel_182876 = $signed({1'h0, add_182776, array_index_182454[0]}) < $signed({1'h0, sel_182778}) ? {add_182776, array_index_182454[0]} : sel_182778;
  assign add_182878 = array_index_182655[11:3] + 9'h0bd;
  assign sel_182881 = $signed({1'h0, add_182780, array_index_182553[2:0]}) < $signed({1'h0, sel_182783}) ? {add_182780, array_index_182553[2:0]} : sel_182783;
  assign add_182883 = array_index_182658[11:3] + 9'h0bd;
  assign sel_182886 = $signed({1'h0, add_182785, array_index_182556[2:0]}) < $signed({1'h0, sel_182788}) ? {add_182785, array_index_182556[2:0]} : sel_182788;
  assign add_182888 = array_index_182757[11:1] + 11'h247;
  assign sel_182891 = $signed({1'h0, add_182790, array_index_182655[0]}) < $signed({1'h0, sel_182793}) ? {add_182790, array_index_182655[0]} : sel_182793;
  assign add_182893 = array_index_182760[11:1] + 11'h247;
  assign sel_182896 = $signed({1'h0, add_182795, array_index_182658[0]}) < $signed({1'h0, sel_182798}) ? {add_182795, array_index_182658[0]} : sel_182798;
  assign add_182944 = array_index_182553[11:1] + 11'h79d;
  assign sel_182946 = $signed({1'h0, add_182862, array_index_182451[0]}) < $signed({1'h0, sel_182864}) ? {add_182862, array_index_182451[0]} : sel_182864;
  assign add_182948 = array_index_182556[11:1] + 11'h79d;
  assign sel_182950 = $signed({1'h0, add_182866, array_index_182454[0]}) < $signed({1'h0, sel_182868}) ? {add_182866, array_index_182454[0]} : sel_182868;
  assign add_182952 = array_index_182655[11:1] + 11'h347;
  assign sel_182954 = $signed({1'h0, add_182870, array_index_182553[0]}) < $signed({1'h0, sel_182872}) ? {add_182870, array_index_182553[0]} : sel_182872;
  assign add_182956 = array_index_182658[11:1] + 11'h347;
  assign sel_182958 = $signed({1'h0, add_182874, array_index_182556[0]}) < $signed({1'h0, sel_182876}) ? {add_182874, array_index_182556[0]} : sel_182876;
  assign add_182960 = array_index_182757[11:3] + 9'h0bd;
  assign sel_182963 = $signed({1'h0, add_182878, array_index_182655[2:0]}) < $signed({1'h0, sel_182881}) ? {add_182878, array_index_182655[2:0]} : sel_182881;
  assign add_182965 = array_index_182760[11:3] + 9'h0bd;
  assign sel_182968 = $signed({1'h0, add_182883, array_index_182658[2:0]}) < $signed({1'h0, sel_182886}) ? {add_182883, array_index_182658[2:0]} : sel_182886;
  assign concat_182971 = {1'h0, ($signed({1'h0, add_182822}) < $signed({1'h0, sel_182824}) ? add_182822 : sel_182824) == ($signed({1'h0, add_182826}) < $signed({1'h0, sel_182828}) ? add_182826 : sel_182828)};
  assign add_182986 = concat_182971 + 2'h1;
  assign add_183006 = array_index_182655[11:1] + 11'h79d;
  assign sel_183008 = $signed({1'h0, add_182944, array_index_182553[0]}) < $signed({1'h0, sel_182946}) ? {add_182944, array_index_182553[0]} : sel_182946;
  assign add_183010 = array_index_182658[11:1] + 11'h79d;
  assign sel_183012 = $signed({1'h0, add_182948, array_index_182556[0]}) < $signed({1'h0, sel_182950}) ? {add_182948, array_index_182556[0]} : sel_182950;
  assign add_183014 = array_index_182757[11:1] + 11'h347;
  assign sel_183016 = $signed({1'h0, add_182952, array_index_182655[0]}) < $signed({1'h0, sel_182954}) ? {add_182952, array_index_182655[0]} : sel_182954;
  assign add_183018 = array_index_182760[11:1] + 11'h347;
  assign sel_183020 = $signed({1'h0, add_182956, array_index_182658[0]}) < $signed({1'h0, sel_182958}) ? {add_182956, array_index_182658[0]} : sel_182958;
  assign concat_183023 = {1'h0, ($signed({1'h0, add_182888, array_index_182757[0]}) < $signed({1'h0, sel_182891}) ? {add_182888, array_index_182757[0]} : sel_182891) == ($signed({1'h0, add_182893, array_index_182760[0]}) < $signed({1'h0, sel_182896}) ? {add_182893, array_index_182760[0]} : sel_182896) ? add_182986 : concat_182971};
  assign add_183034 = concat_183023 + 3'h1;
  assign add_183048 = array_index_182757[11:1] + 11'h79d;
  assign sel_183050 = $signed({1'h0, add_183006, array_index_182655[0]}) < $signed({1'h0, sel_183008}) ? {add_183006, array_index_182655[0]} : sel_183008;
  assign add_183052 = array_index_182760[11:1] + 11'h79d;
  assign sel_183054 = $signed({1'h0, add_183010, array_index_182658[0]}) < $signed({1'h0, sel_183012}) ? {add_183010, array_index_182658[0]} : sel_183012;
  assign concat_183057 = {1'h0, ($signed({1'h0, add_182960, array_index_182757[2:0]}) < $signed({1'h0, sel_182963}) ? {add_182960, array_index_182757[2:0]} : sel_182963) == ($signed({1'h0, add_182965, array_index_182760[2:0]}) < $signed({1'h0, sel_182968}) ? {add_182965, array_index_182760[2:0]} : sel_182968) ? add_183034 : concat_183023};
  assign add_183064 = concat_183057 + 4'h1;
  assign concat_183073 = {1'h0, ($signed({1'h0, add_183014, array_index_182757[0]}) < $signed({1'h0, sel_183016}) ? {add_183014, array_index_182757[0]} : sel_183016) == ($signed({1'h0, add_183018, array_index_182760[0]}) < $signed({1'h0, sel_183020}) ? {add_183018, array_index_182760[0]} : sel_183020) ? add_183064 : concat_183057};
  assign add_183076 = concat_183073 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_183048, array_index_182757[0]}) < $signed({1'h0, sel_183050}) ? {add_183048, array_index_182757[0]} : sel_183050) == ($signed({1'h0, add_183052, array_index_182760[0]}) < $signed({1'h0, sel_183054}) ? {add_183052, array_index_182760[0]} : sel_183054) ? add_183076 : concat_183073}, {set1_unflattened[99], set1_unflattened[98], set1_unflattened[97], set1_unflattened[96], set1_unflattened[95], set1_unflattened[94], set1_unflattened[93], set1_unflattened[92], set1_unflattened[91], set1_unflattened[90], set1_unflattened[89], set1_unflattened[88], set1_unflattened[87], set1_unflattened[86], set1_unflattened[85], set1_unflattened[84], set1_unflattened[83], set1_unflattened[82], set1_unflattened[81], set1_unflattened[80], set1_unflattened[79], set1_unflattened[78], set1_unflattened[77], set1_unflattened[76], set1_unflattened[75], set1_unflattened[74], set1_unflattened[73], set1_unflattened[72], set1_unflattened[71], set1_unflattened[70], set1_unflattened[69], set1_unflattened[68], set1_unflattened[67], set1_unflattened[66], set1_unflattened[65], set1_unflattened[64], set1_unflattened[63], set1_unflattened[62], set1_unflattened[61], set1_unflattened[60], set1_unflattened[59], set1_unflattened[58], set1_unflattened[57], set1_unflattened[56], set1_unflattened[55], set1_unflattened[54], set1_unflattened[53], set1_unflattened[52], set1_unflattened[51], set1_unflattened[50], set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[99], set2_unflattened[98], set2_unflattened[97], set2_unflattened[96], set2_unflattened[95], set2_unflattened[94], set2_unflattened[93], set2_unflattened[92], set2_unflattened[91], set2_unflattened[90], set2_unflattened[89], set2_unflattened[88], set2_unflattened[87], set2_unflattened[86], set2_unflattened[85], set2_unflattened[84], set2_unflattened[83], set2_unflattened[82], set2_unflattened[81], set2_unflattened[80], set2_unflattened[79], set2_unflattened[78], set2_unflattened[77], set2_unflattened[76], set2_unflattened[75], set2_unflattened[74], set2_unflattened[73], set2_unflattened[72], set2_unflattened[71], set2_unflattened[70], set2_unflattened[69], set2_unflattened[68], set2_unflattened[67], set2_unflattened[66], set2_unflattened[65], set2_unflattened[64], set2_unflattened[63], set2_unflattened[62], set2_unflattened[61], set2_unflattened[60], set2_unflattened[59], set2_unflattened[58], set2_unflattened[57], set2_unflattened[56], set2_unflattened[55], set2_unflattened[54], set2_unflattened[53], set2_unflattened[52], set2_unflattened[51], set2_unflattened[50], set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
